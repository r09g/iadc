magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< error_p >>
rect -994 607 -936 887
rect -816 607 -758 887
rect -702 607 -644 887
rect -524 607 -466 887
rect -410 607 -352 887
rect -232 607 -174 887
rect -118 607 -60 887
rect 60 607 118 887
rect 174 607 232 887
rect 352 607 410 887
rect 466 607 524 887
rect 644 607 702 887
rect 758 607 816 887
rect 936 607 994 887
rect -994 109 -936 389
rect -816 109 -758 389
rect -702 109 -644 389
rect -524 109 -466 389
rect -410 109 -352 389
rect -232 109 -174 389
rect -118 109 -60 389
rect 60 109 118 389
rect 174 109 232 389
rect 352 109 410 389
rect 466 109 524 389
rect 644 109 702 389
rect 758 109 816 389
rect 936 109 994 389
rect -994 -389 -936 -109
rect -816 -389 -758 -109
rect -702 -389 -644 -109
rect -524 -389 -466 -109
rect -410 -389 -352 -109
rect -232 -389 -174 -109
rect -118 -389 -60 -109
rect 60 -389 118 -109
rect 174 -389 232 -109
rect 352 -389 410 -109
rect 466 -389 524 -109
rect 644 -389 702 -109
rect 758 -389 816 -109
rect 936 -389 994 -109
rect -994 -887 -936 -607
rect -816 -887 -758 -607
rect -702 -887 -644 -607
rect -524 -887 -466 -607
rect -410 -887 -352 -607
rect -232 -887 -174 -607
rect -118 -887 -60 -607
rect 60 -887 118 -607
rect 174 -887 232 -607
rect 352 -887 410 -607
rect 466 -887 524 -607
rect 644 -887 702 -607
rect 758 -887 816 -607
rect 936 -887 994 -607
<< nmos >>
rect -936 607 -816 887
rect -644 607 -524 887
rect -352 607 -232 887
rect -60 607 60 887
rect 232 607 352 887
rect 524 607 644 887
rect 816 607 936 887
rect -936 109 -816 389
rect -644 109 -524 389
rect -352 109 -232 389
rect -60 109 60 389
rect 232 109 352 389
rect 524 109 644 389
rect 816 109 936 389
rect -936 -389 -816 -109
rect -644 -389 -524 -109
rect -352 -389 -232 -109
rect -60 -389 60 -109
rect 232 -389 352 -109
rect 524 -389 644 -109
rect 816 -389 936 -109
rect -936 -887 -816 -607
rect -644 -887 -524 -607
rect -352 -887 -232 -607
rect -60 -887 60 -607
rect 232 -887 352 -607
rect 524 -887 644 -607
rect 816 -887 936 -607
<< ndiff >>
rect -994 875 -936 887
rect -994 619 -982 875
rect -948 619 -936 875
rect -994 607 -936 619
rect -816 875 -758 887
rect -816 619 -804 875
rect -770 619 -758 875
rect -816 607 -758 619
rect -702 875 -644 887
rect -702 619 -690 875
rect -656 619 -644 875
rect -702 607 -644 619
rect -524 875 -466 887
rect -524 619 -512 875
rect -478 619 -466 875
rect -524 607 -466 619
rect -410 875 -352 887
rect -410 619 -398 875
rect -364 619 -352 875
rect -410 607 -352 619
rect -232 875 -174 887
rect -232 619 -220 875
rect -186 619 -174 875
rect -232 607 -174 619
rect -118 875 -60 887
rect -118 619 -106 875
rect -72 619 -60 875
rect -118 607 -60 619
rect 60 875 118 887
rect 60 619 72 875
rect 106 619 118 875
rect 60 607 118 619
rect 174 875 232 887
rect 174 619 186 875
rect 220 619 232 875
rect 174 607 232 619
rect 352 875 410 887
rect 352 619 364 875
rect 398 619 410 875
rect 352 607 410 619
rect 466 875 524 887
rect 466 619 478 875
rect 512 619 524 875
rect 466 607 524 619
rect 644 875 702 887
rect 644 619 656 875
rect 690 619 702 875
rect 644 607 702 619
rect 758 875 816 887
rect 758 619 770 875
rect 804 619 816 875
rect 758 607 816 619
rect 936 875 994 887
rect 936 619 948 875
rect 982 619 994 875
rect 936 607 994 619
rect -994 377 -936 389
rect -994 121 -982 377
rect -948 121 -936 377
rect -994 109 -936 121
rect -816 377 -758 389
rect -816 121 -804 377
rect -770 121 -758 377
rect -816 109 -758 121
rect -702 377 -644 389
rect -702 121 -690 377
rect -656 121 -644 377
rect -702 109 -644 121
rect -524 377 -466 389
rect -524 121 -512 377
rect -478 121 -466 377
rect -524 109 -466 121
rect -410 377 -352 389
rect -410 121 -398 377
rect -364 121 -352 377
rect -410 109 -352 121
rect -232 377 -174 389
rect -232 121 -220 377
rect -186 121 -174 377
rect -232 109 -174 121
rect -118 377 -60 389
rect -118 121 -106 377
rect -72 121 -60 377
rect -118 109 -60 121
rect 60 377 118 389
rect 60 121 72 377
rect 106 121 118 377
rect 60 109 118 121
rect 174 377 232 389
rect 174 121 186 377
rect 220 121 232 377
rect 174 109 232 121
rect 352 377 410 389
rect 352 121 364 377
rect 398 121 410 377
rect 352 109 410 121
rect 466 377 524 389
rect 466 121 478 377
rect 512 121 524 377
rect 466 109 524 121
rect 644 377 702 389
rect 644 121 656 377
rect 690 121 702 377
rect 644 109 702 121
rect 758 377 816 389
rect 758 121 770 377
rect 804 121 816 377
rect 758 109 816 121
rect 936 377 994 389
rect 936 121 948 377
rect 982 121 994 377
rect 936 109 994 121
rect -994 -121 -936 -109
rect -994 -377 -982 -121
rect -948 -377 -936 -121
rect -994 -389 -936 -377
rect -816 -121 -758 -109
rect -816 -377 -804 -121
rect -770 -377 -758 -121
rect -816 -389 -758 -377
rect -702 -121 -644 -109
rect -702 -377 -690 -121
rect -656 -377 -644 -121
rect -702 -389 -644 -377
rect -524 -121 -466 -109
rect -524 -377 -512 -121
rect -478 -377 -466 -121
rect -524 -389 -466 -377
rect -410 -121 -352 -109
rect -410 -377 -398 -121
rect -364 -377 -352 -121
rect -410 -389 -352 -377
rect -232 -121 -174 -109
rect -232 -377 -220 -121
rect -186 -377 -174 -121
rect -232 -389 -174 -377
rect -118 -121 -60 -109
rect -118 -377 -106 -121
rect -72 -377 -60 -121
rect -118 -389 -60 -377
rect 60 -121 118 -109
rect 60 -377 72 -121
rect 106 -377 118 -121
rect 60 -389 118 -377
rect 174 -121 232 -109
rect 174 -377 186 -121
rect 220 -377 232 -121
rect 174 -389 232 -377
rect 352 -121 410 -109
rect 352 -377 364 -121
rect 398 -377 410 -121
rect 352 -389 410 -377
rect 466 -121 524 -109
rect 466 -377 478 -121
rect 512 -377 524 -121
rect 466 -389 524 -377
rect 644 -121 702 -109
rect 644 -377 656 -121
rect 690 -377 702 -121
rect 644 -389 702 -377
rect 758 -121 816 -109
rect 758 -377 770 -121
rect 804 -377 816 -121
rect 758 -389 816 -377
rect 936 -121 994 -109
rect 936 -377 948 -121
rect 982 -377 994 -121
rect 936 -389 994 -377
rect -994 -619 -936 -607
rect -994 -875 -982 -619
rect -948 -875 -936 -619
rect -994 -887 -936 -875
rect -816 -619 -758 -607
rect -816 -875 -804 -619
rect -770 -875 -758 -619
rect -816 -887 -758 -875
rect -702 -619 -644 -607
rect -702 -875 -690 -619
rect -656 -875 -644 -619
rect -702 -887 -644 -875
rect -524 -619 -466 -607
rect -524 -875 -512 -619
rect -478 -875 -466 -619
rect -524 -887 -466 -875
rect -410 -619 -352 -607
rect -410 -875 -398 -619
rect -364 -875 -352 -619
rect -410 -887 -352 -875
rect -232 -619 -174 -607
rect -232 -875 -220 -619
rect -186 -875 -174 -619
rect -232 -887 -174 -875
rect -118 -619 -60 -607
rect -118 -875 -106 -619
rect -72 -875 -60 -619
rect -118 -887 -60 -875
rect 60 -619 118 -607
rect 60 -875 72 -619
rect 106 -875 118 -619
rect 60 -887 118 -875
rect 174 -619 232 -607
rect 174 -875 186 -619
rect 220 -875 232 -619
rect 174 -887 232 -875
rect 352 -619 410 -607
rect 352 -875 364 -619
rect 398 -875 410 -619
rect 352 -887 410 -875
rect 466 -619 524 -607
rect 466 -875 478 -619
rect 512 -875 524 -619
rect 466 -887 524 -875
rect 644 -619 702 -607
rect 644 -875 656 -619
rect 690 -875 702 -619
rect 644 -887 702 -875
rect 758 -619 816 -607
rect 758 -875 770 -619
rect 804 -875 816 -619
rect 758 -887 816 -875
rect 936 -619 994 -607
rect 936 -875 948 -619
rect 982 -875 994 -619
rect 936 -887 994 -875
<< ndiffc >>
rect -982 619 -948 875
rect -804 619 -770 875
rect -690 619 -656 875
rect -512 619 -478 875
rect -398 619 -364 875
rect -220 619 -186 875
rect -106 619 -72 875
rect 72 619 106 875
rect 186 619 220 875
rect 364 619 398 875
rect 478 619 512 875
rect 656 619 690 875
rect 770 619 804 875
rect 948 619 982 875
rect -982 121 -948 377
rect -804 121 -770 377
rect -690 121 -656 377
rect -512 121 -478 377
rect -398 121 -364 377
rect -220 121 -186 377
rect -106 121 -72 377
rect 72 121 106 377
rect 186 121 220 377
rect 364 121 398 377
rect 478 121 512 377
rect 656 121 690 377
rect 770 121 804 377
rect 948 121 982 377
rect -982 -377 -948 -121
rect -804 -377 -770 -121
rect -690 -377 -656 -121
rect -512 -377 -478 -121
rect -398 -377 -364 -121
rect -220 -377 -186 -121
rect -106 -377 -72 -121
rect 72 -377 106 -121
rect 186 -377 220 -121
rect 364 -377 398 -121
rect 478 -377 512 -121
rect 656 -377 690 -121
rect 770 -377 804 -121
rect 948 -377 982 -121
rect -982 -875 -948 -619
rect -804 -875 -770 -619
rect -690 -875 -656 -619
rect -512 -875 -478 -619
rect -398 -875 -364 -619
rect -220 -875 -186 -619
rect -106 -875 -72 -619
rect 72 -875 106 -619
rect 186 -875 220 -619
rect 364 -875 398 -619
rect 478 -875 512 -619
rect 656 -875 690 -619
rect 770 -875 804 -619
rect 948 -875 982 -619
<< poly >>
rect -918 959 -834 975
rect -918 943 -902 959
rect -936 925 -902 943
rect -850 943 -834 959
rect -626 959 -542 975
rect -626 943 -610 959
rect -850 925 -816 943
rect -936 887 -816 925
rect -644 925 -610 943
rect -558 943 -542 959
rect -334 959 -250 975
rect -334 943 -318 959
rect -558 925 -524 943
rect -644 887 -524 925
rect -352 925 -318 943
rect -266 943 -250 959
rect -42 959 42 975
rect -42 943 -26 959
rect -266 925 -232 943
rect -352 887 -232 925
rect -60 925 -26 943
rect 26 943 42 959
rect 250 959 334 975
rect 250 943 266 959
rect 26 925 60 943
rect -60 887 60 925
rect 232 925 266 943
rect 318 943 334 959
rect 542 959 626 975
rect 542 943 558 959
rect 318 925 352 943
rect 232 887 352 925
rect 524 925 558 943
rect 610 943 626 959
rect 834 959 918 975
rect 834 943 850 959
rect 610 925 644 943
rect 524 887 644 925
rect 816 925 850 943
rect 902 943 918 959
rect 902 925 936 943
rect 816 887 936 925
rect -936 569 -816 607
rect -936 553 -902 569
rect -918 535 -902 553
rect -850 553 -816 569
rect -644 569 -524 607
rect -644 553 -610 569
rect -850 535 -834 553
rect -918 519 -834 535
rect -626 535 -610 553
rect -558 553 -524 569
rect -352 569 -232 607
rect -352 553 -318 569
rect -558 535 -542 553
rect -626 519 -542 535
rect -334 535 -318 553
rect -266 553 -232 569
rect -60 569 60 607
rect -60 553 -26 569
rect -266 535 -250 553
rect -334 519 -250 535
rect -42 535 -26 553
rect 26 553 60 569
rect 232 569 352 607
rect 232 553 266 569
rect 26 535 42 553
rect -42 519 42 535
rect 250 535 266 553
rect 318 553 352 569
rect 524 569 644 607
rect 524 553 558 569
rect 318 535 334 553
rect 250 519 334 535
rect 542 535 558 553
rect 610 553 644 569
rect 816 569 936 607
rect 816 553 850 569
rect 610 535 626 553
rect 542 519 626 535
rect 834 535 850 553
rect 902 553 936 569
rect 902 535 918 553
rect 834 519 918 535
rect -918 461 -834 477
rect -918 445 -902 461
rect -936 427 -902 445
rect -850 445 -834 461
rect -626 461 -542 477
rect -626 445 -610 461
rect -850 427 -816 445
rect -936 389 -816 427
rect -644 427 -610 445
rect -558 445 -542 461
rect -334 461 -250 477
rect -334 445 -318 461
rect -558 427 -524 445
rect -644 389 -524 427
rect -352 427 -318 445
rect -266 445 -250 461
rect -42 461 42 477
rect -42 445 -26 461
rect -266 427 -232 445
rect -352 389 -232 427
rect -60 427 -26 445
rect 26 445 42 461
rect 250 461 334 477
rect 250 445 266 461
rect 26 427 60 445
rect -60 389 60 427
rect 232 427 266 445
rect 318 445 334 461
rect 542 461 626 477
rect 542 445 558 461
rect 318 427 352 445
rect 232 389 352 427
rect 524 427 558 445
rect 610 445 626 461
rect 834 461 918 477
rect 834 445 850 461
rect 610 427 644 445
rect 524 389 644 427
rect 816 427 850 445
rect 902 445 918 461
rect 902 427 936 445
rect 816 389 936 427
rect -936 71 -816 109
rect -936 55 -902 71
rect -918 37 -902 55
rect -850 55 -816 71
rect -644 71 -524 109
rect -644 55 -610 71
rect -850 37 -834 55
rect -918 21 -834 37
rect -626 37 -610 55
rect -558 55 -524 71
rect -352 71 -232 109
rect -352 55 -318 71
rect -558 37 -542 55
rect -626 21 -542 37
rect -334 37 -318 55
rect -266 55 -232 71
rect -60 71 60 109
rect -60 55 -26 71
rect -266 37 -250 55
rect -334 21 -250 37
rect -42 37 -26 55
rect 26 55 60 71
rect 232 71 352 109
rect 232 55 266 71
rect 26 37 42 55
rect -42 21 42 37
rect 250 37 266 55
rect 318 55 352 71
rect 524 71 644 109
rect 524 55 558 71
rect 318 37 334 55
rect 250 21 334 37
rect 542 37 558 55
rect 610 55 644 71
rect 816 71 936 109
rect 816 55 850 71
rect 610 37 626 55
rect 542 21 626 37
rect 834 37 850 55
rect 902 55 936 71
rect 902 37 918 55
rect 834 21 918 37
rect -918 -37 -834 -21
rect -918 -55 -902 -37
rect -936 -71 -902 -55
rect -850 -55 -834 -37
rect -626 -37 -542 -21
rect -626 -55 -610 -37
rect -850 -71 -816 -55
rect -936 -109 -816 -71
rect -644 -71 -610 -55
rect -558 -55 -542 -37
rect -334 -37 -250 -21
rect -334 -55 -318 -37
rect -558 -71 -524 -55
rect -644 -109 -524 -71
rect -352 -71 -318 -55
rect -266 -55 -250 -37
rect -42 -37 42 -21
rect -42 -55 -26 -37
rect -266 -71 -232 -55
rect -352 -109 -232 -71
rect -60 -71 -26 -55
rect 26 -55 42 -37
rect 250 -37 334 -21
rect 250 -55 266 -37
rect 26 -71 60 -55
rect -60 -109 60 -71
rect 232 -71 266 -55
rect 318 -55 334 -37
rect 542 -37 626 -21
rect 542 -55 558 -37
rect 318 -71 352 -55
rect 232 -109 352 -71
rect 524 -71 558 -55
rect 610 -55 626 -37
rect 834 -37 918 -21
rect 834 -55 850 -37
rect 610 -71 644 -55
rect 524 -109 644 -71
rect 816 -71 850 -55
rect 902 -55 918 -37
rect 902 -71 936 -55
rect 816 -109 936 -71
rect -936 -427 -816 -389
rect -936 -445 -902 -427
rect -918 -461 -902 -445
rect -850 -445 -816 -427
rect -644 -427 -524 -389
rect -644 -445 -610 -427
rect -850 -461 -834 -445
rect -918 -477 -834 -461
rect -626 -461 -610 -445
rect -558 -445 -524 -427
rect -352 -427 -232 -389
rect -352 -445 -318 -427
rect -558 -461 -542 -445
rect -626 -477 -542 -461
rect -334 -461 -318 -445
rect -266 -445 -232 -427
rect -60 -427 60 -389
rect -60 -445 -26 -427
rect -266 -461 -250 -445
rect -334 -477 -250 -461
rect -42 -461 -26 -445
rect 26 -445 60 -427
rect 232 -427 352 -389
rect 232 -445 266 -427
rect 26 -461 42 -445
rect -42 -477 42 -461
rect 250 -461 266 -445
rect 318 -445 352 -427
rect 524 -427 644 -389
rect 524 -445 558 -427
rect 318 -461 334 -445
rect 250 -477 334 -461
rect 542 -461 558 -445
rect 610 -445 644 -427
rect 816 -427 936 -389
rect 816 -445 850 -427
rect 610 -461 626 -445
rect 542 -477 626 -461
rect 834 -461 850 -445
rect 902 -445 936 -427
rect 902 -461 918 -445
rect 834 -477 918 -461
rect -918 -535 -834 -519
rect -918 -553 -902 -535
rect -936 -569 -902 -553
rect -850 -553 -834 -535
rect -626 -535 -542 -519
rect -626 -553 -610 -535
rect -850 -569 -816 -553
rect -936 -607 -816 -569
rect -644 -569 -610 -553
rect -558 -553 -542 -535
rect -334 -535 -250 -519
rect -334 -553 -318 -535
rect -558 -569 -524 -553
rect -644 -607 -524 -569
rect -352 -569 -318 -553
rect -266 -553 -250 -535
rect -42 -535 42 -519
rect -42 -553 -26 -535
rect -266 -569 -232 -553
rect -352 -607 -232 -569
rect -60 -569 -26 -553
rect 26 -553 42 -535
rect 250 -535 334 -519
rect 250 -553 266 -535
rect 26 -569 60 -553
rect -60 -607 60 -569
rect 232 -569 266 -553
rect 318 -553 334 -535
rect 542 -535 626 -519
rect 542 -553 558 -535
rect 318 -569 352 -553
rect 232 -607 352 -569
rect 524 -569 558 -553
rect 610 -553 626 -535
rect 834 -535 918 -519
rect 834 -553 850 -535
rect 610 -569 644 -553
rect 524 -607 644 -569
rect 816 -569 850 -553
rect 902 -553 918 -535
rect 902 -569 936 -553
rect 816 -607 936 -569
rect -936 -925 -816 -887
rect -936 -943 -902 -925
rect -918 -959 -902 -943
rect -850 -943 -816 -925
rect -644 -925 -524 -887
rect -644 -943 -610 -925
rect -850 -959 -834 -943
rect -918 -975 -834 -959
rect -626 -959 -610 -943
rect -558 -943 -524 -925
rect -352 -925 -232 -887
rect -352 -943 -318 -925
rect -558 -959 -542 -943
rect -626 -975 -542 -959
rect -334 -959 -318 -943
rect -266 -943 -232 -925
rect -60 -925 60 -887
rect -60 -943 -26 -925
rect -266 -959 -250 -943
rect -334 -975 -250 -959
rect -42 -959 -26 -943
rect 26 -943 60 -925
rect 232 -925 352 -887
rect 232 -943 266 -925
rect 26 -959 42 -943
rect -42 -975 42 -959
rect 250 -959 266 -943
rect 318 -943 352 -925
rect 524 -925 644 -887
rect 524 -943 558 -925
rect 318 -959 334 -943
rect 250 -975 334 -959
rect 542 -959 558 -943
rect 610 -943 644 -925
rect 816 -925 936 -887
rect 816 -943 850 -925
rect 610 -959 626 -943
rect 542 -975 626 -959
rect 834 -959 850 -943
rect 902 -943 936 -925
rect 902 -959 918 -943
rect 834 -975 918 -959
<< polycont >>
rect -902 925 -850 959
rect -610 925 -558 959
rect -318 925 -266 959
rect -26 925 26 959
rect 266 925 318 959
rect 558 925 610 959
rect 850 925 902 959
rect -902 535 -850 569
rect -610 535 -558 569
rect -318 535 -266 569
rect -26 535 26 569
rect 266 535 318 569
rect 558 535 610 569
rect 850 535 902 569
rect -902 427 -850 461
rect -610 427 -558 461
rect -318 427 -266 461
rect -26 427 26 461
rect 266 427 318 461
rect 558 427 610 461
rect 850 427 902 461
rect -902 37 -850 71
rect -610 37 -558 71
rect -318 37 -266 71
rect -26 37 26 71
rect 266 37 318 71
rect 558 37 610 71
rect 850 37 902 71
rect -902 -71 -850 -37
rect -610 -71 -558 -37
rect -318 -71 -266 -37
rect -26 -71 26 -37
rect 266 -71 318 -37
rect 558 -71 610 -37
rect 850 -71 902 -37
rect -902 -461 -850 -427
rect -610 -461 -558 -427
rect -318 -461 -266 -427
rect -26 -461 26 -427
rect 266 -461 318 -427
rect 558 -461 610 -427
rect 850 -461 902 -427
rect -902 -569 -850 -535
rect -610 -569 -558 -535
rect -318 -569 -266 -535
rect -26 -569 26 -535
rect 266 -569 318 -535
rect 558 -569 610 -535
rect 850 -569 902 -535
rect -902 -959 -850 -925
rect -610 -959 -558 -925
rect -318 -959 -266 -925
rect -26 -959 26 -925
rect 266 -959 318 -925
rect 558 -959 610 -925
rect 850 -959 902 -925
<< locali >>
rect -918 925 -902 959
rect -850 925 -834 959
rect -626 925 -610 959
rect -558 925 -542 959
rect -334 925 -318 959
rect -266 925 -250 959
rect -42 925 -26 959
rect 26 925 42 959
rect 250 925 266 959
rect 318 925 334 959
rect 542 925 558 959
rect 610 925 626 959
rect 834 925 850 959
rect 902 925 918 959
rect -982 875 -948 891
rect -982 603 -948 619
rect -804 875 -770 891
rect -804 603 -770 619
rect -690 875 -656 891
rect -690 603 -656 619
rect -512 875 -478 891
rect -512 603 -478 619
rect -398 875 -364 891
rect -398 603 -364 619
rect -220 875 -186 891
rect -220 603 -186 619
rect -106 875 -72 891
rect -106 603 -72 619
rect 72 875 106 891
rect 72 603 106 619
rect 186 875 220 891
rect 186 603 220 619
rect 364 875 398 891
rect 364 603 398 619
rect 478 875 512 891
rect 478 603 512 619
rect 656 875 690 891
rect 656 603 690 619
rect 770 875 804 891
rect 770 603 804 619
rect 948 875 982 891
rect 948 603 982 619
rect -918 535 -902 569
rect -850 535 -834 569
rect -626 535 -610 569
rect -558 535 -542 569
rect -334 535 -318 569
rect -266 535 -250 569
rect -42 535 -26 569
rect 26 535 42 569
rect 250 535 266 569
rect 318 535 334 569
rect 542 535 558 569
rect 610 535 626 569
rect 834 535 850 569
rect 902 535 918 569
rect -918 427 -902 461
rect -850 427 -834 461
rect -626 427 -610 461
rect -558 427 -542 461
rect -334 427 -318 461
rect -266 427 -250 461
rect -42 427 -26 461
rect 26 427 42 461
rect 250 427 266 461
rect 318 427 334 461
rect 542 427 558 461
rect 610 427 626 461
rect 834 427 850 461
rect 902 427 918 461
rect -982 377 -948 393
rect -982 105 -948 121
rect -804 377 -770 393
rect -804 105 -770 121
rect -690 377 -656 393
rect -690 105 -656 121
rect -512 377 -478 393
rect -512 105 -478 121
rect -398 377 -364 393
rect -398 105 -364 121
rect -220 377 -186 393
rect -220 105 -186 121
rect -106 377 -72 393
rect -106 105 -72 121
rect 72 377 106 393
rect 72 105 106 121
rect 186 377 220 393
rect 186 105 220 121
rect 364 377 398 393
rect 364 105 398 121
rect 478 377 512 393
rect 478 105 512 121
rect 656 377 690 393
rect 656 105 690 121
rect 770 377 804 393
rect 770 105 804 121
rect 948 377 982 393
rect 948 105 982 121
rect -918 37 -902 71
rect -850 37 -834 71
rect -626 37 -610 71
rect -558 37 -542 71
rect -334 37 -318 71
rect -266 37 -250 71
rect -42 37 -26 71
rect 26 37 42 71
rect 250 37 266 71
rect 318 37 334 71
rect 542 37 558 71
rect 610 37 626 71
rect 834 37 850 71
rect 902 37 918 71
rect -918 -71 -902 -37
rect -850 -71 -834 -37
rect -626 -71 -610 -37
rect -558 -71 -542 -37
rect -334 -71 -318 -37
rect -266 -71 -250 -37
rect -42 -71 -26 -37
rect 26 -71 42 -37
rect 250 -71 266 -37
rect 318 -71 334 -37
rect 542 -71 558 -37
rect 610 -71 626 -37
rect 834 -71 850 -37
rect 902 -71 918 -37
rect -982 -121 -948 -105
rect -982 -393 -948 -377
rect -804 -121 -770 -105
rect -804 -393 -770 -377
rect -690 -121 -656 -105
rect -690 -393 -656 -377
rect -512 -121 -478 -105
rect -512 -393 -478 -377
rect -398 -121 -364 -105
rect -398 -393 -364 -377
rect -220 -121 -186 -105
rect -220 -393 -186 -377
rect -106 -121 -72 -105
rect -106 -393 -72 -377
rect 72 -121 106 -105
rect 72 -393 106 -377
rect 186 -121 220 -105
rect 186 -393 220 -377
rect 364 -121 398 -105
rect 364 -393 398 -377
rect 478 -121 512 -105
rect 478 -393 512 -377
rect 656 -121 690 -105
rect 656 -393 690 -377
rect 770 -121 804 -105
rect 770 -393 804 -377
rect 948 -121 982 -105
rect 948 -393 982 -377
rect -918 -461 -902 -427
rect -850 -461 -834 -427
rect -626 -461 -610 -427
rect -558 -461 -542 -427
rect -334 -461 -318 -427
rect -266 -461 -250 -427
rect -42 -461 -26 -427
rect 26 -461 42 -427
rect 250 -461 266 -427
rect 318 -461 334 -427
rect 542 -461 558 -427
rect 610 -461 626 -427
rect 834 -461 850 -427
rect 902 -461 918 -427
rect -918 -569 -902 -535
rect -850 -569 -834 -535
rect -626 -569 -610 -535
rect -558 -569 -542 -535
rect -334 -569 -318 -535
rect -266 -569 -250 -535
rect -42 -569 -26 -535
rect 26 -569 42 -535
rect 250 -569 266 -535
rect 318 -569 334 -535
rect 542 -569 558 -535
rect 610 -569 626 -535
rect 834 -569 850 -535
rect 902 -569 918 -535
rect -982 -619 -948 -603
rect -982 -891 -948 -875
rect -804 -619 -770 -603
rect -804 -891 -770 -875
rect -690 -619 -656 -603
rect -690 -891 -656 -875
rect -512 -619 -478 -603
rect -512 -891 -478 -875
rect -398 -619 -364 -603
rect -398 -891 -364 -875
rect -220 -619 -186 -603
rect -220 -891 -186 -875
rect -106 -619 -72 -603
rect -106 -891 -72 -875
rect 72 -619 106 -603
rect 72 -891 106 -875
rect 186 -619 220 -603
rect 186 -891 220 -875
rect 364 -619 398 -603
rect 364 -891 398 -875
rect 478 -619 512 -603
rect 478 -891 512 -875
rect 656 -619 690 -603
rect 656 -891 690 -875
rect 770 -619 804 -603
rect 770 -891 804 -875
rect 948 -619 982 -603
rect 948 -891 982 -875
rect -918 -959 -902 -925
rect -850 -959 -834 -925
rect -626 -959 -610 -925
rect -558 -959 -542 -925
rect -334 -959 -318 -925
rect -266 -959 -250 -925
rect -42 -959 -26 -925
rect 26 -959 42 -925
rect 250 -959 266 -925
rect 318 -959 334 -925
rect 542 -959 558 -925
rect 610 -959 626 -925
rect 834 -959 850 -925
rect 902 -959 918 -925
<< viali >>
rect -902 925 -850 959
rect -610 925 -558 959
rect -318 925 -266 959
rect -26 925 26 959
rect 266 925 318 959
rect 558 925 610 959
rect 850 925 902 959
rect -982 619 -948 875
rect -804 619 -770 875
rect -690 619 -656 875
rect -512 619 -478 875
rect -398 619 -364 875
rect -220 619 -186 875
rect -106 619 -72 875
rect 72 619 106 875
rect 186 619 220 875
rect 364 619 398 875
rect 478 619 512 875
rect 656 619 690 875
rect 770 619 804 875
rect 948 619 982 875
rect -902 535 -850 569
rect -610 535 -558 569
rect -318 535 -266 569
rect -26 535 26 569
rect 266 535 318 569
rect 558 535 610 569
rect 850 535 902 569
rect -902 427 -850 461
rect -610 427 -558 461
rect -318 427 -266 461
rect -26 427 26 461
rect 266 427 318 461
rect 558 427 610 461
rect 850 427 902 461
rect -982 121 -948 377
rect -804 121 -770 377
rect -690 121 -656 377
rect -512 121 -478 377
rect -398 121 -364 377
rect -220 121 -186 377
rect -106 121 -72 377
rect 72 121 106 377
rect 186 121 220 377
rect 364 121 398 377
rect 478 121 512 377
rect 656 121 690 377
rect 770 121 804 377
rect 948 121 982 377
rect -902 37 -850 71
rect -610 37 -558 71
rect -318 37 -266 71
rect -26 37 26 71
rect 266 37 318 71
rect 558 37 610 71
rect 850 37 902 71
rect -902 -71 -850 -37
rect -610 -71 -558 -37
rect -318 -71 -266 -37
rect -26 -71 26 -37
rect 266 -71 318 -37
rect 558 -71 610 -37
rect 850 -71 902 -37
rect -982 -377 -948 -121
rect -804 -377 -770 -121
rect -690 -377 -656 -121
rect -512 -377 -478 -121
rect -398 -377 -364 -121
rect -220 -377 -186 -121
rect -106 -377 -72 -121
rect 72 -377 106 -121
rect 186 -377 220 -121
rect 364 -377 398 -121
rect 478 -377 512 -121
rect 656 -377 690 -121
rect 770 -377 804 -121
rect 948 -377 982 -121
rect -902 -461 -850 -427
rect -610 -461 -558 -427
rect -318 -461 -266 -427
rect -26 -461 26 -427
rect 266 -461 318 -427
rect 558 -461 610 -427
rect 850 -461 902 -427
rect -902 -569 -850 -535
rect -610 -569 -558 -535
rect -318 -569 -266 -535
rect -26 -569 26 -535
rect 266 -569 318 -535
rect 558 -569 610 -535
rect 850 -569 902 -535
rect -982 -875 -948 -619
rect -804 -875 -770 -619
rect -690 -875 -656 -619
rect -512 -875 -478 -619
rect -398 -875 -364 -619
rect -220 -875 -186 -619
rect -106 -875 -72 -619
rect 72 -875 106 -619
rect 186 -875 220 -619
rect 364 -875 398 -619
rect 478 -875 512 -619
rect 656 -875 690 -619
rect 770 -875 804 -619
rect 948 -875 982 -619
rect -902 -959 -850 -925
rect -610 -959 -558 -925
rect -318 -959 -266 -925
rect -26 -959 26 -925
rect 266 -959 318 -925
rect 558 -959 610 -925
rect 850 -959 902 -925
<< metal1 >>
rect -914 963 -838 965
rect -988 959 -764 963
rect -988 925 -902 959
rect -850 925 -764 959
rect -988 917 -764 925
rect -622 959 -546 965
rect -622 925 -610 959
rect -558 925 -546 959
rect -622 919 -546 925
rect -330 959 -254 965
rect -330 925 -318 959
rect -266 925 -254 959
rect -330 919 -254 925
rect -38 959 38 965
rect -38 925 -26 959
rect 26 925 38 959
rect -38 919 38 925
rect 254 959 330 965
rect 254 925 266 959
rect 318 925 330 959
rect 254 919 330 925
rect 546 959 622 965
rect 546 925 558 959
rect 610 925 622 959
rect 546 919 622 925
rect 764 959 988 965
rect 764 925 850 959
rect 902 933 988 959
rect 902 925 992 933
rect 764 919 992 925
rect -988 875 -942 917
rect -988 619 -982 875
rect -948 619 -942 875
rect -988 575 -942 619
rect -810 875 -764 917
rect -810 619 -804 875
rect -770 619 -764 875
rect -810 575 -764 619
rect -696 875 -650 887
rect -696 619 -690 875
rect -656 619 -650 875
rect -696 607 -650 619
rect -518 875 -472 887
rect -518 619 -512 875
rect -478 619 -472 875
rect -518 607 -472 619
rect -404 875 -358 887
rect -404 619 -398 875
rect -364 619 -358 875
rect -404 607 -358 619
rect -226 875 -180 887
rect -226 619 -220 875
rect -186 619 -180 875
rect -226 607 -180 619
rect -112 875 -66 887
rect -112 619 -106 875
rect -72 619 -66 875
rect -112 607 -66 619
rect 66 875 112 887
rect 66 619 72 875
rect 106 619 112 875
rect 66 607 112 619
rect 180 875 226 887
rect 180 619 186 875
rect 220 619 226 875
rect 180 607 226 619
rect 358 875 404 887
rect 358 619 364 875
rect 398 619 404 875
rect 358 607 404 619
rect 472 875 518 887
rect 472 619 478 875
rect 512 619 518 875
rect 472 607 518 619
rect 650 875 696 887
rect 650 619 656 875
rect 690 619 696 875
rect 650 607 696 619
rect 764 875 810 919
rect 764 619 770 875
rect 804 619 810 875
rect 764 575 810 619
rect 942 875 992 919
rect 942 619 948 875
rect 982 619 992 875
rect 942 575 992 619
rect -988 569 -764 575
rect -988 535 -902 569
rect -850 535 -764 569
rect -988 461 -764 535
rect -622 569 -546 575
rect -622 535 -610 569
rect -558 535 -546 569
rect -622 529 -546 535
rect -330 569 -254 575
rect -330 535 -318 569
rect -266 535 -254 569
rect -330 529 -254 535
rect -38 569 38 575
rect -38 535 -26 569
rect 26 535 38 569
rect -38 529 38 535
rect 254 569 330 575
rect 254 535 266 569
rect 318 535 330 569
rect 254 529 330 535
rect 546 569 622 575
rect 546 535 558 569
rect 610 535 622 569
rect 546 529 622 535
rect 764 569 992 575
rect 764 535 850 569
rect 902 535 992 569
rect -988 427 -902 461
rect -850 427 -764 461
rect -988 421 -764 427
rect -622 461 -546 467
rect -622 427 -610 461
rect -558 427 -546 461
rect -622 421 -546 427
rect -330 461 -254 467
rect -330 427 -318 461
rect -266 427 -254 461
rect -330 421 -254 427
rect -38 461 38 467
rect -38 427 -26 461
rect 26 427 38 461
rect -38 421 38 427
rect 254 461 330 467
rect 254 427 266 461
rect 318 427 330 461
rect 254 421 330 427
rect 546 461 622 467
rect 546 427 558 461
rect 610 427 622 461
rect 546 421 622 427
rect 764 461 992 535
rect 764 427 850 461
rect 902 427 992 461
rect 764 423 992 427
rect -988 377 -942 421
rect -988 121 -982 377
rect -948 121 -942 377
rect -988 77 -942 121
rect -810 377 -764 421
rect -810 121 -804 377
rect -770 121 -764 377
rect -810 77 -764 121
rect -696 377 -650 389
rect -696 121 -690 377
rect -656 121 -650 377
rect -696 109 -650 121
rect -518 377 -472 389
rect -518 121 -512 377
rect -478 121 -472 377
rect -518 109 -472 121
rect -404 377 -358 389
rect -404 121 -398 377
rect -364 121 -358 377
rect -404 109 -358 121
rect -226 377 -180 389
rect -226 121 -220 377
rect -186 121 -180 377
rect -226 109 -180 121
rect -112 377 -66 389
rect -112 121 -106 377
rect -72 121 -66 377
rect -112 109 -66 121
rect 66 377 112 389
rect 66 121 72 377
rect 106 121 112 377
rect 66 109 112 121
rect 180 377 226 389
rect 180 121 186 377
rect 220 121 226 377
rect 180 109 226 121
rect 358 377 404 389
rect 358 121 364 377
rect 398 121 404 377
rect 358 109 404 121
rect 472 377 518 389
rect 472 121 478 377
rect 512 121 518 377
rect 472 109 518 121
rect 650 377 696 389
rect 650 121 656 377
rect 690 121 696 377
rect 650 109 696 121
rect 764 377 810 423
rect 838 421 914 423
rect 946 389 992 423
rect 764 121 770 377
rect 804 121 810 377
rect -988 71 -764 77
rect -988 37 -902 71
rect -850 37 -764 71
rect -988 31 -764 37
rect -622 71 -546 77
rect -622 37 -610 71
rect -558 37 -546 71
rect -622 31 -546 37
rect -330 71 -254 77
rect -330 37 -318 71
rect -266 37 -254 71
rect -330 31 -254 37
rect -38 71 38 77
rect -38 37 -26 71
rect 26 37 38 71
rect -38 31 38 37
rect 254 71 330 77
rect 254 37 266 71
rect 318 37 330 71
rect 254 31 330 37
rect 546 71 622 77
rect 546 37 558 71
rect 610 37 622 71
rect 546 31 622 37
rect 764 63 810 121
rect 942 377 992 389
rect 942 121 948 377
rect 982 121 992 377
rect 942 109 992 121
rect 838 71 914 77
rect 838 63 850 71
rect 764 37 850 63
rect 902 63 914 71
rect 946 63 992 109
rect 902 37 992 63
rect -988 -31 -942 31
rect -810 -31 -764 31
rect -988 -37 -764 -31
rect -988 -71 -902 -37
rect -850 -71 -764 -37
rect -988 -77 -764 -71
rect -622 -37 -546 -31
rect -622 -71 -610 -37
rect -558 -71 -546 -37
rect -622 -77 -546 -71
rect -330 -37 -254 -31
rect -330 -71 -318 -37
rect -266 -71 -254 -37
rect -330 -77 -254 -71
rect -38 -37 38 -31
rect -38 -71 -26 -37
rect 26 -71 38 -37
rect -38 -77 38 -71
rect 254 -37 330 -31
rect 254 -71 266 -37
rect 318 -71 330 -37
rect 254 -77 330 -71
rect 546 -37 622 -31
rect 546 -71 558 -37
rect 610 -71 622 -37
rect 546 -77 622 -71
rect 764 -37 992 37
rect 764 -71 850 -37
rect 902 -71 992 -37
rect 764 -75 992 -71
rect -988 -121 -942 -77
rect -988 -377 -982 -121
rect -948 -377 -942 -121
rect -988 -391 -942 -377
rect -810 -121 -764 -77
rect -810 -377 -804 -121
rect -770 -377 -764 -121
rect -810 -391 -764 -377
rect -696 -121 -650 -109
rect -696 -377 -690 -121
rect -656 -377 -650 -121
rect -696 -389 -650 -377
rect -518 -121 -472 -109
rect -518 -377 -512 -121
rect -478 -377 -472 -121
rect -518 -389 -472 -377
rect -404 -121 -358 -109
rect -404 -377 -398 -121
rect -364 -377 -358 -121
rect -404 -389 -358 -377
rect -226 -121 -180 -109
rect -226 -377 -220 -121
rect -186 -377 -180 -121
rect -226 -389 -180 -377
rect -112 -121 -66 -109
rect -112 -377 -106 -121
rect -72 -377 -66 -121
rect -112 -389 -66 -377
rect 66 -121 112 -109
rect 66 -377 72 -121
rect 106 -377 112 -121
rect 66 -389 112 -377
rect 180 -121 226 -109
rect 180 -377 186 -121
rect 220 -377 226 -121
rect 180 -389 226 -377
rect 358 -121 404 -109
rect 358 -377 364 -121
rect 398 -377 404 -121
rect 358 -389 404 -377
rect 472 -121 518 -109
rect 472 -377 478 -121
rect 512 -377 518 -121
rect 472 -389 518 -377
rect 650 -121 696 -109
rect 650 -377 656 -121
rect 690 -377 696 -121
rect 650 -389 696 -377
rect 764 -121 810 -75
rect 838 -77 914 -75
rect 946 -109 992 -75
rect 764 -377 770 -121
rect 804 -377 810 -121
rect -988 -427 -764 -391
rect -988 -461 -902 -427
rect -850 -461 -764 -427
rect -988 -535 -764 -461
rect -622 -427 -546 -421
rect -622 -461 -610 -427
rect -558 -461 -546 -427
rect -622 -467 -546 -461
rect -330 -427 -254 -421
rect -330 -461 -318 -427
rect -266 -461 -254 -427
rect -330 -467 -254 -461
rect -38 -427 38 -421
rect -38 -461 -26 -427
rect 26 -461 38 -427
rect -38 -467 38 -461
rect 254 -427 330 -421
rect 254 -461 266 -427
rect 318 -461 330 -427
rect 254 -467 330 -461
rect 546 -427 622 -421
rect 546 -461 558 -427
rect 610 -461 622 -427
rect 546 -467 622 -461
rect 764 -439 810 -377
rect 942 -121 992 -109
rect 942 -377 948 -121
rect 982 -377 992 -121
rect 942 -389 992 -377
rect 838 -427 914 -421
rect 838 -439 850 -427
rect 764 -461 850 -439
rect 902 -439 914 -427
rect 946 -439 992 -389
rect 902 -461 992 -439
rect -988 -569 -902 -535
rect -850 -569 -764 -535
rect -988 -601 -764 -569
rect -622 -535 -546 -529
rect -622 -569 -610 -535
rect -558 -569 -546 -535
rect -622 -575 -546 -569
rect -330 -535 -254 -529
rect -330 -569 -318 -535
rect -266 -569 -254 -535
rect -330 -575 -254 -569
rect -38 -535 38 -529
rect -38 -569 -26 -535
rect 26 -569 38 -535
rect -38 -575 38 -569
rect 254 -535 330 -529
rect 254 -569 266 -535
rect 318 -569 330 -535
rect 254 -575 330 -569
rect 546 -535 622 -529
rect 546 -569 558 -535
rect 610 -569 622 -535
rect 546 -575 622 -569
rect 764 -535 992 -461
rect 764 -567 850 -535
rect -988 -619 -942 -601
rect -988 -875 -982 -619
rect -948 -875 -942 -619
rect -988 -915 -942 -875
rect -810 -619 -764 -601
rect -810 -875 -804 -619
rect -770 -875 -764 -619
rect -810 -915 -764 -875
rect -696 -619 -650 -607
rect -696 -875 -690 -619
rect -656 -875 -650 -619
rect -696 -887 -650 -875
rect -518 -619 -472 -607
rect -518 -875 -512 -619
rect -478 -875 -472 -619
rect -518 -887 -472 -875
rect -404 -619 -358 -607
rect -404 -875 -398 -619
rect -364 -875 -358 -619
rect -404 -887 -358 -875
rect -226 -619 -180 -607
rect -226 -875 -220 -619
rect -186 -875 -180 -619
rect -226 -887 -180 -875
rect -112 -619 -66 -607
rect -112 -875 -106 -619
rect -72 -875 -66 -619
rect -112 -887 -66 -875
rect 66 -619 112 -607
rect 66 -875 72 -619
rect 106 -875 112 -619
rect 66 -887 112 -875
rect 180 -619 226 -607
rect 180 -875 186 -619
rect 220 -875 226 -619
rect 180 -887 226 -875
rect 358 -619 404 -607
rect 358 -875 364 -619
rect 398 -875 404 -619
rect 358 -887 404 -875
rect 472 -619 518 -607
rect 472 -875 478 -619
rect 512 -875 518 -619
rect 472 -887 518 -875
rect 650 -619 696 -607
rect 650 -875 656 -619
rect 690 -875 696 -619
rect 650 -887 696 -875
rect 764 -619 810 -567
rect 838 -569 850 -567
rect 902 -567 992 -535
rect 902 -569 914 -567
rect 838 -575 914 -569
rect 946 -607 992 -567
rect 764 -875 770 -619
rect 804 -875 810 -619
rect -988 -925 -764 -915
rect 764 -919 810 -875
rect 942 -619 992 -607
rect 942 -875 948 -619
rect 982 -875 992 -619
rect 942 -887 992 -875
rect 946 -919 992 -887
rect -988 -959 -902 -925
rect -850 -959 -764 -925
rect -988 -961 -764 -959
rect -622 -925 -546 -919
rect -622 -959 -610 -925
rect -558 -959 -546 -925
rect -988 -967 -942 -961
rect -914 -965 -838 -961
rect -622 -965 -546 -959
rect -330 -925 -254 -919
rect -330 -959 -318 -925
rect -266 -959 -254 -925
rect -330 -965 -254 -959
rect -38 -925 38 -919
rect -38 -959 -26 -925
rect 26 -959 38 -925
rect -38 -965 38 -959
rect 254 -925 330 -919
rect 254 -959 266 -925
rect 318 -959 330 -925
rect 254 -965 330 -959
rect 546 -925 622 -919
rect 546 -959 558 -925
rect 610 -959 622 -925
rect 546 -965 622 -959
rect 764 -925 992 -919
rect 764 -959 850 -925
rect 902 -959 992 -925
rect 764 -965 992 -959
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 4 nf 7 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
