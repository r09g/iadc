magic
tech sky130A
magscale 1 2
timestamp 1654898484
<< error_p >>
rect -1531 572 -1473 578
rect -1373 572 -1315 578
rect -1215 572 -1157 578
rect -1057 572 -999 578
rect -899 572 -841 578
rect -741 572 -683 578
rect -583 572 -525 578
rect -425 572 -367 578
rect -267 572 -209 578
rect -109 572 -51 578
rect 51 572 109 578
rect 209 572 267 578
rect 367 572 425 578
rect 525 572 583 578
rect 683 572 741 578
rect 841 572 899 578
rect 999 572 1057 578
rect 1157 572 1215 578
rect 1315 572 1373 578
rect 1473 572 1531 578
rect -1531 538 -1519 572
rect -1373 538 -1361 572
rect -1215 538 -1203 572
rect -1057 538 -1045 572
rect -899 538 -887 572
rect -741 538 -729 572
rect -583 538 -571 572
rect -425 538 -413 572
rect -267 538 -255 572
rect -109 538 -97 572
rect 51 538 63 572
rect 209 538 221 572
rect 367 538 379 572
rect 525 538 537 572
rect 683 538 695 572
rect 841 538 853 572
rect 999 538 1011 572
rect 1157 538 1169 572
rect 1315 538 1327 572
rect 1473 538 1485 572
rect -1531 532 -1473 538
rect -1373 532 -1315 538
rect -1215 532 -1157 538
rect -1057 532 -999 538
rect -899 532 -841 538
rect -741 532 -683 538
rect -583 532 -525 538
rect -425 532 -367 538
rect -267 532 -209 538
rect -109 532 -51 538
rect 51 532 109 538
rect 209 532 267 538
rect 367 532 425 538
rect 525 532 583 538
rect 683 532 741 538
rect 841 532 899 538
rect 999 532 1057 538
rect 1157 532 1215 538
rect 1315 532 1373 538
rect 1473 532 1531 538
rect -1531 -538 -1473 -532
rect -1373 -538 -1315 -532
rect -1215 -538 -1157 -532
rect -1057 -538 -999 -532
rect -899 -538 -841 -532
rect -741 -538 -683 -532
rect -583 -538 -525 -532
rect -425 -538 -367 -532
rect -267 -538 -209 -532
rect -109 -538 -51 -532
rect 51 -538 109 -532
rect 209 -538 267 -532
rect 367 -538 425 -532
rect 525 -538 583 -532
rect 683 -538 741 -532
rect 841 -538 899 -532
rect 999 -538 1057 -532
rect 1157 -538 1215 -532
rect 1315 -538 1373 -532
rect 1473 -538 1531 -532
rect -1531 -572 -1519 -538
rect -1373 -572 -1361 -538
rect -1215 -572 -1203 -538
rect -1057 -572 -1045 -538
rect -899 -572 -887 -538
rect -741 -572 -729 -538
rect -583 -572 -571 -538
rect -425 -572 -413 -538
rect -267 -572 -255 -538
rect -109 -572 -97 -538
rect 51 -572 63 -538
rect 209 -572 221 -538
rect 367 -572 379 -538
rect 525 -572 537 -538
rect 683 -572 695 -538
rect 841 -572 853 -538
rect 999 -572 1011 -538
rect 1157 -572 1169 -538
rect 1315 -572 1327 -538
rect 1473 -572 1485 -538
rect -1531 -578 -1473 -572
rect -1373 -578 -1315 -572
rect -1215 -578 -1157 -572
rect -1057 -578 -999 -572
rect -899 -578 -841 -572
rect -741 -578 -683 -572
rect -583 -578 -525 -572
rect -425 -578 -367 -572
rect -267 -578 -209 -572
rect -109 -578 -51 -572
rect 51 -578 109 -572
rect 209 -578 267 -572
rect 367 -578 425 -572
rect 525 -578 583 -572
rect 683 -578 741 -572
rect 841 -578 899 -572
rect 999 -578 1057 -572
rect 1157 -578 1215 -572
rect 1315 -578 1373 -572
rect 1473 -578 1531 -572
<< pwell >>
rect -1779 -758 1779 758
<< mvnmos >>
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
<< mvndiff >>
rect -1609 488 -1551 500
rect -1609 -488 -1597 488
rect -1563 -488 -1551 488
rect -1609 -500 -1551 -488
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
rect 1551 488 1609 500
rect 1551 -488 1563 488
rect 1597 -488 1609 488
rect 1551 -500 1609 -488
<< mvndiffc >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< mvpsubdiff >>
rect -1743 710 1743 722
rect -1743 676 -1635 710
rect 1635 676 1743 710
rect -1743 664 1743 676
rect -1743 614 -1685 664
rect -1743 -614 -1731 614
rect -1697 -614 -1685 614
rect 1685 614 1743 664
rect -1743 -664 -1685 -614
rect 1685 -614 1697 614
rect 1731 -614 1743 614
rect 1685 -664 1743 -614
rect -1743 -676 1743 -664
rect -1743 -710 -1635 -676
rect 1635 -710 1743 -676
rect -1743 -722 1743 -710
<< mvpsubdiffcont >>
rect -1635 676 1635 710
rect -1731 -614 -1697 614
rect 1697 -614 1731 614
rect -1635 -710 1635 -676
<< poly >>
rect -1551 572 -1451 588
rect -1551 538 -1535 572
rect -1467 538 -1451 572
rect -1551 500 -1451 538
rect -1393 572 -1293 588
rect -1393 538 -1377 572
rect -1309 538 -1293 572
rect -1393 500 -1293 538
rect -1235 572 -1135 588
rect -1235 538 -1219 572
rect -1151 538 -1135 572
rect -1235 500 -1135 538
rect -1077 572 -977 588
rect -1077 538 -1061 572
rect -993 538 -977 572
rect -1077 500 -977 538
rect -919 572 -819 588
rect -919 538 -903 572
rect -835 538 -819 572
rect -919 500 -819 538
rect -761 572 -661 588
rect -761 538 -745 572
rect -677 538 -661 572
rect -761 500 -661 538
rect -603 572 -503 588
rect -603 538 -587 572
rect -519 538 -503 572
rect -603 500 -503 538
rect -445 572 -345 588
rect -445 538 -429 572
rect -361 538 -345 572
rect -445 500 -345 538
rect -287 572 -187 588
rect -287 538 -271 572
rect -203 538 -187 572
rect -287 500 -187 538
rect -129 572 -29 588
rect -129 538 -113 572
rect -45 538 -29 572
rect -129 500 -29 538
rect 29 572 129 588
rect 29 538 45 572
rect 113 538 129 572
rect 29 500 129 538
rect 187 572 287 588
rect 187 538 203 572
rect 271 538 287 572
rect 187 500 287 538
rect 345 572 445 588
rect 345 538 361 572
rect 429 538 445 572
rect 345 500 445 538
rect 503 572 603 588
rect 503 538 519 572
rect 587 538 603 572
rect 503 500 603 538
rect 661 572 761 588
rect 661 538 677 572
rect 745 538 761 572
rect 661 500 761 538
rect 819 572 919 588
rect 819 538 835 572
rect 903 538 919 572
rect 819 500 919 538
rect 977 572 1077 588
rect 977 538 993 572
rect 1061 538 1077 572
rect 977 500 1077 538
rect 1135 572 1235 588
rect 1135 538 1151 572
rect 1219 538 1235 572
rect 1135 500 1235 538
rect 1293 572 1393 588
rect 1293 538 1309 572
rect 1377 538 1393 572
rect 1293 500 1393 538
rect 1451 572 1551 588
rect 1451 538 1467 572
rect 1535 538 1551 572
rect 1451 500 1551 538
rect -1551 -538 -1451 -500
rect -1551 -572 -1535 -538
rect -1467 -572 -1451 -538
rect -1551 -588 -1451 -572
rect -1393 -538 -1293 -500
rect -1393 -572 -1377 -538
rect -1309 -572 -1293 -538
rect -1393 -588 -1293 -572
rect -1235 -538 -1135 -500
rect -1235 -572 -1219 -538
rect -1151 -572 -1135 -538
rect -1235 -588 -1135 -572
rect -1077 -538 -977 -500
rect -1077 -572 -1061 -538
rect -993 -572 -977 -538
rect -1077 -588 -977 -572
rect -919 -538 -819 -500
rect -919 -572 -903 -538
rect -835 -572 -819 -538
rect -919 -588 -819 -572
rect -761 -538 -661 -500
rect -761 -572 -745 -538
rect -677 -572 -661 -538
rect -761 -588 -661 -572
rect -603 -538 -503 -500
rect -603 -572 -587 -538
rect -519 -572 -503 -538
rect -603 -588 -503 -572
rect -445 -538 -345 -500
rect -445 -572 -429 -538
rect -361 -572 -345 -538
rect -445 -588 -345 -572
rect -287 -538 -187 -500
rect -287 -572 -271 -538
rect -203 -572 -187 -538
rect -287 -588 -187 -572
rect -129 -538 -29 -500
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect -129 -588 -29 -572
rect 29 -538 129 -500
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 29 -588 129 -572
rect 187 -538 287 -500
rect 187 -572 203 -538
rect 271 -572 287 -538
rect 187 -588 287 -572
rect 345 -538 445 -500
rect 345 -572 361 -538
rect 429 -572 445 -538
rect 345 -588 445 -572
rect 503 -538 603 -500
rect 503 -572 519 -538
rect 587 -572 603 -538
rect 503 -588 603 -572
rect 661 -538 761 -500
rect 661 -572 677 -538
rect 745 -572 761 -538
rect 661 -588 761 -572
rect 819 -538 919 -500
rect 819 -572 835 -538
rect 903 -572 919 -538
rect 819 -588 919 -572
rect 977 -538 1077 -500
rect 977 -572 993 -538
rect 1061 -572 1077 -538
rect 977 -588 1077 -572
rect 1135 -538 1235 -500
rect 1135 -572 1151 -538
rect 1219 -572 1235 -538
rect 1135 -588 1235 -572
rect 1293 -538 1393 -500
rect 1293 -572 1309 -538
rect 1377 -572 1393 -538
rect 1293 -588 1393 -572
rect 1451 -538 1551 -500
rect 1451 -572 1467 -538
rect 1535 -572 1551 -538
rect 1451 -588 1551 -572
<< polycont >>
rect -1535 538 -1467 572
rect -1377 538 -1309 572
rect -1219 538 -1151 572
rect -1061 538 -993 572
rect -903 538 -835 572
rect -745 538 -677 572
rect -587 538 -519 572
rect -429 538 -361 572
rect -271 538 -203 572
rect -113 538 -45 572
rect 45 538 113 572
rect 203 538 271 572
rect 361 538 429 572
rect 519 538 587 572
rect 677 538 745 572
rect 835 538 903 572
rect 993 538 1061 572
rect 1151 538 1219 572
rect 1309 538 1377 572
rect 1467 538 1535 572
rect -1535 -572 -1467 -538
rect -1377 -572 -1309 -538
rect -1219 -572 -1151 -538
rect -1061 -572 -993 -538
rect -903 -572 -835 -538
rect -745 -572 -677 -538
rect -587 -572 -519 -538
rect -429 -572 -361 -538
rect -271 -572 -203 -538
rect -113 -572 -45 -538
rect 45 -572 113 -538
rect 203 -572 271 -538
rect 361 -572 429 -538
rect 519 -572 587 -538
rect 677 -572 745 -538
rect 835 -572 903 -538
rect 993 -572 1061 -538
rect 1151 -572 1219 -538
rect 1309 -572 1377 -538
rect 1467 -572 1535 -538
<< locali >>
rect -1731 676 -1635 710
rect 1635 676 1731 710
rect -1731 614 -1697 676
rect 1697 614 1731 676
rect -1551 538 -1535 572
rect -1467 538 -1451 572
rect -1393 538 -1377 572
rect -1309 538 -1293 572
rect -1235 538 -1219 572
rect -1151 538 -1135 572
rect -1077 538 -1061 572
rect -993 538 -977 572
rect -919 538 -903 572
rect -835 538 -819 572
rect -761 538 -745 572
rect -677 538 -661 572
rect -603 538 -587 572
rect -519 538 -503 572
rect -445 538 -429 572
rect -361 538 -345 572
rect -287 538 -271 572
rect -203 538 -187 572
rect -129 538 -113 572
rect -45 538 -29 572
rect 29 538 45 572
rect 113 538 129 572
rect 187 538 203 572
rect 271 538 287 572
rect 345 538 361 572
rect 429 538 445 572
rect 503 538 519 572
rect 587 538 603 572
rect 661 538 677 572
rect 745 538 761 572
rect 819 538 835 572
rect 903 538 919 572
rect 977 538 993 572
rect 1061 538 1077 572
rect 1135 538 1151 572
rect 1219 538 1235 572
rect 1293 538 1309 572
rect 1377 538 1393 572
rect 1451 538 1467 572
rect 1535 538 1551 572
rect -1597 488 -1563 504
rect -1597 -504 -1563 -488
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect 1563 488 1597 504
rect 1563 -504 1597 -488
rect -1551 -572 -1535 -538
rect -1467 -572 -1451 -538
rect -1393 -572 -1377 -538
rect -1309 -572 -1293 -538
rect -1235 -572 -1219 -538
rect -1151 -572 -1135 -538
rect -1077 -572 -1061 -538
rect -993 -572 -977 -538
rect -919 -572 -903 -538
rect -835 -572 -819 -538
rect -761 -572 -745 -538
rect -677 -572 -661 -538
rect -603 -572 -587 -538
rect -519 -572 -503 -538
rect -445 -572 -429 -538
rect -361 -572 -345 -538
rect -287 -572 -271 -538
rect -203 -572 -187 -538
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 187 -572 203 -538
rect 271 -572 287 -538
rect 345 -572 361 -538
rect 429 -572 445 -538
rect 503 -572 519 -538
rect 587 -572 603 -538
rect 661 -572 677 -538
rect 745 -572 761 -538
rect 819 -572 835 -538
rect 903 -572 919 -538
rect 977 -572 993 -538
rect 1061 -572 1077 -538
rect 1135 -572 1151 -538
rect 1219 -572 1235 -538
rect 1293 -572 1309 -538
rect 1377 -572 1393 -538
rect 1451 -572 1467 -538
rect 1535 -572 1551 -538
rect -1731 -676 -1697 -614
rect 1697 -676 1731 -614
rect -1731 -710 -1635 -676
rect 1635 -710 1731 -676
<< viali >>
rect -1519 538 -1485 572
rect -1361 538 -1327 572
rect -1203 538 -1169 572
rect -1045 538 -1011 572
rect -887 538 -853 572
rect -729 538 -695 572
rect -571 538 -537 572
rect -413 538 -379 572
rect -255 538 -221 572
rect -97 538 -63 572
rect 63 538 97 572
rect 221 538 255 572
rect 379 538 413 572
rect 537 538 571 572
rect 695 538 729 572
rect 853 538 887 572
rect 1011 538 1045 572
rect 1169 538 1203 572
rect 1327 538 1361 572
rect 1485 538 1519 572
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
rect -1519 -572 -1485 -538
rect -1361 -572 -1327 -538
rect -1203 -572 -1169 -538
rect -1045 -572 -1011 -538
rect -887 -572 -853 -538
rect -729 -572 -695 -538
rect -571 -572 -537 -538
rect -413 -572 -379 -538
rect -255 -572 -221 -538
rect -97 -572 -63 -538
rect 63 -572 97 -538
rect 221 -572 255 -538
rect 379 -572 413 -538
rect 537 -572 571 -538
rect 695 -572 729 -538
rect 853 -572 887 -538
rect 1011 -572 1045 -538
rect 1169 -572 1203 -538
rect 1327 -572 1361 -538
rect 1485 -572 1519 -538
<< metal1 >>
rect -1531 572 -1473 578
rect -1531 538 -1519 572
rect -1485 538 -1473 572
rect -1531 532 -1473 538
rect -1373 572 -1315 578
rect -1373 538 -1361 572
rect -1327 538 -1315 572
rect -1373 532 -1315 538
rect -1215 572 -1157 578
rect -1215 538 -1203 572
rect -1169 538 -1157 572
rect -1215 532 -1157 538
rect -1057 572 -999 578
rect -1057 538 -1045 572
rect -1011 538 -999 572
rect -1057 532 -999 538
rect -899 572 -841 578
rect -899 538 -887 572
rect -853 538 -841 572
rect -899 532 -841 538
rect -741 572 -683 578
rect -741 538 -729 572
rect -695 538 -683 572
rect -741 532 -683 538
rect -583 572 -525 578
rect -583 538 -571 572
rect -537 538 -525 572
rect -583 532 -525 538
rect -425 572 -367 578
rect -425 538 -413 572
rect -379 538 -367 572
rect -425 532 -367 538
rect -267 572 -209 578
rect -267 538 -255 572
rect -221 538 -209 572
rect -267 532 -209 538
rect -109 572 -51 578
rect -109 538 -97 572
rect -63 538 -51 572
rect -109 532 -51 538
rect 51 572 109 578
rect 51 538 63 572
rect 97 538 109 572
rect 51 532 109 538
rect 209 572 267 578
rect 209 538 221 572
rect 255 538 267 572
rect 209 532 267 538
rect 367 572 425 578
rect 367 538 379 572
rect 413 538 425 572
rect 367 532 425 538
rect 525 572 583 578
rect 525 538 537 572
rect 571 538 583 572
rect 525 532 583 538
rect 683 572 741 578
rect 683 538 695 572
rect 729 538 741 572
rect 683 532 741 538
rect 841 572 899 578
rect 841 538 853 572
rect 887 538 899 572
rect 841 532 899 538
rect 999 572 1057 578
rect 999 538 1011 572
rect 1045 538 1057 572
rect 999 532 1057 538
rect 1157 572 1215 578
rect 1157 538 1169 572
rect 1203 538 1215 572
rect 1157 532 1215 538
rect 1315 572 1373 578
rect 1315 538 1327 572
rect 1361 538 1373 572
rect 1315 532 1373 538
rect 1473 572 1531 578
rect 1473 538 1485 572
rect 1519 538 1531 572
rect 1473 532 1531 538
rect -1603 488 -1557 500
rect -1603 -488 -1597 488
rect -1563 -488 -1557 488
rect -1603 -500 -1557 -488
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect 1557 488 1603 500
rect 1557 -488 1563 488
rect 1597 -488 1603 488
rect 1557 -500 1603 -488
rect -1531 -538 -1473 -532
rect -1531 -572 -1519 -538
rect -1485 -572 -1473 -538
rect -1531 -578 -1473 -572
rect -1373 -538 -1315 -532
rect -1373 -572 -1361 -538
rect -1327 -572 -1315 -538
rect -1373 -578 -1315 -572
rect -1215 -538 -1157 -532
rect -1215 -572 -1203 -538
rect -1169 -572 -1157 -538
rect -1215 -578 -1157 -572
rect -1057 -538 -999 -532
rect -1057 -572 -1045 -538
rect -1011 -572 -999 -538
rect -1057 -578 -999 -572
rect -899 -538 -841 -532
rect -899 -572 -887 -538
rect -853 -572 -841 -538
rect -899 -578 -841 -572
rect -741 -538 -683 -532
rect -741 -572 -729 -538
rect -695 -572 -683 -538
rect -741 -578 -683 -572
rect -583 -538 -525 -532
rect -583 -572 -571 -538
rect -537 -572 -525 -538
rect -583 -578 -525 -572
rect -425 -538 -367 -532
rect -425 -572 -413 -538
rect -379 -572 -367 -538
rect -425 -578 -367 -572
rect -267 -538 -209 -532
rect -267 -572 -255 -538
rect -221 -572 -209 -538
rect -267 -578 -209 -572
rect -109 -538 -51 -532
rect -109 -572 -97 -538
rect -63 -572 -51 -538
rect -109 -578 -51 -572
rect 51 -538 109 -532
rect 51 -572 63 -538
rect 97 -572 109 -538
rect 51 -578 109 -572
rect 209 -538 267 -532
rect 209 -572 221 -538
rect 255 -572 267 -538
rect 209 -578 267 -572
rect 367 -538 425 -532
rect 367 -572 379 -538
rect 413 -572 425 -538
rect 367 -578 425 -572
rect 525 -538 583 -532
rect 525 -572 537 -538
rect 571 -572 583 -538
rect 525 -578 583 -572
rect 683 -538 741 -532
rect 683 -572 695 -538
rect 729 -572 741 -538
rect 683 -578 741 -572
rect 841 -538 899 -532
rect 841 -572 853 -538
rect 887 -572 899 -538
rect 841 -578 899 -572
rect 999 -538 1057 -532
rect 999 -572 1011 -538
rect 1045 -572 1057 -538
rect 999 -578 1057 -572
rect 1157 -538 1215 -532
rect 1157 -572 1169 -538
rect 1203 -572 1215 -538
rect 1157 -578 1215 -572
rect 1315 -538 1373 -532
rect 1315 -572 1327 -538
rect 1361 -572 1373 -538
rect 1315 -578 1373 -572
rect 1473 -538 1531 -532
rect 1473 -572 1485 -538
rect 1519 -572 1531 -538
rect 1473 -578 1531 -572
<< properties >>
string FIXED_BBOX -1714 -692 1714 692
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
