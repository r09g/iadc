magic
tech sky130A
magscale 1 2
timestamp 1655456512
<< error_p >>
rect -749 181 -691 187
rect -557 181 -499 187
rect -365 181 -307 187
rect -173 181 -115 187
rect 19 181 77 187
rect 211 181 269 187
rect 403 181 461 187
rect 595 181 653 187
rect -749 147 -737 181
rect -557 147 -545 181
rect -365 147 -353 181
rect -173 147 -161 181
rect 19 147 31 181
rect 211 147 223 181
rect 403 147 415 181
rect 595 147 607 181
rect -749 141 -691 147
rect -557 141 -499 147
rect -365 141 -307 147
rect -173 141 -115 147
rect 19 141 77 147
rect 211 141 269 147
rect 403 141 461 147
rect 595 141 653 147
rect -653 -147 -595 -141
rect -461 -147 -403 -141
rect -269 -147 -211 -141
rect -77 -147 -19 -141
rect 115 -147 173 -141
rect 307 -147 365 -141
rect 499 -147 557 -141
rect 691 -147 749 -141
rect -653 -181 -641 -147
rect -461 -181 -449 -147
rect -269 -181 -257 -147
rect -77 -181 -65 -147
rect 115 -181 127 -147
rect 307 -181 319 -147
rect 499 -181 511 -147
rect 691 -181 703 -147
rect -653 -187 -595 -181
rect -461 -187 -403 -181
rect -269 -187 -211 -181
rect -77 -187 -19 -181
rect 115 -187 173 -181
rect 307 -187 365 -181
rect 499 -187 557 -181
rect 691 -187 749 -181
<< nwell >>
rect -1031 -319 1031 319
<< pmos >>
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
<< pdiff >>
rect -893 88 -831 100
rect -893 -88 -881 88
rect -847 -88 -831 88
rect -893 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 893 100
rect 831 -88 847 88
rect 881 -88 893 88
rect 831 -100 893 -88
<< pdiffc >>
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
<< nsubdiff >>
rect -995 249 -899 283
rect 899 249 995 283
rect -995 187 -961 249
rect 961 187 995 249
rect -995 -249 -961 -187
rect 961 -249 995 -187
rect -995 -283 -899 -249
rect 899 -283 995 -249
<< nsubdiffcont >>
rect -899 249 899 283
rect -995 -187 -961 187
rect 961 -187 995 187
rect -899 -283 899 -249
<< poly >>
rect -753 181 -687 197
rect -753 147 -737 181
rect -703 147 -687 181
rect -753 131 -687 147
rect -561 181 -495 197
rect -561 147 -545 181
rect -511 147 -495 181
rect -561 131 -495 147
rect -369 181 -303 197
rect -369 147 -353 181
rect -319 147 -303 181
rect -369 131 -303 147
rect -177 181 -111 197
rect -177 147 -161 181
rect -127 147 -111 181
rect -177 131 -111 147
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect 207 181 273 197
rect 207 147 223 181
rect 257 147 273 181
rect 207 131 273 147
rect 399 181 465 197
rect 399 147 415 181
rect 449 147 465 181
rect 399 131 465 147
rect 591 181 657 197
rect 591 147 607 181
rect 641 147 657 181
rect 591 131 657 147
rect 783 181 849 197
rect 783 147 799 181
rect 833 147 849 181
rect 783 131 849 147
rect -831 100 -801 127
rect -735 100 -705 131
rect -639 100 -609 127
rect -543 100 -513 131
rect -447 100 -417 127
rect -351 100 -321 131
rect -255 100 -225 127
rect -159 100 -129 131
rect -63 100 -33 127
rect 33 100 63 131
rect 129 100 159 127
rect 225 100 255 131
rect 321 100 351 127
rect 417 100 447 131
rect 513 100 543 127
rect 609 100 639 131
rect 705 100 735 127
rect 801 100 831 131
rect -831 -131 -801 -100
rect -735 -127 -705 -100
rect -639 -131 -609 -100
rect -543 -127 -513 -100
rect -447 -131 -417 -100
rect -351 -127 -321 -100
rect -255 -131 -225 -100
rect -159 -127 -129 -100
rect -63 -131 -33 -100
rect 33 -127 63 -100
rect 129 -131 159 -100
rect 225 -127 255 -100
rect 321 -131 351 -100
rect 417 -127 447 -100
rect 513 -131 543 -100
rect 609 -127 639 -100
rect 705 -131 735 -100
rect 801 -127 831 -100
rect -849 -147 -783 -131
rect -849 -181 -833 -147
rect -799 -181 -783 -147
rect -849 -197 -783 -181
rect -657 -147 -591 -131
rect -657 -181 -641 -147
rect -607 -181 -591 -147
rect -657 -197 -591 -181
rect -465 -147 -399 -131
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -465 -197 -399 -181
rect -273 -147 -207 -131
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -273 -197 -207 -181
rect -81 -147 -15 -131
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect -81 -197 -15 -181
rect 111 -147 177 -131
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 111 -197 177 -181
rect 303 -147 369 -131
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 303 -197 369 -181
rect 495 -147 561 -131
rect 495 -181 511 -147
rect 545 -181 561 -147
rect 495 -197 561 -181
rect 687 -147 753 -131
rect 687 -181 703 -147
rect 737 -181 753 -147
rect 687 -197 753 -181
<< polycont >>
rect -737 147 -703 181
rect -545 147 -511 181
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect 607 147 641 181
rect 799 147 833 181
rect -833 -181 -799 -147
rect -641 -181 -607 -147
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
rect 511 -181 545 -147
rect 703 -181 737 -147
<< locali >>
rect -995 249 -899 283
rect 899 249 995 283
rect -995 187 -961 249
rect 847 181 881 249
rect -753 147 -737 181
rect -703 147 -687 181
rect -561 147 -545 181
rect -511 147 -495 181
rect -369 147 -353 181
rect -319 147 -303 181
rect -177 147 -161 181
rect -127 147 -111 181
rect 15 147 31 181
rect 65 147 81 181
rect 207 147 223 181
rect 257 147 273 181
rect 399 147 415 181
rect 449 147 465 181
rect 591 147 607 181
rect 641 147 657 181
rect 783 147 799 181
rect 833 147 881 181
rect -995 -249 -961 -187
rect -881 88 -847 104
rect -881 -147 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 147
rect 847 -104 881 -88
rect 961 187 995 249
rect -881 -181 -833 -147
rect -799 -181 -783 -147
rect -657 -181 -641 -147
rect -607 -181 -591 -147
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 495 -181 511 -147
rect 545 -181 561 -147
rect 687 -181 703 -147
rect 737 -181 753 -147
rect -881 -249 -847 -181
rect 961 -249 995 -187
rect -995 -283 -899 -249
rect 899 -283 995 -249
<< viali >>
rect -737 147 -703 181
rect -545 147 -511 181
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect 607 147 641 181
rect -641 -181 -607 -147
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
rect 511 -181 545 -147
rect 703 -181 737 -147
<< metal1 >>
rect -749 181 -691 187
rect -749 147 -737 181
rect -703 147 -691 181
rect -749 141 -691 147
rect -557 181 -499 187
rect -557 147 -545 181
rect -511 147 -499 181
rect -557 141 -499 147
rect -365 181 -307 187
rect -365 147 -353 181
rect -319 147 -307 181
rect -365 141 -307 147
rect -173 181 -115 187
rect -173 147 -161 181
rect -127 147 -115 181
rect -173 141 -115 147
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect 211 181 269 187
rect 211 147 223 181
rect 257 147 269 181
rect 211 141 269 147
rect 403 181 461 187
rect 403 147 415 181
rect 449 147 461 181
rect 403 141 461 147
rect 595 181 653 187
rect 595 147 607 181
rect 641 147 653 181
rect 595 141 653 147
rect -653 -147 -595 -141
rect -653 -181 -641 -147
rect -607 -181 -595 -147
rect -653 -187 -595 -181
rect -461 -147 -403 -141
rect -461 -181 -449 -147
rect -415 -181 -403 -147
rect -461 -187 -403 -181
rect -269 -147 -211 -141
rect -269 -181 -257 -147
rect -223 -181 -211 -147
rect -269 -187 -211 -181
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
rect 115 -147 173 -141
rect 115 -181 127 -147
rect 161 -181 173 -147
rect 115 -187 173 -181
rect 307 -147 365 -141
rect 307 -181 319 -147
rect 353 -181 365 -147
rect 307 -187 365 -181
rect 499 -147 557 -141
rect 499 -181 511 -147
rect 545 -181 557 -147
rect 499 -187 557 -181
rect 691 -147 749 -141
rect 691 -181 703 -147
rect 737 -181 749 -147
rect 691 -187 749 -181
<< properties >>
string FIXED_BBOX -978 -266 978 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
