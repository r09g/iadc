magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< locali >>
rect 15025 21777 15134 21811
rect 15410 21777 15611 21811
rect 18538 21777 18906 21811
rect 15025 21709 15059 21777
rect 15577 21675 15611 21777
rect 15577 21641 15686 21675
rect 18613 21641 18647 21777
rect 13202 21233 13495 21267
rect 16606 21233 16974 21267
rect 13461 21199 13495 21233
rect 17693 21199 17727 21403
rect 13461 21165 13647 21199
rect 17693 21165 17802 21199
rect 21206 21165 21315 21199
rect 22954 21097 23155 21131
rect 14289 20825 14398 20859
rect 14289 20689 14398 20723
rect 14289 20621 14323 20689
rect 15393 20655 15427 20859
rect 15333 20621 15427 20655
rect 23121 20553 23155 21097
rect 8861 19635 8895 19771
rect 8861 19601 8970 19635
rect 17325 19601 17618 19635
rect 9338 19533 9447 19567
rect 8234 19465 8343 19499
rect 8309 19397 8343 19465
rect 9413 19397 9447 19533
rect 15853 19465 15962 19499
rect 17325 19465 17359 19601
rect 15853 19397 15887 19465
rect 6469 19057 6578 19091
rect 6469 18853 6503 19057
rect 11546 18989 11638 19023
rect 21833 18479 21867 18683
rect 21833 18445 21942 18479
rect 7849 18071 7883 18139
rect 7774 18037 7883 18071
rect 16313 18003 16347 18139
rect 5917 17969 6394 18003
rect 16313 17969 16422 18003
rect 5917 17935 5951 17969
rect 5641 17901 5951 17935
rect 21281 17901 21390 17935
rect 5641 17459 5675 17901
rect 5641 17425 6026 17459
rect 19933 17425 20119 17459
rect 20085 17221 20119 17425
rect 13645 16813 13754 16847
rect 20453 16813 20562 16847
rect 13645 16745 13679 16813
rect 15778 16745 15887 16779
rect 20453 16677 20487 16813
rect 21114 16677 21223 16711
rect 12098 16337 12207 16371
rect 6578 16269 6670 16303
rect 12173 16201 12207 16337
rect 13185 16303 13219 16507
rect 17250 16473 17359 16507
rect 16514 16405 16623 16439
rect 22477 16303 22511 16507
rect 13110 16269 13219 16303
rect 22402 16269 22511 16303
rect 19441 15759 19475 15827
rect 8694 15725 8803 15759
rect 10902 15725 11270 15759
rect 18705 15725 18799 15759
rect 19366 15725 19475 15759
rect 8769 15589 8803 15725
rect 19625 15657 19734 15691
rect 11454 15589 11730 15623
rect 17509 15283 17543 15419
rect 7113 15249 7207 15283
rect 14766 15249 14950 15283
rect 17509 15249 17618 15283
rect 22017 15215 22051 15419
rect 22017 15181 22126 15215
rect 8769 14671 8803 14875
rect 20853 14841 20947 14875
rect 8341 14637 8435 14671
rect 8769 14637 8878 14671
rect 10885 14637 11063 14671
rect 18981 14297 19070 14331
rect 14766 14161 14875 14195
rect 20085 13957 20194 13991
rect 23121 13855 23155 14059
rect 23121 13821 23247 13855
rect 6193 13719 6227 13787
rect 6193 13685 6302 13719
rect 7222 13617 7314 13651
rect 12817 13583 12851 13719
rect 12742 13549 12851 13583
rect 6285 12087 6319 12155
rect 6285 12053 6394 12087
rect 16345 12053 16439 12087
rect 16054 11373 16255 11407
rect 16221 11237 16255 11373
rect 20361 11305 20470 11339
rect 23213 11067 23247 13821
rect 23489 11815 23523 18887
rect 23121 11033 23247 11067
rect 23397 11781 23523 11815
rect 23121 10829 23155 11033
rect 6561 10761 6670 10795
rect 6561 10693 6595 10761
rect 23397 10659 23431 11781
rect 23673 11679 23707 11883
rect 23627 11645 23707 11679
rect 23627 10659 23661 11645
rect 23305 10625 23431 10659
rect 23581 10625 23661 10659
rect 6561 10319 6595 10455
rect 18337 10319 18371 10523
rect 20913 10319 20947 10387
rect 6486 10285 6595 10319
rect 18262 10285 18371 10319
rect 20853 10285 20947 10319
rect 11753 10217 11839 10251
rect 6193 9843 6227 9979
rect 6745 9843 6779 9979
rect 6118 9809 6227 9843
rect 6285 9809 6394 9843
rect 6670 9809 6779 9843
rect 6285 9707 6319 9809
rect 19366 9741 19475 9775
rect 6118 9673 6319 9707
rect 19441 9605 19475 9741
rect 23305 9639 23339 10625
rect 23581 9775 23615 10625
rect 23765 9877 23799 19703
rect 23857 11203 23891 11407
rect 23857 11169 23937 11203
rect 23903 10523 23937 11169
rect 24041 10727 24075 10931
rect 24041 10693 24259 10727
rect 23903 10489 23983 10523
rect 23949 9775 23983 10489
rect 23581 9741 23707 9775
rect 23305 9605 23431 9639
rect 18262 9197 18371 9231
rect 20853 9197 20947 9231
rect 18337 9061 18371 9197
rect 20913 9061 20947 9197
rect 6854 8721 6963 8755
rect 7021 8721 7207 8755
rect 12098 8721 12391 8755
rect 7021 8517 7055 8721
rect 12357 8687 12391 8721
rect 12357 8653 12635 8687
rect 17509 8517 17543 8891
rect 6285 8279 6319 8347
rect 6285 8245 6394 8279
rect 20913 8143 20947 8347
rect 13294 8109 13647 8143
rect 20838 8109 20947 8143
rect 13461 7973 13495 8109
rect 23397 7939 23431 9605
rect 23397 7905 23523 7939
rect 5641 7769 5842 7803
rect 6854 7769 6963 7803
rect 5549 6579 5583 7055
rect 5641 6885 5675 7769
rect 23489 7701 23523 7905
rect 5733 7633 5842 7667
rect 6026 7633 6135 7667
rect 5733 7429 5767 7633
rect 6101 7429 6135 7633
rect 19826 7565 19935 7599
rect 12098 7497 12207 7531
rect 19901 7497 19935 7565
rect 23673 7531 23707 9741
rect 23581 7497 23707 7531
rect 23857 9741 23983 9775
rect 12173 7429 12207 7497
rect 18262 7089 18371 7123
rect 15594 6953 15795 6987
rect 18337 6885 18371 7089
rect 21114 7021 21223 7055
rect 23581 6919 23615 7497
rect 23857 7021 23891 9741
rect 24225 9639 24259 10693
rect 24133 9605 24259 9639
rect 24133 6919 24167 9605
rect 23581 6885 23707 6919
rect 23673 6681 23707 6885
rect 24041 6885 24167 6919
rect 7481 6579 7515 6647
rect 5549 6545 6026 6579
rect 6302 6545 6411 6579
rect 7481 6545 7575 6579
rect 6377 6477 6411 6545
rect 24041 6409 24075 6885
rect 7757 6103 7791 6171
rect 7757 6069 7866 6103
rect 10425 5967 10459 6171
rect 18001 6137 18095 6171
rect 13645 6069 13754 6103
rect 13645 5967 13679 6069
rect 17509 6001 17618 6035
rect 17509 5967 17543 6001
rect 10425 5933 10534 5967
rect 13478 5933 13679 5967
rect 17250 5933 17543 5967
<< metal1 >>
rect 5796 21984 23000 22080
rect 18432 21916 19104 21944
rect 19076 21876 19104 21916
rect 20732 21882 21404 21910
rect 20732 21876 20760 21882
rect 15212 21848 15792 21876
rect 15764 21808 15792 21848
rect 18432 21848 19012 21876
rect 19076 21848 20760 21876
rect 21376 21876 21404 21882
rect 21376 21848 21864 21876
rect 18432 21808 18460 21848
rect 15120 21780 15700 21808
rect 15764 21780 15976 21808
rect 16684 21780 17540 21808
rect 18248 21780 18460 21808
rect 16684 21740 16712 21780
rect 10263 21712 10350 21740
rect 14292 21712 15056 21740
rect 16500 21712 16712 21740
rect 17512 21740 17540 21780
rect 17512 21712 19748 21740
rect 20272 21672 20300 21808
rect 20548 21780 20576 21848
rect 21836 21808 21864 21848
rect 21008 21780 21312 21808
rect 21836 21780 22692 21808
rect 22756 21780 22876 21808
rect 20364 21712 20484 21740
rect 20548 21712 20944 21740
rect 21100 21712 21772 21740
rect 21947 21712 22034 21740
rect 20548 21672 20576 21712
rect 10079 21644 10166 21672
rect 15856 21644 16344 21672
rect 18432 21644 18644 21672
rect 19536 21644 20116 21672
rect 20272 21644 20576 21672
rect 20916 21672 20944 21712
rect 20916 21644 22784 21672
rect 15856 21604 15884 21644
rect 16316 21638 16344 21644
rect 16316 21610 17264 21638
rect 10447 21576 10534 21604
rect 15396 21576 15516 21604
rect 15672 21576 15884 21604
rect 17236 21604 17264 21610
rect 17236 21576 17448 21604
rect 19095 21576 19182 21604
rect 19831 21576 19918 21604
rect 19996 21576 20760 21604
rect 21560 21576 21680 21604
rect 22315 21576 22402 21604
rect 5796 21440 23000 21536
rect 10079 21372 10166 21400
rect 15875 21372 15962 21400
rect 17144 21372 17724 21400
rect 18156 21372 18276 21400
rect 19812 21372 20024 21400
rect 21468 21372 22048 21400
rect 17144 21304 17172 21372
rect 19812 21332 19840 21372
rect 19168 21304 19288 21332
rect 19720 21304 19840 21332
rect 22204 21304 22523 21332
rect 13372 21236 14044 21264
rect 15672 21236 16528 21264
rect 17347 21236 18000 21264
rect 19076 21236 19656 21264
rect 21468 21236 21758 21264
rect 10980 21168 13124 21196
rect 13372 21168 13400 21236
rect 15672 21196 15700 21236
rect 13832 21128 13860 21196
rect 14108 21168 14504 21196
rect 15120 21168 15700 21196
rect 15764 21168 15976 21196
rect 17144 21168 17356 21196
rect 17972 21168 18000 21236
rect 19812 21168 20116 21196
rect 21284 21168 21666 21196
rect 17328 21128 17356 21168
rect 13832 21100 14320 21128
rect 15503 21100 16160 21128
rect 17328 21100 18460 21128
rect 19996 21100 20096 21128
rect 19996 21060 20024 21100
rect 9968 21032 10088 21060
rect 12636 21032 12848 21060
rect 14311 21032 14398 21060
rect 14752 21032 15884 21060
rect 16151 21032 16238 21060
rect 17696 21032 18092 21060
rect 18819 21032 18906 21060
rect 19352 21032 20024 21060
rect 5796 20896 23000 20992
rect 10885 20761 10949 20868
rect 12603 20761 12667 20868
rect 14219 20828 14306 20856
rect 15396 20828 15516 20856
rect 20456 20828 20668 20856
rect 20640 20788 20668 20828
rect 21284 20828 21496 20856
rect 21284 20788 21312 20828
rect 13096 20760 14688 20788
rect 16151 20760 16252 20788
rect 18831 20760 18935 20788
rect 19904 20760 20377 20788
rect 20640 20760 21312 20788
rect 14660 20720 14688 20760
rect 7503 20692 7604 20720
rect 10888 20692 11192 20720
rect 12360 20692 12664 20720
rect 7227 20624 7314 20652
rect 13372 20624 14504 20652
rect 13372 20584 13400 20624
rect 11532 20556 12020 20584
rect 11992 20516 12020 20556
rect 13280 20556 13400 20584
rect 13280 20516 13308 20556
rect 14568 20516 14596 20720
rect 14660 20692 15148 20720
rect 21928 20692 22600 20720
rect 15875 20624 15962 20652
rect 19095 20624 19182 20652
rect 20015 20624 20102 20652
rect 21744 20624 22048 20652
rect 21560 20556 23152 20584
rect 8680 20488 9168 20516
rect 9784 20488 9996 20516
rect 11992 20488 13308 20516
rect 13372 20488 14596 20516
rect 14936 20488 15516 20516
rect 17144 20488 17356 20516
rect 17696 20488 17816 20516
rect 5796 20352 23000 20448
rect 10336 20284 11100 20312
rect 6767 20148 6854 20176
rect 10520 20148 10732 20176
rect 22867 20148 22954 20176
rect 12452 20080 16252 20108
rect 20088 20080 20208 20108
rect 20364 20080 21404 20108
rect 6932 20012 7129 20040
rect 7300 20012 8064 20040
rect 10183 20012 10287 20040
rect 12191 20012 12388 20040
rect 15319 20012 15516 20040
rect 16316 20012 16513 20040
rect 16684 20012 17448 20040
rect 7300 19972 7328 20012
rect 6748 19944 7328 19972
rect 8036 19972 8064 20012
rect 16684 19972 16712 20012
rect 8036 19944 8800 19972
rect 8956 19944 9168 19972
rect 13464 19944 14780 19972
rect 16040 19944 16712 19972
rect 17420 19972 17448 20012
rect 18064 20012 18644 20040
rect 18892 20012 19947 20040
rect 18064 19972 18092 20012
rect 17420 19944 17632 19972
rect 17880 19944 18092 19972
rect 18616 19972 18644 20012
rect 20364 19972 20392 20080
rect 18616 19944 18828 19972
rect 20180 19944 20392 19972
rect 21376 19972 21404 20080
rect 22679 20012 22968 20040
rect 21376 19944 21588 19972
rect 5796 19808 23000 19904
rect 7576 19740 7880 19768
rect 8864 19740 8984 19768
rect 9067 19740 9154 19768
rect 10244 19740 10364 19768
rect 15488 19740 16160 19768
rect 16243 19740 16330 19768
rect 16776 19740 16988 19768
rect 16960 19734 16988 19740
rect 17880 19740 18920 19768
rect 21100 19740 21312 19768
rect 17880 19734 17908 19740
rect 16960 19706 17908 19734
rect 21284 19700 21312 19740
rect 21836 19740 22048 19768
rect 21836 19700 21864 19740
rect 8772 19672 9076 19700
rect 12728 19672 13109 19700
rect 13280 19672 15056 19700
rect 21284 19672 21864 19700
rect 22219 19672 23796 19700
rect 13280 19632 13308 19672
rect 7024 19604 10548 19632
rect 11992 19604 12204 19632
rect 12360 19604 12572 19632
rect 12636 19604 12848 19632
rect 12912 19604 13308 19632
rect 15028 19632 15056 19672
rect 15028 19604 16896 19632
rect 17696 19604 17986 19632
rect 12544 19564 12572 19604
rect 12912 19564 12940 19604
rect 12544 19536 12940 19564
rect 22480 19536 22784 19564
rect 8128 19502 8892 19530
rect 8128 19496 8156 19502
rect 7944 19468 8156 19496
rect 8864 19496 8892 19502
rect 13924 19502 14964 19530
rect 13924 19496 13952 19502
rect 8864 19468 9076 19496
rect 10336 19468 10732 19496
rect 11992 19468 12388 19496
rect 13740 19468 13952 19496
rect 14936 19496 14964 19502
rect 14936 19468 15148 19496
rect 16408 19468 17356 19496
rect 13740 19428 13768 19468
rect 18041 19428 18069 19496
rect 8312 19400 8800 19428
rect 9416 19400 9996 19428
rect 11808 19400 11928 19428
rect 13188 19400 13768 19428
rect 14127 19400 14214 19428
rect 14568 19400 15884 19428
rect 17604 19400 18069 19428
rect 19076 19400 19288 19428
rect 5796 19264 23000 19360
rect 6859 19196 6946 19224
rect 10263 19196 10350 19224
rect 15948 19196 16344 19224
rect 10520 19128 11284 19156
rect 12084 19128 12365 19156
rect 13004 19128 13400 19156
rect 14200 19088 14228 19156
rect 14826 19116 14956 19168
rect 16316 19156 16344 19196
rect 17052 19196 17632 19224
rect 21100 19196 21312 19224
rect 17052 19156 17080 19196
rect 21284 19156 21312 19196
rect 21744 19196 22232 19224
rect 21744 19156 21772 19196
rect 16316 19128 17080 19156
rect 19260 19128 20093 19156
rect 21284 19128 21772 19156
rect 8956 19060 9720 19088
rect 9895 19060 9982 19088
rect 11348 19060 11744 19088
rect 11919 19060 12006 19088
rect 13110 19060 14228 19088
rect 14495 19060 14582 19088
rect 15686 19060 16160 19088
rect 11348 19020 11376 19060
rect 6748 18992 6960 19020
rect 10244 18992 11008 19020
rect 11256 18992 11376 19020
rect 11551 18992 11638 19020
rect 11808 18952 11836 19020
rect 13202 18992 13400 19020
rect 15778 18992 17172 19020
rect 17236 18992 17356 19020
rect 17497 18992 17908 19020
rect 22756 18992 22876 19020
rect 5736 18924 6316 18952
rect 11440 18924 11836 18952
rect 22587 18924 23520 18952
rect 5736 18680 5764 18924
rect 6288 18884 6316 18924
rect 6288 18856 6500 18884
rect 9508 18856 9996 18884
rect 10888 18856 11008 18884
rect 17788 18856 18644 18884
rect 19720 18856 20944 18884
rect 21284 18856 21496 18884
rect 23492 18856 23520 18924
rect 5796 18720 23000 18816
rect 5736 18652 6132 18680
rect 8312 18652 8800 18680
rect 12084 18652 12204 18680
rect 12544 18652 13216 18680
rect 19812 18652 20116 18680
rect 20916 18652 21864 18680
rect 22296 18652 22968 18680
rect 14016 18584 14872 18612
rect 16132 18584 17095 18612
rect 17604 18584 17724 18612
rect 17802 18584 17889 18612
rect 20180 18584 20377 18612
rect 7852 18550 8984 18578
rect 7852 18544 7880 18550
rect 6675 18516 6762 18544
rect 7668 18516 7880 18544
rect 8956 18544 8984 18550
rect 20548 18550 21128 18578
rect 20548 18544 20576 18550
rect 8956 18516 9168 18544
rect 10907 18516 11008 18544
rect 15580 18516 17540 18544
rect 17807 18516 17894 18544
rect 19352 18516 20576 18544
rect 21100 18544 21128 18550
rect 21652 18544 21680 18612
rect 21100 18516 21680 18544
rect 22112 18516 22968 18544
rect 6656 18408 6684 18476
rect 7944 18448 8248 18476
rect 8680 18448 8800 18476
rect 8975 18448 9062 18476
rect 10631 18448 10718 18476
rect 13662 18448 14596 18476
rect 17328 18448 17724 18476
rect 19628 18448 19840 18476
rect 19904 18448 20116 18476
rect 8220 18408 8248 18448
rect 6656 18380 7512 18408
rect 8220 18380 8616 18408
rect 12889 18380 13032 18408
rect 19812 18340 19840 18448
rect 6564 18312 6960 18340
rect 8864 18312 9444 18340
rect 15764 18312 15976 18340
rect 18064 18312 18460 18340
rect 18892 18312 19012 18340
rect 19812 18312 20392 18340
rect 21468 18312 21864 18340
rect 5796 18176 23000 18272
rect 7852 18108 8064 18136
rect 8036 18068 8064 18108
rect 8680 18108 8892 18136
rect 9048 18108 9720 18136
rect 13280 18108 15148 18136
rect 8680 18068 8708 18108
rect 12176 18074 12848 18102
rect 12176 18068 12204 18074
rect 6748 18040 7512 18068
rect 8036 18040 8708 18068
rect 11992 18040 12204 18068
rect 12820 18068 12848 18074
rect 15120 18068 15148 18108
rect 15856 18108 16344 18136
rect 21192 18108 26464 18136
rect 15856 18068 15884 18108
rect 12820 18040 13055 18068
rect 15120 18040 15884 18068
rect 16040 18040 16528 18068
rect 17623 18040 17710 18068
rect 9982 17972 10069 18000
rect 10428 17972 11192 18000
rect 11348 17972 11836 18000
rect 11900 17972 12112 18000
rect 10428 17932 10456 17972
rect 6564 17904 9628 17932
rect 9784 17904 9904 17932
rect 10244 17904 10456 17932
rect 11164 17932 11192 17972
rect 16592 17932 16620 18000
rect 22680 17972 22770 18000
rect 11164 17904 11652 17932
rect 14016 17904 14412 17932
rect 15488 17904 15608 17932
rect 15691 17904 15778 17932
rect 15870 17904 15957 17932
rect 16040 17904 16620 17932
rect 19736 17904 19826 17932
rect 20073 17904 20300 17932
rect 14384 17864 14412 17904
rect 20272 17864 20300 17904
rect 20824 17904 21496 17932
rect 22419 17904 22523 17932
rect 20824 17864 20852 17904
rect 14219 17836 14320 17864
rect 14384 17836 14504 17864
rect 15672 17836 16344 17864
rect 20272 17836 20852 17864
rect 7116 17768 7420 17796
rect 10336 17768 10548 17796
rect 10980 17768 11468 17796
rect 13299 17768 13386 17796
rect 14844 17768 15424 17796
rect 21192 17768 21496 17796
rect 5796 17632 23000 17728
rect 9600 17564 10456 17592
rect 12176 17564 12940 17592
rect 14752 17564 14964 17592
rect 9416 17496 10180 17524
rect 7208 17428 7328 17456
rect 7411 17428 7512 17456
rect 8864 17428 9168 17456
rect 9232 17388 9260 17456
rect 10152 17428 10180 17496
rect 10428 17428 10456 17564
rect 12912 17524 12940 17564
rect 14936 17524 14964 17564
rect 20272 17564 20760 17592
rect 11256 17496 11928 17524
rect 12912 17496 13661 17524
rect 14108 17496 14596 17524
rect 14936 17496 15424 17524
rect 18340 17496 18920 17524
rect 19734 17496 19821 17524
rect 11256 17456 11284 17496
rect 10704 17428 10824 17456
rect 11057 17428 11284 17456
rect 11900 17456 11928 17496
rect 14568 17456 14596 17496
rect 18340 17456 18368 17496
rect 11900 17428 12112 17456
rect 12084 17388 12112 17428
rect 12728 17428 12940 17456
rect 13004 17428 13124 17456
rect 13372 17428 14504 17456
rect 14568 17428 15332 17456
rect 15488 17428 15608 17456
rect 15686 17428 15773 17456
rect 15948 17428 16988 17456
rect 17696 17428 17908 17456
rect 18141 17428 18368 17456
rect 12728 17388 12756 17428
rect 6491 17360 6578 17388
rect 6656 17360 7236 17388
rect 7208 17252 7236 17360
rect 8864 17360 9260 17388
rect 10244 17360 10364 17388
rect 12084 17360 12756 17388
rect 8864 17252 8892 17360
rect 13280 17292 13400 17320
rect 15304 17252 15332 17428
rect 15580 17388 15608 17428
rect 15948 17388 15976 17428
rect 15580 17360 15976 17388
rect 16960 17388 16988 17428
rect 18892 17388 18920 17496
rect 20272 17456 20300 17564
rect 20732 17524 20760 17564
rect 21376 17564 21864 17592
rect 21376 17524 21404 17564
rect 20732 17496 21404 17524
rect 19463 17428 19550 17456
rect 19628 17428 20300 17456
rect 22143 17428 22247 17456
rect 22480 17428 22784 17456
rect 16960 17360 17172 17388
rect 18892 17360 19472 17388
rect 19444 17354 19472 17360
rect 19444 17326 20576 17354
rect 20548 17320 20576 17326
rect 16132 17292 16712 17320
rect 19076 17292 19288 17320
rect 20548 17292 21128 17320
rect 16132 17252 16160 17292
rect 6767 17224 6854 17252
rect 7208 17224 8892 17252
rect 9048 17224 9168 17252
rect 10336 17224 10640 17252
rect 14752 17224 15148 17252
rect 15304 17224 16160 17252
rect 16684 17252 16712 17292
rect 17052 17258 17724 17286
rect 17052 17252 17080 17258
rect 16684 17224 17080 17252
rect 17696 17252 17724 17258
rect 17696 17224 17908 17252
rect 18616 17224 19380 17252
rect 20088 17224 20208 17252
rect 5796 17088 23000 17184
rect 9508 17020 10180 17048
rect 11275 17020 11362 17048
rect 11919 17020 12006 17048
rect 14292 17020 15332 17048
rect 16316 17020 16804 17048
rect 19720 17020 20208 17048
rect 12084 16952 13047 16980
rect 10815 16884 10902 16912
rect 11716 16884 11928 16912
rect 11900 16844 11928 16884
rect 14016 16884 14320 16912
rect 18083 16884 18828 16912
rect 20088 16884 23520 16912
rect 10336 16816 10655 16844
rect 11532 16816 11652 16844
rect 11735 16816 11822 16844
rect 11900 16816 12190 16844
rect 13280 16816 13952 16844
rect 14016 16816 14044 16884
rect 14122 16816 14209 16844
rect 14384 16816 14504 16844
rect 14587 16816 14688 16844
rect 15396 16816 15608 16844
rect 16040 16816 16528 16844
rect 18432 16816 19089 16844
rect 20843 16816 20930 16844
rect 15396 16776 15424 16816
rect 16040 16776 16068 16816
rect 13648 16748 15424 16776
rect 15856 16748 16068 16776
rect 16500 16776 16528 16816
rect 16500 16748 16712 16776
rect 17788 16748 17923 16776
rect 20659 16748 20746 16776
rect 20824 16748 21496 16776
rect 13096 16680 13400 16708
rect 20088 16680 20484 16708
rect 21008 16680 21220 16708
rect 5796 16544 23000 16640
rect 8772 16476 8892 16504
rect 11624 16476 11836 16504
rect 13096 16476 13216 16504
rect 13280 16476 13400 16504
rect 15764 16476 16068 16504
rect 16684 16476 16988 16504
rect 17328 16476 17816 16504
rect 19904 16476 20760 16504
rect 21468 16476 21680 16504
rect 22020 16476 22232 16504
rect 22388 16476 22508 16504
rect 10603 16436 10631 16446
rect 7024 16408 7681 16436
rect 7944 16408 9168 16436
rect 10603 16408 11008 16436
rect 6123 16340 6210 16368
rect 6840 16340 6960 16368
rect 7300 16340 7420 16368
rect 8975 16340 9062 16368
rect 9140 16340 9168 16408
rect 12820 16368 12848 16436
rect 14491 16408 14872 16436
rect 15323 16408 15424 16436
rect 16040 16368 16068 16476
rect 16592 16408 16896 16436
rect 16960 16408 16988 16476
rect 18616 16408 18813 16436
rect 20291 16408 20392 16436
rect 10336 16340 10640 16368
rect 11624 16340 11836 16368
rect 11900 16340 12020 16368
rect 12820 16340 13400 16368
rect 14752 16340 15976 16368
rect 16040 16340 16712 16368
rect 16868 16340 17080 16368
rect 19904 16340 20116 16368
rect 6288 16272 6776 16300
rect 8791 16272 8878 16300
rect 9416 16272 9996 16300
rect 16868 16272 16896 16340
rect 17972 16272 18552 16300
rect 22204 16272 22968 16300
rect 6748 16232 6776 16272
rect 6748 16204 7420 16232
rect 9159 16204 9246 16232
rect 9784 16204 10272 16232
rect 11716 16204 12204 16232
rect 7392 16164 7420 16204
rect 7392 16136 8800 16164
rect 9048 16136 9168 16164
rect 9600 16136 10088 16164
rect 10152 16136 11008 16164
rect 12655 16136 12742 16164
rect 21284 16136 21496 16164
rect 5796 16000 23000 16096
rect 6932 15932 8064 15960
rect 8588 15932 8892 15960
rect 9416 15932 11192 15960
rect 11735 15932 11822 15960
rect 13004 15932 14044 15960
rect 8036 15892 8064 15932
rect 8036 15864 8616 15892
rect 8975 15864 9062 15892
rect 8588 15756 8616 15864
rect 6932 15728 7236 15756
rect 7484 15679 7512 15756
rect 7944 15728 8524 15756
rect 8588 15728 9260 15756
rect 9435 15728 9522 15756
rect 9769 15728 10088 15756
rect 10796 15728 11008 15756
rect 11348 15728 11652 15756
rect 12084 15728 12388 15756
rect 11348 15688 11376 15728
rect 14016 15688 14044 15932
rect 16868 15864 17816 15892
rect 17788 15824 17816 15864
rect 18432 15864 18828 15892
rect 18432 15824 18460 15864
rect 16611 15796 16698 15824
rect 17788 15796 18460 15824
rect 18800 15756 18828 15864
rect 19444 15796 20116 15824
rect 22683 15796 22770 15824
rect 14384 15728 14504 15756
rect 16500 15728 16988 15756
rect 17420 15688 17448 15742
rect 18616 15728 18736 15756
rect 18800 15728 19012 15756
rect 19090 15728 19177 15756
rect 20839 15728 21036 15756
rect 21100 15728 21496 15756
rect 7199 15651 7512 15679
rect 10428 15660 11376 15688
rect 12345 15660 12480 15688
rect 14016 15660 14673 15688
rect 14844 15660 15608 15688
rect 17328 15660 17448 15688
rect 14844 15620 14872 15660
rect 8312 15592 8800 15620
rect 10244 15592 11376 15620
rect 14292 15592 14872 15620
rect 15580 15620 15608 15660
rect 18984 15620 19012 15728
rect 19168 15660 19656 15688
rect 21928 15660 22523 15688
rect 15580 15592 15792 15620
rect 17715 15592 17802 15620
rect 18984 15592 19104 15620
rect 21376 15592 21772 15620
rect 5796 15456 23000 15552
rect 6104 15388 6224 15416
rect 9232 15388 9996 15416
rect 16316 15348 16344 15416
rect 16960 15388 17540 15416
rect 18984 15388 19196 15416
rect 19168 15348 19196 15388
rect 20916 15388 21404 15416
rect 20916 15348 20944 15388
rect 21376 15348 21404 15388
rect 21836 15388 22048 15416
rect 21836 15348 21864 15388
rect 8327 15320 9076 15348
rect 12084 15320 12204 15348
rect 14016 15320 15225 15348
rect 16316 15320 16712 15348
rect 19168 15320 20944 15348
rect 21100 15320 21235 15348
rect 21376 15320 21864 15348
rect 14016 15280 14044 15320
rect 6564 15252 6868 15280
rect 6932 15252 7972 15280
rect 8588 15252 8708 15280
rect 8864 15252 8984 15280
rect 10152 15252 10272 15280
rect 10336 15252 10994 15280
rect 12636 15252 14044 15280
rect 14306 15252 14780 15280
rect 15672 15252 16436 15280
rect 16500 15252 16620 15280
rect 16776 15252 16896 15280
rect 18616 15252 18813 15280
rect 6932 15212 6960 15252
rect 16500 15212 16528 15252
rect 6288 15184 6960 15212
rect 10442 15184 10529 15212
rect 10631 15184 10718 15212
rect 13115 15184 13202 15212
rect 16040 15184 16528 15212
rect 17972 15184 18552 15212
rect 21395 15184 21482 15212
rect 22223 15184 22310 15212
rect 6932 15116 7696 15144
rect 7668 15076 7696 15116
rect 8588 15116 8708 15144
rect 8588 15076 8616 15116
rect 7668 15048 8616 15076
rect 11057 15076 11085 15144
rect 13188 15116 13400 15144
rect 14403 15116 14490 15144
rect 19812 15116 20116 15144
rect 13188 15076 13216 15116
rect 13556 15082 14228 15110
rect 13556 15076 13584 15082
rect 11057 15048 11376 15076
rect 12820 15048 13584 15076
rect 14200 15076 14228 15082
rect 14200 15048 16344 15076
rect 16960 15048 17356 15076
rect 19904 15048 20024 15076
rect 22407 15048 22494 15076
rect 5796 14912 23000 15008
rect 8772 14844 10180 14872
rect 10336 14844 10456 14872
rect 10704 14844 10916 14872
rect 10888 14804 10916 14844
rect 11348 14844 12480 14872
rect 17420 14844 17632 14872
rect 20916 14844 21036 14872
rect 11348 14804 11376 14844
rect 9048 14776 9329 14804
rect 10888 14776 11376 14804
rect 12452 14804 12480 14844
rect 12452 14776 13676 14804
rect 20364 14776 21404 14804
rect 6859 14708 6946 14736
rect 8404 14708 9154 14736
rect 6748 14640 7221 14668
rect 8404 14640 8432 14708
rect 10166 14640 10916 14668
rect 10980 14640 11468 14668
rect 11440 14600 11468 14640
rect 11992 14640 12219 14668
rect 12360 14640 12480 14668
rect 13372 14640 13860 14668
rect 14403 14640 14490 14668
rect 16151 14640 16238 14668
rect 16427 14640 16528 14668
rect 17328 14640 18092 14668
rect 11992 14600 12020 14640
rect 17328 14600 17356 14640
rect 7392 14572 8156 14600
rect 11440 14572 12020 14600
rect 14568 14572 14765 14600
rect 15212 14572 16068 14600
rect 7392 14566 7420 14572
rect 6748 14538 7420 14566
rect 6748 14532 6776 14538
rect 6564 14504 6776 14532
rect 8128 14532 8156 14572
rect 8128 14504 8340 14532
rect 13464 14504 14044 14532
rect 14568 14504 14596 14572
rect 16040 14566 16068 14572
rect 16592 14572 17356 14600
rect 18064 14600 18092 14640
rect 18230 14631 18294 14748
rect 18727 14708 18814 14736
rect 20456 14708 20576 14736
rect 22680 14708 22770 14736
rect 20088 14640 20392 14668
rect 20548 14640 20576 14708
rect 18064 14572 18644 14600
rect 16592 14566 16620 14572
rect 16040 14538 16620 14566
rect 18966 14560 19099 14612
rect 19996 14572 20484 14600
rect 15783 14504 15870 14532
rect 20107 14504 20194 14532
rect 20640 14504 20668 14651
rect 22419 14640 22523 14668
rect 5796 14368 23000 14464
rect 10612 14300 10824 14328
rect 11808 14300 12020 14328
rect 11992 14294 12020 14300
rect 12820 14300 14596 14328
rect 17144 14300 17540 14328
rect 18911 14300 18998 14328
rect 21928 14300 22048 14328
rect 12820 14294 12848 14300
rect 11992 14266 12848 14294
rect 12989 14232 13492 14260
rect 14292 14232 14504 14260
rect 6491 14164 6578 14192
rect 7300 14164 7880 14192
rect 7944 14164 8141 14192
rect 11164 14164 12848 14192
rect 14200 14124 14228 14192
rect 14311 14164 14398 14192
rect 14495 14164 14582 14192
rect 14844 14164 15240 14192
rect 16776 14164 16988 14192
rect 18555 14164 18659 14192
rect 18800 14164 18920 14192
rect 19076 14164 19288 14192
rect 6656 14096 6960 14124
rect 12176 14096 12756 14124
rect 14200 14096 14412 14124
rect 14384 14056 14412 14096
rect 15212 14096 15608 14124
rect 16606 14096 16693 14124
rect 15212 14056 15240 14096
rect 14384 14028 15240 14056
rect 15415 14028 15502 14056
rect 19352 13988 19380 14192
rect 19444 14124 19472 14192
rect 19628 14164 20392 14192
rect 21223 14164 21327 14192
rect 21468 14164 21588 14192
rect 22204 14164 22324 14192
rect 19444 14096 19932 14124
rect 22388 14028 23152 14056
rect 5736 13960 6316 13988
rect 9140 13960 9260 13988
rect 10796 13960 11836 13988
rect 19352 13960 22968 13988
rect 5736 13784 5764 13960
rect 5796 13824 23000 13920
rect 5736 13756 6224 13784
rect 6656 13756 6776 13784
rect 7668 13756 7972 13784
rect 9048 13756 9352 13784
rect 11256 13756 11376 13784
rect 14384 13756 14596 13784
rect 10244 13688 10387 13716
rect 10796 13688 12319 13716
rect 12820 13688 13860 13716
rect 14568 13648 14596 13756
rect 16040 13756 16252 13784
rect 18267 13756 18354 13784
rect 20180 13756 21772 13784
rect 16040 13648 16068 13756
rect 19812 13688 20300 13716
rect 6380 13620 6776 13648
rect 6840 13620 9591 13648
rect 12466 13620 12572 13648
rect 12728 13620 12940 13648
rect 14568 13620 16068 13648
rect 17604 13620 18000 13648
rect 18724 13620 18814 13648
rect 6472 13444 6500 13580
rect 6840 13512 6868 13620
rect 6932 13552 7052 13580
rect 6748 13484 6868 13512
rect 7484 13444 7512 13580
rect 10980 13552 11454 13580
rect 12636 13552 14044 13580
rect 17788 13552 18184 13580
rect 12636 13444 12664 13552
rect 19812 13512 19840 13688
rect 20456 13654 20944 13682
rect 20456 13648 20484 13654
rect 19904 13620 20484 13648
rect 20916 13648 20944 13654
rect 21376 13648 21404 13716
rect 20916 13620 21404 13648
rect 22680 13620 22770 13648
rect 20383 13552 20470 13580
rect 20732 13552 20852 13580
rect 22419 13552 22523 13580
rect 17144 13484 17371 13512
rect 19061 13484 19840 13512
rect 20475 13484 20562 13512
rect 20640 13444 20668 13512
rect 6196 13416 7512 13444
rect 10631 13416 10718 13444
rect 11624 13416 12664 13444
rect 13004 13416 13308 13444
rect 13464 13416 14228 13444
rect 20180 13416 20668 13444
rect 5796 13280 23000 13376
rect 6656 13212 6960 13240
rect 8680 13212 8892 13240
rect 8864 13172 8892 13212
rect 9324 13212 9720 13240
rect 9324 13172 9352 13212
rect 9692 13206 9720 13212
rect 10428 13212 10916 13240
rect 12544 13212 14228 13240
rect 15948 13212 16068 13240
rect 17328 13212 17448 13240
rect 20088 13212 20576 13240
rect 21744 13212 21956 13240
rect 10428 13206 10456 13212
rect 9692 13178 10456 13206
rect 7760 13144 8432 13172
rect 8864 13144 9352 13172
rect 10612 13144 10824 13172
rect 7760 13104 7788 13144
rect 6380 13076 6592 13104
rect 6675 13076 6762 13104
rect 7561 13076 7788 13104
rect 8404 13104 8432 13144
rect 8404 13076 8616 13104
rect 8588 13036 8616 13076
rect 9876 13076 10088 13104
rect 10888 13090 10916 13212
rect 17420 13172 17448 13212
rect 12176 13144 12756 13172
rect 13081 13144 13492 13172
rect 14568 13144 15424 13172
rect 15488 13144 16160 13172
rect 17420 13144 18659 13172
rect 21215 13144 21680 13172
rect 21928 13144 21956 13212
rect 13372 13076 13860 13104
rect 15231 13076 15318 13104
rect 15580 13076 15700 13104
rect 17067 13076 17264 13104
rect 17328 13076 17540 13104
rect 18800 13076 18920 13104
rect 20456 13076 21772 13104
rect 21850 13076 21937 13104
rect 22020 13076 22140 13104
rect 9876 13036 9904 13076
rect 13832 13036 13860 13076
rect 7227 13008 7314 13036
rect 8588 13008 9904 13036
rect 10060 13008 10272 13036
rect 10428 13008 10732 13036
rect 11914 13008 12020 13036
rect 12360 13008 12848 13036
rect 13832 13008 14780 13036
rect 21395 13008 21482 13036
rect 10060 12940 10088 13008
rect 14752 12968 14780 13008
rect 14936 12974 15792 13002
rect 14936 12968 14964 12974
rect 10796 12940 11767 12968
rect 14752 12940 14964 12968
rect 15764 12968 15792 12974
rect 15764 12940 16436 12968
rect 16408 12900 16436 12940
rect 15120 12872 15700 12900
rect 16408 12872 17080 12900
rect 17439 12872 17526 12900
rect 20180 12872 21588 12900
rect 5796 12736 23000 12832
rect 8772 12668 8984 12696
rect 8956 12662 8984 12668
rect 9600 12668 10272 12696
rect 11900 12668 13676 12696
rect 16776 12668 16988 12696
rect 17071 12668 17158 12696
rect 21652 12668 22968 12696
rect 9600 12662 9628 12668
rect 8956 12634 9628 12662
rect 9807 12600 10456 12628
rect 13648 12560 13676 12668
rect 16040 12600 16620 12628
rect 16040 12560 16068 12600
rect 7484 12532 9062 12560
rect 13207 12532 13294 12560
rect 13648 12532 13768 12560
rect 15856 12532 16068 12560
rect 16592 12560 16620 12600
rect 16592 12532 16896 12560
rect 7484 12492 7512 12532
rect 13740 12492 13768 12532
rect 6380 12464 6500 12492
rect 6578 12464 6665 12492
rect 7116 12464 7512 12492
rect 8864 12464 8970 12492
rect 12943 12464 13047 12492
rect 13464 12464 13676 12492
rect 13740 12464 13937 12492
rect 15580 12464 16620 12492
rect 16868 12464 16896 12532
rect 16960 12492 16988 12668
rect 18616 12532 18828 12560
rect 16960 12464 17172 12492
rect 19168 12464 19932 12492
rect 20107 12464 20194 12492
rect 21027 12464 21404 12492
rect 22480 12464 23060 12492
rect 6472 12424 6500 12464
rect 6472 12396 6960 12424
rect 18355 12396 19012 12424
rect 15212 12362 16620 12390
rect 15212 12356 15240 12362
rect 5736 12328 6500 12356
rect 10152 12328 10272 12356
rect 15028 12328 15240 12356
rect 16592 12356 16620 12362
rect 19168 12356 19196 12464
rect 19904 12390 19932 12464
rect 22480 12424 22508 12464
rect 21579 12396 21680 12424
rect 21836 12396 22508 12424
rect 19904 12362 20944 12390
rect 16592 12328 16804 12356
rect 17236 12328 19196 12356
rect 20916 12356 20944 12362
rect 21836 12356 21864 12396
rect 20916 12328 21864 12356
rect 23032 12356 23060 12464
rect 23032 12328 28764 12356
rect 5736 12152 5764 12328
rect 5796 12192 23000 12288
rect 5736 12124 6316 12152
rect 6564 12124 6776 12152
rect 8791 12124 9076 12152
rect 9048 12084 9076 12124
rect 10428 12124 10916 12152
rect 14568 12124 14780 12152
rect 16776 12124 17080 12152
rect 21560 12124 21680 12152
rect 10428 12118 10456 12124
rect 9508 12090 10456 12118
rect 9508 12084 9536 12090
rect 7944 12056 8524 12084
rect 9048 12056 9536 12084
rect 10612 12056 10824 12084
rect 7944 12016 7972 12056
rect 6564 11988 6684 12016
rect 7745 11988 7972 12016
rect 8496 12016 8524 12056
rect 8496 11988 8708 12016
rect 8680 11948 8708 11988
rect 9692 11988 9904 12016
rect 10888 12002 10916 12124
rect 11900 12056 12296 12084
rect 9692 11948 9720 11988
rect 7300 11920 7512 11948
rect 8680 11920 9720 11948
rect 9987 11920 10074 11948
rect 10171 11920 10258 11948
rect 11900 11934 11928 12056
rect 12268 12016 12296 12056
rect 13096 12056 13661 12084
rect 15197 12056 15700 12084
rect 16408 12056 16988 12084
rect 17052 12056 17080 12124
rect 17512 12056 17908 12084
rect 17986 12056 18073 12084
rect 18785 12056 20116 12084
rect 13096 12016 13124 12056
rect 12268 11988 13124 12016
rect 13372 11988 13492 12016
rect 14936 11988 15516 12016
rect 15580 11988 16804 12016
rect 17071 11988 17816 12016
rect 11992 11920 12112 11948
rect 16500 11880 16528 11988
rect 18156 11880 18184 12016
rect 21131 11988 21235 12016
rect 18451 11920 18538 11948
rect 21395 11920 21482 11948
rect 21744 11920 22232 11948
rect 22388 11920 23060 11948
rect 22388 11880 22416 11920
rect 10612 11852 10824 11880
rect 10796 11846 10824 11852
rect 11532 11852 11767 11880
rect 16500 11852 16804 11880
rect 17255 11852 17342 11880
rect 17420 11852 18276 11880
rect 21928 11852 22416 11880
rect 23032 11880 23060 11920
rect 23032 11852 23704 11880
rect 11532 11846 11560 11852
rect 10796 11818 11560 11846
rect 16776 11812 16804 11852
rect 17420 11812 17448 11852
rect 6307 11784 6394 11812
rect 16776 11784 17448 11812
rect 17531 11784 17618 11812
rect 19904 11784 20024 11812
rect 20088 11784 21772 11812
rect 5796 11648 23000 11744
rect 7944 11580 8340 11608
rect 10428 11580 10640 11608
rect 13280 11580 13492 11608
rect 6380 11512 6500 11540
rect 8864 11512 9605 11540
rect 11440 11512 12020 11540
rect 20180 11512 21680 11540
rect 9416 11404 9444 11458
rect 13943 11444 14030 11472
rect 22683 11444 22770 11472
rect 6196 11376 6684 11404
rect 6932 11376 7236 11404
rect 8680 11376 9444 11404
rect 10442 11376 10548 11404
rect 11551 11376 11638 11404
rect 12084 11376 12388 11404
rect 14277 11376 14596 11404
rect 15415 11376 15502 11404
rect 15783 11376 15870 11404
rect 16795 11376 16882 11404
rect 17129 11376 17632 11404
rect 18064 11376 18552 11404
rect 18727 11376 18814 11404
rect 20456 11376 20668 11404
rect 21008 11376 21220 11404
rect 22495 11376 23888 11404
rect 18064 11336 18092 11376
rect 6840 11308 7216 11336
rect 11808 11308 12368 11336
rect 15672 11268 15700 11336
rect 15778 11308 15865 11336
rect 17880 11308 18092 11336
rect 18524 11336 18552 11376
rect 18524 11308 19089 11336
rect 19168 11308 20392 11336
rect 20456 11308 20484 11376
rect 20548 11308 20760 11336
rect 20838 11308 20925 11336
rect 16408 11274 17172 11302
rect 16408 11268 16436 11274
rect 9048 11240 9260 11268
rect 15396 11240 15700 11268
rect 16224 11240 16436 11268
rect 17144 11268 17172 11274
rect 17144 11240 17356 11268
rect 17880 11240 17908 11308
rect 18064 11240 18276 11268
rect 21303 11240 21390 11268
rect 5796 11104 23000 11200
rect 11348 11036 11928 11064
rect 14752 11036 14964 11064
rect 14936 10996 14964 11036
rect 15488 11036 15792 11064
rect 19720 11036 19932 11064
rect 15488 10996 15516 11036
rect 19904 11030 19932 11036
rect 20640 11036 20852 11064
rect 20640 11030 20668 11036
rect 19904 11002 20668 11030
rect 10428 10968 10640 10996
rect 13280 10968 13661 10996
rect 14936 10968 15516 10996
rect 18800 10968 19380 10996
rect 21100 10968 21404 10996
rect 22296 10968 23244 10996
rect 6656 10900 6868 10928
rect 7024 10900 7589 10928
rect 9140 10900 10088 10928
rect 10520 10900 10718 10928
rect 13280 10860 13308 10968
rect 18800 10928 18828 10968
rect 13372 10900 13492 10928
rect 15948 10900 16359 10928
rect 18340 10900 18460 10928
rect 18601 10900 18828 10928
rect 19352 10928 19380 10968
rect 22296 10928 22324 10968
rect 19352 10900 20208 10928
rect 22112 10900 22324 10928
rect 23216 10928 23244 10968
rect 23216 10900 24072 10928
rect 7227 10832 7314 10860
rect 8956 10832 9076 10860
rect 11730 10832 13308 10860
rect 16592 10832 16896 10860
rect 21395 10832 21482 10860
rect 21928 10832 22048 10860
rect 22480 10832 23152 10860
rect 5736 10764 6408 10792
rect 10888 10764 11583 10792
rect 14476 10764 15240 10792
rect 5736 10520 5764 10764
rect 6380 10724 6408 10764
rect 6380 10696 6592 10724
rect 8607 10696 8694 10724
rect 9048 10696 9352 10724
rect 14476 10696 14504 10764
rect 21560 10730 23060 10758
rect 21560 10724 21588 10730
rect 20088 10696 21588 10724
rect 23032 10724 23060 10730
rect 23032 10696 26280 10724
rect 5796 10560 23000 10656
rect 5736 10492 6684 10520
rect 10520 10492 10640 10520
rect 13280 10492 13492 10520
rect 14016 10492 14596 10520
rect 16132 10492 16252 10520
rect 18248 10492 20208 10520
rect 20286 10492 20373 10520
rect 20180 10452 20208 10492
rect 6564 10424 7328 10452
rect 7300 10384 7328 10424
rect 8496 10424 8708 10452
rect 11275 10424 11362 10452
rect 17623 10424 17710 10452
rect 20180 10424 20944 10452
rect 8496 10384 8524 10424
rect 20916 10384 20944 10424
rect 6380 10356 6960 10384
rect 7300 10356 8524 10384
rect 11532 10356 11652 10384
rect 6380 10316 6408 10356
rect 6932 10316 6960 10356
rect 17972 10316 18000 10384
rect 18724 10356 18814 10384
rect 20916 10356 21312 10384
rect 5736 10288 6408 10316
rect 5736 9976 5764 10288
rect 6840 10248 6868 10316
rect 6932 10288 7144 10316
rect 9140 10288 9260 10316
rect 12084 10288 12388 10316
rect 13280 10288 14228 10316
rect 14384 10288 14504 10316
rect 14568 10288 15332 10316
rect 16040 10288 17632 10316
rect 17880 10288 18000 10316
rect 18078 10288 18165 10316
rect 20364 10288 20484 10316
rect 20567 10288 20654 10316
rect 21376 10288 21496 10316
rect 21560 10288 23244 10316
rect 21560 10248 21588 10288
rect 6380 10220 6868 10248
rect 9048 10220 9521 10248
rect 11808 10220 12368 10248
rect 14292 10180 14320 10248
rect 15779 10220 16160 10248
rect 17267 10220 17371 10248
rect 17512 10220 18000 10248
rect 18524 10220 19089 10248
rect 20548 10220 21588 10248
rect 21637 10220 21956 10248
rect 17512 10180 17540 10220
rect 18524 10180 18552 10220
rect 14292 10152 14596 10180
rect 14660 10152 14964 10180
rect 17236 10152 17540 10180
rect 18156 10152 18552 10180
rect 20180 10152 20852 10180
rect 22683 10152 22770 10180
rect 5796 10016 23000 10112
rect 5736 9948 6040 9976
rect 6196 9948 6776 9976
rect 8864 9948 9076 9976
rect 17328 9948 17540 9976
rect 17991 9948 18078 9976
rect 18156 9948 18276 9976
rect 20640 9948 21496 9976
rect 22407 9948 22494 9976
rect 9048 9908 9076 9948
rect 6012 9880 6224 9908
rect 6012 9840 6040 9880
rect 5920 9812 6040 9840
rect 6196 9840 6224 9880
rect 6564 9880 6868 9908
rect 9048 9880 9352 9908
rect 14936 9880 15516 9908
rect 16209 9880 16436 9908
rect 6564 9840 6592 9880
rect 18156 9840 18184 9948
rect 22020 9880 22508 9908
rect 22480 9840 22508 9880
rect 23032 9880 23796 9908
rect 23032 9840 23060 9880
rect 6196 9812 6592 9840
rect 7024 9812 8064 9840
rect 9062 9812 10902 9840
rect 12563 9812 12664 9840
rect 15231 9812 15318 9840
rect 15507 9812 15594 9840
rect 7852 9744 7972 9772
rect 8036 9758 8064 9812
rect 15672 9772 15700 9840
rect 15948 9812 16068 9840
rect 16776 9812 18184 9840
rect 19352 9812 20116 9840
rect 20180 9812 20377 9840
rect 20824 9812 22324 9840
rect 22480 9812 23060 9840
rect 10060 9744 10180 9772
rect 12287 9744 12374 9772
rect 14292 9744 15792 9772
rect 7944 9636 7972 9744
rect 8147 9676 8248 9704
rect 9600 9676 9996 9704
rect 10704 9676 10916 9704
rect 11072 9676 11767 9704
rect 15856 9676 15976 9704
rect 17604 9676 18184 9704
rect 19095 9676 19182 9704
rect 21579 9676 21666 9704
rect 22112 9676 22232 9704
rect 9600 9670 9628 9676
rect 8404 9642 9628 9670
rect 8404 9636 8432 9642
rect 17604 9636 17632 9676
rect 18156 9670 18184 9676
rect 18156 9642 18920 9670
rect 5736 9608 6408 9636
rect 7944 9608 8432 9636
rect 10263 9608 10350 9636
rect 12061 9608 13032 9636
rect 13740 9608 14320 9636
rect 17052 9608 17632 9636
rect 18892 9636 18920 9642
rect 18892 9608 19472 9636
rect 5736 9296 5764 9608
rect 5796 9472 23000 9568
rect 8239 9404 8326 9432
rect 10631 9404 10718 9432
rect 11348 9404 11560 9432
rect 11624 9404 13124 9432
rect 14568 9404 15056 9432
rect 16132 9404 16252 9432
rect 20180 9404 20300 9432
rect 21560 9404 21680 9432
rect 22020 9404 22416 9432
rect 6288 9336 6500 9364
rect 6288 9296 6316 9336
rect 5736 9268 6316 9296
rect 6583 9268 6670 9296
rect 9140 9268 9352 9296
rect 10336 9228 10364 9364
rect 12931 9336 13018 9364
rect 13096 9296 13124 9404
rect 19996 9336 20668 9364
rect 13096 9268 13216 9296
rect 13464 9268 13676 9296
rect 6932 9200 7236 9228
rect 9585 9200 10364 9228
rect 12544 9200 12940 9228
rect 15856 9200 16436 9228
rect 16703 9200 16790 9228
rect 17696 9200 18015 9228
rect 18708 9200 18828 9228
rect 20364 9200 20484 9228
rect 20640 9200 20668 9336
rect 20824 9268 21312 9296
rect 22020 9268 22048 9404
rect 22388 9364 22416 9404
rect 23032 9404 23428 9432
rect 23032 9364 23060 9404
rect 22388 9336 23060 9364
rect 22112 9268 22232 9296
rect 12544 9160 12572 9200
rect 20824 9160 20852 9268
rect 21284 9228 21312 9268
rect 21284 9200 21864 9228
rect 6840 9132 7221 9160
rect 11716 9132 12296 9160
rect 12452 9132 12572 9160
rect 12651 9132 13400 9160
rect 13464 9132 13937 9160
rect 16427 9132 16514 9160
rect 16592 9132 16896 9160
rect 18524 9132 18644 9160
rect 19061 9132 20024 9160
rect 20180 9132 20852 9160
rect 21836 9160 21864 9200
rect 21836 9132 22048 9160
rect 11716 9092 11744 9132
rect 11532 9064 11744 9092
rect 12268 9092 12296 9132
rect 13464 9092 13492 9132
rect 12268 9064 13492 9092
rect 16868 9064 16896 9132
rect 18616 9092 18644 9132
rect 18340 9064 19380 9092
rect 20180 9064 20208 9132
rect 20916 9064 21220 9092
rect 21836 9064 22416 9092
rect 5796 8928 23000 9024
rect 8128 8860 8892 8888
rect 10796 8860 11100 8888
rect 12636 8860 13032 8888
rect 13188 8860 13308 8888
rect 14752 8860 15424 8888
rect 16500 8860 16896 8888
rect 17512 8860 19564 8888
rect 20180 8860 21588 8888
rect 10796 8820 10824 8860
rect 19536 8820 19564 8860
rect 6840 8792 7328 8820
rect 10520 8792 10824 8820
rect 11808 8792 12572 8820
rect 6840 8752 6868 8792
rect 6472 8724 6868 8752
rect 6932 8724 7880 8752
rect 9338 8724 10810 8752
rect 11808 8670 11836 8792
rect 12544 8786 12572 8792
rect 13004 8792 14320 8820
rect 16960 8792 17448 8820
rect 13004 8786 13032 8792
rect 12544 8758 13032 8786
rect 17420 8786 17448 8792
rect 18156 8792 19012 8820
rect 19536 8792 20116 8820
rect 18156 8786 18184 8792
rect 17420 8758 18184 8786
rect 18984 8752 19012 8792
rect 13207 8724 13294 8752
rect 13372 8724 13492 8752
rect 15415 8724 15502 8752
rect 15749 8724 16252 8752
rect 18340 8724 18722 8752
rect 18984 8724 19840 8752
rect 19996 8724 20378 8752
rect 7208 8588 8156 8616
rect 7208 8548 7236 8588
rect 5736 8520 6408 8548
rect 6748 8520 7236 8548
rect 8128 8548 8156 8588
rect 8312 8548 8340 8670
rect 12820 8656 13124 8684
rect 14476 8656 15240 8684
rect 8481 8588 10456 8616
rect 11647 8588 12756 8616
rect 12728 8582 12756 8588
rect 12728 8554 13400 8582
rect 13372 8548 13400 8554
rect 14476 8548 14504 8656
rect 8128 8520 8340 8548
rect 8680 8520 9536 8548
rect 13372 8520 14504 8548
rect 15212 8548 15240 8656
rect 16776 8656 18828 8684
rect 16776 8616 16804 8656
rect 18800 8616 18828 8656
rect 16684 8588 16804 8616
rect 18451 8588 18538 8616
rect 18800 8588 19656 8616
rect 19996 8548 20024 8724
rect 20272 8656 20470 8684
rect 20180 8588 20392 8616
rect 20364 8582 20392 8588
rect 21008 8588 21243 8616
rect 21008 8582 21036 8588
rect 20364 8554 21036 8582
rect 15212 8520 17540 8548
rect 17604 8520 20024 8548
rect 5736 8344 5764 8520
rect 5796 8384 23000 8480
rect 5736 8316 6316 8344
rect 8239 8316 8326 8344
rect 10631 8316 10718 8344
rect 13188 8316 13308 8344
rect 16316 8316 16896 8344
rect 17163 8316 17250 8344
rect 18248 8316 18644 8344
rect 18984 8316 20300 8344
rect 20916 8316 21220 8344
rect 22756 8316 23244 8344
rect 16316 8310 16344 8316
rect 13832 8282 16344 8310
rect 13832 8276 13860 8282
rect 12452 8248 13860 8276
rect 16500 8248 16804 8276
rect 16500 8208 16528 8248
rect 10704 8180 11100 8208
rect 13740 8180 16528 8208
rect 16868 8208 16896 8316
rect 17328 8248 17632 8276
rect 17328 8208 17356 8248
rect 16868 8180 17356 8208
rect 18616 8180 18644 8316
rect 6564 8112 6684 8140
rect 6932 8112 7236 8140
rect 9140 8112 9352 8140
rect 11808 8112 13124 8140
rect 14219 8112 14306 8140
rect 15028 8112 15148 8140
rect 15304 8112 15332 8180
rect 18064 8112 18383 8140
rect 18524 8112 18828 8140
rect 19003 8112 19104 8140
rect 20364 8112 20484 8140
rect 20562 8112 20649 8140
rect 21376 8112 21496 8140
rect 6748 8044 7216 8072
rect 9416 8044 9613 8072
rect 11333 8044 11437 8072
rect 14844 8044 14964 8072
rect 15212 8044 20024 8072
rect 20640 8004 20668 8072
rect 20732 8044 21680 8072
rect 11992 7976 12480 8004
rect 13391 7976 13478 8004
rect 14476 7976 15148 8004
rect 20180 7976 20668 8004
rect 5796 7840 23000 7936
rect 6932 7772 7497 7800
rect 9232 7772 9444 7800
rect 10060 7772 11008 7800
rect 11256 7772 11376 7800
rect 13740 7772 13952 7800
rect 7116 7704 7420 7732
rect 7469 7704 7497 7772
rect 10980 7732 11008 7772
rect 13924 7766 13952 7772
rect 14568 7772 15240 7800
rect 15967 7772 16054 7800
rect 18984 7772 19196 7800
rect 14568 7766 14596 7772
rect 13924 7738 14596 7766
rect 19168 7732 19196 7772
rect 19812 7772 21588 7800
rect 19812 7732 19840 7772
rect 7576 7704 10088 7732
rect 10980 7704 11468 7732
rect 11716 7704 12649 7732
rect 13280 7704 13400 7732
rect 19168 7704 19840 7732
rect 20088 7704 20208 7732
rect 22296 7704 22600 7732
rect 7116 7664 7144 7704
rect 7392 7664 7420 7704
rect 7576 7664 7604 7704
rect 10060 7698 10088 7704
rect 10060 7670 10732 7698
rect 6583 7636 7144 7664
rect 7208 7636 7328 7664
rect 7392 7636 7604 7664
rect 10704 7664 10732 7670
rect 11440 7664 11468 7704
rect 10704 7636 10931 7664
rect 11440 7636 12940 7664
rect 13372 7596 13400 7704
rect 22572 7664 22600 7704
rect 23032 7704 23520 7732
rect 23032 7664 23060 7704
rect 14016 7636 14136 7664
rect 14200 7636 14504 7664
rect 14752 7636 18368 7664
rect 18616 7636 18920 7664
rect 19996 7636 20378 7664
rect 22388 7596 22416 7664
rect 22572 7636 23060 7664
rect 8791 7568 8878 7596
rect 9048 7568 10088 7596
rect 11164 7568 12388 7596
rect 13372 7568 14412 7596
rect 17158 7568 17245 7596
rect 17328 7568 17448 7596
rect 18064 7568 20470 7596
rect 21560 7568 22416 7596
rect 5920 7460 5948 7528
rect 6380 7500 6500 7528
rect 9784 7500 9812 7568
rect 11551 7500 11638 7528
rect 14292 7500 16620 7528
rect 19812 7500 19932 7528
rect 21008 7500 21243 7528
rect 21928 7500 22048 7528
rect 21008 7494 21036 7500
rect 18340 7466 19656 7494
rect 18340 7460 18368 7466
rect 5736 7432 5948 7460
rect 6104 7432 9168 7460
rect 12176 7432 12572 7460
rect 13096 7432 13768 7460
rect 18156 7432 18368 7460
rect 19628 7460 19656 7466
rect 20364 7466 21036 7494
rect 20364 7460 20392 7466
rect 19628 7432 20392 7460
rect 5736 7120 5764 7432
rect 5796 7296 23000 7392
rect 6012 7228 6132 7256
rect 6307 7228 6394 7256
rect 13188 7228 14688 7256
rect 14752 7228 15056 7256
rect 16960 7228 17632 7256
rect 17807 7228 17894 7256
rect 18800 7228 19012 7256
rect 20272 7228 20668 7256
rect 21192 7228 21588 7256
rect 12123 7160 12227 7188
rect 5552 7092 5948 7120
rect 6859 7092 6946 7120
rect 10980 7092 11454 7120
rect 12471 7092 12558 7120
rect 5552 7024 5580 7092
rect 6196 6916 6224 7052
rect 9248 7024 9338 7052
rect 10980 6984 11008 7092
rect 14660 7052 14688 7228
rect 15212 7160 15700 7188
rect 18800 7160 18828 7228
rect 21192 7120 21220 7228
rect 16151 7092 16238 7120
rect 19187 7092 19274 7120
rect 20659 7092 20746 7120
rect 20916 7092 21220 7120
rect 21303 7092 21390 7120
rect 12282 7024 13124 7052
rect 13575 7024 13662 7052
rect 14660 7024 16712 7052
rect 16684 6984 16712 7024
rect 17236 7024 19012 7052
rect 21192 7024 23888 7052
rect 17236 6984 17264 7024
rect 7024 6956 7221 6984
rect 7668 6956 8156 6984
rect 7668 6916 7696 6956
rect 5644 6888 6500 6916
rect 6564 6888 6868 6916
rect 7484 6888 7696 6916
rect 8128 6916 8156 6956
rect 8496 6956 9076 6984
rect 10171 6956 10258 6984
rect 10428 6956 11008 6984
rect 11072 6956 11284 6984
rect 13280 6956 14044 6984
rect 15764 6956 16513 6984
rect 16684 6956 17264 6984
rect 19168 6956 19549 6984
rect 21579 6956 21680 6984
rect 8496 6916 8524 6956
rect 8128 6888 8524 6916
rect 9048 6916 9076 6956
rect 10428 6916 10456 6956
rect 9048 6888 10456 6916
rect 13280 6888 13308 6956
rect 18340 6888 19012 6916
rect 22480 6888 22784 6916
rect 5796 6752 23000 6848
rect 6196 6684 6776 6712
rect 6748 6644 6776 6684
rect 7668 6684 8156 6712
rect 11624 6684 12112 6712
rect 13280 6684 13768 6712
rect 20180 6684 20760 6712
rect 22296 6684 23704 6712
rect 7668 6644 7696 6684
rect 6031 6616 6118 6644
rect 6748 6616 7512 6644
rect 7595 6616 7696 6644
rect 7779 6616 7866 6644
rect 6748 6548 6776 6616
rect 6840 6548 7052 6576
rect 7576 6548 7972 6576
rect 8128 6556 8156 6684
rect 10428 6616 10640 6644
rect 13832 6616 14044 6644
rect 14016 6576 14044 6616
rect 14476 6616 15225 6644
rect 21744 6616 22232 6644
rect 14476 6576 14504 6616
rect 21744 6576 21772 6616
rect 22204 6576 22232 6616
rect 22756 6616 22968 6644
rect 22756 6576 22784 6616
rect 8423 6548 8524 6576
rect 11822 6548 12020 6576
rect 12287 6548 12374 6576
rect 12452 6548 12649 6576
rect 14016 6548 14504 6576
rect 14660 6548 14964 6576
rect 18267 6548 18354 6576
rect 20824 6548 21036 6576
rect 21652 6548 21772 6576
rect 21836 6548 21956 6576
rect 22204 6548 22784 6576
rect 12452 6508 12480 6548
rect 6380 6480 7512 6508
rect 7852 6480 8064 6508
rect 8234 6480 8321 6508
rect 9876 6480 10994 6508
rect 11992 6480 12480 6508
rect 18543 6480 18630 6508
rect 19812 6480 20576 6508
rect 9876 6440 9904 6480
rect 9600 6412 9904 6440
rect 11256 6412 11767 6440
rect 10152 6378 11100 6406
rect 10152 6372 10180 6378
rect 6491 6344 6578 6372
rect 7760 6344 7880 6372
rect 9968 6344 10180 6372
rect 11072 6372 11100 6378
rect 11992 6372 12020 6480
rect 21192 6446 21956 6474
rect 21192 6440 21220 6446
rect 21008 6412 21220 6440
rect 21928 6440 21956 6446
rect 21928 6412 24072 6440
rect 11072 6344 12020 6372
rect 16224 6344 16344 6372
rect 21468 6344 21864 6372
rect 5796 6208 23000 6304
rect 6932 6140 7052 6168
rect 7687 6140 7774 6168
rect 8220 6140 8432 6168
rect 9140 6100 9168 6168
rect 10336 6140 10456 6168
rect 12268 6140 12388 6168
rect 13188 6140 13860 6168
rect 18064 6140 18828 6168
rect 18911 6140 18998 6168
rect 19739 6140 19826 6168
rect 21100 6140 21956 6168
rect 22020 6140 22416 6168
rect 21928 6100 21956 6140
rect 9140 6072 10272 6100
rect 10244 6066 10272 6072
rect 12360 6072 13492 6100
rect 10244 6038 10824 6066
rect 10796 6032 10824 6038
rect 12360 6032 12388 6072
rect 6491 6004 6578 6032
rect 7668 6004 8156 6032
rect 10796 6004 12388 6032
rect 12544 6004 12572 6072
rect 8128 5964 8156 6004
rect 6748 5936 8064 5964
rect 8128 5936 10640 5964
rect 12728 5896 12756 6032
rect 12820 6004 13400 6032
rect 13464 5964 13492 6072
rect 13924 6072 14504 6100
rect 13924 5964 13952 6072
rect 14476 6032 14504 6072
rect 16040 6072 16344 6100
rect 16408 6072 16712 6100
rect 16040 6032 16068 6072
rect 14219 6004 14306 6032
rect 14476 6004 16068 6032
rect 16316 6032 16344 6072
rect 16684 6032 16712 6072
rect 19536 6072 20300 6100
rect 20732 6072 21588 6100
rect 21928 6072 22232 6100
rect 16316 6004 16620 6032
rect 16684 6004 18184 6032
rect 19536 6004 19564 6072
rect 20088 6004 20484 6032
rect 20732 6004 20760 6072
rect 21284 6004 21772 6032
rect 21850 6004 21937 6032
rect 12912 5936 13032 5964
rect 13207 5936 13294 5964
rect 13464 5936 13768 5964
rect 13832 5936 13952 5964
rect 13832 5896 13860 5936
rect 12728 5868 12940 5896
rect 12912 5862 12940 5868
rect 13648 5868 13860 5896
rect 13648 5862 13676 5868
rect 12912 5834 13676 5862
rect 14090 5856 14154 5973
rect 16795 5936 16882 5964
rect 17715 5936 17802 5964
rect 19628 5936 20392 5964
rect 5796 5664 23000 5760
rect 10888 4168 19196 4196
rect 19168 4100 19196 4168
rect 32 156 2636 184
rect 2608 116 2636 156
rect 13464 116 13492 184
rect 2608 88 13492 116
<< metal2 >>
rect 32 14760 60 27744
rect 18616 21808 18644 27720
rect 10152 21372 10180 21672
rect 7300 20176 7328 20652
rect 6840 20148 7328 20176
rect 6748 19768 6776 19972
rect 6656 19740 6776 19768
rect 6656 18748 6684 19740
rect 6932 19196 6960 20040
rect 6932 18816 6960 19020
rect 7024 18816 7052 19632
rect 6932 18788 7052 18816
rect 6656 18720 6776 18748
rect 6748 18516 6776 18720
rect 6564 17360 6592 18340
rect 6840 17048 6868 17252
rect 6656 17020 6868 17048
rect 6196 15388 6224 16368
rect 6656 15824 6684 17020
rect 6932 15932 6960 18788
rect 7116 15980 7144 17796
rect 6656 15796 6868 15824
rect 6840 15252 6868 15796
rect 7208 15552 7236 15756
rect 7300 15552 7328 20148
rect 7576 19740 7604 20720
rect 8772 19672 8800 19972
rect 7484 17428 7512 18068
rect 7944 16408 7972 19496
rect 8772 18652 8800 19428
rect 8956 19060 8984 19972
rect 9140 18516 9168 20516
rect 9968 19060 9996 21060
rect 10336 20176 10364 21740
rect 10520 20856 10548 21604
rect 10520 20828 10931 20856
rect 10704 20692 10916 20720
rect 10336 20148 10548 20176
rect 10244 19740 10272 20040
rect 10520 19604 10548 20148
rect 10336 19196 10364 19496
rect 8680 17524 8708 18476
rect 8864 18108 8892 18340
rect 9048 18108 9076 18476
rect 9968 17972 9996 18884
rect 9600 17564 9628 17932
rect 8588 17496 8708 17524
rect 9784 17496 9812 17932
rect 10244 17864 10272 19020
rect 9968 17836 10272 17864
rect 8588 16776 8616 17496
rect 8588 16748 8708 16776
rect 7484 15728 7512 16008
rect 8680 15960 8708 16748
rect 8864 16476 8892 17456
rect 9048 16340 9076 17252
rect 9968 16504 9996 17836
rect 10152 17020 10180 17456
rect 10336 17360 10364 17796
rect 10336 16816 10364 17252
rect 10704 16912 10732 20692
rect 10980 18992 11008 21196
rect 12636 20856 12664 21060
rect 12621 20828 12664 20856
rect 13096 20760 13124 21196
rect 11532 19060 11560 20584
rect 10980 18516 11008 18884
rect 10704 16884 10916 16912
rect 9876 16476 9996 16504
rect 8680 15932 8800 15960
rect 8864 15932 8892 16300
rect 9876 16272 9904 16476
rect 9140 16204 9260 16232
rect 7208 15524 7328 15552
rect 7300 14872 7328 15524
rect 7944 15252 7972 15756
rect 8680 15252 8708 15764
rect 8772 15592 8800 15932
rect 9048 15864 9076 16164
rect 9140 15960 9168 16204
rect 9140 15932 9260 15960
rect 8956 15252 8984 15756
rect 9232 15388 9260 15932
rect 9968 15892 9996 16476
rect 10704 16368 10732 16884
rect 10980 16408 11008 17796
rect 11348 17020 11376 18000
rect 11624 16476 11652 19020
rect 11808 18992 11836 19428
rect 11992 19060 12020 19496
rect 12176 19428 12204 19632
rect 12360 19604 12388 20040
rect 12636 19604 12664 20720
rect 13372 20108 13400 21196
rect 14292 20828 14320 21740
rect 13280 20080 13400 20108
rect 13280 19632 13308 20080
rect 13464 19768 13492 19972
rect 13464 19740 13584 19768
rect 13556 19632 13584 19740
rect 13280 19604 13400 19632
rect 13556 19604 13676 19632
rect 12176 19400 12296 19428
rect 12084 18884 12112 19156
rect 12268 18884 12296 19400
rect 12728 19360 12756 19564
rect 12728 19332 12848 19360
rect 12820 19224 12848 19332
rect 11992 18856 12112 18884
rect 12176 18856 12296 18884
rect 12636 19196 12848 19224
rect 11992 18272 12020 18856
rect 11992 18244 12112 18272
rect 11992 17020 12020 18068
rect 12084 17972 12112 18244
rect 12176 17904 12204 18856
rect 12636 18272 12664 19196
rect 13004 18380 13032 19156
rect 13188 18652 13216 19428
rect 13372 18992 13400 19604
rect 13648 19088 13676 19604
rect 13556 19060 13676 19088
rect 13556 18952 13584 19060
rect 13464 18924 13584 18952
rect 14200 18952 14228 19428
rect 14384 18952 14412 21060
rect 14476 20624 14504 21196
rect 14752 19944 14780 21060
rect 15120 20692 15148 21196
rect 15488 20828 15516 21604
rect 15948 21372 15976 21808
rect 16500 21236 16528 21740
rect 15488 20012 15516 20516
rect 15948 20080 15976 21196
rect 16040 19632 16068 19972
rect 16132 19740 16160 21128
rect 16224 20760 16252 21060
rect 16316 19740 16344 20040
rect 16040 19604 16160 19632
rect 14568 19060 14596 19428
rect 14200 18924 14320 18952
rect 14384 18924 14596 18952
rect 13464 18516 13492 18924
rect 12636 18244 12848 18272
rect 12268 17564 12296 18000
rect 12820 17456 12848 18244
rect 13188 18108 13308 18136
rect 12820 17428 13032 17456
rect 10612 16340 10732 16368
rect 9876 15864 9996 15892
rect 9508 15728 9536 15764
rect 9876 15144 9904 15864
rect 10060 15728 10088 16164
rect 10244 15824 10272 16232
rect 10152 15796 10272 15824
rect 9876 15116 9996 15144
rect 6932 14844 7328 14872
rect 6932 14708 6960 14844
rect 6564 14164 6592 14532
rect 5828 13648 5856 13812
rect 6748 13756 6776 14668
rect 5828 13620 5948 13648
rect 5920 7500 5948 13620
rect 6196 11376 6224 13444
rect 6380 12328 6408 13648
rect 6748 13076 6776 13512
rect 6932 13212 6960 14124
rect 6564 11880 6592 12492
rect 6748 12124 6776 12424
rect 6564 11852 6868 11880
rect 6380 11512 6408 11812
rect 6656 10724 6684 11404
rect 6840 11268 6868 11852
rect 7300 11404 7328 14844
rect 7944 13756 7972 14192
rect 9048 13756 9076 14804
rect 9140 13620 9168 13988
rect 9508 13212 9536 13580
rect 9968 13240 9996 15116
rect 10152 14844 10180 15796
rect 10704 15736 10732 16340
rect 10244 15252 10272 15620
rect 10428 14844 10456 15688
rect 10796 15252 10824 15756
rect 10704 14844 10732 15212
rect 10612 14300 10640 14788
rect 10888 13920 10916 14668
rect 10980 14640 11008 16164
rect 11164 15756 11192 15960
rect 11164 15728 11284 15756
rect 11624 15728 11652 16368
rect 11808 15932 11836 16844
rect 11900 16204 11928 16844
rect 12084 16776 12112 16980
rect 12084 16748 12296 16776
rect 11992 15824 12020 16368
rect 12268 15960 12296 16748
rect 12820 16408 12848 17428
rect 12912 16884 13032 16912
rect 11900 15796 12020 15824
rect 12084 15932 12296 15960
rect 11256 15280 11284 15728
rect 11164 15252 11284 15280
rect 11900 15252 11928 15796
rect 12084 15320 12112 15932
rect 11164 14164 11192 15252
rect 11348 14872 11376 15076
rect 11348 14844 11468 14872
rect 11440 14056 11468 14844
rect 11808 14300 11836 15212
rect 11348 14028 11468 14056
rect 10888 13892 11008 13920
rect 9968 13212 10088 13240
rect 10060 12628 10088 13212
rect 10244 12668 10272 13716
rect 10704 13008 10732 13444
rect 10796 13144 10824 13716
rect 10980 13552 11008 13892
rect 11348 13756 11376 14028
rect 11624 13240 11652 13444
rect 11532 13212 11652 13240
rect 9968 12600 10088 12628
rect 7944 11580 7972 12560
rect 8864 12124 8892 12492
rect 9968 12152 9996 12600
rect 9968 12124 10088 12152
rect 7208 11376 7328 11404
rect 6840 11240 6960 11268
rect 6564 10696 6684 10724
rect 6564 10248 6592 10696
rect 6932 10520 6960 11240
rect 6840 10492 6960 10520
rect 6840 10288 6868 10492
rect 6564 10220 6684 10248
rect 6472 9772 6500 9976
rect 6380 9744 6500 9772
rect 6380 8956 6408 9744
rect 6380 8928 6500 8956
rect 6472 8724 6500 8928
rect 6104 6616 6132 7460
rect 6380 7228 6408 7528
rect 6656 6440 6684 10220
rect 7300 9228 7328 11376
rect 8680 10424 8708 11404
rect 8864 9948 8892 11540
rect 9048 10832 9076 11268
rect 9048 10220 9076 10724
rect 7208 9200 7328 9228
rect 7300 8140 7328 9200
rect 8220 9160 8248 9704
rect 8312 9404 8340 9772
rect 8220 9132 8708 9160
rect 7208 8112 7328 8140
rect 7300 7120 7328 8112
rect 6932 7092 7328 7120
rect 6840 6548 6868 6916
rect 6656 6412 6776 6440
rect 6564 6004 6592 6372
rect 6748 5936 6776 6412
rect 7024 6140 7052 6984
rect 7300 6586 7328 7092
rect 7484 6480 7512 6916
rect 7668 6004 7696 6644
rect 7852 6480 7880 8752
rect 8312 8316 8340 8548
rect 8680 8520 8708 9132
rect 8864 7568 8892 8888
rect 9140 7684 9168 10316
rect 9416 7772 9444 8072
rect 10060 7568 10088 12124
rect 10244 11920 10272 12356
rect 10428 11580 10456 12628
rect 10796 12056 10824 12968
rect 10612 11676 10640 11880
rect 10612 11648 10732 11676
rect 10520 10492 10548 11404
rect 10704 11200 10732 11648
rect 11532 11608 11560 13212
rect 11532 11580 11652 11608
rect 10612 11172 10732 11200
rect 10612 10968 10640 11172
rect 10336 9336 10364 9636
rect 10704 9404 10732 9840
rect 10888 9676 10916 10792
rect 11348 10424 11376 11064
rect 11072 8860 11100 9704
rect 11348 9404 11376 9772
rect 11624 9404 11652 11580
rect 11808 11336 11836 13988
rect 11992 12668 12020 13036
rect 11992 11512 12020 11948
rect 11808 11308 11928 11336
rect 11900 9296 11928 11308
rect 11808 9268 11928 9296
rect 7760 6140 7788 6372
rect 8220 6342 8248 6508
rect 8496 6440 8524 6576
rect 8404 6412 8524 6440
rect 8404 6140 8432 6412
rect 9140 6140 9168 7460
rect 9306 6929 9370 7064
rect 10244 6586 10272 6984
rect 10428 6616 10456 8616
rect 10704 8316 10732 8752
rect 10704 7684 10732 8208
rect 11808 8112 11836 9268
rect 12360 9160 12388 15756
rect 12728 15688 12756 16164
rect 13004 15932 13032 16884
rect 13096 16476 13124 16708
rect 12452 15660 12756 15688
rect 12544 15252 12664 15280
rect 12544 13212 12572 15252
rect 12820 14164 12848 15076
rect 13188 15008 13216 18108
rect 14292 17836 14320 18924
rect 14568 18272 14596 18924
rect 14844 18584 14872 19156
rect 16132 18584 16160 19604
rect 16868 19152 16896 19632
rect 17144 18992 17172 21332
rect 17420 21236 17448 21604
rect 18248 21372 18276 21808
rect 18616 21780 18736 21808
rect 18432 21100 18460 21672
rect 18708 21264 18736 21780
rect 19168 21304 19196 21604
rect 18616 21236 18736 21264
rect 19628 21236 19656 21740
rect 17696 19604 17724 21060
rect 17604 19196 17632 19428
rect 14568 18244 14688 18272
rect 13372 17292 13400 17796
rect 13280 16476 13308 16844
rect 14108 16816 14136 17524
rect 14292 16884 14320 17472
rect 13372 16164 13400 16368
rect 13372 16136 13492 16164
rect 13464 15688 13492 16136
rect 13096 14980 13216 15008
rect 13372 15660 13492 15688
rect 13096 13648 13124 14980
rect 12728 13144 12756 13648
rect 13096 13620 13216 13648
rect 13004 12464 13032 13444
rect 13188 13104 13216 13620
rect 13372 13552 13400 15660
rect 14292 15348 14320 15620
rect 14200 15320 14320 15348
rect 14200 14600 14228 15320
rect 14476 14640 14504 17864
rect 14660 16816 14688 18244
rect 14844 17444 14872 17796
rect 15580 17456 15608 18544
rect 17328 18448 17356 19020
rect 17880 18992 17908 19972
rect 17604 18408 17632 18612
rect 17788 18584 17816 18884
rect 18616 18856 18644 21236
rect 18892 20760 18920 21060
rect 19904 20760 19932 21604
rect 19996 21372 20024 21604
rect 20364 21400 20392 21864
rect 20364 21372 20484 21400
rect 19168 20128 19196 20652
rect 20088 20080 20116 21196
rect 20456 20584 20484 21372
rect 20364 20556 20484 20584
rect 20364 20108 20392 20556
rect 20364 20080 20484 20108
rect 18892 19740 18920 20040
rect 20180 19768 20208 19972
rect 20088 19740 20208 19768
rect 19076 19496 19104 19668
rect 18984 19468 19104 19496
rect 18984 19020 19012 19468
rect 19260 19128 19288 19428
rect 20088 19292 20116 19740
rect 20456 19496 20484 20080
rect 20364 19468 20484 19496
rect 20088 19264 20208 19292
rect 18984 18992 19104 19020
rect 17512 18380 17632 18408
rect 15764 17904 15792 18340
rect 15580 17428 15700 17456
rect 14752 17048 14780 17252
rect 14752 17020 14872 17048
rect 14844 16408 14872 17020
rect 15304 16776 15332 17048
rect 15304 16748 15424 16776
rect 15396 16408 15424 16748
rect 15580 16504 15608 17428
rect 15856 17224 15884 17932
rect 16040 16504 16068 17932
rect 16500 17864 16528 18068
rect 16316 17020 16344 17864
rect 16500 17836 16620 17864
rect 16592 16980 16620 17836
rect 15580 16476 15792 16504
rect 15856 16476 16068 16504
rect 16500 16952 16620 16980
rect 15580 15892 15608 16476
rect 15856 15960 15884 16476
rect 15948 16340 16252 16368
rect 15856 15932 15976 15960
rect 15488 15864 15608 15892
rect 15488 15416 15516 15864
rect 15488 15388 15608 15416
rect 15580 15280 15608 15388
rect 14200 14572 14320 14600
rect 13464 14232 13492 14532
rect 14292 14232 14320 14572
rect 14568 14300 14596 14532
rect 14384 13756 14412 14192
rect 14568 13662 14596 14192
rect 13464 13144 13492 13444
rect 13188 13076 13400 13104
rect 14568 12968 14596 13172
rect 14476 12940 14596 12968
rect 13280 12532 13308 12592
rect 13280 11580 13308 12084
rect 13280 10492 13308 10860
rect 12360 9132 12480 9160
rect 11348 7772 11376 8072
rect 9968 6168 9996 6372
rect 9600 6140 9996 6168
rect 10336 6140 10364 6508
rect 32 0 60 184
rect 9600 0 9628 6140
rect 10888 4168 10916 7664
rect 11256 6412 11284 6984
rect 11624 6684 11652 7528
rect 11992 7324 12020 8004
rect 11900 7296 12020 7324
rect 11900 6780 11928 7296
rect 11900 6752 12020 6780
rect 11992 6548 12020 6752
rect 12176 6576 12204 7188
rect 12176 6548 12296 6576
rect 12360 6548 12388 9132
rect 12636 8860 12664 9840
rect 13004 9336 13032 9636
rect 13096 8480 13124 9296
rect 13280 8860 13308 10316
rect 13004 8452 13124 8480
rect 13004 7868 13032 8452
rect 13004 7840 13124 7868
rect 13096 7664 13124 7840
rect 13280 7704 13308 8752
rect 13464 8724 13492 12492
rect 14476 12356 14504 12940
rect 14476 12328 14596 12356
rect 14568 12124 14596 12328
rect 14016 11444 14044 11982
rect 14200 10288 14320 10316
rect 14476 10288 14504 10724
rect 14568 10492 14596 11404
rect 14292 9744 14320 10288
rect 14292 8792 14320 9636
rect 14568 9404 14596 10180
rect 12912 7460 12940 7664
rect 13096 7636 13216 7664
rect 12544 7092 12572 7460
rect 12820 7432 12940 7460
rect 12820 6916 12848 7432
rect 13096 7024 13124 7460
rect 13188 7228 13216 7636
rect 12820 6888 12940 6916
rect 12268 5976 12296 6548
rect 12912 5936 12940 6888
rect 13280 6684 13308 6916
rect 13280 5936 13308 6004
rect 13464 156 13492 8004
rect 13648 7024 13676 7712
rect 14016 6956 14044 7664
rect 13832 6140 13860 6644
rect 14292 6004 14320 8140
rect 14752 8072 14780 15280
rect 15580 15252 15700 15280
rect 15212 14164 15240 14600
rect 15580 14096 15608 15252
rect 15764 14150 15792 15886
rect 15948 15048 15976 15932
rect 15304 12930 15332 13690
rect 15488 11954 15516 14056
rect 15580 11880 15608 13104
rect 15672 12056 15700 12900
rect 15856 12532 15884 14532
rect 16040 13212 16068 15212
rect 16224 14638 16252 16340
rect 15488 11852 15608 11880
rect 15488 10520 15516 11852
rect 15764 11036 15792 11336
rect 15856 10928 15884 12348
rect 15304 10492 15516 10520
rect 15764 10900 15884 10928
rect 14936 9880 14964 10180
rect 15304 9812 15332 10492
rect 15580 9432 15608 9840
rect 15764 9568 15792 10900
rect 15948 9676 15976 10928
rect 16132 10492 16160 13172
rect 15764 9540 15884 9568
rect 15396 9404 15608 9432
rect 15396 8860 15424 9404
rect 15488 8724 15516 8810
rect 14752 8044 14872 8072
rect 14476 7636 14504 8004
rect 14660 6548 14688 7712
rect 14752 7636 14780 8044
rect 15028 7528 15056 8140
rect 15212 7772 15240 8072
rect 14752 7500 15056 7528
rect 14752 7228 14780 7500
rect 15672 7160 15700 9420
rect 15856 9200 15884 9540
rect 16040 7772 16068 9840
rect 16132 9404 16160 10248
rect 16316 9636 16344 15076
rect 16500 14640 16528 16952
rect 16684 16476 16712 16776
rect 16684 16300 16712 16374
rect 16684 14464 16712 15824
rect 16868 15252 16896 17252
rect 16592 14436 16712 14464
rect 16408 9296 16436 9908
rect 16362 9268 16436 9296
rect 16592 9296 16620 14436
rect 16960 13648 16988 15756
rect 17144 14300 17172 17388
rect 17328 15660 17356 17932
rect 17512 15824 17540 18380
rect 17696 17428 17724 18476
rect 17880 18340 17908 18544
rect 17880 18312 18000 18340
rect 17972 17660 18000 18312
rect 17880 17632 18000 17660
rect 17880 17224 17908 17632
rect 17972 16884 18184 16912
rect 17788 16476 17816 16776
rect 17420 15796 17540 15824
rect 17328 14668 17356 15076
rect 17420 14844 17448 15796
rect 17328 14640 17448 14668
rect 17420 14192 17448 14640
rect 16868 13620 16988 13648
rect 17328 14164 17448 14192
rect 16868 13172 16896 13620
rect 16868 13144 16942 13172
rect 16776 12668 16804 12958
rect 16776 12464 16804 12592
rect 16776 12124 16804 12356
rect 16914 11608 16942 13144
rect 17052 11812 17080 12900
rect 17144 12668 17172 13512
rect 17328 13212 17356 14164
rect 17788 13552 17816 15620
rect 17972 14872 18000 16884
rect 18432 16816 18460 18340
rect 18892 18136 18920 18340
rect 18800 18108 18920 18136
rect 18800 17456 18828 18108
rect 18800 17428 18920 17456
rect 18616 16408 18644 17252
rect 18616 15252 18644 15756
rect 18892 15416 18920 17428
rect 19076 16436 19104 18992
rect 19812 17838 19840 17932
rect 19904 17838 19932 18476
rect 19812 17810 19932 17838
rect 19536 16834 19564 17472
rect 19720 17020 19748 17524
rect 19076 16408 19196 16436
rect 19168 15960 19196 16408
rect 19904 16340 19932 17810
rect 20088 16884 20116 18680
rect 20180 18584 20208 19264
rect 20364 18992 20392 19468
rect 20916 18652 20944 18884
rect 19076 15932 19196 15960
rect 19076 15728 19104 15932
rect 18892 15388 19012 15416
rect 18524 14872 18552 15154
rect 17972 14844 18552 14872
rect 17972 13620 18000 14844
rect 18248 13920 18276 14736
rect 18524 14640 18552 14844
rect 18616 14164 18644 14600
rect 18248 13892 18368 13920
rect 18340 13756 18368 13892
rect 17236 13076 17356 13104
rect 17512 13076 17540 13202
rect 17144 11988 17172 12492
rect 17328 11852 17356 13076
rect 17512 12564 17540 12900
rect 17512 11880 17540 12084
rect 17972 12056 18000 12356
rect 17466 11852 17540 11880
rect 17052 11784 17172 11812
rect 16914 11580 16988 11608
rect 16868 10288 16896 11404
rect 16960 10112 16988 11580
rect 17144 10384 17172 11784
rect 17466 11268 17494 11852
rect 17604 11376 17632 11812
rect 16914 10084 16988 10112
rect 17098 10356 17172 10384
rect 16592 9268 16666 9296
rect 16362 8752 16390 9268
rect 16500 8860 16528 9160
rect 16638 8820 16666 9268
rect 16592 8792 16666 8820
rect 16224 8538 16252 8752
rect 16362 8724 16436 8752
rect 16224 7092 16252 7712
rect 16224 6072 16252 6372
rect 16408 6168 16436 8724
rect 16592 8616 16620 8792
rect 16592 8588 16712 8616
rect 16592 7500 16620 8588
rect 16776 8248 16804 9840
rect 16914 9500 16942 10084
rect 17098 9840 17126 10356
rect 17328 10220 17356 11268
rect 17466 11240 17540 11268
rect 17052 9812 17126 9840
rect 17052 9608 17080 9812
rect 16914 9472 16988 9500
rect 16960 8792 16988 9472
rect 17052 8072 17080 8566
rect 17236 8316 17264 10180
rect 17512 9948 17540 11240
rect 16868 8044 17080 8072
rect 16868 7460 16896 8044
rect 17144 7568 17172 7956
rect 17420 7568 17448 9636
rect 17696 9200 17724 10452
rect 17604 8248 17632 8548
rect 17880 8072 17908 11268
rect 17972 10322 18000 10396
rect 18064 10288 18092 11268
rect 18156 10124 18184 10180
rect 18064 8344 18092 9976
rect 18248 9948 18276 11880
rect 18524 10928 18552 11948
rect 18432 10900 18552 10928
rect 18064 8316 18276 8344
rect 17788 8044 17908 8072
rect 17788 7460 17816 8044
rect 18064 7568 18092 8140
rect 16868 7432 16988 7460
rect 17788 7432 17908 7460
rect 16960 7228 16988 7432
rect 17880 7228 17908 7432
rect 18156 7052 18184 7460
rect 16408 6140 16896 6168
rect 16868 5936 16896 6140
rect 17788 5936 17816 7052
rect 18064 7024 18184 7052
rect 18064 6440 18092 7024
rect 18340 6548 18368 9840
rect 18524 8112 18552 10900
rect 18616 6480 18644 12592
rect 18800 12532 18828 14736
rect 18984 14300 19012 14600
rect 19076 13662 19104 15620
rect 19812 14600 19840 15144
rect 19812 14572 19932 14600
rect 19996 14572 20024 15076
rect 20088 14640 20116 16708
rect 20180 16680 20208 17252
rect 20364 14776 20392 18340
rect 21100 18068 21128 21740
rect 21284 21168 21312 21808
rect 21468 20992 21496 21264
rect 21376 20964 21496 20992
rect 21376 19088 21404 20964
rect 21376 19060 21496 19088
rect 21008 18040 21128 18068
rect 21008 17524 21036 18040
rect 21008 17496 21128 17524
rect 21100 17292 21128 17496
rect 20916 16788 20944 16862
rect 20732 16476 20760 16776
rect 21008 16232 21036 16708
rect 21284 16346 21312 18884
rect 21468 17904 21496 19060
rect 21652 18584 21680 21604
rect 21468 16748 21496 17796
rect 21652 17388 21680 17716
rect 21836 17564 21864 25280
rect 22756 21780 22784 21864
rect 22020 21372 22048 21740
rect 22388 21400 22416 21604
rect 22388 21372 22508 21400
rect 22020 19904 22048 20652
rect 22204 19972 22232 21332
rect 22480 20924 22508 21372
rect 22388 20896 22508 20924
rect 22204 19944 22278 19972
rect 22020 19876 22140 19904
rect 22020 19564 22048 19768
rect 21974 19536 22048 19564
rect 21974 19020 22002 19536
rect 22112 19088 22140 19876
rect 22250 19428 22278 19944
rect 22204 19400 22278 19428
rect 22204 19196 22232 19400
rect 22112 19060 22232 19088
rect 21974 18992 22048 19020
rect 22020 18340 22048 18992
rect 22204 18516 22232 19060
rect 22020 18312 22140 18340
rect 22112 17660 22140 18312
rect 22020 17632 22140 17660
rect 21652 17360 21772 17388
rect 21744 16708 21772 17360
rect 21652 16680 21772 16708
rect 21652 16476 21680 16680
rect 21008 16204 21128 16232
rect 21100 15960 21128 16204
rect 21008 15932 21128 15960
rect 21008 15728 21036 15932
rect 21100 14872 21128 15348
rect 21008 14844 21128 14872
rect 19904 14096 19932 14572
rect 18708 8782 18736 9228
rect 18800 7684 18828 11404
rect 18984 8316 19012 12424
rect 19904 12084 19932 13648
rect 20180 13416 20208 14532
rect 20364 13784 20392 14668
rect 20456 14516 20484 14736
rect 20640 14504 20668 14788
rect 21284 14516 21312 16164
rect 21468 15126 21496 15756
rect 22020 15688 22048 17632
rect 22204 16476 22232 17456
rect 22388 16476 22416 20896
rect 22572 18136 22600 20720
rect 22480 18108 22600 18136
rect 22756 20040 22784 20156
rect 22848 20148 22968 20176
rect 22848 20040 22876 20148
rect 22756 20012 22876 20040
rect 22480 17904 22508 18108
rect 21284 14164 21312 14300
rect 20364 13756 20760 13784
rect 20456 13104 20484 13690
rect 20364 13076 20484 13104
rect 20180 12696 20208 12900
rect 19812 12056 19932 12084
rect 20088 12668 20208 12696
rect 20088 12056 20116 12668
rect 20180 12464 20208 12592
rect 19812 11948 19840 12056
rect 19720 11920 19840 11948
rect 19720 11472 19748 11920
rect 19996 11608 20024 11812
rect 19996 11580 20116 11608
rect 19720 11444 19840 11472
rect 19812 11336 19840 11444
rect 19076 11308 19196 11336
rect 19812 11308 19932 11336
rect 19076 11064 19104 11308
rect 19904 11064 19932 11308
rect 20088 11132 20116 11580
rect 19076 11036 19196 11064
rect 19168 10928 19196 11036
rect 19812 11036 19932 11064
rect 19996 11104 20116 11132
rect 20364 11336 20392 13076
rect 20548 12930 20576 13512
rect 20732 13376 20760 13756
rect 20732 13348 20852 13376
rect 20824 13174 20852 13348
rect 21100 12442 21128 12492
rect 21192 11954 21220 12016
rect 21284 11880 21312 13202
rect 21192 11852 21312 11880
rect 20364 11308 20484 11336
rect 19812 10928 19840 11036
rect 19168 10900 19288 10928
rect 19260 10384 19288 10900
rect 19168 10356 19288 10384
rect 19720 10900 19840 10928
rect 19720 10384 19748 10900
rect 19720 10356 19840 10384
rect 19168 10248 19196 10356
rect 19076 10220 19196 10248
rect 19812 10248 19840 10356
rect 19812 10220 19932 10248
rect 19076 8820 19104 10220
rect 19904 9976 19932 10220
rect 19812 9948 19932 9976
rect 19812 9840 19840 9948
rect 19168 9636 19196 9704
rect 19352 9064 19380 9840
rect 19720 9812 19840 9840
rect 19720 9364 19748 9812
rect 19720 9336 19840 9364
rect 19996 9336 20024 11104
rect 20180 10520 20208 10928
rect 20180 10492 20300 10520
rect 20180 9404 20208 9840
rect 19812 9132 19840 9336
rect 19996 8820 20024 9160
rect 20180 8860 20208 9298
rect 19076 8792 19196 8820
rect 19168 8344 19196 8792
rect 19076 8316 19196 8344
rect 19904 8792 20024 8820
rect 19076 8112 19104 8316
rect 19904 8208 19932 8792
rect 19904 8180 20116 8208
rect 18984 7228 19012 7800
rect 19260 7092 19288 7712
rect 19812 7500 19840 7712
rect 19996 7636 20024 8072
rect 18064 6412 18184 6440
rect 18156 6004 18184 6412
rect 18800 6140 18828 6492
rect 18984 6140 19012 6916
rect 19812 6140 19840 6508
rect 20088 6004 20116 8180
rect 20180 7704 20208 8616
rect 20272 8538 20300 8684
rect 20364 8112 20392 11308
rect 20548 10696 20576 11336
rect 20824 11036 20852 11336
rect 21192 11064 21220 11852
rect 21192 11036 21312 11064
rect 20640 9948 20668 10316
rect 20824 9812 20852 10180
rect 21100 9364 21128 10996
rect 21008 9336 21128 9364
rect 21008 9228 21036 9336
rect 21284 9296 21312 11036
rect 21376 10968 21404 11268
rect 20916 9200 21036 9228
rect 21192 9268 21312 9296
rect 20916 8752 20944 9200
rect 20916 8724 21036 8752
rect 21008 8616 21036 8724
rect 21008 8588 21128 8616
rect 21100 8276 21128 8588
rect 21192 8316 21220 9268
rect 21008 8248 21128 8276
rect 20548 8050 20576 8140
rect 20272 7228 20300 7596
rect 20732 7528 20760 8072
rect 20364 7500 20760 7528
rect 21008 7528 21036 8248
rect 21008 7500 21128 7528
rect 20364 5936 20392 7500
rect 21100 7256 21128 7500
rect 21008 7228 21128 7256
rect 20732 6684 20760 7120
rect 21008 6548 21036 7228
rect 21284 6004 21312 8322
rect 21468 8112 21496 14192
rect 21744 13920 21772 15620
rect 21928 14300 21956 15688
rect 22020 15660 22140 15688
rect 21744 13892 21956 13920
rect 21744 13212 21772 13784
rect 21652 12668 21680 13172
rect 21836 12696 21864 13104
rect 21790 12668 21864 12696
rect 21652 12124 21680 12424
rect 21790 12016 21818 12668
rect 21744 11988 21818 12016
rect 21744 11608 21772 11988
rect 21744 11580 21818 11608
rect 21652 10248 21680 11540
rect 21790 10384 21818 11580
rect 21790 10356 21864 10384
rect 21652 10220 21772 10248
rect 21836 10246 21864 10356
rect 21928 10220 21956 13892
rect 22020 13076 22048 13202
rect 22112 12220 22140 15660
rect 22066 12192 22140 12220
rect 22066 11676 22094 12192
rect 22296 12152 22324 16300
rect 22480 14640 22508 15076
rect 22204 12124 22324 12152
rect 22204 11744 22232 12124
rect 22204 11716 22324 11744
rect 22066 11648 22140 11676
rect 21744 9840 21772 10220
rect 22112 10044 22140 11648
rect 22296 10044 22324 11716
rect 22480 11268 22508 13580
rect 22756 11444 22784 20012
rect 22940 19836 22968 20040
rect 22940 19808 23060 19836
rect 23032 18884 23060 19808
rect 22940 18856 23060 18884
rect 22940 18652 22968 18856
rect 22940 18340 22968 18544
rect 22940 18312 23060 18340
rect 23032 16504 23060 18312
rect 26436 18108 26464 22718
rect 22940 16476 23060 16504
rect 22940 16272 22968 16476
rect 22940 15076 22968 15276
rect 22940 15048 23060 15076
rect 23032 14192 23060 15048
rect 22940 14164 23060 14192
rect 22940 13960 22968 14164
rect 22940 12492 22968 12696
rect 22940 12464 23060 12492
rect 23032 11336 23060 12464
rect 22940 11308 23060 11336
rect 22480 11240 22600 11268
rect 22572 10384 22600 11240
rect 22020 10016 22140 10044
rect 22204 10016 22324 10044
rect 22480 10356 22600 10384
rect 21744 9812 21864 9840
rect 21652 9404 21680 9704
rect 21836 9296 21864 9812
rect 22020 9500 22048 10016
rect 22204 9840 22232 10016
rect 22480 9948 22508 10356
rect 22204 9812 22324 9840
rect 22020 9472 22140 9500
rect 21652 9268 21864 9296
rect 22112 9268 22140 9472
rect 21652 8044 21680 9268
rect 21376 7092 21404 7712
rect 21560 7228 21588 7596
rect 21652 6464 21680 6984
rect 21836 6548 21864 9092
rect 22020 7684 22048 9160
rect 21836 6004 21864 6372
rect 22020 6140 22048 7528
rect 22204 6072 22232 9704
rect 22296 9432 22324 9812
rect 22296 9404 22508 9432
rect 22480 7868 22508 9404
rect 22756 8050 22784 10180
rect 22388 7840 22508 7868
rect 22388 7636 22416 7840
rect 22480 6220 22508 6916
rect 22940 6616 22968 11308
rect 14108 5868 14320 5896
rect 14292 120 14320 5868
rect 23216 5244 23244 10316
rect 23492 9432 23520 16912
rect 28736 12328 28764 27744
rect 23400 9404 23520 9432
rect 19168 0 19196 4128
rect 26252 2682 26280 10724
rect 28552 120 28580 8078
rect 28736 0 28764 392
<< metal3 >>
rect 18600 27676 28796 27736
rect 21820 25236 28796 25296
rect 26420 22674 28796 22734
rect 20348 21820 22800 21880
rect 23016 20234 28796 20294
rect 15932 20112 22800 20172
rect 23016 19684 23076 20234
rect 19060 19624 23076 19684
rect 16852 19136 22156 19196
rect 17680 17794 19856 17854
rect 21636 17672 28796 17732
rect 14276 17428 14888 17488
rect 17864 17428 19580 17488
rect 19520 16818 20960 16878
rect 16668 16330 20132 16390
rect 21176 16330 21298 16390
rect 7100 15964 7528 16024
rect 15748 15842 17372 15902
rect 7284 15720 10748 15780
rect 22924 15232 28796 15292
rect 18508 15110 21512 15170
rect 16 14744 10656 14804
rect 19060 14744 20684 14804
rect 16208 14622 18016 14682
rect 20440 14500 21328 14560
rect 21268 14256 22156 14316
rect 14736 14134 15808 14194
rect 0 13768 5872 13828
rect 14552 13646 15348 13706
rect 19060 13646 20500 13706
rect 15472 13158 18844 13218
rect 20808 13158 22064 13218
rect 15288 12914 16820 12974
rect 20532 12914 22524 12974
rect 12344 12548 13324 12608
rect 15840 12304 15900 12914
rect 22464 12730 22524 12914
rect 22464 12670 28796 12730
rect 16760 12548 17556 12608
rect 18600 12548 20224 12608
rect 21084 12426 22800 12486
rect 14000 11938 15532 11998
rect 21173 11935 21336 12001
rect 16852 10596 18568 10656
rect 15748 10352 18292 10412
rect 18232 10290 18292 10352
rect 10044 10230 14428 10290
rect 18232 10230 20408 10290
rect 21820 10230 28796 10290
rect 14368 10168 14428 10230
rect 14368 10108 18200 10168
rect 18048 9864 21512 9924
rect 16300 9620 19212 9680
rect 17128 9498 17188 9620
rect 15656 9376 16636 9436
rect 16576 9314 16636 9376
rect 16576 9254 20224 9314
rect 13448 8766 18752 8826
rect 16208 8522 17464 8582
rect 17404 8338 17464 8522
rect 19980 8522 20316 8582
rect 19980 8338 20040 8522
rect 17404 8278 20040 8338
rect 21176 8278 21298 8338
rect 20532 8034 28596 8094
rect 17036 7912 17158 7972
rect 9124 7668 21420 7728
rect 22004 7668 28796 7728
rect 9308 6936 18660 6996
rect 7284 6570 10288 6630
rect 8480 6386 8540 6570
rect 18784 6448 21696 6508
rect 8204 6326 8540 6386
rect 22464 6020 22524 6264
rect 12252 5960 13324 6020
rect 16852 5960 22524 6020
rect 23200 5228 28796 5288
rect 26236 2666 28796 2726
rect 28352 348 28780 408
rect 28352 164 28412 348
rect 14276 104 28412 164
rect 28536 104 28796 164
<< metal4 >>
rect 3936 0 4556 27744
rect 5176 0 5796 27744
rect 8000 3852 8620 23892
rect 9240 5092 9860 22652
rect 13600 3852 14220 23892
rect 14840 5092 15460 22652
rect 17128 7912 17188 9558
rect 19200 3852 19820 23892
rect 20440 5092 21060 22652
rect 21268 16024 21328 16390
rect 21268 15964 21604 16024
rect 21544 12364 21604 15964
rect 21268 12304 21604 12364
rect 21268 11632 21328 12304
rect 21268 11572 21466 11632
rect 21406 8704 21466 11572
rect 21268 8644 21466 8704
rect 21268 8278 21328 8644
rect 23000 0 23620 27744
rect 24240 0 24860 27744
<< metal5 >>
rect 0 23272 28796 23892
rect 0 22032 28796 22652
rect 0 5092 28796 5712
rect 0 3852 28796 4472
use L1M1_PR  L1M1_PR_0
timestamp 1655484843
transform 1 0 18262 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1
timestamp 1655484843
transform 1 0 18078 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_2
timestamp 1655484843
transform 1 0 16882 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_3
timestamp 1655484843
transform 1 0 16606 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_4
timestamp 1655484843
transform 1 0 15502 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_5
timestamp 1655484843
transform 1 0 14674 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_6
timestamp 1655484843
transform 1 0 15226 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_7
timestamp 1655484843
transform 1 0 14398 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_8
timestamp 1655484843
transform 1 0 15686 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_9
timestamp 1655484843
transform 1 0 15410 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_10
timestamp 1655484843
transform 1 0 16238 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_11
timestamp 1655484843
transform 1 0 15502 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_12
timestamp 1655484843
transform 1 0 16974 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_13
timestamp 1655484843
transform 1 0 16422 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_14
timestamp 1655484843
transform 1 0 16606 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_15
timestamp 1655484843
transform 1 0 15962 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_16
timestamp 1655484843
transform 1 0 17526 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_17
timestamp 1655484843
transform 1 0 16790 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_18
timestamp 1655484843
transform 1 0 16238 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_19
timestamp 1655484843
transform 1 0 14398 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_20
timestamp 1655484843
transform 1 0 17526 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_21
timestamp 1655484843
transform 1 0 15502 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_22
timestamp 1655484843
transform 1 0 13938 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_23
timestamp 1655484843
transform 1 0 13386 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_24
timestamp 1655484843
transform 1 0 16882 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_25
timestamp 1655484843
transform 1 0 16606 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_26
timestamp 1655484843
transform 1 0 16790 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_27
timestamp 1655484843
transform 1 0 15686 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_28
timestamp 1655484843
transform 1 0 17710 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_29
timestamp 1655484843
transform 1 0 17618 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_30
timestamp 1655484843
transform 1 0 20194 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_31
timestamp 1655484843
transform 1 0 19734 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_32
timestamp 1655484843
transform 1 0 20746 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_33
timestamp 1655484843
transform 1 0 19918 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_34
timestamp 1655484843
transform 1 0 19642 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_35
timestamp 1655484843
transform 1 0 19182 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_36
timestamp 1655484843
transform 1 0 20470 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_37
timestamp 1655484843
transform 1 0 19918 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_38
timestamp 1655484843
transform 1 0 20102 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_39
timestamp 1655484843
transform 1 0 19458 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_40
timestamp 1655484843
transform 1 0 20654 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_41
timestamp 1655484843
transform 1 0 20194 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_42
timestamp 1655484843
transform 1 0 21942 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_43
timestamp 1655484843
transform 1 0 20194 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_44
timestamp 1655484843
transform 1 0 20654 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_45
timestamp 1655484843
transform 1 0 19918 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_46
timestamp 1655484843
transform 1 0 21482 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_47
timestamp 1655484843
transform 1 0 20654 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_48
timestamp 1655484843
transform 1 0 20838 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_49
timestamp 1655484843
transform 1 0 19734 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_50
timestamp 1655484843
transform 1 0 20654 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_51
timestamp 1655484843
transform 1 0 20194 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_52
timestamp 1655484843
transform 1 0 14122 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_53
timestamp 1655484843
transform 1 0 13923 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_54
timestamp 1655484843
transform 1 0 13754 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_55
timestamp 1655484843
transform 1 0 15134 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_56
timestamp 1655484843
transform 1 0 15042 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_57
timestamp 1655484843
transform 1 0 21758 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_58
timestamp 1655484843
transform 1 0 20930 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_59
timestamp 1655484843
transform 1 0 20654 0 1 14637
box -29 -23 29 23
use L1M1_PR  L1M1_PR_60
timestamp 1655484843
transform 1 0 20654 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_61
timestamp 1655484843
transform 1 0 20470 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_62
timestamp 1655484843
transform 1 0 20470 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_63
timestamp 1655484843
transform 1 0 20470 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_64
timestamp 1655484843
transform 1 0 20470 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_65
timestamp 1655484843
transform 1 0 19550 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_66
timestamp 1655484843
transform 1 0 19274 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_67
timestamp 1655484843
transform 1 0 18998 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_68
timestamp 1655484843
transform 1 0 17894 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_69
timestamp 1655484843
transform 1 0 17894 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_70
timestamp 1655484843
transform 1 0 17802 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_71
timestamp 1655484843
transform 1 0 17158 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_72
timestamp 1655484843
transform 1 0 17066 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_73
timestamp 1655484843
transform 1 0 16974 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_74
timestamp 1655484843
transform 1 0 16790 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_75
timestamp 1655484843
transform 1 0 16422 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_76
timestamp 1655484843
transform 1 0 15870 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_77
timestamp 1655484843
transform 1 0 15870 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_78
timestamp 1655484843
transform 1 0 15686 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_79
timestamp 1655484843
transform 1 0 15318 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_80
timestamp 1655484843
transform 1 0 15318 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_81
timestamp 1655484843
transform 1 0 14582 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_82
timestamp 1655484843
transform 1 0 14214 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_83
timestamp 1655484843
transform 1 0 14122 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_84
timestamp 1655484843
transform 1 0 13202 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_85
timestamp 1655484843
transform 1 0 22126 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_86
timestamp 1655484843
transform 1 0 21022 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_87
timestamp 1655484843
transform 1 0 20930 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_88
timestamp 1655484843
transform 1 0 20930 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_89
timestamp 1655484843
transform 1 0 20930 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_90
timestamp 1655484843
transform 1 0 20838 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_91
timestamp 1655484843
transform 1 0 20470 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_92
timestamp 1655484843
transform 1 0 20274 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_93
timestamp 1655484843
transform 1 0 20102 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_94
timestamp 1655484843
transform 1 0 19642 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_95
timestamp 1655484843
transform 1 0 19458 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_96
timestamp 1655484843
transform 1 0 18354 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_97
timestamp 1655484843
transform 1 0 18170 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_98
timestamp 1655484843
transform 1 0 17526 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_99
timestamp 1655484843
transform 1 0 16790 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_100
timestamp 1655484843
transform 1 0 16790 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_101
timestamp 1655484843
transform 1 0 16698 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_102
timestamp 1655484843
transform 1 0 16606 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_103
timestamp 1655484843
transform 1 0 16422 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_104
timestamp 1655484843
transform 1 0 15686 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_105
timestamp 1655484843
transform 1 0 15686 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_106
timestamp 1655484843
transform 1 0 15502 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_107
timestamp 1655484843
transform 1 0 15502 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_108
timestamp 1655484843
transform 1 0 15318 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_109
timestamp 1655484843
transform 1 0 15318 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_110
timestamp 1655484843
transform 1 0 14582 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_111
timestamp 1655484843
transform 1 0 14214 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_112
timestamp 1655484843
transform 1 0 13754 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_113
timestamp 1655484843
transform 1 0 13662 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_114
timestamp 1655484843
transform 1 0 15134 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_115
timestamp 1655484843
transform 1 0 14214 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_116
timestamp 1655484843
transform 1 0 14398 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_117
timestamp 1655484843
transform 1 0 13294 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_118
timestamp 1655484843
transform 1 0 13202 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_119
timestamp 1655484843
transform 1 0 19826 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_120
timestamp 1655484843
transform 1 0 17526 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_121
timestamp 1655484843
transform 1 0 16790 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_122
timestamp 1655484843
transform 1 0 16514 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_123
timestamp 1655484843
transform 1 0 20286 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_124
timestamp 1655484843
transform 1 0 18369 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_125
timestamp 1655484843
transform 1 0 20378 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_126
timestamp 1655484843
transform 1 0 19075 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_127
timestamp 1655484843
transform 1 0 20286 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_128
timestamp 1655484843
transform 1 0 18615 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_129
timestamp 1655484843
transform 1 0 20363 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_130
timestamp 1655484843
transform 1 0 20286 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_131
timestamp 1655484843
transform 1 0 21574 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_132
timestamp 1655484843
transform 1 0 18799 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_133
timestamp 1655484843
transform 1 0 20286 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_134
timestamp 1655484843
transform 1 0 19075 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_135
timestamp 1655484843
transform 1 0 19070 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_136
timestamp 1655484843
transform 1 0 18998 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_137
timestamp 1655484843
transform 1 0 21221 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_138
timestamp 1655484843
transform 1 0 20930 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_139
timestamp 1655484843
transform 1 0 18799 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_140
timestamp 1655484843
transform 1 0 18722 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_141
timestamp 1655484843
transform 1 0 21206 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_142
timestamp 1655484843
transform 1 0 20853 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_143
timestamp 1655484843
transform 1 0 19366 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_144
timestamp 1655484843
transform 1 0 18799 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_145
timestamp 1655484843
transform 1 0 19075 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_146
timestamp 1655484843
transform 1 0 18078 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_147
timestamp 1655484843
transform 1 0 16499 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_148
timestamp 1655484843
transform 1 0 16054 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_149
timestamp 1655484843
transform 1 0 17909 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_150
timestamp 1655484843
transform 1 0 17342 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_151
timestamp 1655484843
transform 1 0 15395 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_152
timestamp 1655484843
transform 1 0 14306 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_153
timestamp 1655484843
transform 1 0 15134 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_154
timestamp 1655484843
transform 1 0 14505 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_155
timestamp 1655484843
transform 1 0 18645 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_156
timestamp 1655484843
transform 1 0 14858 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_157
timestamp 1655484843
transform 1 0 17357 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_158
timestamp 1655484843
transform 1 0 17158 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_159
timestamp 1655484843
transform 1 0 18645 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_160
timestamp 1655484843
transform 1 0 16974 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_161
timestamp 1655484843
transform 1 0 17342 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_162
timestamp 1655484843
transform 1 0 17081 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_163
timestamp 1655484843
transform 1 0 15211 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_164
timestamp 1655484843
transform 1 0 15134 0 1 12886
box -29 -23 29 23
use L1M1_PR  L1M1_PR_165
timestamp 1655484843
transform 1 0 17357 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_166
timestamp 1655484843
transform 1 0 16238 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_167
timestamp 1655484843
transform 1 0 14291 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_168
timestamp 1655484843
transform 1 0 14030 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_169
timestamp 1655484843
transform 1 0 16345 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_170
timestamp 1655484843
transform 1 0 15870 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_171
timestamp 1655484843
transform 1 0 16238 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_172
timestamp 1655484843
transform 1 0 15793 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_173
timestamp 1655484843
transform 1 0 18001 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_174
timestamp 1655484843
transform 1 0 17710 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_175
timestamp 1655484843
transform 1 0 17618 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_176
timestamp 1655484843
transform 1 0 17143 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_177
timestamp 1655484843
transform 1 0 19642 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_178
timestamp 1655484843
transform 1 0 16698 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_179
timestamp 1655484843
transform 1 0 16606 0 1 14110
box -29 -23 29 23
use L1M1_PR  L1M1_PR_180
timestamp 1655484843
transform 1 0 14306 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_181
timestamp 1655484843
transform 1 0 18906 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_182
timestamp 1655484843
transform 1 0 18906 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_183
timestamp 1655484843
transform 1 0 18814 0 1 14722
box -29 -23 29 23
use L1M1_PR  L1M1_PR_184
timestamp 1655484843
transform 1 0 18814 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_185
timestamp 1655484843
transform 1 0 18630 0 1 12546
box -29 -23 29 23
use L1M1_PR  L1M1_PR_186
timestamp 1655484843
transform 1 0 17342 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_187
timestamp 1655484843
transform 1 0 15502 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_188
timestamp 1655484843
transform 1 0 14950 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_189
timestamp 1655484843
transform 1 0 14030 0 1 11458
box -29 -23 29 23
use L1M1_PR  L1M1_PR_190
timestamp 1655484843
transform 1 0 20102 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_191
timestamp 1655484843
transform 1 0 18814 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_192
timestamp 1655484843
transform 1 0 18538 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_193
timestamp 1655484843
transform 1 0 18538 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_194
timestamp 1655484843
transform 1 0 18354 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_195
timestamp 1655484843
transform 1 0 18354 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_196
timestamp 1655484843
transform 1 0 17618 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_197
timestamp 1655484843
transform 1 0 16882 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_198
timestamp 1655484843
transform 1 0 16606 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_199
timestamp 1655484843
transform 1 0 16054 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_200
timestamp 1655484843
transform 1 0 21482 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_201
timestamp 1655484843
transform 1 0 21114 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_202
timestamp 1655484843
transform 1 0 18814 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_203
timestamp 1655484843
transform 1 0 18538 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_204
timestamp 1655484843
transform 1 0 18538 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_205
timestamp 1655484843
transform 1 0 18538 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_206
timestamp 1655484843
transform 1 0 18170 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_207
timestamp 1655484843
transform 1 0 17618 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_208
timestamp 1655484843
transform 1 0 16238 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_209
timestamp 1655484843
transform 1 0 15134 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_210
timestamp 1655484843
transform 1 0 14766 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_211
timestamp 1655484843
transform 1 0 18354 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_212
timestamp 1655484843
transform 1 0 18262 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_213
timestamp 1655484843
transform 1 0 18170 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_214
timestamp 1655484843
transform 1 0 17802 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_215
timestamp 1655484843
transform 1 0 6854 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_216
timestamp 1655484843
transform 1 0 6578 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_217
timestamp 1655484843
transform 1 0 6946 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_218
timestamp 1655484843
transform 1 0 6578 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_219
timestamp 1655484843
transform 1 0 7498 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_220
timestamp 1655484843
transform 1 0 6670 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_221
timestamp 1655484843
transform 1 0 8602 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_222
timestamp 1655484843
transform 1 0 7958 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_223
timestamp 1655484843
transform 1 0 9706 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_224
timestamp 1655484843
transform 1 0 9062 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_225
timestamp 1655484843
transform 1 0 9982 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_226
timestamp 1655484843
transform 1 0 9522 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_227
timestamp 1655484843
transform 1 0 6210 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_228
timestamp 1655484843
transform 1 0 6118 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_229
timestamp 1655484843
transform 1 0 10074 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_230
timestamp 1655484843
transform 1 0 9982 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_231
timestamp 1655484843
transform 1 0 9798 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_232
timestamp 1655484843
transform 1 0 9430 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_233
timestamp 1655484843
transform 1 0 9706 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_234
timestamp 1655484843
transform 1 0 9154 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_235
timestamp 1655484843
transform 1 0 8878 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_236
timestamp 1655484843
transform 1 0 9890 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_237
timestamp 1655484843
transform 1 0 9522 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_238
timestamp 1655484843
transform 1 0 9430 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_239
timestamp 1655484843
transform 1 0 8786 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_240
timestamp 1655484843
transform 1 0 8786 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_241
timestamp 1655484843
transform 1 0 8326 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_242
timestamp 1655484843
transform 1 0 9154 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_243
timestamp 1655484843
transform 1 0 8694 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_244
timestamp 1655484843
transform 1 0 7682 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_245
timestamp 1655484843
transform 1 0 9062 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_246
timestamp 1655484843
transform 1 0 8234 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_247
timestamp 1655484843
transform 1 0 6762 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_248
timestamp 1655484843
transform 1 0 9246 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_249
timestamp 1655484843
transform 1 0 8602 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_250
timestamp 1655484843
transform 1 0 6670 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_251
timestamp 1655484843
transform 1 0 8510 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_252
timestamp 1655484843
transform 1 0 7130 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_253
timestamp 1655484843
transform 1 0 6302 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_254
timestamp 1655484843
transform 1 0 9154 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_255
timestamp 1655484843
transform 1 0 8786 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_256
timestamp 1655484843
transform 1 0 8786 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_257
timestamp 1655484843
transform 1 0 6302 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_258
timestamp 1655484843
transform 1 0 8878 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_259
timestamp 1655484843
transform 1 0 8602 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_260
timestamp 1655484843
transform 1 0 9154 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_261
timestamp 1655484843
transform 1 0 9062 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_262
timestamp 1655484843
transform 1 0 9154 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_263
timestamp 1655484843
transform 1 0 9062 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_264
timestamp 1655484843
transform 1 0 7667 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_265
timestamp 1655484843
transform 1 0 7038 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_266
timestamp 1655484843
transform 1 0 9062 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_267
timestamp 1655484843
transform 1 0 8341 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_268
timestamp 1655484843
transform 1 0 7483 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_269
timestamp 1655484843
transform 1 0 6762 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_270
timestamp 1655484843
transform 1 0 7115 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_271
timestamp 1655484843
transform 1 0 6946 0 1 19210
box -29 -23 29 23
use L1M1_PR  L1M1_PR_272
timestamp 1655484843
transform 1 0 7866 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_273
timestamp 1655484843
transform 1 0 7575 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_274
timestamp 1655484843
transform 1 0 7406 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_275
timestamp 1655484843
transform 1 0 7213 0 1 15665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_276
timestamp 1655484843
transform 1 0 10641 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_277
timestamp 1655484843
transform 1 0 10626 0 1 17238
box -29 -23 29 23
use L1M1_PR  L1M1_PR_278
timestamp 1655484843
transform 1 0 10350 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_279
timestamp 1655484843
transform 1 0 10273 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_280
timestamp 1655484843
transform 1 0 10917 0 1 20784
box -29 -23 29 23
use L1M1_PR  L1M1_PR_281
timestamp 1655484843
transform 1 0 10534 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_282
timestamp 1655484843
transform 1 0 19182 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_283
timestamp 1655484843
transform 1 0 17158 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_284
timestamp 1655484843
transform 1 0 16606 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_285
timestamp 1655484843
transform 1 0 13386 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_286
timestamp 1655484843
transform 1 0 11929 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_287
timestamp 1655484843
transform 1 0 9430 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_288
timestamp 1655484843
transform 1 0 19458 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_289
timestamp 1655484843
transform 1 0 17342 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_290
timestamp 1655484843
transform 1 0 16330 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_291
timestamp 1655484843
transform 1 0 14766 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_292
timestamp 1655484843
transform 1 0 13202 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_293
timestamp 1655484843
transform 1 0 9154 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_294
timestamp 1655484843
transform 1 0 9062 0 1 15878
box -29 -23 29 23
use L1M1_PR  L1M1_PR_295
timestamp 1655484843
transform 1 0 8694 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_296
timestamp 1655484843
transform 1 0 6946 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_297
timestamp 1655484843
transform 1 0 6486 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_298
timestamp 1655484843
transform 1 0 6118 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_299
timestamp 1655484843
transform 1 0 8326 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_300
timestamp 1655484843
transform 1 0 8326 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_301
timestamp 1655484843
transform 1 0 9430 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_302
timestamp 1655484843
transform 1 0 7866 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_303
timestamp 1655484843
transform 1 0 10534 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_304
timestamp 1655484843
transform 1 0 10258 0 1 17374
box -29 -23 29 23
use L1M1_PR  L1M1_PR_305
timestamp 1655484843
transform 1 0 10718 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_306
timestamp 1655484843
transform 1 0 10350 0 1 19210
box -29 -23 29 23
use L1M1_PR  L1M1_PR_307
timestamp 1655484843
transform 1 0 10166 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_308
timestamp 1655484843
transform 1 0 10166 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_309
timestamp 1655484843
transform 1 0 18814 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_310
timestamp 1655484843
transform 1 0 16054 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_311
timestamp 1655484843
transform 1 0 15962 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_312
timestamp 1655484843
transform 1 0 15502 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_313
timestamp 1655484843
transform 1 0 13662 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_314
timestamp 1655484843
transform 1 0 13662 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_315
timestamp 1655484843
transform 1 0 13386 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_316
timestamp 1655484843
transform 1 0 13386 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_317
timestamp 1655484843
transform 1 0 13386 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_318
timestamp 1655484843
transform 1 0 14490 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_319
timestamp 1655484843
transform 1 0 14490 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_320
timestamp 1655484843
transform 1 0 14398 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_321
timestamp 1655484843
transform 1 0 14398 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_322
timestamp 1655484843
transform 1 0 14030 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_323
timestamp 1655484843
transform 1 0 13386 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_324
timestamp 1655484843
transform 1 0 21574 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_325
timestamp 1655484843
transform 1 0 21482 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_326
timestamp 1655484843
transform 1 0 21482 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_327
timestamp 1655484843
transform 1 0 21482 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_328
timestamp 1655484843
transform 1 0 21390 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_329
timestamp 1655484843
transform 1 0 21390 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_330
timestamp 1655484843
transform 1 0 18630 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_331
timestamp 1655484843
transform 1 0 18078 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_332
timestamp 1655484843
transform 1 0 20102 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_333
timestamp 1655484843
transform 1 0 20102 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_334
timestamp 1655484843
transform 1 0 19826 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_335
timestamp 1655484843
transform 1 0 17894 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_336
timestamp 1655484843
transform 1 0 17710 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_337
timestamp 1655484843
transform 1 0 17342 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_338
timestamp 1655484843
transform 1 0 17250 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_339
timestamp 1655484843
transform 1 0 20562 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_340
timestamp 1655484843
transform 1 0 19826 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_341
timestamp 1655484843
transform 1 0 20286 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_342
timestamp 1655484843
transform 1 0 19550 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_343
timestamp 1655484843
transform 1 0 21574 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_344
timestamp 1655484843
transform 1 0 20746 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_345
timestamp 1655484843
transform 1 0 21850 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_346
timestamp 1655484843
transform 1 0 21482 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_347
timestamp 1655484843
transform 1 0 22402 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_348
timestamp 1655484843
transform 1 0 21942 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_349
timestamp 1655484843
transform 1 0 22034 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_350
timestamp 1655484843
transform 1 0 19826 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_351
timestamp 1655484843
transform 1 0 21574 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_352
timestamp 1655484843
transform 1 0 19366 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_353
timestamp 1655484843
transform 1 0 22034 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_354
timestamp 1655484843
transform 1 0 21482 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_355
timestamp 1655484843
transform 1 0 22509 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_356
timestamp 1655484843
transform 1 0 21114 0 1 19210
box -29 -23 29 23
use L1M1_PR  L1M1_PR_357
timestamp 1655484843
transform 1 0 20079 0 1 19142
box -29 -23 29 23
use L1M1_PR  L1M1_PR_358
timestamp 1655484843
transform 1 0 19090 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_359
timestamp 1655484843
transform 1 0 18055 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_360
timestamp 1655484843
transform 1 0 15962 0 1 19210
box -29 -23 29 23
use L1M1_PR  L1M1_PR_361
timestamp 1655484843
transform 1 0 14927 0 1 19142
box -29 -23 29 23
use L1M1_PR  L1M1_PR_362
timestamp 1655484843
transform 1 0 14030 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_363
timestamp 1655484843
transform 1 0 13386 0 1 19142
box -29 -23 29 23
use L1M1_PR  L1M1_PR_364
timestamp 1655484843
transform 1 0 12903 0 1 18394
box -29 -23 29 23
use L1M1_PR  L1M1_PR_365
timestamp 1655484843
transform 1 0 12351 0 1 19142
box -29 -23 29 23
use L1M1_PR  L1M1_PR_366
timestamp 1655484843
transform 1 0 11914 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_367
timestamp 1655484843
transform 1 0 13041 0 1 18054
box -29 -23 29 23
use L1M1_PR  L1M1_PR_368
timestamp 1655484843
transform 1 0 12006 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_369
timestamp 1655484843
transform 1 0 13033 0 1 16966
box -29 -23 29 23
use L1M1_PR  L1M1_PR_370
timestamp 1655484843
transform 1 0 12190 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_371
timestamp 1655484843
transform 1 0 11270 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_372
timestamp 1655484843
transform 1 0 11071 0 1 15130
box -29 -23 29 23
use L1M1_PR  L1M1_PR_373
timestamp 1655484843
transform 1 0 12305 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_374
timestamp 1655484843
transform 1 0 10626 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_375
timestamp 1655484843
transform 1 0 11753 0 1 12954
box -29 -23 29 23
use L1M1_PR  L1M1_PR_376
timestamp 1655484843
transform 1 0 10626 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_377
timestamp 1655484843
transform 1 0 11753 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_378
timestamp 1655484843
transform 1 0 10442 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_379
timestamp 1655484843
transform 1 0 11569 0 1 10778
box -29 -23 29 23
use L1M1_PR  L1M1_PR_380
timestamp 1655484843
transform 1 0 10718 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_381
timestamp 1655484843
transform 1 0 11753 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_382
timestamp 1655484843
transform 1 0 10534 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_383
timestamp 1655484843
transform 1 0 20102 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_384
timestamp 1655484843
transform 1 0 17526 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_385
timestamp 1655484843
transform 1 0 17526 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_386
timestamp 1655484843
transform 1 0 11661 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_387
timestamp 1655484843
transform 1 0 21229 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_388
timestamp 1655484843
transform 1 0 20102 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_389
timestamp 1655484843
transform 1 0 21229 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_390
timestamp 1655484843
transform 1 0 16422 0 1 6086
box -29 -23 29 23
use L1M1_PR  L1M1_PR_391
timestamp 1655484843
transform 1 0 24058 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_392
timestamp 1655484843
transform 1 0 24058 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_393
timestamp 1655484843
transform 1 0 22126 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_394
timestamp 1655484843
transform 1 0 21022 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_395
timestamp 1655484843
transform 1 0 22509 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_396
timestamp 1655484843
transform 1 0 22034 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_397
timestamp 1655484843
transform 1 0 23874 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_398
timestamp 1655484843
transform 1 0 23874 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_399
timestamp 1655484843
transform 1 0 22509 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_400
timestamp 1655484843
transform 1 0 21206 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_401
timestamp 1655484843
transform 1 0 19075 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_402
timestamp 1655484843
transform 1 0 17894 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_403
timestamp 1655484843
transform 1 0 22509 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_404
timestamp 1655484843
transform 1 0 22494 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_405
timestamp 1655484843
transform 1 0 23506 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_406
timestamp 1655484843
transform 1 0 23506 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_407
timestamp 1655484843
transform 1 0 22601 0 1 18938
box -29 -23 29 23
use L1M1_PR  L1M1_PR_408
timestamp 1655484843
transform 1 0 22310 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_409
timestamp 1655484843
transform 1 0 21651 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_410
timestamp 1655484843
transform 1 0 21574 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_411
timestamp 1655484843
transform 1 0 23782 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_412
timestamp 1655484843
transform 1 0 23782 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_413
timestamp 1655484843
transform 1 0 22233 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_414
timestamp 1655484843
transform 1 0 22034 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_415
timestamp 1655484843
transform 1 0 22509 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_416
timestamp 1655484843
transform 1 0 22494 0 1 15062
box -29 -23 29 23
use L1M1_PR  L1M1_PR_417
timestamp 1655484843
transform 1 0 22233 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_418
timestamp 1655484843
transform 1 0 22034 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_419
timestamp 1655484843
transform 1 0 22509 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_420
timestamp 1655484843
transform 1 0 21942 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_421
timestamp 1655484843
transform 1 0 22693 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_422
timestamp 1655484843
transform 1 0 22310 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_423
timestamp 1655484843
transform 1 0 19933 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_424
timestamp 1655484843
transform 1 0 16790 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_425
timestamp 1655484843
transform 1 0 16499 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_426
timestamp 1655484843
transform 1 0 16330 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_427
timestamp 1655484843
transform 1 0 15517 0 1 21114
box -29 -23 29 23
use L1M1_PR  L1M1_PR_428
timestamp 1655484843
transform 1 0 15502 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_429
timestamp 1655484843
transform 1 0 13095 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_430
timestamp 1655484843
transform 1 0 12742 0 1 19686
box -29 -23 29 23
use L1M1_PR  L1M1_PR_431
timestamp 1655484843
transform 1 0 12926 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_432
timestamp 1655484843
transform 1 0 11071 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_433
timestamp 1655484843
transform 1 0 12742 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_434
timestamp 1655484843
transform 1 0 12359 0 1 15665
box -29 -23 29 23
use L1M1_PR  L1M1_PR_435
timestamp 1655484843
transform 1 0 14030 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_436
timestamp 1655484843
transform 1 0 13003 0 1 14246
box -29 -23 29 23
use L1M1_PR  L1M1_PR_437
timestamp 1655484843
transform 1 0 14214 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_438
timestamp 1655484843
transform 1 0 13095 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_439
timestamp 1655484843
transform 1 0 13294 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_440
timestamp 1655484843
transform 1 0 13033 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_441
timestamp 1655484843
transform 1 0 12354 0 1 11313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_442
timestamp 1655484843
transform 1 0 11822 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_443
timestamp 1655484843
transform 1 0 12354 0 1 10225
box -29 -23 29 23
use L1M1_PR  L1M1_PR_444
timestamp 1655484843
transform 1 0 11822 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_445
timestamp 1655484843
transform 1 0 13386 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_446
timestamp 1655484843
transform 1 0 12665 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_447
timestamp 1655484843
transform 1 0 13018 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_448
timestamp 1655484843
transform 1 0 12635 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_449
timestamp 1655484843
transform 1 0 16499 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_450
timestamp 1655484843
transform 1 0 15778 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_451
timestamp 1655484843
transform 1 0 19535 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_452
timestamp 1655484843
transform 1 0 19182 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_453
timestamp 1655484843
transform 1 0 21651 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_454
timestamp 1655484843
transform 1 0 18078 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_455
timestamp 1655484843
transform 1 0 23138 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_456
timestamp 1655484843
transform 1 0 23138 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_457
timestamp 1655484843
transform 1 0 22494 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_458
timestamp 1655484843
transform 1 0 22402 0 1 14042
box -29 -23 29 23
use L1M1_PR  L1M1_PR_459
timestamp 1655484843
transform 1 0 20746 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_460
timestamp 1655484843
transform 1 0 20194 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_461
timestamp 1655484843
transform 1 0 18998 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_462
timestamp 1655484843
transform 1 0 18354 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_463
timestamp 1655484843
transform 1 0 22126 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_464
timestamp 1655484843
transform 1 0 21114 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_465
timestamp 1655484843
transform 1 0 22402 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_466
timestamp 1655484843
transform 1 0 21942 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_467
timestamp 1655484843
transform 1 0 23690 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_468
timestamp 1655484843
transform 1 0 23690 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_469
timestamp 1655484843
transform 1 0 22310 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_470
timestamp 1655484843
transform 1 0 21942 0 1 11866
box -29 -23 29 23
use L1M1_PR  L1M1_PR_471
timestamp 1655484843
transform 1 0 21666 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_472
timestamp 1655484843
transform 1 0 21574 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_473
timestamp 1655484843
transform 1 0 22034 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_474
timestamp 1655484843
transform 1 0 18998 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_475
timestamp 1655484843
transform 1 0 22494 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_476
timestamp 1655484843
transform 1 0 22402 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_477
timestamp 1655484843
transform 1 0 23138 0 1 20570
box -29 -23 29 23
use L1M1_PR  L1M1_PR_478
timestamp 1655484843
transform 1 0 21574 0 1 20570
box -29 -23 29 23
use L1M1_PR  L1M1_PR_479
timestamp 1655484843
transform 1 0 21850 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_480
timestamp 1655484843
transform 1 0 19734 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_481
timestamp 1655484843
transform 1 0 17342 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_482
timestamp 1655484843
transform 1 0 16422 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_483
timestamp 1655484843
transform 1 0 15870 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_484
timestamp 1655484843
transform 1 0 14582 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_485
timestamp 1655484843
transform 1 0 15134 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_486
timestamp 1655484843
transform 1 0 12558 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_487
timestamp 1655484843
transform 1 0 12374 0 1 19482
box -29 -23 29 23
use L1M1_PR  L1M1_PR_488
timestamp 1655484843
transform 1 0 12006 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_489
timestamp 1655484843
transform 1 0 13386 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_490
timestamp 1655484843
transform 1 0 13294 0 1 17306
box -29 -23 29 23
use L1M1_PR  L1M1_PR_491
timestamp 1655484843
transform 1 0 13386 0 1 16694
box -29 -23 29 23
use L1M1_PR  L1M1_PR_492
timestamp 1655484843
transform 1 0 13202 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_493
timestamp 1655484843
transform 1 0 13662 0 1 14790
box -29 -23 29 23
use L1M1_PR  L1M1_PR_494
timestamp 1655484843
transform 1 0 10718 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_495
timestamp 1655484843
transform 1 0 13846 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_496
timestamp 1655484843
transform 1 0 12834 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_497
timestamp 1655484843
transform 1 0 12926 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_498
timestamp 1655484843
transform 1 0 12190 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_499
timestamp 1655484843
transform 1 0 12098 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_500
timestamp 1655484843
transform 1 0 11454 0 1 11526
box -29 -23 29 23
use L1M1_PR  L1M1_PR_501
timestamp 1655484843
transform 1 0 11914 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_502
timestamp 1655484843
transform 1 0 11362 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_503
timestamp 1655484843
transform 1 0 13018 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_504
timestamp 1655484843
transform 1 0 12075 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_505
timestamp 1655484843
transform 1 0 21574 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_506
timestamp 1655484843
transform 1 0 15226 0 1 7174
box -29 -23 29 23
use L1M1_PR  L1M1_PR_507
timestamp 1655484843
transform 1 0 21574 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_508
timestamp 1655484843
transform 1 0 18814 0 1 7174
box -29 -23 29 23
use L1M1_PR  L1M1_PR_509
timestamp 1655484843
transform 1 0 22678 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_510
timestamp 1655484843
transform 1 0 20562 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_511
timestamp 1655484843
transform 1 0 19182 0 1 21862
box -29 -23 29 23
use L1M1_PR  L1M1_PR_512
timestamp 1655484843
transform 1 0 18446 0 1 21930
box -29 -23 29 23
use L1M1_PR  L1M1_PR_513
timestamp 1655484843
transform 1 0 22770 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_514
timestamp 1655484843
transform 1 0 20930 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_515
timestamp 1655484843
transform 1 0 20286 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_516
timestamp 1655484843
transform 1 0 18998 0 1 21862
box -29 -23 29 23
use L1M1_PR  L1M1_PR_517
timestamp 1655484843
transform 1 0 18354 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_518
timestamp 1655484843
transform 1 0 18170 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_519
timestamp 1655484843
transform 1 0 18630 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_520
timestamp 1655484843
transform 1 0 17894 0 1 21114
box -29 -23 29 23
use L1M1_PR  L1M1_PR_521
timestamp 1655484843
transform 1 0 17158 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_522
timestamp 1655484843
transform 1 0 17986 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_523
timestamp 1655484843
transform 1 0 17434 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_524
timestamp 1655484843
transform 1 0 15686 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_525
timestamp 1655484843
transform 1 0 15962 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_526
timestamp 1655484843
transform 1 0 15870 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_527
timestamp 1655484843
transform 1 0 15226 0 1 21862
box -29 -23 29 23
use L1M1_PR  L1M1_PR_528
timestamp 1655484843
transform 1 0 15686 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_529
timestamp 1655484843
transform 1 0 15134 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_530
timestamp 1655484843
transform 1 0 15042 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_531
timestamp 1655484843
transform 1 0 14306 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_532
timestamp 1655484843
transform 1 0 13846 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_533
timestamp 1655484843
transform 1 0 14306 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_534
timestamp 1655484843
transform 1 0 14122 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_535
timestamp 1655484843
transform 1 0 11730 0 1 19074
box -29 -23 29 23
use L1M1_PR  L1M1_PR_536
timestamp 1655484843
transform 1 0 11270 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_537
timestamp 1655484843
transform 1 0 11914 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_538
timestamp 1655484843
transform 1 0 11822 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_539
timestamp 1655484843
transform 1 0 11454 0 1 18938
box -29 -23 29 23
use L1M1_PR  L1M1_PR_540
timestamp 1655484843
transform 1 0 11822 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_541
timestamp 1655484843
transform 1 0 11638 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_542
timestamp 1655484843
transform 1 0 11546 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_543
timestamp 1655484843
transform 1 0 11822 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_544
timestamp 1655484843
transform 1 0 11822 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_545
timestamp 1655484843
transform 1 0 11362 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_546
timestamp 1655484843
transform 1 0 10166 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_547
timestamp 1655484843
transform 1 0 11822 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_548
timestamp 1655484843
transform 1 0 11454 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_549
timestamp 1655484843
transform 1 0 10442 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_550
timestamp 1655484843
transform 1 0 10350 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_551
timestamp 1655484843
transform 1 0 9338 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_552
timestamp 1655484843
transform 1 0 9315 0 1 14790
box -29 -23 29 23
use L1M1_PR  L1M1_PR_553
timestamp 1655484843
transform 1 0 10373 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_554
timestamp 1655484843
transform 1 0 8786 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_555
timestamp 1655484843
transform 1 0 10626 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_556
timestamp 1655484843
transform 1 0 9821 0 1 12614
box -29 -23 29 23
use L1M1_PR  L1M1_PR_557
timestamp 1655484843
transform 1 0 9591 0 1 11526
box -29 -23 29 23
use L1M1_PR  L1M1_PR_558
timestamp 1655484843
transform 1 0 9338 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_559
timestamp 1655484843
transform 1 0 9522 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_560
timestamp 1655484843
transform 1 0 8211 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_561
timestamp 1655484843
transform 1 0 10626 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_562
timestamp 1655484843
transform 1 0 8495 0 1 8602
box -29 -23 29 23
use L1M1_PR  L1M1_PR_563
timestamp 1655484843
transform 1 0 11753 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_564
timestamp 1655484843
transform 1 0 11086 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_565
timestamp 1655484843
transform 1 0 13294 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_566
timestamp 1655484843
transform 1 0 12374 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_567
timestamp 1655484843
transform 1 0 12213 0 1 7174
box -29 -23 29 23
use L1M1_PR  L1M1_PR_568
timestamp 1655484843
transform 1 0 15211 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_569
timestamp 1655484843
transform 1 0 13202 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_570
timestamp 1655484843
transform 1 0 12635 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_571
timestamp 1655484843
transform 1 0 11730 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_572
timestamp 1655484843
transform 1 0 11347 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_573
timestamp 1655484843
transform 1 0 11270 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_574
timestamp 1655484843
transform 1 0 9599 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_575
timestamp 1655484843
transform 1 0 9246 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_576
timestamp 1655484843
transform 1 0 10350 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_577
timestamp 1655484843
transform 1 0 9599 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_578
timestamp 1655484843
transform 1 0 9507 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_579
timestamp 1655484843
transform 1 0 9338 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_580
timestamp 1655484843
transform 1 0 9890 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_581
timestamp 1655484843
transform 1 0 7759 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_582
timestamp 1655484843
transform 1 0 10074 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_583
timestamp 1655484843
transform 1 0 7575 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_584
timestamp 1655484843
transform 1 0 12205 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_585
timestamp 1655484843
transform 1 0 10166 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_586
timestamp 1655484843
transform 1 0 9783 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_587
timestamp 1655484843
transform 1 0 9614 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_588
timestamp 1655484843
transform 1 0 11454 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_589
timestamp 1655484843
transform 1 0 10617 0 1 16432
box -29 -23 29 23
use L1M1_PR  L1M1_PR_590
timestamp 1655484843
transform 1 0 10979 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_591
timestamp 1655484843
transform 1 0 10902 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_592
timestamp 1655484843
transform 1 0 12834 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_593
timestamp 1655484843
transform 1 0 12635 0 1 20784
box -29 -23 29 23
use L1M1_PR  L1M1_PR_594
timestamp 1655484843
transform 1 0 15333 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_595
timestamp 1655484843
transform 1 0 14950 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_596
timestamp 1655484843
transform 1 0 16238 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_597
timestamp 1655484843
transform 1 0 16223 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_598
timestamp 1655484843
transform 1 0 18921 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_599
timestamp 1655484843
transform 1 0 18906 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_600
timestamp 1655484843
transform 1 0 20082 0 1 21105
box -29 -23 29 23
use L1M1_PR  L1M1_PR_601
timestamp 1655484843
transform 1 0 19366 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_602
timestamp 1655484843
transform 1 0 20363 0 1 20774
box -29 -23 29 23
use L1M1_PR  L1M1_PR_603
timestamp 1655484843
transform 1 0 19918 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_604
timestamp 1655484843
transform 1 0 20746 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_605
timestamp 1655484843
transform 1 0 19734 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_606
timestamp 1655484843
transform 1 0 20102 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_607
timestamp 1655484843
transform 1 0 19550 0 1 21658
box -29 -23 29 23
use L1M1_PR  L1M1_PR_608
timestamp 1655484843
transform 1 0 19274 0 1 21318
box -29 -23 29 23
use L1M1_PR  L1M1_PR_609
timestamp 1655484843
transform 1 0 19182 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_610
timestamp 1655484843
transform 1 0 15410 0 1 21590
box -29 -23 29 23
use L1M1_PR  L1M1_PR_611
timestamp 1655484843
transform 1 0 15410 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_612
timestamp 1655484843
transform 1 0 11270 0 1 19142
box -29 -23 29 23
use L1M1_PR  L1M1_PR_613
timestamp 1655484843
transform 1 0 10534 0 1 19142
box -29 -23 29 23
use L1M1_PR  L1M1_PR_614
timestamp 1655484843
transform 1 0 11822 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_615
timestamp 1655484843
transform 1 0 11362 0 1 17034
box -29 -23 29 23
use L1M1_PR  L1M1_PR_616
timestamp 1655484843
transform 1 0 9982 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_617
timestamp 1655484843
transform 1 0 9246 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_618
timestamp 1655484843
transform 1 0 9798 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_619
timestamp 1655484843
transform 1 0 8786 0 1 14858
box -29 -23 29 23
use L1M1_PR  L1M1_PR_620
timestamp 1655484843
transform 1 0 10718 0 1 13430
box -29 -23 29 23
use L1M1_PR  L1M1_PR_621
timestamp 1655484843
transform 1 0 10442 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_622
timestamp 1655484843
transform 1 0 10258 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_623
timestamp 1655484843
transform 1 0 10166 0 1 12342
box -29 -23 29 23
use L1M1_PR  L1M1_PR_624
timestamp 1655484843
transform 1 0 9246 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_625
timestamp 1655484843
transform 1 0 8970 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_626
timestamp 1655484843
transform 1 0 9982 0 1 9690
box -29 -23 29 23
use L1M1_PR  L1M1_PR_627
timestamp 1655484843
transform 1 0 7866 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_628
timestamp 1655484843
transform 1 0 8878 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_629
timestamp 1655484843
transform 1 0 8142 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_630
timestamp 1655484843
transform 1 0 12098 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_631
timestamp 1655484843
transform 1 0 11638 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_632
timestamp 1655484843
transform 1 0 12558 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_633
timestamp 1655484843
transform 1 0 12190 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_634
timestamp 1655484843
transform 1 0 13386 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_635
timestamp 1655484843
transform 1 0 12834 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_636
timestamp 1655484843
transform 1 0 6762 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_637
timestamp 1655484843
transform 1 0 6578 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_638
timestamp 1655484843
transform 1 0 6486 0 1 12342
box -29 -23 29 23
use L1M1_PR  L1M1_PR_639
timestamp 1655484843
transform 1 0 6302 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_640
timestamp 1655484843
transform 1 0 7038 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_641
timestamp 1655484843
transform 1 0 6670 0 1 14110
box -29 -23 29 23
use L1M1_PR  L1M1_PR_642
timestamp 1655484843
transform 1 0 6670 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_643
timestamp 1655484843
transform 1 0 6946 0 1 12410
box -29 -23 29 23
use L1M1_PR  L1M1_PR_644
timestamp 1655484843
transform 1 0 6578 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_645
timestamp 1655484843
transform 1 0 6394 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_646
timestamp 1655484843
transform 1 0 6854 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_647
timestamp 1655484843
transform 1 0 6670 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_648
timestamp 1655484843
transform 1 0 6578 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_649
timestamp 1655484843
transform 1 0 6394 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_650
timestamp 1655484843
transform 1 0 7130 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_651
timestamp 1655484843
transform 1 0 6302 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_652
timestamp 1655484843
transform 1 0 6026 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_653
timestamp 1655484843
transform 1 0 6854 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_654
timestamp 1655484843
transform 1 0 6578 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_655
timestamp 1655484843
transform 1 0 5934 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_656
timestamp 1655484843
transform 1 0 7314 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_657
timestamp 1655484843
transform 1 0 6762 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_658
timestamp 1655484843
transform 1 0 6578 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_659
timestamp 1655484843
transform 1 0 6210 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_660
timestamp 1655484843
transform 1 0 8050 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_661
timestamp 1655484843
transform 1 0 7866 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_662
timestamp 1655484843
transform 1 0 7406 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_663
timestamp 1655484843
transform 1 0 6946 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_664
timestamp 1655484843
transform 1 0 10626 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_665
timestamp 1655484843
transform 1 0 8142 0 1 6570
box -29 -23 29 23
use L1M1_PR  L1M1_PR_666
timestamp 1655484843
transform 1 0 7682 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_667
timestamp 1655484843
transform 1 0 7958 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_668
timestamp 1655484843
transform 1 0 7590 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_669
timestamp 1655484843
transform 1 0 7498 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_670
timestamp 1655484843
transform 1 0 6762 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_671
timestamp 1655484843
transform 1 0 6210 0 1 6698
box -29 -23 29 23
use L1M1_PR  L1M1_PR_672
timestamp 1655484843
transform 1 0 7038 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_673
timestamp 1655484843
transform 1 0 6578 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_674
timestamp 1655484843
transform 1 0 6486 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_675
timestamp 1655484843
transform 1 0 6210 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_676
timestamp 1655484843
transform 1 0 5658 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_677
timestamp 1655484843
transform 1 0 7483 0 1 7718
box -29 -23 29 23
use L1M1_PR  L1M1_PR_678
timestamp 1655484843
transform 1 0 6946 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_679
timestamp 1655484843
transform 1 0 7207 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_680
timestamp 1655484843
transform 1 0 6946 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_681
timestamp 1655484843
transform 1 0 8495 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_682
timestamp 1655484843
transform 1 0 8234 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_683
timestamp 1655484843
transform 1 0 7202 0 1 8049
box -29 -23 29 23
use L1M1_PR  L1M1_PR_684
timestamp 1655484843
transform 1 0 6762 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_685
timestamp 1655484843
transform 1 0 7207 0 1 9137
box -29 -23 29 23
use L1M1_PR  L1M1_PR_686
timestamp 1655484843
transform 1 0 6854 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_687
timestamp 1655484843
transform 1 0 7575 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_688
timestamp 1655484843
transform 1 0 7038 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_689
timestamp 1655484843
transform 1 0 7202 0 1 11313
box -29 -23 29 23
use L1M1_PR  L1M1_PR_690
timestamp 1655484843
transform 1 0 6854 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_691
timestamp 1655484843
transform 1 0 7207 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_692
timestamp 1655484843
transform 1 0 6670 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_693
timestamp 1655484843
transform 1 0 8127 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_694
timestamp 1655484843
transform 1 0 7682 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_695
timestamp 1655484843
transform 1 0 6302 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_696
timestamp 1655484843
transform 1 0 6210 0 1 13770
box -29 -23 29 23
use L1M1_PR  L1M1_PR_697
timestamp 1655484843
transform 1 0 6486 0 1 11526
box -29 -23 29 23
use L1M1_PR  L1M1_PR_698
timestamp 1655484843
transform 1 0 6394 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_699
timestamp 1655484843
transform 1 0 6670 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_700
timestamp 1655484843
transform 1 0 6578 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_701
timestamp 1655484843
transform 1 0 6486 0 1 9350
box -29 -23 29 23
use L1M1_PR  L1M1_PR_702
timestamp 1655484843
transform 1 0 6394 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_703
timestamp 1655484843
transform 1 0 6394 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_704
timestamp 1655484843
transform 1 0 6302 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_705
timestamp 1655484843
transform 1 0 7866 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_706
timestamp 1655484843
transform 1 0 7774 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_707
timestamp 1655484843
transform 1 0 6578 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_708
timestamp 1655484843
transform 1 0 6578 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_709
timestamp 1655484843
transform 1 0 6486 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_710
timestamp 1655484843
transform 1 0 6394 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_711
timestamp 1655484843
transform 1 0 22770 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_712
timestamp 1655484843
transform 1 0 16882 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_713
timestamp 1655484843
transform 1 0 16223 0 1 9894
box -29 -23 29 23
use L1M1_PR  L1M1_PR_714
timestamp 1655484843
transform 1 0 20654 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_715
timestamp 1655484843
transform 1 0 18369 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_716
timestamp 1655484843
transform 1 0 17618 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_717
timestamp 1655484843
transform 1 0 15763 0 1 8738
box -29 -23 29 23
use L1M1_PR  L1M1_PR_718
timestamp 1655484843
transform 1 0 13754 0 1 9622
box -29 -23 29 23
use L1M1_PR  L1M1_PR_719
timestamp 1655484843
transform 1 0 13647 0 1 8806
box -29 -23 29 23
use L1M1_PR  L1M1_PR_720
timestamp 1655484843
transform 1 0 13923 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_721
timestamp 1655484843
transform 1 0 11546 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_722
timestamp 1655484843
transform 1 0 11546 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_723
timestamp 1655484843
transform 1 0 13647 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_724
timestamp 1655484843
transform 1 0 13478 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_725
timestamp 1655484843
transform 1 0 13647 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_726
timestamp 1655484843
transform 1 0 13478 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_727
timestamp 1655484843
transform 1 0 13923 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_728
timestamp 1655484843
transform 1 0 11914 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_729
timestamp 1655484843
transform 1 0 15211 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_730
timestamp 1655484843
transform 1 0 14214 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_731
timestamp 1655484843
transform 1 0 14751 0 1 14586
box -29 -23 29 23
use L1M1_PR  L1M1_PR_732
timestamp 1655484843
transform 1 0 14122 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_733
timestamp 1655484843
transform 1 0 14659 0 1 15674
box -29 -23 29 23
use L1M1_PR  L1M1_PR_734
timestamp 1655484843
transform 1 0 13478 0 1 15946
box -29 -23 29 23
use L1M1_PR  L1M1_PR_735
timestamp 1655484843
transform 1 0 13647 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_736
timestamp 1655484843
transform 1 0 12190 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_737
timestamp 1655484843
transform 1 0 14291 0 1 17850
box -29 -23 29 23
use L1M1_PR  L1M1_PR_738
timestamp 1655484843
transform 1 0 14214 0 1 19414
box -29 -23 29 23
use L1M1_PR  L1M1_PR_739
timestamp 1655484843
transform 1 0 14659 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_740
timestamp 1655484843
transform 1 0 14398 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_741
timestamp 1655484843
transform 1 0 17618 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_742
timestamp 1655484843
transform 1 0 17081 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_743
timestamp 1655484843
transform 1 0 18814 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_744
timestamp 1655484843
transform 1 0 17511 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_745
timestamp 1655484843
transform 1 0 21574 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_746
timestamp 1655484843
transform 1 0 20363 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_747
timestamp 1655484843
transform 1 0 21298 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_748
timestamp 1655484843
transform 1 0 20087 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_749
timestamp 1655484843
transform 1 0 21758 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_750
timestamp 1655484843
transform 1 0 21114 0 1 17306
box -29 -23 29 23
use L1M1_PR  L1M1_PR_751
timestamp 1655484843
transform 1 0 18155 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_752
timestamp 1655484843
transform 1 0 21390 0 1 14790
box -29 -23 29 23
use L1M1_PR  L1M1_PR_753
timestamp 1655484843
transform 1 0 20363 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_754
timestamp 1655484843
transform 1 0 19642 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_755
timestamp 1655484843
transform 1 0 22218 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_756
timestamp 1655484843
transform 1 0 21313 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_757
timestamp 1655484843
transform 1 0 21114 0 1 19754
box -29 -23 29 23
use L1M1_PR  L1M1_PR_758
timestamp 1655484843
transform 1 0 22770 0 1 12682
box -29 -23 29 23
use L1M1_PR  L1M1_PR_759
timestamp 1655484843
transform 1 0 21666 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_760
timestamp 1655484843
transform 1 0 21229 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_761
timestamp 1655484843
transform 1 0 21758 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_762
timestamp 1655484843
transform 1 0 21482 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_763
timestamp 1655484843
transform 1 0 21221 0 1 12002
box -29 -23 29 23
use L1M1_PR  L1M1_PR_764
timestamp 1655484843
transform 1 0 21390 0 1 13702
box -29 -23 29 23
use L1M1_PR  L1M1_PR_765
timestamp 1655484843
transform 1 0 20470 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_766
timestamp 1655484843
transform 1 0 19075 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_767
timestamp 1655484843
transform 1 0 21651 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_768
timestamp 1655484843
transform 1 0 20194 0 1 11526
box -29 -23 29 23
use L1M1_PR  L1M1_PR_769
timestamp 1655484843
transform 1 0 19642 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_770
timestamp 1655484843
transform 1 0 21390 0 1 11254
box -29 -23 29 23
use L1M1_PR  L1M1_PR_771
timestamp 1655484843
transform 1 0 21229 0 1 10982
box -29 -23 29 23
use L1M1_PR  L1M1_PR_772
timestamp 1655484843
transform 1 0 20838 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_773
timestamp 1655484843
transform 1 0 22034 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_774
timestamp 1655484843
transform 1 0 21651 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_775
timestamp 1655484843
transform 1 0 21390 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_776
timestamp 1655484843
transform 1 0 16606 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_777
timestamp 1655484843
transform 1 0 16330 0 1 6358
box -29 -23 29 23
use L1M1_PR  L1M1_PR_778
timestamp 1655484843
transform 1 0 13938 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_779
timestamp 1655484843
transform 1 0 12742 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_780
timestamp 1655484843
transform 1 0 13754 0 1 7786
box -29 -23 29 23
use L1M1_PR  L1M1_PR_781
timestamp 1655484843
transform 1 0 13754 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_782
timestamp 1655484843
transform 1 0 12466 0 1 8262
box -29 -23 29 23
use L1M1_PR  L1M1_PR_783
timestamp 1655484843
transform 1 0 12466 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_784
timestamp 1655484843
transform 1 0 10718 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_785
timestamp 1655484843
transform 1 0 10718 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_786
timestamp 1655484843
transform 1 0 10626 0 1 10506
box -29 -23 29 23
use L1M1_PR  L1M1_PR_787
timestamp 1655484843
transform 1 0 8878 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_788
timestamp 1655484843
transform 1 0 8694 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_789
timestamp 1655484843
transform 1 0 10902 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_790
timestamp 1655484843
transform 1 0 11914 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_791
timestamp 1655484843
transform 1 0 10994 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_792
timestamp 1655484843
transform 1 0 10350 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_793
timestamp 1655484843
transform 1 0 12190 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_794
timestamp 1655484843
transform 1 0 11730 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_795
timestamp 1655484843
transform 1 0 11730 0 1 16218
box -29 -23 29 23
use L1M1_PR  L1M1_PR_796
timestamp 1655484843
transform 1 0 12098 0 1 18666
box -29 -23 29 23
use L1M1_PR  L1M1_PR_797
timestamp 1655484843
transform 1 0 12006 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_798
timestamp 1655484843
transform 1 0 14582 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_799
timestamp 1655484843
transform 1 0 14030 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_800
timestamp 1655484843
transform 1 0 13754 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_801
timestamp 1655484843
transform 1 0 15870 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_802
timestamp 1655484843
transform 1 0 14214 0 1 19958
box -29 -23 29 23
use L1M1_PR  L1M1_PR_803
timestamp 1655484843
transform 1 0 17710 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_804
timestamp 1655484843
transform 1 0 17342 0 1 21386
box -29 -23 29 23
use L1M1_PR  L1M1_PR_805
timestamp 1655484843
transform 1 0 17342 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_806
timestamp 1655484843
transform 1 0 18078 0 1 21046
box -29 -23 29 23
use L1M1_PR  L1M1_PR_807
timestamp 1655484843
transform 1 0 17802 0 1 20502
box -29 -23 29 23
use L1M1_PR  L1M1_PR_808
timestamp 1655484843
transform 1 0 22862 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_809
timestamp 1655484843
transform 1 0 21482 0 1 20842
box -29 -23 29 23
use L1M1_PR  L1M1_PR_810
timestamp 1655484843
transform 1 0 20470 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_811
timestamp 1655484843
transform 1 0 21298 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_812
timestamp 1655484843
transform 1 0 21022 0 1 21794
box -29 -23 29 23
use L1M1_PR  L1M1_PR_813
timestamp 1655484843
transform 1 0 13754 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_814
timestamp 1655484843
transform 1 0 12558 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_815
timestamp 1655484843
transform 1 0 8602 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_816
timestamp 1655484843
transform 1 0 6118 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_817
timestamp 1655484843
transform 1 0 6118 0 1 6630
box -29 -23 29 23
use L1M1_PR  L1M1_PR_818
timestamp 1655484843
transform 1 0 6026 0 1 7242
box -29 -23 29 23
use L1M1_PR  L1M1_PR_819
timestamp 1655484843
transform 1 0 8326 0 1 6902
box -29 -23 29 23
use L1M1_PR  L1M1_PR_820
timestamp 1655484843
transform 1 0 6946 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_821
timestamp 1655484843
transform 1 0 6394 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_822
timestamp 1655484843
transform 1 0 10442 0 1 6154
box -29 -23 29 23
use L1M1_PR  L1M1_PR_823
timestamp 1655484843
transform 1 0 9614 0 1 6426
box -29 -23 29 23
use L1M1_PR  L1M1_PR_824
timestamp 1655484843
transform 1 0 8326 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_825
timestamp 1655484843
transform 1 0 7038 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_826
timestamp 1655484843
transform 1 0 6762 0 1 8534
box -29 -23 29 23
use L1M1_PR  L1M1_PR_827
timestamp 1655484843
transform 1 0 8326 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_828
timestamp 1655484843
transform 1 0 7038 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_829
timestamp 1655484843
transform 1 0 8694 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_830
timestamp 1655484843
transform 1 0 7038 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_831
timestamp 1655484843
transform 1 0 6578 0 1 10438
box -29 -23 29 23
use L1M1_PR  L1M1_PR_832
timestamp 1655484843
transform 1 0 8326 0 1 11594
box -29 -23 29 23
use L1M1_PR  L1M1_PR_833
timestamp 1655484843
transform 1 0 7130 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_834
timestamp 1655484843
transform 1 0 9246 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_835
timestamp 1655484843
transform 1 0 6854 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_836
timestamp 1655484843
transform 1 0 6762 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_837
timestamp 1655484843
transform 1 0 8418 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_838
timestamp 1655484843
transform 1 0 8326 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_839
timestamp 1655484843
transform 1 0 6578 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_840
timestamp 1655484843
transform 1 0 17894 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_841
timestamp 1655484843
transform 1 0 17342 0 1 9962
box -29 -23 29 23
use L1M1_PR  L1M1_PR_842
timestamp 1655484843
transform 1 0 17986 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_843
timestamp 1655484843
transform 1 0 17250 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_844
timestamp 1655484843
transform 1 0 16882 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_845
timestamp 1655484843
transform 1 0 16514 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_846
timestamp 1655484843
transform 1 0 15594 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_847
timestamp 1655484843
transform 1 0 14766 0 1 8874
box -29 -23 29 23
use L1M1_PR  L1M1_PR_848
timestamp 1655484843
transform 1 0 15042 0 1 9418
box -29 -23 29 23
use L1M1_PR  L1M1_PR_849
timestamp 1655484843
transform 1 0 14306 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_850
timestamp 1655484843
transform 1 0 15778 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_851
timestamp 1655484843
transform 1 0 14766 0 1 11050
box -29 -23 29 23
use L1M1_PR  L1M1_PR_852
timestamp 1655484843
transform 1 0 15410 0 1 13158
box -29 -23 29 23
use L1M1_PR  L1M1_PR_853
timestamp 1655484843
transform 1 0 14766 0 1 12138
box -29 -23 29 23
use L1M1_PR  L1M1_PR_854
timestamp 1655484843
transform 1 0 17066 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_855
timestamp 1655484843
transform 1 0 15042 0 1 12342
box -29 -23 29 23
use L1M1_PR  L1M1_PR_856
timestamp 1655484843
transform 1 0 16698 0 1 15334
box -29 -23 29 23
use L1M1_PR  L1M1_PR_857
timestamp 1655484843
transform 1 0 16330 0 1 15402
box -29 -23 29 23
use L1M1_PR  L1M1_PR_858
timestamp 1655484843
transform 1 0 16882 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_859
timestamp 1655484843
transform 1 0 15870 0 1 14518
box -29 -23 29 23
use L1M1_PR  L1M1_PR_860
timestamp 1655484843
transform 1 0 15778 0 1 15606
box -29 -23 29 23
use L1M1_PR  L1M1_PR_861
timestamp 1655484843
transform 1 0 14490 0 1 14246
box -29 -23 29 23
use L1M1_PR  L1M1_PR_862
timestamp 1655484843
transform 1 0 15410 0 1 17510
box -29 -23 29 23
use L1M1_PR  L1M1_PR_863
timestamp 1655484843
transform 1 0 14766 0 1 17578
box -29 -23 29 23
use L1M1_PR  L1M1_PR_864
timestamp 1655484843
transform 1 0 15410 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_865
timestamp 1655484843
transform 1 0 14030 0 1 16830
box -29 -23 29 23
use L1M1_PR  L1M1_PR_866
timestamp 1655484843
transform 1 0 16974 0 1 16422
box -29 -23 29 23
use L1M1_PR  L1M1_PR_867
timestamp 1655484843
transform 1 0 15870 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_868
timestamp 1655484843
transform 1 0 15962 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_869
timestamp 1655484843
transform 1 0 15778 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_870
timestamp 1655484843
transform 1 0 11086 0 1 20298
box -29 -23 29 23
use L1M1_PR  L1M1_PR_871
timestamp 1655484843
transform 1 0 10534 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_872
timestamp 1655484843
transform 1 0 10442 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_873
timestamp 1655484843
transform 1 0 10350 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_874
timestamp 1655484843
transform 1 0 9246 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_875
timestamp 1655484843
transform 1 0 8878 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_876
timestamp 1655484843
transform 1 0 8050 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_877
timestamp 1655484843
transform 1 0 7590 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_878
timestamp 1655484843
transform 1 0 6854 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_879
timestamp 1655484843
transform 1 0 6762 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_880
timestamp 1655484843
transform 1 0 6578 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_881
timestamp 1655484843
transform 1 0 22310 0 1 15198
box -29 -23 29 23
use L1M1_PR  L1M1_PR_882
timestamp 1655484843
transform 1 0 22310 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_883
timestamp 1655484843
transform 1 0 22218 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_884
timestamp 1655484843
transform 1 0 22218 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_885
timestamp 1655484843
transform 1 0 22126 0 1 18530
box -29 -23 29 23
use L1M1_PR  L1M1_PR_886
timestamp 1655484843
transform 1 0 22126 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_887
timestamp 1655484843
transform 1 0 21850 0 1 9826
box -29 -23 29 23
use L1M1_PR  L1M1_PR_888
timestamp 1655484843
transform 1 0 21758 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_889
timestamp 1655484843
transform 1 0 21758 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_890
timestamp 1655484843
transform 1 0 20930 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_891
timestamp 1655484843
transform 1 0 20194 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_892
timestamp 1655484843
transform 1 0 18998 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_893
timestamp 1655484843
transform 1 0 18078 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_894
timestamp 1655484843
transform 1 0 17802 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_895
timestamp 1655484843
transform 1 0 16606 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_896
timestamp 1655484843
transform 1 0 16146 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_897
timestamp 1655484843
transform 1 0 15410 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_898
timestamp 1655484843
transform 1 0 15318 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_899
timestamp 1655484843
transform 1 0 14030 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_900
timestamp 1655484843
transform 1 0 13846 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_901
timestamp 1655484843
transform 1 0 13202 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_902
timestamp 1655484843
transform 1 0 13110 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_903
timestamp 1655484843
transform 1 0 13110 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_904
timestamp 1655484843
transform 1 0 12926 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_905
timestamp 1655484843
transform 1 0 12834 0 1 8670
box -29 -23 29 23
use L1M1_PR  L1M1_PR_906
timestamp 1655484843
transform 1 0 12558 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_907
timestamp 1655484843
transform 1 0 12205 0 1 20026
box -29 -23 29 23
use L1M1_PR  L1M1_PR_908
timestamp 1655484843
transform 1 0 11638 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_909
timestamp 1655484843
transform 1 0 11546 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_910
timestamp 1655484843
transform 1 0 19734 0 1 21726
box -29 -23 29 23
use L1M1_PR  L1M1_PR_911
timestamp 1655484843
transform 1 0 19550 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_912
timestamp 1655484843
transform 1 0 19090 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_913
timestamp 1655484843
transform 1 0 19075 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_914
timestamp 1655484843
transform 1 0 16422 0 1 21250
box -29 -23 29 23
use L1M1_PR  L1M1_PR_915
timestamp 1655484843
transform 1 0 15134 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_916
timestamp 1655484843
transform 1 0 13018 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_917
timestamp 1655484843
transform 1 0 13018 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_918
timestamp 1655484843
transform 1 0 11914 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_919
timestamp 1655484843
transform 1 0 11638 0 1 17918
box -29 -23 29 23
use L1M1_PR  L1M1_PR_920
timestamp 1655484843
transform 1 0 11454 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_921
timestamp 1655484843
transform 1 0 10718 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_922
timestamp 1655484843
transform 1 0 10258 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_923
timestamp 1655484843
transform 1 0 10166 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_924
timestamp 1655484843
transform 1 0 10074 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_925
timestamp 1655484843
transform 1 0 9982 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_926
timestamp 1655484843
transform 1 0 9798 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_927
timestamp 1655484843
transform 1 0 9430 0 1 16286
box -29 -23 29 23
use L1M1_PR  L1M1_PR_928
timestamp 1655484843
transform 1 0 9154 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_929
timestamp 1655484843
transform 1 0 9062 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_930
timestamp 1655484843
transform 1 0 11178 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_931
timestamp 1655484843
transform 1 0 10902 0 1 16898
box -29 -23 29 23
use L1M1_PR  L1M1_PR_932
timestamp 1655484843
transform 1 0 10810 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_933
timestamp 1655484843
transform 1 0 10718 0 1 18462
box -29 -23 29 23
use L1M1_PR  L1M1_PR_934
timestamp 1655484843
transform 1 0 10534 0 1 20162
box -29 -23 29 23
use L1M1_PR  L1M1_PR_935
timestamp 1655484843
transform 1 0 10350 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_936
timestamp 1655484843
transform 1 0 10258 0 1 6970
box -29 -23 29 23
use L1M1_PR  L1M1_PR_937
timestamp 1655484843
transform 1 0 9522 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_938
timestamp 1655484843
transform 1 0 8602 0 1 15266
box -29 -23 29 23
use L1M1_PR  L1M1_PR_939
timestamp 1655484843
transform 1 0 8234 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_940
timestamp 1655484843
transform 1 0 7866 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_941
timestamp 1655484843
transform 1 0 7498 0 1 11934
box -29 -23 29 23
use L1M1_PR  L1M1_PR_942
timestamp 1655484843
transform 1 0 7406 0 1 16354
box -29 -23 29 23
use L1M1_PR  L1M1_PR_943
timestamp 1655484843
transform 1 0 7314 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_944
timestamp 1655484843
transform 1 0 7314 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_945
timestamp 1655484843
transform 1 0 7314 0 1 10846
box -29 -23 29 23
use L1M1_PR  L1M1_PR_946
timestamp 1655484843
transform 1 0 7222 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_947
timestamp 1655484843
transform 1 0 7222 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_948
timestamp 1655484843
transform 1 0 6946 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_949
timestamp 1655484843
transform 1 0 6946 0 1 14722
box -29 -23 29 23
use L1M1_PR  L1M1_PR_950
timestamp 1655484843
transform 1 0 6946 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_951
timestamp 1655484843
transform 1 0 6946 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_952
timestamp 1655484843
transform 1 0 6946 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_953
timestamp 1655484843
transform 1 0 6946 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_954
timestamp 1655484843
transform 1 0 6854 0 1 20162
box -29 -23 29 23
use L1M1_PR  L1M1_PR_955
timestamp 1655484843
transform 1 0 21390 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_956
timestamp 1655484843
transform 1 0 19918 0 1 7514
box -29 -23 29 23
use L1M1_PR  L1M1_PR_957
timestamp 1655484843
transform 1 0 19274 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_958
timestamp 1655484843
transform 1 0 18814 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_959
timestamp 1655484843
transform 1 0 18814 0 1 10370
box -29 -23 29 23
use L1M1_PR  L1M1_PR_960
timestamp 1655484843
transform 1 0 16238 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_961
timestamp 1655484843
transform 1 0 14950 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_962
timestamp 1655484843
transform 1 0 13662 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_963
timestamp 1655484843
transform 1 0 13294 0 1 12546
box -29 -23 29 23
use L1M1_PR  L1M1_PR_964
timestamp 1655484843
transform 1 0 12926 0 1 9214
box -29 -23 29 23
use L1M1_PR  L1M1_PR_965
timestamp 1655484843
transform 1 0 12834 0 1 13022
box -29 -23 29 23
use L1M1_PR  L1M1_PR_966
timestamp 1655484843
transform 1 0 12742 0 1 14110
box -29 -23 29 23
use L1M1_PR  L1M1_PR_967
timestamp 1655484843
transform 1 0 12466 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_968
timestamp 1655484843
transform 1 0 12374 0 1 9758
box -29 -23 29 23
use L1M1_PR  L1M1_PR_969
timestamp 1655484843
transform 1 0 12374 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_970
timestamp 1655484843
transform 1 0 12374 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_971
timestamp 1655484843
transform 1 0 12190 0 1 14110
box -29 -23 29 23
use L1M1_PR  L1M1_PR_972
timestamp 1655484843
transform 1 0 12098 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_973
timestamp 1655484843
transform 1 0 12098 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_974
timestamp 1655484843
transform 1 0 12098 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_975
timestamp 1655484843
transform 1 0 11178 0 1 7582
box -29 -23 29 23
use L1M1_PR  L1M1_PR_976
timestamp 1655484843
transform 1 0 11086 0 1 8194
box -29 -23 29 23
use L1M1_PR  L1M1_PR_977
timestamp 1655484843
transform 1 0 9338 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_978
timestamp 1655484843
transform 1 0 9338 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_979
timestamp 1655484843
transform 1 0 9246 0 1 10302
box -29 -23 29 23
use L1M1_PR  L1M1_PR_980
timestamp 1655484843
transform 1 0 22954 0 1 20162
box -29 -23 29 23
use L1M1_PR  L1M1_PR_981
timestamp 1655484843
transform 1 0 22862 0 1 19006
box -29 -23 29 23
use L1M1_PR  L1M1_PR_982
timestamp 1655484843
transform 1 0 22770 0 1 17986
box -29 -23 29 23
use L1M1_PR  L1M1_PR_983
timestamp 1655484843
transform 1 0 22770 0 1 15810
box -29 -23 29 23
use L1M1_PR  L1M1_PR_984
timestamp 1655484843
transform 1 0 22770 0 1 14722
box -29 -23 29 23
use L1M1_PR  L1M1_PR_985
timestamp 1655484843
transform 1 0 22770 0 1 13634
box -29 -23 29 23
use L1M1_PR  L1M1_PR_986
timestamp 1655484843
transform 1 0 22770 0 1 11458
box -29 -23 29 23
use L1M1_PR  L1M1_PR_987
timestamp 1655484843
transform 1 0 22494 0 1 19550
box -29 -23 29 23
use L1M1_PR  L1M1_PR_988
timestamp 1655484843
transform 1 0 22494 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_989
timestamp 1655484843
transform 1 0 21390 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_990
timestamp 1655484843
transform 1 0 21114 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_991
timestamp 1655484843
transform 1 0 20194 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_992
timestamp 1655484843
transform 1 0 20102 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_993
timestamp 1655484843
transform 1 0 19826 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_994
timestamp 1655484843
transform 1 0 19182 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_995
timestamp 1655484843
transform 1 0 16238 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_996
timestamp 1655484843
transform 1 0 15962 0 1 20638
box -29 -23 29 23
use L1M1_PR  L1M1_PR_997
timestamp 1655484843
transform 1 0 15778 0 1 21182
box -29 -23 29 23
use L1M1_PR  L1M1_PR_998
timestamp 1655484843
transform 1 0 15594 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_999
timestamp 1655484843
transform 1 0 12834 0 1 19618
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1000
timestamp 1655484843
transform 1 0 12466 0 1 20094
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1001
timestamp 1655484843
transform 1 0 12374 0 1 20706
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1002
timestamp 1655484843
transform 1 0 20194 0 1 12478
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1003
timestamp 1655484843
transform 1 0 18906 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1004
timestamp 1655484843
transform 1 0 18630 0 1 6494
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1005
timestamp 1655484843
transform 1 0 9338 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1006
timestamp 1655484843
transform 1 0 18354 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1007
timestamp 1655484843
transform 1 0 14950 0 1 8058
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1008
timestamp 1655484843
transform 1 0 14306 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1009
timestamp 1655484843
transform 1 0 14306 0 1 6018
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1010
timestamp 1655484843
transform 1 0 17986 0 1 12070
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1011
timestamp 1655484843
transform 1 0 17250 0 1 12342
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1012
timestamp 1655484843
transform 1 0 13110 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1013
timestamp 1655484843
transform 1 0 10810 0 1 14314
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1014
timestamp 1655484843
transform 1 0 10810 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1015
timestamp 1655484843
transform 1 0 18630 0 1 18870
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1016
timestamp 1655484843
transform 1 0 17802 0 1 18598
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1017
timestamp 1655484843
transform 1 0 21482 0 1 18326
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1018
timestamp 1655484843
transform 1 0 19642 0 1 17442
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1019
timestamp 1655484843
transform 1 0 21206 0 1 18122
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1020
timestamp 1655484843
transform 1 0 21206 0 1 17782
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1021
timestamp 1655484843
transform 1 0 20838 0 1 16762
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1022
timestamp 1655484843
transform 1 0 19274 0 1 17306
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1023
timestamp 1655484843
transform 1 0 19090 0 1 15742
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1024
timestamp 1655484843
transform 1 0 21482 0 1 16490
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1025
timestamp 1655484843
transform 1 0 21482 0 1 16150
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1026
timestamp 1655484843
transform 1 0 20562 0 1 14654
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1027
timestamp 1655484843
transform 1 0 20102 0 1 13974
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1028
timestamp 1655484843
transform 1 0 19366 0 1 14178
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1029
timestamp 1655484843
transform 1 0 20562 0 1 13498
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1030
timestamp 1655484843
transform 1 0 20102 0 1 13226
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1031
timestamp 1655484843
transform 1 0 21850 0 1 13090
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1032
timestamp 1655484843
transform 1 0 20102 0 1 11798
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1033
timestamp 1655484843
transform 1 0 20562 0 1 9146
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1034
timestamp 1655484843
transform 1 0 20194 0 1 9078
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1035
timestamp 1655484843
transform 1 0 22770 0 1 8330
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1036
timestamp 1655484843
transform 1 0 20562 0 1 10234
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1037
timestamp 1655484843
transform 1 0 20746 0 1 11322
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1038
timestamp 1655484843
transform 1 0 20102 0 1 10710
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1039
timestamp 1655484843
transform 1 0 22770 0 1 10166
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1040
timestamp 1655484843
transform 1 0 20562 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1041
timestamp 1655484843
transform 1 0 5934 0 1 7106
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1042
timestamp 1655484843
transform 1 0 5750 0 1 7446
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1043
timestamp 1655484843
transform 1 0 5566 0 1 7038
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1044
timestamp 1655484843
transform 1 0 13478 0 1 7990
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1045
timestamp 1655484843
transform 1 0 12635 0 1 6562
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1046
timestamp 1655484843
transform 1 0 10917 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1047
timestamp 1655484843
transform 1 0 8050 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1048
timestamp 1655484843
transform 1 0 7498 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1049
timestamp 1655484843
transform 1 0 6854 0 1 10914
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1050
timestamp 1655484843
transform 1 0 6762 0 1 5950
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1051
timestamp 1655484843
transform 1 0 6670 0 1 11390
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1052
timestamp 1655484843
transform 1 0 6670 0 1 9282
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1053
timestamp 1655484843
transform 1 0 6670 0 1 7650
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1054
timestamp 1655484843
transform 1 0 6578 0 1 8126
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1055
timestamp 1655484843
transform 1 0 6486 0 1 13566
box -29 -23 29 23
use L1M1_PR  L1M1_PR_1056
timestamp 1655484843
transform 1 0 14122 0 1 5950
box -29 -23 29 23
use M1M2_PR  M1M2_PR_0
timestamp 1655484843
transform 1 0 18078 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_1
timestamp 1655484843
transform 1 0 18078 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_2
timestamp 1655484843
transform 1 0 14950 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_3
timestamp 1655484843
transform 1 0 14950 0 1 9894
box -32 -32 32 32
use M1M2_PR  M1M2_PR_4
timestamp 1655484843
transform 1 0 14490 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_5
timestamp 1655484843
transform 1 0 14490 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_6
timestamp 1655484843
transform 1 0 16146 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_7
timestamp 1655484843
transform 1 0 16146 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_8
timestamp 1655484843
transform 1 0 16054 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_9
timestamp 1655484843
transform 1 0 17526 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_10
timestamp 1655484843
transform 1 0 16790 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_11
timestamp 1655484843
transform 1 0 14398 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_12
timestamp 1655484843
transform 1 0 14398 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_13
timestamp 1655484843
transform 1 0 17158 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_14
timestamp 1655484843
transform 1 0 17158 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_15
timestamp 1655484843
transform 1 0 13294 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_16
timestamp 1655484843
transform 1 0 13294 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_17
timestamp 1655484843
transform 1 0 16330 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_18
timestamp 1655484843
transform 1 0 16330 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_19
timestamp 1655484843
transform 1 0 17618 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_20
timestamp 1655484843
transform 1 0 17434 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_21
timestamp 1655484843
transform 1 0 19734 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_22
timestamp 1655484843
transform 1 0 19734 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_23
timestamp 1655484843
transform 1 0 20746 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_24
timestamp 1655484843
transform 1 0 20746 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_25
timestamp 1655484843
transform 1 0 20010 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_26
timestamp 1655484843
transform 1 0 20010 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_27
timestamp 1655484843
transform 1 0 19918 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_28
timestamp 1655484843
transform 1 0 19826 0 1 15130
box -32 -32 32 32
use M1M2_PR  M1M2_PR_29
timestamp 1655484843
transform 1 0 20194 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_30
timestamp 1655484843
transform 1 0 20194 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_31
timestamp 1655484843
transform 1 0 21758 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_32
timestamp 1655484843
transform 1 0 21758 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_33
timestamp 1655484843
transform 1 0 20010 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_34
timestamp 1655484843
transform 1 0 20010 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_35
timestamp 1655484843
transform 1 0 20654 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_36
timestamp 1655484843
transform 1 0 20654 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_37
timestamp 1655484843
transform 1 0 20838 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_38
timestamp 1655484843
transform 1 0 20838 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_39
timestamp 1655484843
transform 1 0 14030 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_40
timestamp 1655484843
transform 1 0 14030 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_41
timestamp 1655484843
transform 1 0 13294 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_42
timestamp 1655484843
transform 1 0 13294 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_43
timestamp 1655484843
transform 1 0 15042 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_44
timestamp 1655484843
transform 1 0 14766 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_45
timestamp 1655484843
transform 1 0 20930 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_46
timestamp 1655484843
transform 1 0 20654 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_47
timestamp 1655484843
transform 1 0 20470 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_48
timestamp 1655484843
transform 1 0 20470 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_49
timestamp 1655484843
transform 1 0 20470 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_50
timestamp 1655484843
transform 1 0 20378 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_51
timestamp 1655484843
transform 1 0 20378 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_52
timestamp 1655484843
transform 1 0 20378 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_53
timestamp 1655484843
transform 1 0 19550 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_54
timestamp 1655484843
transform 1 0 19090 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_55
timestamp 1655484843
transform 1 0 19090 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_56
timestamp 1655484843
transform 1 0 17986 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_57
timestamp 1655484843
transform 1 0 17894 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_58
timestamp 1655484843
transform 1 0 17894 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_59
timestamp 1655484843
transform 1 0 17158 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_60
timestamp 1655484843
transform 1 0 17158 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_61
timestamp 1655484843
transform 1 0 16882 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_62
timestamp 1655484843
transform 1 0 16882 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_63
timestamp 1655484843
transform 1 0 16882 0 1 15878
box -32 -32 32 32
use M1M2_PR  M1M2_PR_64
timestamp 1655484843
transform 1 0 16882 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_65
timestamp 1655484843
transform 1 0 16790 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_66
timestamp 1655484843
transform 1 0 15870 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_67
timestamp 1655484843
transform 1 0 15870 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_68
timestamp 1655484843
transform 1 0 15870 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_69
timestamp 1655484843
transform 1 0 15870 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_70
timestamp 1655484843
transform 1 0 15778 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_71
timestamp 1655484843
transform 1 0 15318 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_72
timestamp 1655484843
transform 1 0 14582 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_73
timestamp 1655484843
transform 1 0 14306 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_74
timestamp 1655484843
transform 1 0 14214 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_75
timestamp 1655484843
transform 1 0 14122 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_76
timestamp 1655484843
transform 1 0 14122 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_77
timestamp 1655484843
transform 1 0 13294 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_78
timestamp 1655484843
transform 1 0 13294 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_79
timestamp 1655484843
transform 1 0 22034 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_80
timestamp 1655484843
transform 1 0 21298 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_81
timestamp 1655484843
transform 1 0 21206 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_82
timestamp 1655484843
transform 1 0 21206 0 1 9078
box -32 -32 32 32
use M1M2_PR  M1M2_PR_83
timestamp 1655484843
transform 1 0 21206 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_84
timestamp 1655484843
transform 1 0 20746 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_85
timestamp 1655484843
transform 1 0 20378 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_86
timestamp 1655484843
transform 1 0 20194 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_87
timestamp 1655484843
transform 1 0 20194 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_88
timestamp 1655484843
transform 1 0 20102 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_89
timestamp 1655484843
transform 1 0 20102 0 1 15810
box -32 -32 32 32
use M1M2_PR  M1M2_PR_90
timestamp 1655484843
transform 1 0 18262 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_91
timestamp 1655484843
transform 1 0 18262 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_92
timestamp 1655484843
transform 1 0 18262 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_93
timestamp 1655484843
transform 1 0 16790 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_94
timestamp 1655484843
transform 1 0 16790 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_95
timestamp 1655484843
transform 1 0 16790 0 1 8262
box -32 -32 32 32
use M1M2_PR  M1M2_PR_96
timestamp 1655484843
transform 1 0 16698 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_97
timestamp 1655484843
transform 1 0 15778 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_98
timestamp 1655484843
transform 1 0 15686 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_99
timestamp 1655484843
transform 1 0 15686 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_100
timestamp 1655484843
transform 1 0 15594 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_101
timestamp 1655484843
transform 1 0 15594 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_102
timestamp 1655484843
transform 1 0 15594 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_103
timestamp 1655484843
transform 1 0 15594 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_104
timestamp 1655484843
transform 1 0 15594 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_105
timestamp 1655484843
transform 1 0 15594 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_106
timestamp 1655484843
transform 1 0 15594 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_107
timestamp 1655484843
transform 1 0 15502 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_108
timestamp 1655484843
transform 1 0 15318 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_109
timestamp 1655484843
transform 1 0 15318 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_110
timestamp 1655484843
transform 1 0 14490 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_111
timestamp 1655484843
transform 1 0 14490 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_112
timestamp 1655484843
transform 1 0 13294 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_113
timestamp 1655484843
transform 1 0 13294 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_114
timestamp 1655484843
transform 1 0 13294 0 1 7718
box -32 -32 32 32
use M1M2_PR  M1M2_PR_115
timestamp 1655484843
transform 1 0 16974 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_116
timestamp 1655484843
transform 1 0 16974 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_117
timestamp 1655484843
transform 1 0 16974 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_118
timestamp 1655484843
transform 1 0 16974 0 1 8806
box -32 -32 32 32
use M1M2_PR  M1M2_PR_119
timestamp 1655484843
transform 1 0 18998 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_120
timestamp 1655484843
transform 1 0 18998 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_121
timestamp 1655484843
transform 1 0 19182 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_122
timestamp 1655484843
transform 1 0 19090 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_123
timestamp 1655484843
transform 1 0 20286 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_124
timestamp 1655484843
transform 1 0 20194 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_125
timestamp 1655484843
transform 1 0 20194 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_126
timestamp 1655484843
transform 1 0 20194 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_127
timestamp 1655484843
transform 1 0 20194 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_128
timestamp 1655484843
transform 1 0 20102 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_129
timestamp 1655484843
transform 1 0 18998 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_130
timestamp 1655484843
transform 1 0 18998 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_131
timestamp 1655484843
transform 1 0 21114 0 1 15334
box -32 -32 32 32
use M1M2_PR  M1M2_PR_132
timestamp 1655484843
transform 1 0 18630 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_133
timestamp 1655484843
transform 1 0 18630 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_134
timestamp 1655484843
transform 1 0 21022 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_135
timestamp 1655484843
transform 1 0 21022 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_136
timestamp 1655484843
transform 1 0 18630 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_137
timestamp 1655484843
transform 1 0 18630 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_138
timestamp 1655484843
transform 1 0 18446 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_139
timestamp 1655484843
transform 1 0 18446 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_140
timestamp 1655484843
transform 1 0 16514 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_141
timestamp 1655484843
transform 1 0 16514 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_142
timestamp 1655484843
transform 1 0 17802 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_143
timestamp 1655484843
transform 1 0 17802 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_144
timestamp 1655484843
transform 1 0 15410 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_145
timestamp 1655484843
transform 1 0 14858 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_146
timestamp 1655484843
transform 1 0 14766 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_147
timestamp 1655484843
transform 1 0 18630 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_148
timestamp 1655484843
transform 1 0 18630 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_149
timestamp 1655484843
transform 1 0 15226 0 1 14586
box -32 -32 32 32
use M1M2_PR  M1M2_PR_150
timestamp 1655484843
transform 1 0 15226 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_151
timestamp 1655484843
transform 1 0 17158 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_152
timestamp 1655484843
transform 1 0 17158 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_153
timestamp 1655484843
transform 1 0 17342 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_154
timestamp 1655484843
transform 1 0 17342 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_155
timestamp 1655484843
transform 1 0 17342 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_156
timestamp 1655484843
transform 1 0 17250 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_157
timestamp 1655484843
transform 1 0 15686 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_158
timestamp 1655484843
transform 1 0 15686 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_159
timestamp 1655484843
transform 1 0 17342 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_160
timestamp 1655484843
transform 1 0 17342 0 1 10234
box -32 -32 32 32
use M1M2_PR  M1M2_PR_161
timestamp 1655484843
transform 1 0 14582 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_162
timestamp 1655484843
transform 1 0 14582 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_163
timestamp 1655484843
transform 1 0 15962 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_164
timestamp 1655484843
transform 1 0 15962 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_165
timestamp 1655484843
transform 1 0 16146 0 1 10234
box -32 -32 32 32
use M1M2_PR  M1M2_PR_166
timestamp 1655484843
transform 1 0 16146 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_167
timestamp 1655484843
transform 1 0 17710 0 1 10438
box -32 -32 32 32
use M1M2_PR  M1M2_PR_168
timestamp 1655484843
transform 1 0 17710 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_169
timestamp 1655484843
transform 1 0 17618 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_170
timestamp 1655484843
transform 1 0 17618 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_171
timestamp 1655484843
transform 1 0 16698 0 1 15810
box -32 -32 32 32
use M1M2_PR  M1M2_PR_172
timestamp 1655484843
transform 1 0 16698 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_173
timestamp 1655484843
transform 1 0 16606 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_174
timestamp 1655484843
transform 1 0 16606 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_175
timestamp 1655484843
transform 1 0 18814 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_176
timestamp 1655484843
transform 1 0 18814 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_177
timestamp 1655484843
transform 1 0 18814 0 1 12546
box -32 -32 32 32
use M1M2_PR  M1M2_PR_178
timestamp 1655484843
transform 1 0 17526 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_179
timestamp 1655484843
transform 1 0 15502 0 1 14042
box -32 -32 32 32
use M1M2_PR  M1M2_PR_180
timestamp 1655484843
transform 1 0 15502 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_181
timestamp 1655484843
transform 1 0 14030 0 1 11458
box -32 -32 32 32
use M1M2_PR  M1M2_PR_182
timestamp 1655484843
transform 1 0 19366 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_183
timestamp 1655484843
transform 1 0 18538 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_184
timestamp 1655484843
transform 1 0 18538 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_185
timestamp 1655484843
transform 1 0 18538 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_186
timestamp 1655484843
transform 1 0 18446 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_187
timestamp 1655484843
transform 1 0 16882 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_188
timestamp 1655484843
transform 1 0 16882 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_189
timestamp 1655484843
transform 1 0 16882 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_190
timestamp 1655484843
transform 1 0 21482 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_191
timestamp 1655484843
transform 1 0 21482 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_192
timestamp 1655484843
transform 1 0 18538 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_193
timestamp 1655484843
transform 1 0 18170 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_194
timestamp 1655484843
transform 1 0 17986 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_195
timestamp 1655484843
transform 1 0 17986 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_196
timestamp 1655484843
transform 1 0 17986 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_197
timestamp 1655484843
transform 1 0 16238 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_198
timestamp 1655484843
transform 1 0 15962 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_199
timestamp 1655484843
transform 1 0 18354 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_200
timestamp 1655484843
transform 1 0 18262 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_201
timestamp 1655484843
transform 1 0 17802 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_202
timestamp 1655484843
transform 1 0 17802 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_203
timestamp 1655484843
transform 1 0 6854 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_204
timestamp 1655484843
transform 1 0 6854 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_205
timestamp 1655484843
transform 1 0 6578 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_206
timestamp 1655484843
transform 1 0 6578 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_207
timestamp 1655484843
transform 1 0 9062 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_208
timestamp 1655484843
transform 1 0 9062 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_209
timestamp 1655484843
transform 1 0 9982 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_210
timestamp 1655484843
transform 1 0 9982 0 1 17986
box -32 -32 32 32
use M1M2_PR  M1M2_PR_211
timestamp 1655484843
transform 1 0 6210 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_212
timestamp 1655484843
transform 1 0 6210 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_213
timestamp 1655484843
transform 1 0 9982 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_214
timestamp 1655484843
transform 1 0 9982 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_215
timestamp 1655484843
transform 1 0 9982 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_216
timestamp 1655484843
transform 1 0 9982 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_217
timestamp 1655484843
transform 1 0 8970 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_218
timestamp 1655484843
transform 1 0 8970 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_219
timestamp 1655484843
transform 1 0 8970 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_220
timestamp 1655484843
transform 1 0 10166 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_221
timestamp 1655484843
transform 1 0 10166 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_222
timestamp 1655484843
transform 1 0 9798 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_223
timestamp 1655484843
transform 1 0 9798 0 1 17510
box -32 -32 32 32
use M1M2_PR  M1M2_PR_224
timestamp 1655484843
transform 1 0 8786 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_225
timestamp 1655484843
transform 1 0 8694 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_226
timestamp 1655484843
transform 1 0 9154 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_227
timestamp 1655484843
transform 1 0 9154 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_228
timestamp 1655484843
transform 1 0 9154 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_229
timestamp 1655484843
transform 1 0 8786 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_230
timestamp 1655484843
transform 1 0 8786 0 1 19686
box -32 -32 32 32
use M1M2_PR  M1M2_PR_231
timestamp 1655484843
transform 1 0 6762 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_232
timestamp 1655484843
transform 1 0 6762 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_233
timestamp 1655484843
transform 1 0 7958 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_234
timestamp 1655484843
transform 1 0 7958 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_235
timestamp 1655484843
transform 1 0 8878 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_236
timestamp 1655484843
transform 1 0 8878 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_237
timestamp 1655484843
transform 1 0 8878 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_238
timestamp 1655484843
transform 1 0 8878 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_239
timestamp 1655484843
transform 1 0 9062 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_240
timestamp 1655484843
transform 1 0 9062 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_241
timestamp 1655484843
transform 1 0 7958 0 1 19482
box -32 -32 32 32
use M1M2_PR  M1M2_PR_242
timestamp 1655484843
transform 1 0 7958 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_243
timestamp 1655484843
transform 1 0 7498 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_244
timestamp 1655484843
transform 1 0 7498 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_245
timestamp 1655484843
transform 1 0 6946 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_246
timestamp 1655484843
transform 1 0 6946 0 1 19210
box -32 -32 32 32
use M1M2_PR  M1M2_PR_247
timestamp 1655484843
transform 1 0 7590 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_248
timestamp 1655484843
transform 1 0 7590 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_249
timestamp 1655484843
transform 1 0 7498 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_250
timestamp 1655484843
transform 1 0 7130 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_251
timestamp 1655484843
transform 1 0 10350 0 1 17238
box -32 -32 32 32
use M1M2_PR  M1M2_PR_252
timestamp 1655484843
transform 1 0 10350 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_253
timestamp 1655484843
transform 1 0 10258 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_254
timestamp 1655484843
transform 1 0 10258 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_255
timestamp 1655484843
transform 1 0 10917 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_256
timestamp 1655484843
transform 1 0 10534 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_257
timestamp 1655484843
transform 1 0 19182 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_258
timestamp 1655484843
transform 1 0 17158 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_259
timestamp 1655484843
transform 1 0 16330 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_260
timestamp 1655484843
transform 1 0 16054 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_261
timestamp 1655484843
transform 1 0 15962 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_262
timestamp 1655484843
transform 1 0 12834 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_263
timestamp 1655484843
transform 1 0 12834 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_264
timestamp 1655484843
transform 1 0 11178 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_265
timestamp 1655484843
transform 1 0 11178 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_266
timestamp 1655484843
transform 1 0 17434 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_267
timestamp 1655484843
transform 1 0 17434 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_268
timestamp 1655484843
transform 1 0 17066 0 1 12886
box -32 -32 32 32
use M1M2_PR  M1M2_PR_269
timestamp 1655484843
transform 1 0 17066 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_270
timestamp 1655484843
transform 1 0 13386 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_271
timestamp 1655484843
transform 1 0 13294 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_272
timestamp 1655484843
transform 1 0 13202 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_273
timestamp 1655484843
transform 1 0 9062 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_274
timestamp 1655484843
transform 1 0 9062 0 1 15878
box -32 -32 32 32
use M1M2_PR  M1M2_PR_275
timestamp 1655484843
transform 1 0 8786 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_276
timestamp 1655484843
transform 1 0 8786 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_277
timestamp 1655484843
transform 1 0 8878 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_278
timestamp 1655484843
transform 1 0 8878 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_279
timestamp 1655484843
transform 1 0 10350 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_280
timestamp 1655484843
transform 1 0 10350 0 1 17374
box -32 -32 32 32
use M1M2_PR  M1M2_PR_281
timestamp 1655484843
transform 1 0 10350 0 1 19482
box -32 -32 32 32
use M1M2_PR  M1M2_PR_282
timestamp 1655484843
transform 1 0 10350 0 1 19210
box -32 -32 32 32
use M1M2_PR  M1M2_PR_283
timestamp 1655484843
transform 1 0 10166 0 1 21658
box -32 -32 32 32
use M1M2_PR  M1M2_PR_284
timestamp 1655484843
transform 1 0 10166 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_285
timestamp 1655484843
transform 1 0 18722 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_286
timestamp 1655484843
transform 1 0 16054 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_287
timestamp 1655484843
transform 1 0 16054 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_288
timestamp 1655484843
transform 1 0 15502 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_289
timestamp 1655484843
transform 1 0 13478 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_290
timestamp 1655484843
transform 1 0 13478 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_291
timestamp 1655484843
transform 1 0 13478 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_292
timestamp 1655484843
transform 1 0 13478 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_293
timestamp 1655484843
transform 1 0 14490 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_294
timestamp 1655484843
transform 1 0 14490 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_295
timestamp 1655484843
transform 1 0 14490 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_296
timestamp 1655484843
transform 1 0 14490 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_297
timestamp 1655484843
transform 1 0 14490 0 1 15130
box -32 -32 32 32
use M1M2_PR  M1M2_PR_298
timestamp 1655484843
transform 1 0 14490 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_299
timestamp 1655484843
transform 1 0 21482 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_300
timestamp 1655484843
transform 1 0 21482 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_301
timestamp 1655484843
transform 1 0 21482 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_302
timestamp 1655484843
transform 1 0 21482 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_303
timestamp 1655484843
transform 1 0 21482 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_304
timestamp 1655484843
transform 1 0 21482 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_305
timestamp 1655484843
transform 1 0 18262 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_306
timestamp 1655484843
transform 1 0 18078 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_307
timestamp 1655484843
transform 1 0 19918 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_308
timestamp 1655484843
transform 1 0 19918 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_309
timestamp 1655484843
transform 1 0 17710 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_310
timestamp 1655484843
transform 1 0 17710 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_311
timestamp 1655484843
transform 1 0 17710 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_312
timestamp 1655484843
transform 1 0 17342 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_313
timestamp 1655484843
transform 1 0 17342 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_314
timestamp 1655484843
transform 1 0 19826 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_315
timestamp 1655484843
transform 1 0 19826 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_316
timestamp 1655484843
transform 1 0 21850 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_317
timestamp 1655484843
transform 1 0 21850 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_318
timestamp 1655484843
transform 1 0 21850 0 1 9078
box -32 -32 32 32
use M1M2_PR  M1M2_PR_319
timestamp 1655484843
transform 1 0 21850 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_320
timestamp 1655484843
transform 1 0 23506 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_321
timestamp 1655484843
transform 1 0 23414 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_322
timestamp 1655484843
transform 1 0 20102 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_323
timestamp 1655484843
transform 1 0 20102 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_324
timestamp 1655484843
transform 1 0 21666 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_325
timestamp 1655484843
transform 1 0 21666 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_326
timestamp 1655484843
transform 1 0 22034 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_327
timestamp 1655484843
transform 1 0 22034 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_328
timestamp 1655484843
transform 1 0 22218 0 1 21318
box -32 -32 32 32
use M1M2_PR  M1M2_PR_329
timestamp 1655484843
transform 1 0 22218 0 1 19210
box -32 -32 32 32
use M1M2_PR  M1M2_PR_330
timestamp 1655484843
transform 1 0 19274 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_331
timestamp 1655484843
transform 1 0 19274 0 1 19142
box -32 -32 32 32
use M1M2_PR  M1M2_PR_332
timestamp 1655484843
transform 1 0 17618 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_333
timestamp 1655484843
transform 1 0 17618 0 1 19210
box -32 -32 32 32
use M1M2_PR  M1M2_PR_334
timestamp 1655484843
transform 1 0 14858 0 1 19142
box -32 -32 32 32
use M1M2_PR  M1M2_PR_335
timestamp 1655484843
transform 1 0 14858 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_336
timestamp 1655484843
transform 1 0 13018 0 1 19142
box -32 -32 32 32
use M1M2_PR  M1M2_PR_337
timestamp 1655484843
transform 1 0 13018 0 1 18394
box -32 -32 32 32
use M1M2_PR  M1M2_PR_338
timestamp 1655484843
transform 1 0 12098 0 1 19142
box -32 -32 32 32
use M1M2_PR  M1M2_PR_339
timestamp 1655484843
transform 1 0 12098 0 1 17986
box -32 -32 32 32
use M1M2_PR  M1M2_PR_340
timestamp 1655484843
transform 1 0 12006 0 1 18054
box -32 -32 32 32
use M1M2_PR  M1M2_PR_341
timestamp 1655484843
transform 1 0 12006 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_342
timestamp 1655484843
transform 1 0 12098 0 1 16966
box -32 -32 32 32
use M1M2_PR  M1M2_PR_343
timestamp 1655484843
transform 1 0 12098 0 1 15334
box -32 -32 32 32
use M1M2_PR  M1M2_PR_344
timestamp 1655484843
transform 1 0 11362 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_345
timestamp 1655484843
transform 1 0 11362 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_346
timestamp 1655484843
transform 1 0 10810 0 1 13702
box -32 -32 32 32
use M1M2_PR  M1M2_PR_347
timestamp 1655484843
transform 1 0 10810 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_348
timestamp 1655484843
transform 1 0 10810 0 1 12954
box -32 -32 32 32
use M1M2_PR  M1M2_PR_349
timestamp 1655484843
transform 1 0 10810 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_350
timestamp 1655484843
transform 1 0 10626 0 1 11866
box -32 -32 32 32
use M1M2_PR  M1M2_PR_351
timestamp 1655484843
transform 1 0 10626 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_352
timestamp 1655484843
transform 1 0 10902 0 1 10778
box -32 -32 32 32
use M1M2_PR  M1M2_PR_353
timestamp 1655484843
transform 1 0 10902 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_354
timestamp 1655484843
transform 1 0 11086 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_355
timestamp 1655484843
transform 1 0 11086 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_356
timestamp 1655484843
transform 1 0 20194 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_357
timestamp 1655484843
transform 1 0 20194 0 1 7718
box -32 -32 32 32
use M1M2_PR  M1M2_PR_358
timestamp 1655484843
transform 1 0 18170 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_359
timestamp 1655484843
transform 1 0 18170 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_360
timestamp 1655484843
transform 1 0 21942 0 1 15674
box -32 -32 32 32
use M1M2_PR  M1M2_PR_361
timestamp 1655484843
transform 1 0 21942 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_362
timestamp 1655484843
transform 1 0 17894 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_363
timestamp 1655484843
transform 1 0 17894 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_364
timestamp 1655484843
transform 1 0 22494 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_365
timestamp 1655484843
transform 1 0 22494 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_366
timestamp 1655484843
transform 1 0 21666 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_367
timestamp 1655484843
transform 1 0 21666 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_368
timestamp 1655484843
transform 1 0 22494 0 1 15062
box -32 -32 32 32
use M1M2_PR  M1M2_PR_369
timestamp 1655484843
transform 1 0 22494 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_370
timestamp 1655484843
transform 1 0 22218 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_371
timestamp 1655484843
transform 1 0 22218 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_372
timestamp 1655484843
transform 1 0 22586 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_373
timestamp 1655484843
transform 1 0 22494 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_374
timestamp 1655484843
transform 1 0 22954 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_375
timestamp 1655484843
transform 1 0 22954 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_376
timestamp 1655484843
transform 1 0 18906 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_377
timestamp 1655484843
transform 1 0 18906 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_378
timestamp 1655484843
transform 1 0 16330 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_379
timestamp 1655484843
transform 1 0 16330 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_380
timestamp 1655484843
transform 1 0 16146 0 1 21114
box -32 -32 32 32
use M1M2_PR  M1M2_PR_381
timestamp 1655484843
transform 1 0 16146 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_382
timestamp 1655484843
transform 1 0 12742 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_383
timestamp 1655484843
transform 1 0 12466 0 1 15674
box -32 -32 32 32
use M1M2_PR  M1M2_PR_384
timestamp 1655484843
transform 1 0 13478 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_385
timestamp 1655484843
transform 1 0 13478 0 1 14246
box -32 -32 32 32
use M1M2_PR  M1M2_PR_386
timestamp 1655484843
transform 1 0 13478 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_387
timestamp 1655484843
transform 1 0 13478 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_388
timestamp 1655484843
transform 1 0 13018 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_389
timestamp 1655484843
transform 1 0 13018 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_390
timestamp 1655484843
transform 1 0 12650 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_391
timestamp 1655484843
transform 1 0 12650 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_392
timestamp 1655484843
transform 1 0 21666 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_393
timestamp 1655484843
transform 1 0 18814 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_394
timestamp 1655484843
transform 1 0 20746 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_395
timestamp 1655484843
transform 1 0 20746 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_396
timestamp 1655484843
transform 1 0 18998 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_397
timestamp 1655484843
transform 1 0 18998 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_398
timestamp 1655484843
transform 1 0 22218 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_399
timestamp 1655484843
transform 1 0 22218 0 1 6086
box -32 -32 32 32
use M1M2_PR  M1M2_PR_400
timestamp 1655484843
transform 1 0 22034 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_401
timestamp 1655484843
transform 1 0 22034 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_402
timestamp 1655484843
transform 1 0 21666 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_403
timestamp 1655484843
transform 1 0 21666 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_404
timestamp 1655484843
transform 1 0 18998 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_405
timestamp 1655484843
transform 1 0 18906 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_406
timestamp 1655484843
transform 1 0 22402 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_407
timestamp 1655484843
transform 1 0 22402 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_408
timestamp 1655484843
transform 1 0 20930 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_409
timestamp 1655484843
transform 1 0 20930 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_410
timestamp 1655484843
transform 1 0 14582 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_411
timestamp 1655484843
transform 1 0 14582 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_412
timestamp 1655484843
transform 1 0 13202 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_413
timestamp 1655484843
transform 1 0 13202 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_414
timestamp 1655484843
transform 1 0 12006 0 1 19482
box -32 -32 32 32
use M1M2_PR  M1M2_PR_415
timestamp 1655484843
transform 1 0 12006 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_416
timestamp 1655484843
transform 1 0 13386 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_417
timestamp 1655484843
transform 1 0 13386 0 1 17306
box -32 -32 32 32
use M1M2_PR  M1M2_PR_418
timestamp 1655484843
transform 1 0 13110 0 1 16694
box -32 -32 32 32
use M1M2_PR  M1M2_PR_419
timestamp 1655484843
transform 1 0 13110 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_420
timestamp 1655484843
transform 1 0 10718 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_421
timestamp 1655484843
transform 1 0 10718 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_422
timestamp 1655484843
transform 1 0 12742 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_423
timestamp 1655484843
transform 1 0 12742 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_424
timestamp 1655484843
transform 1 0 12006 0 1 11526
box -32 -32 32 32
use M1M2_PR  M1M2_PR_425
timestamp 1655484843
transform 1 0 11362 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_426
timestamp 1655484843
transform 1 0 11362 0 1 10438
box -32 -32 32 32
use M1M2_PR  M1M2_PR_427
timestamp 1655484843
transform 1 0 13018 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_428
timestamp 1655484843
transform 1 0 13018 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_429
timestamp 1655484843
transform 1 0 20194 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_430
timestamp 1655484843
transform 1 0 15686 0 1 7174
box -32 -32 32 32
use M1M2_PR  M1M2_PR_431
timestamp 1655484843
transform 1 0 18998 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_432
timestamp 1655484843
transform 1 0 18262 0 1 21794
box -32 -32 32 32
use M1M2_PR  M1M2_PR_433
timestamp 1655484843
transform 1 0 18262 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_434
timestamp 1655484843
transform 1 0 18446 0 1 21658
box -32 -32 32 32
use M1M2_PR  M1M2_PR_435
timestamp 1655484843
transform 1 0 18446 0 1 21114
box -32 -32 32 32
use M1M2_PR  M1M2_PR_436
timestamp 1655484843
transform 1 0 17434 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_437
timestamp 1655484843
transform 1 0 17434 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_438
timestamp 1655484843
transform 1 0 15962 0 1 21794
box -32 -32 32 32
use M1M2_PR  M1M2_PR_439
timestamp 1655484843
transform 1 0 15962 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_440
timestamp 1655484843
transform 1 0 14306 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_441
timestamp 1655484843
transform 1 0 14306 0 1 21114
box -32 -32 32 32
use M1M2_PR  M1M2_PR_442
timestamp 1655484843
transform 1 0 14306 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_443
timestamp 1655484843
transform 1 0 14490 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_444
timestamp 1655484843
transform 1 0 14490 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_445
timestamp 1655484843
transform 1 0 11546 0 1 20570
box -32 -32 32 32
use M1M2_PR  M1M2_PR_446
timestamp 1655484843
transform 1 0 11546 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_447
timestamp 1655484843
transform 1 0 11822 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_448
timestamp 1655484843
transform 1 0 11822 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_449
timestamp 1655484843
transform 1 0 11638 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_450
timestamp 1655484843
transform 1 0 11638 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_451
timestamp 1655484843
transform 1 0 11638 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_452
timestamp 1655484843
transform 1 0 11822 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_453
timestamp 1655484843
transform 1 0 11822 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_454
timestamp 1655484843
transform 1 0 10258 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_455
timestamp 1655484843
transform 1 0 10258 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_456
timestamp 1655484843
transform 1 0 11638 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_457
timestamp 1655484843
transform 1 0 11638 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_458
timestamp 1655484843
transform 1 0 10442 0 1 15674
box -32 -32 32 32
use M1M2_PR  M1M2_PR_459
timestamp 1655484843
transform 1 0 10442 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_460
timestamp 1655484843
transform 1 0 10442 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_461
timestamp 1655484843
transform 1 0 9062 0 1 14790
box -32 -32 32 32
use M1M2_PR  M1M2_PR_462
timestamp 1655484843
transform 1 0 9062 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_463
timestamp 1655484843
transform 1 0 10258 0 1 13702
box -32 -32 32 32
use M1M2_PR  M1M2_PR_464
timestamp 1655484843
transform 1 0 10258 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_465
timestamp 1655484843
transform 1 0 10442 0 1 12614
box -32 -32 32 32
use M1M2_PR  M1M2_PR_466
timestamp 1655484843
transform 1 0 10442 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_467
timestamp 1655484843
transform 1 0 8878 0 1 11526
box -32 -32 32 32
use M1M2_PR  M1M2_PR_468
timestamp 1655484843
transform 1 0 8878 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_469
timestamp 1655484843
transform 1 0 8694 0 1 8534
box -32 -32 32 32
use M1M2_PR  M1M2_PR_470
timestamp 1655484843
transform 1 0 8234 0 1 9690
box -32 -32 32 32
use M1M2_PR  M1M2_PR_471
timestamp 1655484843
transform 1 0 10442 0 1 8602
box -32 -32 32 32
use M1M2_PR  M1M2_PR_472
timestamp 1655484843
transform 1 0 10442 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_473
timestamp 1655484843
transform 1 0 11270 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_474
timestamp 1655484843
transform 1 0 11270 0 1 6426
box -32 -32 32 32
use M1M2_PR  M1M2_PR_475
timestamp 1655484843
transform 1 0 13294 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_476
timestamp 1655484843
transform 1 0 12282 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_477
timestamp 1655484843
transform 1 0 12190 0 1 7174
box -32 -32 32 32
use M1M2_PR  M1M2_PR_478
timestamp 1655484843
transform 1 0 13846 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_479
timestamp 1655484843
transform 1 0 13846 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_480
timestamp 1655484843
transform 1 0 11362 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_481
timestamp 1655484843
transform 1 0 11362 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_482
timestamp 1655484843
transform 1 0 9430 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_483
timestamp 1655484843
transform 1 0 9430 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_484
timestamp 1655484843
transform 1 0 10350 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_485
timestamp 1655484843
transform 1 0 10350 0 1 9350
box -32 -32 32 32
use M1M2_PR  M1M2_PR_486
timestamp 1655484843
transform 1 0 9062 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_487
timestamp 1655484843
transform 1 0 9062 0 1 10234
box -32 -32 32 32
use M1M2_PR  M1M2_PR_488
timestamp 1655484843
transform 1 0 10994 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_489
timestamp 1655484843
transform 1 0 10994 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_490
timestamp 1655484843
transform 1 0 10074 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_491
timestamp 1655484843
transform 1 0 10074 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_492
timestamp 1655484843
transform 1 0 10994 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_493
timestamp 1655484843
transform 1 0 10994 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_494
timestamp 1655484843
transform 1 0 10994 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_495
timestamp 1655484843
transform 1 0 10994 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_496
timestamp 1655484843
transform 1 0 12650 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_497
timestamp 1655484843
transform 1 0 12635 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_498
timestamp 1655484843
transform 1 0 15502 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_499
timestamp 1655484843
transform 1 0 16238 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_500
timestamp 1655484843
transform 1 0 16238 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_501
timestamp 1655484843
transform 1 0 18906 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_502
timestamp 1655484843
transform 1 0 18906 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_503
timestamp 1655484843
transform 1 0 19918 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_504
timestamp 1655484843
transform 1 0 19918 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_505
timestamp 1655484843
transform 1 0 20010 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_506
timestamp 1655484843
transform 1 0 20010 0 1 21386
box -32 -32 32 32
use M1M2_PR  M1M2_PR_507
timestamp 1655484843
transform 1 0 19182 0 1 21590
box -32 -32 32 32
use M1M2_PR  M1M2_PR_508
timestamp 1655484843
transform 1 0 19182 0 1 21318
box -32 -32 32 32
use M1M2_PR  M1M2_PR_509
timestamp 1655484843
transform 1 0 15502 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_510
timestamp 1655484843
transform 1 0 11362 0 1 17986
box -32 -32 32 32
use M1M2_PR  M1M2_PR_511
timestamp 1655484843
transform 1 0 11362 0 1 17034
box -32 -32 32 32
use M1M2_PR  M1M2_PR_512
timestamp 1655484843
transform 1 0 9246 0 1 16218
box -32 -32 32 32
use M1M2_PR  M1M2_PR_513
timestamp 1655484843
transform 1 0 9246 0 1 15402
box -32 -32 32 32
use M1M2_PR  M1M2_PR_514
timestamp 1655484843
transform 1 0 10258 0 1 16218
box -32 -32 32 32
use M1M2_PR  M1M2_PR_515
timestamp 1655484843
transform 1 0 10166 0 1 14858
box -32 -32 32 32
use M1M2_PR  M1M2_PR_516
timestamp 1655484843
transform 1 0 10718 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_517
timestamp 1655484843
transform 1 0 10718 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_518
timestamp 1655484843
transform 1 0 10258 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_519
timestamp 1655484843
transform 1 0 10258 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_520
timestamp 1655484843
transform 1 0 9062 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_521
timestamp 1655484843
transform 1 0 9062 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_522
timestamp 1655484843
transform 1 0 8878 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_523
timestamp 1655484843
transform 1 0 8878 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_524
timestamp 1655484843
transform 1 0 11638 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_525
timestamp 1655484843
transform 1 0 11638 0 1 6698
box -32 -32 32 32
use M1M2_PR  M1M2_PR_526
timestamp 1655484843
transform 1 0 12558 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_527
timestamp 1655484843
transform 1 0 12558 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_528
timestamp 1655484843
transform 1 0 6394 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_529
timestamp 1655484843
transform 1 0 6394 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_530
timestamp 1655484843
transform 1 0 6394 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_531
timestamp 1655484843
transform 1 0 6946 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_532
timestamp 1655484843
transform 1 0 6946 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_533
timestamp 1655484843
transform 1 0 6946 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_534
timestamp 1655484843
transform 1 0 6762 0 1 12410
box -32 -32 32 32
use M1M2_PR  M1M2_PR_535
timestamp 1655484843
transform 1 0 6762 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_536
timestamp 1655484843
transform 1 0 6854 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_537
timestamp 1655484843
transform 1 0 6578 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_538
timestamp 1655484843
transform 1 0 6578 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_539
timestamp 1655484843
transform 1 0 6486 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_540
timestamp 1655484843
transform 1 0 6486 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_541
timestamp 1655484843
transform 1 0 7866 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_542
timestamp 1655484843
transform 1 0 7866 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_543
timestamp 1655484843
transform 1 0 7866 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_544
timestamp 1655484843
transform 1 0 7682 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_545
timestamp 1655484843
transform 1 0 7682 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_546
timestamp 1655484843
transform 1 0 6854 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_547
timestamp 1655484843
transform 1 0 6854 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_548
timestamp 1655484843
transform 1 0 7038 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_549
timestamp 1655484843
transform 1 0 7038 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_550
timestamp 1655484843
transform 1 0 8510 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_551
timestamp 1655484843
transform 1 0 8418 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_552
timestamp 1655484843
transform 1 0 6762 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_553
timestamp 1655484843
transform 1 0 6762 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_554
timestamp 1655484843
transform 1 0 7958 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_555
timestamp 1655484843
transform 1 0 7958 0 1 13770
box -32 -32 32 32
use M1M2_PR  M1M2_PR_556
timestamp 1655484843
transform 1 0 6394 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_557
timestamp 1655484843
transform 1 0 6394 0 1 11526
box -32 -32 32 32
use M1M2_PR  M1M2_PR_558
timestamp 1655484843
transform 1 0 7774 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_559
timestamp 1655484843
transform 1 0 7774 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_560
timestamp 1655484843
transform 1 0 6578 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_561
timestamp 1655484843
transform 1 0 6578 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_562
timestamp 1655484843
transform 1 0 6394 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_563
timestamp 1655484843
transform 1 0 6394 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_564
timestamp 1655484843
transform 1 0 22494 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_565
timestamp 1655484843
transform 1 0 16882 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_566
timestamp 1655484843
transform 1 0 16422 0 1 9894
box -32 -32 32 32
use M1M2_PR  M1M2_PR_567
timestamp 1655484843
transform 1 0 20286 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_568
timestamp 1655484843
transform 1 0 20286 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_569
timestamp 1655484843
transform 1 0 18078 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_570
timestamp 1655484843
transform 1 0 18078 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_571
timestamp 1655484843
transform 1 0 20286 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_572
timestamp 1655484843
transform 1 0 16974 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_573
timestamp 1655484843
transform 1 0 16238 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_574
timestamp 1655484843
transform 1 0 14306 0 1 9622
box -32 -32 32 32
use M1M2_PR  M1M2_PR_575
timestamp 1655484843
transform 1 0 14306 0 1 8806
box -32 -32 32 32
use M1M2_PR  M1M2_PR_576
timestamp 1655484843
transform 1 0 11362 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_577
timestamp 1655484843
transform 1 0 11362 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_578
timestamp 1655484843
transform 1 0 13294 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_579
timestamp 1655484843
transform 1 0 13294 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_580
timestamp 1655484843
transform 1 0 13294 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_581
timestamp 1655484843
transform 1 0 13294 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_582
timestamp 1655484843
transform 1 0 12006 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_583
timestamp 1655484843
transform 1 0 12650 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_584
timestamp 1655484843
transform 1 0 12558 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_585
timestamp 1655484843
transform 1 0 14582 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_586
timestamp 1655484843
transform 1 0 14582 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_587
timestamp 1655484843
transform 1 0 11822 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_588
timestamp 1655484843
transform 1 0 11822 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_589
timestamp 1655484843
transform 1 0 13018 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_590
timestamp 1655484843
transform 1 0 12926 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_591
timestamp 1655484843
transform 1 0 12282 0 1 17986
box -32 -32 32 32
use M1M2_PR  M1M2_PR_592
timestamp 1655484843
transform 1 0 12282 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_593
timestamp 1655484843
transform 1 0 14306 0 1 17850
box -32 -32 32 32
use M1M2_PR  M1M2_PR_594
timestamp 1655484843
transform 1 0 14214 0 1 19414
box -32 -32 32 32
use M1M2_PR  M1M2_PR_595
timestamp 1655484843
transform 1 0 14214 0 1 19142
box -32 -32 32 32
use M1M2_PR  M1M2_PR_596
timestamp 1655484843
transform 1 0 14674 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_597
timestamp 1655484843
transform 1 0 14582 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_598
timestamp 1655484843
transform 1 0 14398 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_599
timestamp 1655484843
transform 1 0 16146 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_600
timestamp 1655484843
transform 1 0 16146 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_601
timestamp 1655484843
transform 1 0 16054 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_602
timestamp 1655484843
transform 1 0 17894 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_603
timestamp 1655484843
transform 1 0 17894 0 1 19550
box -32 -32 32 32
use M1M2_PR  M1M2_PR_604
timestamp 1655484843
transform 1 0 17894 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_605
timestamp 1655484843
transform 1 0 20194 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_606
timestamp 1655484843
transform 1 0 20194 0 1 19074
box -32 -32 32 32
use M1M2_PR  M1M2_PR_607
timestamp 1655484843
transform 1 0 20194 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_608
timestamp 1655484843
transform 1 0 21482 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_609
timestamp 1655484843
transform 1 0 21482 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_610
timestamp 1655484843
transform 1 0 21114 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_611
timestamp 1655484843
transform 1 0 21114 0 1 17306
box -32 -32 32 32
use M1M2_PR  M1M2_PR_612
timestamp 1655484843
transform 1 0 20378 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_613
timestamp 1655484843
transform 1 0 20378 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_614
timestamp 1655484843
transform 1 0 20378 0 1 14790
box -32 -32 32 32
use M1M2_PR  M1M2_PR_615
timestamp 1655484843
transform 1 0 22126 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_616
timestamp 1655484843
transform 1 0 22034 0 1 19754
box -32 -32 32 32
use M1M2_PR  M1M2_PR_617
timestamp 1655484843
transform 1 0 21298 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_618
timestamp 1655484843
transform 1 0 22954 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_619
timestamp 1655484843
transform 1 0 22954 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_620
timestamp 1655484843
transform 1 0 21666 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_621
timestamp 1655484843
transform 1 0 21666 0 1 12682
box -32 -32 32 32
use M1M2_PR  M1M2_PR_622
timestamp 1655484843
transform 1 0 21298 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_623
timestamp 1655484843
transform 1 0 21298 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_624
timestamp 1655484843
transform 1 0 21206 0 1 12002
box -32 -32 32 32
use M1M2_PR  M1M2_PR_625
timestamp 1655484843
transform 1 0 20102 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_626
timestamp 1655484843
transform 1 0 20010 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_627
timestamp 1655484843
transform 1 0 19918 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_628
timestamp 1655484843
transform 1 0 19826 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_629
timestamp 1655484843
transform 1 0 21666 0 1 11526
box -32 -32 32 32
use M1M2_PR  M1M2_PR_630
timestamp 1655484843
transform 1 0 21666 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_631
timestamp 1655484843
transform 1 0 20746 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_632
timestamp 1655484843
transform 1 0 20378 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_633
timestamp 1655484843
transform 1 0 21390 0 1 11254
box -32 -32 32 32
use M1M2_PR  M1M2_PR_634
timestamp 1655484843
transform 1 0 21390 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_635
timestamp 1655484843
transform 1 0 21114 0 1 10982
box -32 -32 32 32
use M1M2_PR  M1M2_PR_636
timestamp 1655484843
transform 1 0 21022 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_637
timestamp 1655484843
transform 1 0 21942 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_638
timestamp 1655484843
transform 1 0 21942 0 1 10234
box -32 -32 32 32
use M1M2_PR  M1M2_PR_639
timestamp 1655484843
transform 1 0 21758 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_640
timestamp 1655484843
transform 1 0 16238 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_641
timestamp 1655484843
transform 1 0 16238 0 1 6086
box -32 -32 32 32
use M1M2_PR  M1M2_PR_642
timestamp 1655484843
transform 1 0 20010 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_643
timestamp 1655484843
transform 1 0 20010 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_644
timestamp 1655484843
transform 1 0 15226 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_645
timestamp 1655484843
transform 1 0 15226 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_646
timestamp 1655484843
transform 1 0 13110 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_647
timestamp 1655484843
transform 1 0 13110 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_648
timestamp 1655484843
transform 1 0 17618 0 1 8534
box -32 -32 32 32
use M1M2_PR  M1M2_PR_649
timestamp 1655484843
transform 1 0 17618 0 1 8262
box -32 -32 32 32
use M1M2_PR  M1M2_PR_650
timestamp 1655484843
transform 1 0 12006 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_651
timestamp 1655484843
transform 1 0 12006 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_652
timestamp 1655484843
transform 1 0 10718 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_653
timestamp 1655484843
transform 1 0 10718 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_654
timestamp 1655484843
transform 1 0 10718 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_655
timestamp 1655484843
transform 1 0 10718 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_656
timestamp 1655484843
transform 1 0 10534 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_657
timestamp 1655484843
transform 1 0 10534 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_658
timestamp 1655484843
transform 1 0 10534 0 1 10506
box -32 -32 32 32
use M1M2_PR  M1M2_PR_659
timestamp 1655484843
transform 1 0 8878 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_660
timestamp 1655484843
transform 1 0 8878 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_661
timestamp 1655484843
transform 1 0 9522 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_662
timestamp 1655484843
transform 1 0 9522 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_663
timestamp 1655484843
transform 1 0 10994 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_664
timestamp 1655484843
transform 1 0 10902 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_665
timestamp 1655484843
transform 1 0 12006 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_666
timestamp 1655484843
transform 1 0 11914 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_667
timestamp 1655484843
transform 1 0 10810 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_668
timestamp 1655484843
transform 1 0 10810 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_669
timestamp 1655484843
transform 1 0 11914 0 1 16830
box -32 -32 32 32
use M1M2_PR  M1M2_PR_670
timestamp 1655484843
transform 1 0 11914 0 1 16218
box -32 -32 32 32
use M1M2_PR  M1M2_PR_671
timestamp 1655484843
transform 1 0 12190 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_672
timestamp 1655484843
transform 1 0 12190 0 1 18666
box -32 -32 32 32
use M1M2_PR  M1M2_PR_673
timestamp 1655484843
transform 1 0 12190 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_674
timestamp 1655484843
transform 1 0 13386 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_675
timestamp 1655484843
transform 1 0 13386 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_676
timestamp 1655484843
transform 1 0 13386 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_677
timestamp 1655484843
transform 1 0 14766 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_678
timestamp 1655484843
transform 1 0 14766 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_679
timestamp 1655484843
transform 1 0 13478 0 1 19958
box -32 -32 32 32
use M1M2_PR  M1M2_PR_680
timestamp 1655484843
transform 1 0 13478 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_681
timestamp 1655484843
transform 1 0 17158 0 1 21318
box -32 -32 32 32
use M1M2_PR  M1M2_PR_682
timestamp 1655484843
transform 1 0 17158 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_683
timestamp 1655484843
transform 1 0 17158 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_684
timestamp 1655484843
transform 1 0 17710 0 1 21046
box -32 -32 32 32
use M1M2_PR  M1M2_PR_685
timestamp 1655484843
transform 1 0 17710 0 1 20502
box -32 -32 32 32
use M1M2_PR  M1M2_PR_686
timestamp 1655484843
transform 1 0 17710 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_687
timestamp 1655484843
transform 1 0 22770 0 1 21794
box -32 -32 32 32
use M1M2_PR  M1M2_PR_688
timestamp 1655484843
transform 1 0 20470 0 1 20842
box -32 -32 32 32
use M1M2_PR  M1M2_PR_689
timestamp 1655484843
transform 1 0 20378 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_690
timestamp 1655484843
transform 1 0 20378 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_691
timestamp 1655484843
transform 1 0 21298 0 1 21794
box -32 -32 32 32
use M1M2_PR  M1M2_PR_692
timestamp 1655484843
transform 1 0 21298 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_693
timestamp 1655484843
transform 1 0 9154 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_694
timestamp 1655484843
transform 1 0 9154 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_695
timestamp 1655484843
transform 1 0 6118 0 1 7446
box -32 -32 32 32
use M1M2_PR  M1M2_PR_696
timestamp 1655484843
transform 1 0 6118 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_697
timestamp 1655484843
transform 1 0 6118 0 1 6630
box -32 -32 32 32
use M1M2_PR  M1M2_PR_698
timestamp 1655484843
transform 1 0 7498 0 1 6902
box -32 -32 32 32
use M1M2_PR  M1M2_PR_699
timestamp 1655484843
transform 1 0 7498 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_700
timestamp 1655484843
transform 1 0 10350 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_701
timestamp 1655484843
transform 1 0 10350 0 1 6154
box -32 -32 32 32
use M1M2_PR  M1M2_PR_702
timestamp 1655484843
transform 1 0 8326 0 1 8534
box -32 -32 32 32
use M1M2_PR  M1M2_PR_703
timestamp 1655484843
transform 1 0 8326 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_704
timestamp 1655484843
transform 1 0 8326 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_705
timestamp 1655484843
transform 1 0 8326 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_706
timestamp 1655484843
transform 1 0 8694 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_707
timestamp 1655484843
transform 1 0 8694 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_708
timestamp 1655484843
transform 1 0 8694 0 1 10438
box -32 -32 32 32
use M1M2_PR  M1M2_PR_709
timestamp 1655484843
transform 1 0 7958 0 1 12546
box -32 -32 32 32
use M1M2_PR  M1M2_PR_710
timestamp 1655484843
transform 1 0 7958 0 1 11594
box -32 -32 32 32
use M1M2_PR  M1M2_PR_711
timestamp 1655484843
transform 1 0 9154 0 1 13974
box -32 -32 32 32
use M1M2_PR  M1M2_PR_712
timestamp 1655484843
transform 1 0 9154 0 1 13634
box -32 -32 32 32
use M1M2_PR  M1M2_PR_713
timestamp 1655484843
transform 1 0 6762 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_714
timestamp 1655484843
transform 1 0 6762 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_715
timestamp 1655484843
transform 1 0 6578 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_716
timestamp 1655484843
transform 1 0 6578 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_717
timestamp 1655484843
transform 1 0 17526 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_718
timestamp 1655484843
transform 1 0 17526 0 1 9962
box -32 -32 32 32
use M1M2_PR  M1M2_PR_719
timestamp 1655484843
transform 1 0 17250 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_720
timestamp 1655484843
transform 1 0 17250 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_721
timestamp 1655484843
transform 1 0 16514 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_722
timestamp 1655484843
transform 1 0 16514 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_723
timestamp 1655484843
transform 1 0 15594 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_724
timestamp 1655484843
transform 1 0 15410 0 1 8874
box -32 -32 32 32
use M1M2_PR  M1M2_PR_725
timestamp 1655484843
transform 1 0 14582 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_726
timestamp 1655484843
transform 1 0 14582 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_727
timestamp 1655484843
transform 1 0 15778 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_728
timestamp 1655484843
transform 1 0 15778 0 1 11050
box -32 -32 32 32
use M1M2_PR  M1M2_PR_729
timestamp 1655484843
transform 1 0 14582 0 1 13158
box -32 -32 32 32
use M1M2_PR  M1M2_PR_730
timestamp 1655484843
transform 1 0 14582 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_731
timestamp 1655484843
transform 1 0 16790 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_732
timestamp 1655484843
transform 1 0 16790 0 1 12138
box -32 -32 32 32
use M1M2_PR  M1M2_PR_733
timestamp 1655484843
transform 1 0 15870 0 1 14518
box -32 -32 32 32
use M1M2_PR  M1M2_PR_734
timestamp 1655484843
transform 1 0 15870 0 1 12546
box -32 -32 32 32
use M1M2_PR  M1M2_PR_735
timestamp 1655484843
transform 1 0 14306 0 1 15606
box -32 -32 32 32
use M1M2_PR  M1M2_PR_736
timestamp 1655484843
transform 1 0 14306 0 1 14246
box -32 -32 32 32
use M1M2_PR  M1M2_PR_737
timestamp 1655484843
transform 1 0 14858 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_738
timestamp 1655484843
transform 1 0 14306 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_739
timestamp 1655484843
transform 1 0 16698 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_740
timestamp 1655484843
transform 1 0 16698 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_741
timestamp 1655484843
transform 1 0 15778 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_742
timestamp 1655484843
transform 1 0 15778 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_743
timestamp 1655484843
transform 1 0 10534 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_744
timestamp 1655484843
transform 1 0 10350 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_745
timestamp 1655484843
transform 1 0 10350 0 1 20298
box -32 -32 32 32
use M1M2_PR  M1M2_PR_746
timestamp 1655484843
transform 1 0 9614 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_747
timestamp 1655484843
transform 1 0 9614 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_748
timestamp 1655484843
transform 1 0 8970 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_749
timestamp 1655484843
transform 1 0 8970 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_750
timestamp 1655484843
transform 1 0 7038 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_751
timestamp 1655484843
transform 1 0 6946 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_752
timestamp 1655484843
transform 1 0 6946 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_753
timestamp 1655484843
transform 1 0 6946 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_754
timestamp 1655484843
transform 1 0 6946 0 1 15946
box -32 -32 32 32
use M1M2_PR  M1M2_PR_755
timestamp 1655484843
transform 1 0 22954 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_756
timestamp 1655484843
transform 1 0 22954 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_757
timestamp 1655484843
transform 1 0 22402 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_758
timestamp 1655484843
transform 1 0 22310 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_759
timestamp 1655484843
transform 1 0 22310 0 1 15198
box -32 -32 32 32
use M1M2_PR  M1M2_PR_760
timestamp 1655484843
transform 1 0 22310 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_761
timestamp 1655484843
transform 1 0 22218 0 1 18530
box -32 -32 32 32
use M1M2_PR  M1M2_PR_762
timestamp 1655484843
transform 1 0 22218 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_763
timestamp 1655484843
transform 1 0 22218 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_764
timestamp 1655484843
transform 1 0 22034 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_765
timestamp 1655484843
transform 1 0 21574 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_766
timestamp 1655484843
transform 1 0 21574 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_767
timestamp 1655484843
transform 1 0 20838 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_768
timestamp 1655484843
transform 1 0 20838 0 1 9826
box -32 -32 32 32
use M1M2_PR  M1M2_PR_769
timestamp 1655484843
transform 1 0 17802 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_770
timestamp 1655484843
transform 1 0 17802 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_771
timestamp 1655484843
transform 1 0 16882 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_772
timestamp 1655484843
transform 1 0 13386 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_773
timestamp 1655484843
transform 1 0 13386 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_774
timestamp 1655484843
transform 1 0 13386 0 1 13566
box -32 -32 32 32
use M1M2_PR  M1M2_PR_775
timestamp 1655484843
transform 1 0 13202 0 1 7242
box -32 -32 32 32
use M1M2_PR  M1M2_PR_776
timestamp 1655484843
transform 1 0 13110 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_777
timestamp 1655484843
transform 1 0 13110 0 1 8670
box -32 -32 32 32
use M1M2_PR  M1M2_PR_778
timestamp 1655484843
transform 1 0 13018 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_779
timestamp 1655484843
transform 1 0 12834 0 1 16422
box -32 -32 32 32
use M1M2_PR  M1M2_PR_780
timestamp 1655484843
transform 1 0 12742 0 1 19550
box -32 -32 32 32
use M1M2_PR  M1M2_PR_781
timestamp 1655484843
transform 1 0 12374 0 1 20026
box -32 -32 32 32
use M1M2_PR  M1M2_PR_782
timestamp 1655484843
transform 1 0 12374 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_783
timestamp 1655484843
transform 1 0 11638 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_784
timestamp 1655484843
transform 1 0 11638 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_785
timestamp 1655484843
transform 1 0 11638 0 1 10370
box -32 -32 32 32
use M1M2_PR  M1M2_PR_786
timestamp 1655484843
transform 1 0 11638 0 1 9418
box -32 -32 32 32
use M1M2_PR  M1M2_PR_787
timestamp 1655484843
transform 1 0 19642 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_788
timestamp 1655484843
transform 1 0 19642 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_789
timestamp 1655484843
transform 1 0 18170 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_790
timestamp 1655484843
transform 1 0 16514 0 1 21726
box -32 -32 32 32
use M1M2_PR  M1M2_PR_791
timestamp 1655484843
transform 1 0 16514 0 1 21250
box -32 -32 32 32
use M1M2_PR  M1M2_PR_792
timestamp 1655484843
transform 1 0 15134 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_793
timestamp 1655484843
transform 1 0 15134 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_794
timestamp 1655484843
transform 1 0 13110 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_795
timestamp 1655484843
transform 1 0 13110 0 1 20774
box -32 -32 32 32
use M1M2_PR  M1M2_PR_796
timestamp 1655484843
transform 1 0 12926 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_797
timestamp 1655484843
transform 1 0 12926 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_798
timestamp 1655484843
transform 1 0 10994 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_799
timestamp 1655484843
transform 1 0 10994 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_800
timestamp 1655484843
transform 1 0 10258 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_801
timestamp 1655484843
transform 1 0 10074 0 1 12954
box -32 -32 32 32
use M1M2_PR  M1M2_PR_802
timestamp 1655484843
transform 1 0 10074 0 1 11934
box -32 -32 32 32
use M1M2_PR  M1M2_PR_803
timestamp 1655484843
transform 1 0 10074 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_804
timestamp 1655484843
transform 1 0 10074 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_805
timestamp 1655484843
transform 1 0 10074 0 1 7786
box -32 -32 32 32
use M1M2_PR  M1M2_PR_806
timestamp 1655484843
transform 1 0 10074 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_807
timestamp 1655484843
transform 1 0 9890 0 1 16286
box -32 -32 32 32
use M1M2_PR  M1M2_PR_808
timestamp 1655484843
transform 1 0 10902 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_809
timestamp 1655484843
transform 1 0 10902 0 1 16898
box -32 -32 32 32
use M1M2_PR  M1M2_PR_810
timestamp 1655484843
transform 1 0 10718 0 1 18462
box -32 -32 32 32
use M1M2_PR  M1M2_PR_811
timestamp 1655484843
transform 1 0 10718 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_812
timestamp 1655484843
transform 1 0 10626 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_813
timestamp 1655484843
transform 1 0 10258 0 1 6970
box -32 -32 32 32
use M1M2_PR  M1M2_PR_814
timestamp 1655484843
transform 1 0 9522 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_815
timestamp 1655484843
transform 1 0 8694 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_816
timestamp 1655484843
transform 1 0 8234 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_817
timestamp 1655484843
transform 1 0 7314 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_818
timestamp 1655484843
transform 1 0 7314 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_819
timestamp 1655484843
transform 1 0 7314 0 1 16354
box -32 -32 32 32
use M1M2_PR  M1M2_PR_820
timestamp 1655484843
transform 1 0 7314 0 1 14178
box -32 -32 32 32
use M1M2_PR  M1M2_PR_821
timestamp 1655484843
transform 1 0 7314 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_822
timestamp 1655484843
transform 1 0 7314 0 1 10846
box -32 -32 32 32
use M1M2_PR  M1M2_PR_823
timestamp 1655484843
transform 1 0 7314 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_824
timestamp 1655484843
transform 1 0 7222 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_825
timestamp 1655484843
transform 1 0 7222 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_826
timestamp 1655484843
transform 1 0 7222 0 1 9214
box -32 -32 32 32
use M1M2_PR  M1M2_PR_827
timestamp 1655484843
transform 1 0 7222 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_828
timestamp 1655484843
transform 1 0 6946 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_829
timestamp 1655484843
transform 1 0 6946 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_830
timestamp 1655484843
transform 1 0 6854 0 1 20162
box -32 -32 32 32
use M1M2_PR  M1M2_PR_831
timestamp 1655484843
transform 1 0 21390 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_832
timestamp 1655484843
transform 1 0 19826 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_833
timestamp 1655484843
transform 1 0 19274 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_834
timestamp 1655484843
transform 1 0 18814 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_835
timestamp 1655484843
transform 1 0 16238 0 1 7106
box -32 -32 32 32
use M1M2_PR  M1M2_PR_836
timestamp 1655484843
transform 1 0 14674 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_837
timestamp 1655484843
transform 1 0 13662 0 1 7038
box -32 -32 32 32
use M1M2_PR  M1M2_PR_838
timestamp 1655484843
transform 1 0 13294 0 1 12546
box -32 -32 32 32
use M1M2_PR  M1M2_PR_839
timestamp 1655484843
transform 1 0 12466 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_840
timestamp 1655484843
transform 1 0 12374 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_841
timestamp 1655484843
transform 1 0 12374 0 1 14654
box -32 -32 32 32
use M1M2_PR  M1M2_PR_842
timestamp 1655484843
transform 1 0 12374 0 1 14110
box -32 -32 32 32
use M1M2_PR  M1M2_PR_843
timestamp 1655484843
transform 1 0 12374 0 1 13022
box -32 -32 32 32
use M1M2_PR  M1M2_PR_844
timestamp 1655484843
transform 1 0 12374 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_845
timestamp 1655484843
transform 1 0 12374 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_846
timestamp 1655484843
transform 1 0 12374 0 1 9758
box -32 -32 32 32
use M1M2_PR  M1M2_PR_847
timestamp 1655484843
transform 1 0 12374 0 1 7582
box -32 -32 32 32
use M1M2_PR  M1M2_PR_848
timestamp 1655484843
transform 1 0 12374 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_849
timestamp 1655484843
transform 1 0 10718 0 1 8194
box -32 -32 32 32
use M1M2_PR  M1M2_PR_850
timestamp 1655484843
transform 1 0 9154 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_851
timestamp 1655484843
transform 1 0 9154 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_852
timestamp 1655484843
transform 1 0 9154 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_853
timestamp 1655484843
transform 1 0 22954 0 1 20162
box -32 -32 32 32
use M1M2_PR  M1M2_PR_854
timestamp 1655484843
transform 1 0 22770 0 1 19550
box -32 -32 32 32
use M1M2_PR  M1M2_PR_855
timestamp 1655484843
transform 1 0 22770 0 1 19006
box -32 -32 32 32
use M1M2_PR  M1M2_PR_856
timestamp 1655484843
transform 1 0 22770 0 1 17442
box -32 -32 32 32
use M1M2_PR  M1M2_PR_857
timestamp 1655484843
transform 1 0 22770 0 1 15810
box -32 -32 32 32
use M1M2_PR  M1M2_PR_858
timestamp 1655484843
transform 1 0 22770 0 1 11458
box -32 -32 32 32
use M1M2_PR  M1M2_PR_859
timestamp 1655484843
transform 1 0 21114 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_860
timestamp 1655484843
transform 1 0 20102 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_861
timestamp 1655484843
transform 1 0 20102 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_862
timestamp 1655484843
transform 1 0 20102 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_863
timestamp 1655484843
transform 1 0 19182 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_864
timestamp 1655484843
transform 1 0 15962 0 1 21182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_865
timestamp 1655484843
transform 1 0 15962 0 1 20638
box -32 -32 32 32
use M1M2_PR  M1M2_PR_866
timestamp 1655484843
transform 1 0 15962 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_867
timestamp 1655484843
transform 1 0 12650 0 1 20706
box -32 -32 32 32
use M1M2_PR  M1M2_PR_868
timestamp 1655484843
transform 1 0 12650 0 1 20094
box -32 -32 32 32
use M1M2_PR  M1M2_PR_869
timestamp 1655484843
transform 1 0 12650 0 1 19618
box -32 -32 32 32
use M1M2_PR  M1M2_PR_870
timestamp 1655484843
transform 1 0 20194 0 1 12478
box -32 -32 32 32
use M1M2_PR  M1M2_PR_871
timestamp 1655484843
transform 1 0 18630 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_872
timestamp 1655484843
transform 1 0 18630 0 1 6494
box -32 -32 32 32
use M1M2_PR  M1M2_PR_873
timestamp 1655484843
transform 1 0 18354 0 1 8738
box -32 -32 32 32
use M1M2_PR  M1M2_PR_874
timestamp 1655484843
transform 1 0 18354 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_875
timestamp 1655484843
transform 1 0 18354 0 1 6562
box -32 -32 32 32
use M1M2_PR  M1M2_PR_876
timestamp 1655484843
transform 1 0 17342 0 1 17918
box -32 -32 32 32
use M1M2_PR  M1M2_PR_877
timestamp 1655484843
transform 1 0 14858 0 1 8058
box -32 -32 32 32
use M1M2_PR  M1M2_PR_878
timestamp 1655484843
transform 1 0 14766 0 1 15266
box -32 -32 32 32
use M1M2_PR  M1M2_PR_879
timestamp 1655484843
transform 1 0 14766 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_880
timestamp 1655484843
transform 1 0 14306 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_881
timestamp 1655484843
transform 1 0 14306 0 1 6018
box -32 -32 32 32
use M1M2_PR  M1M2_PR_882
timestamp 1655484843
transform 1 0 28750 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_883
timestamp 1655484843
transform 1 0 17986 0 1 12342
box -32 -32 32 32
use M1M2_PR  M1M2_PR_884
timestamp 1655484843
transform 1 0 17986 0 1 12070
box -32 -32 32 32
use M1M2_PR  M1M2_PR_885
timestamp 1655484843
transform 1 0 11822 0 1 13974
box -32 -32 32 32
use M1M2_PR  M1M2_PR_886
timestamp 1655484843
transform 1 0 11822 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_887
timestamp 1655484843
transform 1 0 10626 0 1 14314
box -32 -32 32 32
use M1M2_PR  M1M2_PR_888
timestamp 1655484843
transform 1 0 18630 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_889
timestamp 1655484843
transform 1 0 17802 0 1 18870
box -32 -32 32 32
use M1M2_PR  M1M2_PR_890
timestamp 1655484843
transform 1 0 17802 0 1 18598
box -32 -32 32 32
use M1M2_PR  M1M2_PR_891
timestamp 1655484843
transform 1 0 21850 0 1 18326
box -32 -32 32 32
use M1M2_PR  M1M2_PR_892
timestamp 1655484843
transform 1 0 21850 0 1 17578
box -32 -32 32 32
use M1M2_PR  M1M2_PR_893
timestamp 1655484843
transform 1 0 26450 0 1 18122
box -32 -32 32 32
use M1M2_PR  M1M2_PR_894
timestamp 1655484843
transform 1 0 21482 0 1 17782
box -32 -32 32 32
use M1M2_PR  M1M2_PR_895
timestamp 1655484843
transform 1 0 21482 0 1 16762
box -32 -32 32 32
use M1M2_PR  M1M2_PR_896
timestamp 1655484843
transform 1 0 19090 0 1 17306
box -32 -32 32 32
use M1M2_PR  M1M2_PR_897
timestamp 1655484843
transform 1 0 19090 0 1 15742
box -32 -32 32 32
use M1M2_PR  M1M2_PR_898
timestamp 1655484843
transform 1 0 21666 0 1 16490
box -32 -32 32 32
use M1M2_PR  M1M2_PR_899
timestamp 1655484843
transform 1 0 21298 0 1 16150
box -32 -32 32 32
use M1M2_PR  M1M2_PR_900
timestamp 1655484843
transform 1 0 20470 0 1 14722
box -32 -32 32 32
use M1M2_PR  M1M2_PR_901
timestamp 1655484843
transform 1 0 22954 0 1 13974
box -32 -32 32 32
use M1M2_PR  M1M2_PR_902
timestamp 1655484843
transform 1 0 20562 0 1 13498
box -32 -32 32 32
use M1M2_PR  M1M2_PR_903
timestamp 1655484843
transform 1 0 20562 0 1 13226
box -32 -32 32 32
use M1M2_PR  M1M2_PR_904
timestamp 1655484843
transform 1 0 21850 0 1 13090
box -32 -32 32 32
use M1M2_PR  M1M2_PR_905
timestamp 1655484843
transform 1 0 21758 0 1 11798
box -32 -32 32 32
use M1M2_PR  M1M2_PR_906
timestamp 1655484843
transform 1 0 22034 0 1 9146
box -32 -32 32 32
use M1M2_PR  M1M2_PR_907
timestamp 1655484843
transform 1 0 23230 0 1 10302
box -32 -32 32 32
use M1M2_PR  M1M2_PR_908
timestamp 1655484843
transform 1 0 23230 0 1 8330
box -32 -32 32 32
use M1M2_PR  M1M2_PR_909
timestamp 1655484843
transform 1 0 26266 0 1 10710
box -32 -32 32 32
use M1M2_PR  M1M2_PR_910
timestamp 1655484843
transform 1 0 20562 0 1 11322
box -32 -32 32 32
use M1M2_PR  M1M2_PR_911
timestamp 1655484843
transform 1 0 22770 0 1 10166
box -32 -32 32 32
use M1M2_PR  M1M2_PR_912
timestamp 1655484843
transform 1 0 20562 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_913
timestamp 1655484843
transform 1 0 5934 0 1 7514
box -32 -32 32 32
use M1M2_PR  M1M2_PR_914
timestamp 1655484843
transform 1 0 13478 0 1 7990
box -32 -32 32 32
use M1M2_PR  M1M2_PR_915
timestamp 1655484843
transform 1 0 13478 0 1 170
box -32 -32 32 32
use M1M2_PR  M1M2_PR_916
timestamp 1655484843
transform 1 0 46 0 1 170
box -32 -32 32 32
use M1M2_PR  M1M2_PR_917
timestamp 1655484843
transform 1 0 9982 0 1 6358
box -32 -32 32 32
use M1M2_PR  M1M2_PR_918
timestamp 1655484843
transform 1 0 19182 0 1 4114
box -32 -32 32 32
use M1M2_PR  M1M2_PR_919
timestamp 1655484843
transform 1 0 10902 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_920
timestamp 1655484843
transform 1 0 10902 0 1 4182
box -32 -32 32 32
use M1M2_PR  M1M2_PR_921
timestamp 1655484843
transform 1 0 6762 0 1 5950
box -32 -32 32 32
use M1M2_PR  M1M2_PR_922
timestamp 1655484843
transform 1 0 6670 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_923
timestamp 1655484843
transform 1 0 6670 0 1 10914
box -32 -32 32 32
use M1M2_PR  M1M2_PR_924
timestamp 1655484843
transform 1 0 6670 0 1 9282
box -32 -32 32 32
use M1M2_PR  M1M2_PR_925
timestamp 1655484843
transform 1 0 6670 0 1 8126
box -32 -32 32 32
use M1M2_PR  M1M2_PR_926
timestamp 1655484843
transform 1 0 6670 0 1 7650
box -32 -32 32 32
use M1M2_PR  M1M2_PR_927
timestamp 1655484843
transform 1 0 6210 0 1 13430
box -32 -32 32 32
use M1M2_PR  M1M2_PR_928
timestamp 1655484843
transform 1 0 6210 0 1 11390
box -32 -32 32 32
use M1M2_PR  M1M2_PR_929
timestamp 1655484843
transform 1 0 14122 0 1 5882
box -32 -32 32 32
use M1M2_PR_MR  M1M2_PR_MR_0
timestamp 1655484843
transform 1 0 12006 0 1 11934
box -26 -32 26 32
use M1M2_PR_MR  M1M2_PR_MR_1
timestamp 1655484843
transform 1 0 12006 0 1 13022
box -26 -32 26 32
use M1M2_PR_MR  M1M2_PR_MR_2
timestamp 1655484843
transform 1 0 12558 0 1 13634
box -26 -32 26 32
use M1M2_PR_MR  M1M2_PR_MR_3
timestamp 1655484843
transform 1 0 18354 0 1 9826
box -26 -32 26 32
use M1M2_PR_MR  M1M2_PR_MR_4
timestamp 1655484843
transform 1 0 15778 0 1 14178
box -26 -32 26 32
use M1M2_PR_M  M1M2_PR_M_0
timestamp 1655484843
transform 1 0 16054 0 1 13226
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_1
timestamp 1655484843
transform 1 0 20378 0 1 14654
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_2
timestamp 1655484843
transform 1 0 20102 0 1 14654
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_3
timestamp 1655484843
transform 1 0 21022 0 1 14858
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_4
timestamp 1655484843
transform 1 0 15318 0 1 17034
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_5
timestamp 1655484843
transform 1 0 18814 0 1 14722
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_6
timestamp 1655484843
transform 1 0 19366 0 1 9078
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_7
timestamp 1655484843
transform 1 0 18538 0 1 9146
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_8
timestamp 1655484843
transform 1 0 13478 0 1 9282
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_9
timestamp 1655484843
transform 1 0 18998 0 1 7242
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_10
timestamp 1655484843
transform 1 0 15502 0 1 20502
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_11
timestamp 1655484843
transform 1 0 15502 0 1 21590
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_12
timestamp 1655484843
transform 1 0 10258 0 1 17918
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_13
timestamp 1655484843
transform 1 0 10718 0 1 20162
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_14
timestamp 1655484843
transform 1 0 7314 0 1 11934
box -32 -26 32 26
use M1M2_PR_M  M1M2_PR_M_15
timestamp 1655484843
transform 1 0 20562 0 1 10710
box -32 -26 32 26
use M1M2_PR_R  M1M2_PR_R_0
timestamp 1655484843
transform 1 0 18814 0 1 13634
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_1
timestamp 1655484843
transform 1 0 19826 0 1 17918
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_2
timestamp 1655484843
transform 1 0 18814 0 1 10370
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_3
timestamp 1655484843
transform 1 0 22770 0 1 17986
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_4
timestamp 1655484843
transform 1 0 22770 0 1 14722
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_5
timestamp 1655484843
transform 1 0 22770 0 1 13634
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_6
timestamp 1655484843
transform 1 0 9338 0 1 7038
box -32 -32 32 32
use M1M2_PR_R  M1M2_PR_R_7
timestamp 1655484843
transform 1 0 17342 0 1 15674
box -32 -32 32 32
use M2M3_PR  M2M3_PR_0
timestamp 1655484843
transform 1 0 17526 0 1 12578
box -33 -37 33 37
use M2M3_PR  M2M3_PR_1
timestamp 1655484843
transform 1 0 16790 0 1 12578
box -33 -37 33 37
use M2M3_PR  M2M3_PR_2
timestamp 1655484843
transform 1 0 20930 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_3
timestamp 1655484843
transform 1 0 20654 0 1 14774
box -33 -37 33 37
use M2M3_PR  M2M3_PR_4
timestamp 1655484843
transform 1 0 20470 0 1 13676
box -33 -37 33 37
use M2M3_PR  M2M3_PR_5
timestamp 1655484843
transform 1 0 20378 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_6
timestamp 1655484843
transform 1 0 19550 0 1 17458
box -33 -37 33 37
use M2M3_PR  M2M3_PR_7
timestamp 1655484843
transform 1 0 19550 0 1 16848
box -33 -37 33 37
use M2M3_PR  M2M3_PR_8
timestamp 1655484843
transform 1 0 19090 0 1 14774
box -33 -37 33 37
use M2M3_PR  M2M3_PR_9
timestamp 1655484843
transform 1 0 19090 0 1 13676
box -33 -37 33 37
use M2M3_PR  M2M3_PR_10
timestamp 1655484843
transform 1 0 17986 0 1 10382
box -33 -37 33 37
use M2M3_PR  M2M3_PR_11
timestamp 1655484843
transform 1 0 17894 0 1 17458
box -33 -37 33 37
use M2M3_PR  M2M3_PR_12
timestamp 1655484843
transform 1 0 16790 0 1 12944
box -33 -37 33 37
use M2M3_PR  M2M3_PR_13
timestamp 1655484843
transform 1 0 15870 0 1 12334
box -33 -37 33 37
use M2M3_PR  M2M3_PR_14
timestamp 1655484843
transform 1 0 15778 0 1 10382
box -33 -37 33 37
use M2M3_PR  M2M3_PR_15
timestamp 1655484843
transform 1 0 15318 0 1 13676
box -33 -37 33 37
use M2M3_PR  M2M3_PR_16
timestamp 1655484843
transform 1 0 15318 0 1 12944
box -33 -37 33 37
use M2M3_PR  M2M3_PR_17
timestamp 1655484843
transform 1 0 14582 0 1 13676
box -33 -37 33 37
use M2M3_PR  M2M3_PR_18
timestamp 1655484843
transform 1 0 22034 0 1 13188
box -33 -37 33 37
use M2M3_PR  M2M3_PR_19
timestamp 1655484843
transform 1 0 21298 0 1 13188
box -33 -37 33 37
use M2M3_PR  M2M3_PR_20
timestamp 1655484843
transform 1 0 20838 0 1 13188
box -33 -37 33 37
use M2M3_PR  M2M3_PR_21
timestamp 1655484843
transform 1 0 20102 0 1 16360
box -33 -37 33 37
use M2M3_PR  M2M3_PR_22
timestamp 1655484843
transform 1 0 16698 0 1 16360
box -33 -37 33 37
use M2M3_PR  M2M3_PR_23
timestamp 1655484843
transform 1 0 18814 0 1 13188
box -33 -37 33 37
use M2M3_PR  M2M3_PR_24
timestamp 1655484843
transform 1 0 17526 0 1 13188
box -33 -37 33 37
use M2M3_PR  M2M3_PR_25
timestamp 1655484843
transform 1 0 15502 0 1 13188
box -33 -37 33 37
use M2M3_PR  M2M3_PR_26
timestamp 1655484843
transform 1 0 15502 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_27
timestamp 1655484843
transform 1 0 14030 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_28
timestamp 1655484843
transform 1 0 18538 0 1 10626
box -33 -37 33 37
use M2M3_PR  M2M3_PR_29
timestamp 1655484843
transform 1 0 16882 0 1 10626
box -33 -37 33 37
use M2M3_PR  M2M3_PR_30
timestamp 1655484843
transform 1 0 21482 0 1 15140
box -33 -37 33 37
use M2M3_PR  M2M3_PR_31
timestamp 1655484843
transform 1 0 18538 0 1 15140
box -33 -37 33 37
use M2M3_PR  M2M3_PR_32
timestamp 1655484843
transform 1 0 17986 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_33
timestamp 1655484843
transform 1 0 16238 0 1 14652
box -33 -37 33 37
use M2M3_PR  M2M3_PR_34
timestamp 1655484843
transform 1 0 7498 0 1 15994
box -33 -37 33 37
use M2M3_PR  M2M3_PR_35
timestamp 1655484843
transform 1 0 7130 0 1 15994
box -33 -37 33 37
use M2M3_PR  M2M3_PR_36
timestamp 1655484843
transform 1 0 19182 0 1 9650
box -33 -37 33 37
use M2M3_PR  M2M3_PR_37
timestamp 1655484843
transform 1 0 17158 0 1 7942
box -33 -37 33 37
use M2M3_PR  M2M3_PR_38
timestamp 1655484843
transform 1 0 16330 0 1 9650
box -33 -37 33 37
use M2M3_PR  M2M3_PR_39
timestamp 1655484843
transform 1 0 18722 0 1 8796
box -33 -37 33 37
use M2M3_PR  M2M3_PR_40
timestamp 1655484843
transform 1 0 16054 0 1 8796
box -33 -37 33 37
use M2M3_PR  M2M3_PR_41
timestamp 1655484843
transform 1 0 15502 0 1 8796
box -33 -37 33 37
use M2M3_PR  M2M3_PR_42
timestamp 1655484843
transform 1 0 13478 0 1 8796
box -33 -37 33 37
use M2M3_PR  M2M3_PR_43
timestamp 1655484843
transform 1 0 21482 0 1 9894
box -33 -37 33 37
use M2M3_PR  M2M3_PR_44
timestamp 1655484843
transform 1 0 18078 0 1 9894
box -33 -37 33 37
use M2M3_PR  M2M3_PR_45
timestamp 1655484843
transform 1 0 19826 0 1 17824
box -33 -37 33 37
use M2M3_PR  M2M3_PR_46
timestamp 1655484843
transform 1 0 17710 0 1 17824
box -33 -37 33 37
use M2M3_PR  M2M3_PR_47
timestamp 1655484843
transform 1 0 21666 0 1 6478
box -33 -37 33 37
use M2M3_PR  M2M3_PR_48
timestamp 1655484843
transform 1 0 18814 0 1 6478
box -33 -37 33 37
use M2M3_PR  M2M3_PR_49
timestamp 1655484843
transform 1 0 20194 0 1 9284
box -33 -37 33 37
use M2M3_PR  M2M3_PR_50
timestamp 1655484843
transform 1 0 15686 0 1 9406
box -33 -37 33 37
use M2M3_PR  M2M3_PR_51
timestamp 1655484843
transform 1 0 13294 0 1 5990
box -33 -37 33 37
use M2M3_PR  M2M3_PR_52
timestamp 1655484843
transform 1 0 12282 0 1 5990
box -33 -37 33 37
use M2M3_PR  M2M3_PR_53
timestamp 1655484843
transform 1 0 22494 0 1 6234
box -33 -37 33 37
use M2M3_PR  M2M3_PR_54
timestamp 1655484843
transform 1 0 16882 0 1 5990
box -33 -37 33 37
use M2M3_PR  M2M3_PR_55
timestamp 1655484843
transform 1 0 20286 0 1 8552
box -33 -37 33 37
use M2M3_PR  M2M3_PR_56
timestamp 1655484843
transform 1 0 17066 0 1 8552
box -33 -37 33 37
use M2M3_PR  M2M3_PR_57
timestamp 1655484843
transform 1 0 16238 0 1 8552
box -33 -37 33 37
use M2M3_PR  M2M3_PR_58
timestamp 1655484843
transform 1 0 22126 0 1 14286
box -33 -37 33 37
use M2M3_PR  M2M3_PR_59
timestamp 1655484843
transform 1 0 21298 0 1 14286
box -33 -37 33 37
use M2M3_PR  M2M3_PR_60
timestamp 1655484843
transform 1 0 21298 0 1 16360
box -33 -37 33 37
use M2M3_PR  M2M3_PR_61
timestamp 1655484843
transform 1 0 21298 0 1 8308
box -33 -37 33 37
use M2M3_PR  M2M3_PR_62
timestamp 1655484843
transform 1 0 21206 0 1 11968
box -33 -37 33 37
use M2M3_PR  M2M3_PR_63
timestamp 1655484843
transform 1 0 22770 0 1 21850
box -33 -37 33 37
use M2M3_PR  M2M3_PR_64
timestamp 1655484843
transform 1 0 20378 0 1 21850
box -33 -37 33 37
use M2M3_PR  M2M3_PR_65
timestamp 1655484843
transform 1 0 14858 0 1 17458
box -33 -37 33 37
use M2M3_PR  M2M3_PR_66
timestamp 1655484843
transform 1 0 14306 0 1 17458
box -33 -37 33 37
use M2M3_PR  M2M3_PR_67
timestamp 1655484843
transform 1 0 22126 0 1 19166
box -33 -37 33 37
use M2M3_PR  M2M3_PR_68
timestamp 1655484843
transform 1 0 16882 0 1 19166
box -33 -37 33 37
use M2M3_PR  M2M3_PR_69
timestamp 1655484843
transform 1 0 18170 0 1 10138
box -33 -37 33 37
use M2M3_PR  M2M3_PR_70
timestamp 1655484843
transform 1 0 10074 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_71
timestamp 1655484843
transform 1 0 10718 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_72
timestamp 1655484843
transform 1 0 10258 0 1 6600
box -33 -37 33 37
use M2M3_PR  M2M3_PR_73
timestamp 1655484843
transform 1 0 9522 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_74
timestamp 1655484843
transform 1 0 8694 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_75
timestamp 1655484843
transform 1 0 8234 0 1 6356
box -33 -37 33 37
use M2M3_PR  M2M3_PR_76
timestamp 1655484843
transform 1 0 7314 0 1 15750
box -33 -37 33 37
use M2M3_PR  M2M3_PR_77
timestamp 1655484843
transform 1 0 7314 0 1 6600
box -33 -37 33 37
use M2M3_PR  M2M3_PR_78
timestamp 1655484843
transform 1 0 21390 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_79
timestamp 1655484843
transform 1 0 19826 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_80
timestamp 1655484843
transform 1 0 19274 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_81
timestamp 1655484843
transform 1 0 18814 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_82
timestamp 1655484843
transform 1 0 16238 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_83
timestamp 1655484843
transform 1 0 14674 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_84
timestamp 1655484843
transform 1 0 13662 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_85
timestamp 1655484843
transform 1 0 13294 0 1 12578
box -33 -37 33 37
use M2M3_PR  M2M3_PR_86
timestamp 1655484843
transform 1 0 12374 0 1 12578
box -33 -37 33 37
use M2M3_PR  M2M3_PR_87
timestamp 1655484843
transform 1 0 12374 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_88
timestamp 1655484843
transform 1 0 10718 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_89
timestamp 1655484843
transform 1 0 9154 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_90
timestamp 1655484843
transform 1 0 22770 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_91
timestamp 1655484843
transform 1 0 22770 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_92
timestamp 1655484843
transform 1 0 21114 0 1 12456
box -33 -37 33 37
use M2M3_PR  M2M3_PR_93
timestamp 1655484843
transform 1 0 20102 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_94
timestamp 1655484843
transform 1 0 19182 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_95
timestamp 1655484843
transform 1 0 15962 0 1 20142
box -33 -37 33 37
use M2M3_PR  M2M3_PR_96
timestamp 1655484843
transform 1 0 20194 0 1 12578
box -33 -37 33 37
use M2M3_PR  M2M3_PR_97
timestamp 1655484843
transform 1 0 18630 0 1 12578
box -33 -37 33 37
use M2M3_PR  M2M3_PR_98
timestamp 1655484843
transform 1 0 18630 0 1 6966
box -33 -37 33 37
use M2M3_PR  M2M3_PR_99
timestamp 1655484843
transform 1 0 9338 0 1 6966
box -33 -37 33 37
use M2M3_PR  M2M3_PR_100
timestamp 1655484843
transform 1 0 17342 0 1 15872
box -33 -37 33 37
use M2M3_PR  M2M3_PR_101
timestamp 1655484843
transform 1 0 15778 0 1 15872
box -33 -37 33 37
use M2M3_PR  M2M3_PR_102
timestamp 1655484843
transform 1 0 15778 0 1 14164
box -33 -37 33 37
use M2M3_PR  M2M3_PR_103
timestamp 1655484843
transform 1 0 14766 0 1 14164
box -33 -37 33 37
use M2M3_PR  M2M3_PR_104
timestamp 1655484843
transform 1 0 10626 0 1 14774
box -33 -37 33 37
use M2M3_PR  M2M3_PR_105
timestamp 1655484843
transform 1 0 46 0 1 14774
box -33 -37 33 37
use M2M3_PR  M2M3_PR_106
timestamp 1655484843
transform 1 0 18630 0 1 27706
box -33 -37 33 37
use M2M3_PR  M2M3_PR_107
timestamp 1655484843
transform 1 0 21850 0 1 25266
box -33 -37 33 37
use M2M3_PR  M2M3_PR_108
timestamp 1655484843
transform 1 0 26450 0 1 22704
box -33 -37 33 37
use M2M3_PR  M2M3_PR_109
timestamp 1655484843
transform 1 0 19090 0 1 19654
box -33 -37 33 37
use M2M3_PR  M2M3_PR_110
timestamp 1655484843
transform 1 0 21666 0 1 17702
box -33 -37 33 37
use M2M3_PR  M2M3_PR_111
timestamp 1655484843
transform 1 0 21298 0 1 14530
box -33 -37 33 37
use M2M3_PR  M2M3_PR_112
timestamp 1655484843
transform 1 0 20470 0 1 14530
box -33 -37 33 37
use M2M3_PR  M2M3_PR_113
timestamp 1655484843
transform 1 0 22954 0 1 15262
box -33 -37 33 37
use M2M3_PR  M2M3_PR_114
timestamp 1655484843
transform 1 0 20562 0 1 12944
box -33 -37 33 37
use M2M3_PR  M2M3_PR_115
timestamp 1655484843
transform 1 0 21850 0 1 10260
box -33 -37 33 37
use M2M3_PR  M2M3_PR_116
timestamp 1655484843
transform 1 0 22034 0 1 7698
box -33 -37 33 37
use M2M3_PR  M2M3_PR_117
timestamp 1655484843
transform 1 0 23230 0 1 5258
box -33 -37 33 37
use M2M3_PR  M2M3_PR_118
timestamp 1655484843
transform 1 0 26266 0 1 2696
box -33 -37 33 37
use M2M3_PR  M2M3_PR_119
timestamp 1655484843
transform 1 0 28566 0 1 8064
box -33 -37 33 37
use M2M3_PR  M2M3_PR_120
timestamp 1655484843
transform 1 0 28566 0 1 134
box -33 -37 33 37
use M2M3_PR  M2M3_PR_121
timestamp 1655484843
transform 1 0 22770 0 1 8064
box -33 -37 33 37
use M2M3_PR  M2M3_PR_122
timestamp 1655484843
transform 1 0 20562 0 1 8064
box -33 -37 33 37
use M2M3_PR  M2M3_PR_123
timestamp 1655484843
transform 1 0 5842 0 1 13798
box -33 -37 33 37
use M2M3_PR  M2M3_PR_124
timestamp 1655484843
transform 1 0 28750 0 1 378
box -33 -37 33 37
use M2M3_PR  M2M3_PR_125
timestamp 1655484843
transform 1 0 14306 0 1 134
box -33 -37 33 37
use M3M4_PR  M3M4_PR_0
timestamp 1655484843
transform 1 0 17158 0 1 9528
box -38 -33 38 33
use M3M4_PR  M3M4_PR_1
timestamp 1655484843
transform 1 0 17158 0 1 7942
box -38 -33 38 33
use M3M4_PR  M3M4_PR_2
timestamp 1655484843
transform 1 0 21298 0 1 16360
box -38 -33 38 33
use M3M4_PR  M3M4_PR_3
timestamp 1655484843
transform 1 0 21298 0 1 11968
box -38 -33 38 33
use M3M4_PR  M3M4_PR_4
timestamp 1655484843
transform 1 0 21298 0 1 8308
box -38 -33 38 33
use digital_filter_VIA0  digital_filter_VIA0_0
timestamp 1655484843
transform 1 0 20750 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_1
timestamp 1655484843
transform 1 0 15150 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_2
timestamp 1655484843
transform 1 0 9550 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_3
timestamp 1655484843
transform 1 0 20750 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_4
timestamp 1655484843
transform 1 0 15150 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_5
timestamp 1655484843
transform 1 0 9550 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_6
timestamp 1655484843
transform 1 0 23310 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_7
timestamp 1655484843
transform 1 0 23310 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_8
timestamp 1655484843
transform 1 0 5486 0 1 22342
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_9
timestamp 1655484843
transform 1 0 5486 0 1 5402
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_10
timestamp 1655484843
transform 1 0 19510 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_11
timestamp 1655484843
transform 1 0 13910 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_12
timestamp 1655484843
transform 1 0 8310 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_13
timestamp 1655484843
transform 1 0 19510 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_14
timestamp 1655484843
transform 1 0 13910 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_15
timestamp 1655484843
transform 1 0 8310 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_16
timestamp 1655484843
transform 1 0 24550 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_17
timestamp 1655484843
transform 1 0 24550 0 1 4162
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_18
timestamp 1655484843
transform 1 0 4246 0 1 23582
box -310 -310 310 310
use digital_filter_VIA0  digital_filter_VIA0_19
timestamp 1655484843
transform 1 0 4246 0 1 4162
box -310 -310 310 310
use digital_filter_VIA1  digital_filter_VIA1_0
timestamp 1655484843
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_1
timestamp 1655484843
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_2
timestamp 1655484843
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_3
timestamp 1655484843
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_4
timestamp 1655484843
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_5
timestamp 1655484843
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_6
timestamp 1655484843
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_7
timestamp 1655484843
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_8
timestamp 1655484843
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_9
timestamp 1655484843
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_10
timestamp 1655484843
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_11
timestamp 1655484843
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_12
timestamp 1655484843
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_13
timestamp 1655484843
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_14
timestamp 1655484843
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_15
timestamp 1655484843
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_16
timestamp 1655484843
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_17
timestamp 1655484843
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_18
timestamp 1655484843
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_19
timestamp 1655484843
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_20
timestamp 1655484843
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_21
timestamp 1655484843
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_22
timestamp 1655484843
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_23
timestamp 1655484843
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_24
timestamp 1655484843
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_25
timestamp 1655484843
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_26
timestamp 1655484843
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_27
timestamp 1655484843
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_28
timestamp 1655484843
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_29
timestamp 1655484843
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_30
timestamp 1655484843
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_31
timestamp 1655484843
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_32
timestamp 1655484843
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_33
timestamp 1655484843
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_34
timestamp 1655484843
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_35
timestamp 1655484843
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_36
timestamp 1655484843
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_37
timestamp 1655484843
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_38
timestamp 1655484843
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_39
timestamp 1655484843
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_40
timestamp 1655484843
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_41
timestamp 1655484843
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_42
timestamp 1655484843
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_43
timestamp 1655484843
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_44
timestamp 1655484843
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_45
timestamp 1655484843
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_46
timestamp 1655484843
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_47
timestamp 1655484843
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_48
timestamp 1655484843
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_49
timestamp 1655484843
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_50
timestamp 1655484843
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_51
timestamp 1655484843
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_52
timestamp 1655484843
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_53
timestamp 1655484843
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_54
timestamp 1655484843
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_55
timestamp 1655484843
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_56
timestamp 1655484843
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_57
timestamp 1655484843
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_58
timestamp 1655484843
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_59
timestamp 1655484843
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_60
timestamp 1655484843
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_61
timestamp 1655484843
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_62
timestamp 1655484843
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_63
timestamp 1655484843
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_64
timestamp 1655484843
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_65
timestamp 1655484843
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_66
timestamp 1655484843
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_67
timestamp 1655484843
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_68
timestamp 1655484843
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_69
timestamp 1655484843
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_70
timestamp 1655484843
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_71
timestamp 1655484843
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_72
timestamp 1655484843
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_73
timestamp 1655484843
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_74
timestamp 1655484843
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_75
timestamp 1655484843
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_76
timestamp 1655484843
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_77
timestamp 1655484843
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_78
timestamp 1655484843
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_79
timestamp 1655484843
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_80
timestamp 1655484843
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_81
timestamp 1655484843
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_82
timestamp 1655484843
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_83
timestamp 1655484843
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_84
timestamp 1655484843
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_85
timestamp 1655484843
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_86
timestamp 1655484843
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_87
timestamp 1655484843
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_88
timestamp 1655484843
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_89
timestamp 1655484843
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_90
timestamp 1655484843
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_91
timestamp 1655484843
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA1  digital_filter_VIA1_92
timestamp 1655484843
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_0
timestamp 1655484843
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_1
timestamp 1655484843
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_2
timestamp 1655484843
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_3
timestamp 1655484843
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_4
timestamp 1655484843
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_5
timestamp 1655484843
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_6
timestamp 1655484843
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_7
timestamp 1655484843
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_8
timestamp 1655484843
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_9
timestamp 1655484843
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_10
timestamp 1655484843
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_11
timestamp 1655484843
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_12
timestamp 1655484843
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_13
timestamp 1655484843
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_14
timestamp 1655484843
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_15
timestamp 1655484843
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_16
timestamp 1655484843
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_17
timestamp 1655484843
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_18
timestamp 1655484843
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_19
timestamp 1655484843
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_20
timestamp 1655484843
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_21
timestamp 1655484843
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_22
timestamp 1655484843
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_23
timestamp 1655484843
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_24
timestamp 1655484843
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_25
timestamp 1655484843
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_26
timestamp 1655484843
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_27
timestamp 1655484843
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_28
timestamp 1655484843
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_29
timestamp 1655484843
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_30
timestamp 1655484843
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_31
timestamp 1655484843
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_32
timestamp 1655484843
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_33
timestamp 1655484843
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_34
timestamp 1655484843
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_35
timestamp 1655484843
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_36
timestamp 1655484843
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_37
timestamp 1655484843
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_38
timestamp 1655484843
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_39
timestamp 1655484843
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_40
timestamp 1655484843
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_41
timestamp 1655484843
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_42
timestamp 1655484843
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_43
timestamp 1655484843
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_44
timestamp 1655484843
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_45
timestamp 1655484843
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_46
timestamp 1655484843
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_47
timestamp 1655484843
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_48
timestamp 1655484843
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_49
timestamp 1655484843
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_50
timestamp 1655484843
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_51
timestamp 1655484843
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_52
timestamp 1655484843
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_53
timestamp 1655484843
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_54
timestamp 1655484843
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_55
timestamp 1655484843
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_56
timestamp 1655484843
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_57
timestamp 1655484843
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_58
timestamp 1655484843
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_59
timestamp 1655484843
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_60
timestamp 1655484843
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_61
timestamp 1655484843
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_62
timestamp 1655484843
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_63
timestamp 1655484843
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_64
timestamp 1655484843
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_65
timestamp 1655484843
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_66
timestamp 1655484843
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_67
timestamp 1655484843
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_68
timestamp 1655484843
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_69
timestamp 1655484843
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_70
timestamp 1655484843
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_71
timestamp 1655484843
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_72
timestamp 1655484843
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_73
timestamp 1655484843
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_74
timestamp 1655484843
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_75
timestamp 1655484843
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_76
timestamp 1655484843
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_77
timestamp 1655484843
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_78
timestamp 1655484843
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_79
timestamp 1655484843
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_80
timestamp 1655484843
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_81
timestamp 1655484843
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_82
timestamp 1655484843
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_83
timestamp 1655484843
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_84
timestamp 1655484843
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_85
timestamp 1655484843
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_86
timestamp 1655484843
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_87
timestamp 1655484843
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_88
timestamp 1655484843
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_89
timestamp 1655484843
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_90
timestamp 1655484843
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_91
timestamp 1655484843
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA2  digital_filter_VIA2_92
timestamp 1655484843
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_0
timestamp 1655484843
transform 1 0 20750 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_1
timestamp 1655484843
transform 1 0 20750 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_2
timestamp 1655484843
transform 1 0 20750 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_3
timestamp 1655484843
transform 1 0 20750 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_4
timestamp 1655484843
transform 1 0 20750 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_5
timestamp 1655484843
transform 1 0 20750 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_6
timestamp 1655484843
transform 1 0 20750 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_7
timestamp 1655484843
transform 1 0 20750 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_8
timestamp 1655484843
transform 1 0 20750 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_9
timestamp 1655484843
transform 1 0 20750 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_10
timestamp 1655484843
transform 1 0 20750 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_11
timestamp 1655484843
transform 1 0 20750 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_12
timestamp 1655484843
transform 1 0 20750 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_13
timestamp 1655484843
transform 1 0 20750 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_14
timestamp 1655484843
transform 1 0 20750 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_15
timestamp 1655484843
transform 1 0 15150 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_16
timestamp 1655484843
transform 1 0 15150 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_17
timestamp 1655484843
transform 1 0 15150 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_18
timestamp 1655484843
transform 1 0 15150 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_19
timestamp 1655484843
transform 1 0 15150 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_20
timestamp 1655484843
transform 1 0 15150 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_21
timestamp 1655484843
transform 1 0 15150 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_22
timestamp 1655484843
transform 1 0 15150 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_23
timestamp 1655484843
transform 1 0 15150 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_24
timestamp 1655484843
transform 1 0 15150 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_25
timestamp 1655484843
transform 1 0 15150 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_26
timestamp 1655484843
transform 1 0 15150 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_27
timestamp 1655484843
transform 1 0 15150 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_28
timestamp 1655484843
transform 1 0 15150 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_29
timestamp 1655484843
transform 1 0 15150 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_30
timestamp 1655484843
transform 1 0 9550 0 1 21488
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_31
timestamp 1655484843
transform 1 0 9550 0 1 20400
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_32
timestamp 1655484843
transform 1 0 9550 0 1 19312
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_33
timestamp 1655484843
transform 1 0 9550 0 1 18224
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_34
timestamp 1655484843
transform 1 0 9550 0 1 17136
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_35
timestamp 1655484843
transform 1 0 9550 0 1 16048
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_36
timestamp 1655484843
transform 1 0 9550 0 1 14960
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_37
timestamp 1655484843
transform 1 0 9550 0 1 13872
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_38
timestamp 1655484843
transform 1 0 9550 0 1 12784
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_39
timestamp 1655484843
transform 1 0 9550 0 1 11696
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_40
timestamp 1655484843
transform 1 0 9550 0 1 10608
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_41
timestamp 1655484843
transform 1 0 9550 0 1 9520
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_42
timestamp 1655484843
transform 1 0 9550 0 1 8432
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_43
timestamp 1655484843
transform 1 0 9550 0 1 7344
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_44
timestamp 1655484843
transform 1 0 9550 0 1 6256
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_45
timestamp 1655484843
transform 1 0 19510 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_46
timestamp 1655484843
transform 1 0 19510 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_47
timestamp 1655484843
transform 1 0 19510 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_48
timestamp 1655484843
transform 1 0 19510 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_49
timestamp 1655484843
transform 1 0 19510 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_50
timestamp 1655484843
transform 1 0 19510 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_51
timestamp 1655484843
transform 1 0 19510 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_52
timestamp 1655484843
transform 1 0 19510 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_53
timestamp 1655484843
transform 1 0 19510 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_54
timestamp 1655484843
transform 1 0 19510 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_55
timestamp 1655484843
transform 1 0 19510 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_56
timestamp 1655484843
transform 1 0 19510 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_57
timestamp 1655484843
transform 1 0 19510 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_58
timestamp 1655484843
transform 1 0 19510 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_59
timestamp 1655484843
transform 1 0 19510 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_60
timestamp 1655484843
transform 1 0 19510 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_61
timestamp 1655484843
transform 1 0 13910 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_62
timestamp 1655484843
transform 1 0 13910 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_63
timestamp 1655484843
transform 1 0 13910 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_64
timestamp 1655484843
transform 1 0 13910 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_65
timestamp 1655484843
transform 1 0 13910 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_66
timestamp 1655484843
transform 1 0 13910 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_67
timestamp 1655484843
transform 1 0 13910 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_68
timestamp 1655484843
transform 1 0 13910 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_69
timestamp 1655484843
transform 1 0 13910 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_70
timestamp 1655484843
transform 1 0 13910 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_71
timestamp 1655484843
transform 1 0 13910 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_72
timestamp 1655484843
transform 1 0 13910 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_73
timestamp 1655484843
transform 1 0 13910 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_74
timestamp 1655484843
transform 1 0 13910 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_75
timestamp 1655484843
transform 1 0 13910 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_76
timestamp 1655484843
transform 1 0 13910 0 1 5712
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_77
timestamp 1655484843
transform 1 0 8310 0 1 22032
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_78
timestamp 1655484843
transform 1 0 8310 0 1 20944
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_79
timestamp 1655484843
transform 1 0 8310 0 1 19856
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_80
timestamp 1655484843
transform 1 0 8310 0 1 18768
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_81
timestamp 1655484843
transform 1 0 8310 0 1 17680
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_82
timestamp 1655484843
transform 1 0 8310 0 1 16592
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_83
timestamp 1655484843
transform 1 0 8310 0 1 15504
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_84
timestamp 1655484843
transform 1 0 8310 0 1 14416
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_85
timestamp 1655484843
transform 1 0 8310 0 1 13328
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_86
timestamp 1655484843
transform 1 0 8310 0 1 12240
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_87
timestamp 1655484843
transform 1 0 8310 0 1 11152
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_88
timestamp 1655484843
transform 1 0 8310 0 1 10064
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_89
timestamp 1655484843
transform 1 0 8310 0 1 8976
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_90
timestamp 1655484843
transform 1 0 8310 0 1 7888
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_91
timestamp 1655484843
transform 1 0 8310 0 1 6800
box -310 -48 310 48
use digital_filter_VIA3  digital_filter_VIA3_92
timestamp 1655484843
transform 1 0 8310 0 1 5712
box -310 -48 310 48
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 19228 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_1
timestamp 1655484843
transform -1 0 15456 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_2
timestamp 1655484843
transform 1 0 11224 0 1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_3
timestamp 1655484843
transform 1 0 6348 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_4
timestamp 1655484843
transform 1 0 6348 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  sky130_fd_sc_hd__a21oi_1_5
timestamp 1655484843
transform -1 0 7912 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 20884 0 1 7888
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_1
timestamp 1655484843
transform -1 0 21068 0 1 11152
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_2
timestamp 1655484843
transform -1 0 20884 0 1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_3
timestamp 1655484843
transform -1 0 20884 0 1 8976
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_4
timestamp 1655484843
transform -1 0 22172 0 -1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_5
timestamp 1655484843
transform -1 0 20884 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_6
timestamp 1655484843
transform -1 0 19688 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_7
timestamp 1655484843
transform 1 0 20240 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_8
timestamp 1655484843
transform -1 0 19412 0 1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_9
timestamp 1655484843
transform 1 0 20516 0 1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_10
timestamp 1655484843
transform -1 0 19964 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_11
timestamp 1655484843
transform 1 0 17480 0 -1 18768
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_12
timestamp 1655484843
transform 1 0 15456 0 1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_13
timestamp 1655484843
transform 1 0 16652 0 -1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_14
timestamp 1655484843
transform 1 0 13708 0 1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_15
timestamp 1655484843
transform -1 0 15732 0 -1 17680
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_16
timestamp 1655484843
transform 1 0 14168 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_17
timestamp 1655484843
transform 1 0 16560 0 1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_18
timestamp 1655484843
transform 1 0 16376 0 -1 15504
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_19
timestamp 1655484843
transform 1 0 16744 0 -1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_20
timestamp 1655484843
transform -1 0 15732 0 -1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_21
timestamp 1655484843
transform 1 0 15456 0 1 11152
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_22
timestamp 1655484843
transform -1 0 14628 0 1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_23
timestamp 1655484843
transform 1 0 15272 0 -1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_24
timestamp 1655484843
transform -1 0 16836 0 1 8976
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_25
timestamp 1655484843
transform -1 0 18308 0 1 10064
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  sky130_fd_sc_hd__a22o_1_26
timestamp 1655484843
transform -1 0 18216 0 -1 12240
box -38 -48 682 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 10120 0 -1 22032
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_1
timestamp 1655484843
transform 1 0 9016 0 1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_2
timestamp 1655484843
transform -1 0 10764 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_3
timestamp 1655484843
transform 1 0 10212 0 -1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_4
timestamp 1655484843
transform -1 0 7820 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_5
timestamp 1655484843
transform -1 0 8280 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_6
timestamp 1655484843
transform 1 0 6532 0 1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_7
timestamp 1655484843
transform 1 0 6348 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_8
timestamp 1655484843
transform 1 0 8648 0 -1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_9
timestamp 1655484843
transform 1 0 6624 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_10
timestamp 1655484843
transform 1 0 17572 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_11
timestamp 1655484843
transform 1 0 18768 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_12
timestamp 1655484843
transform 1 0 15180 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_13
timestamp 1655484843
transform 1 0 12604 0 -1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_14
timestamp 1655484843
transform 1 0 12972 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_15
timestamp 1655484843
transform 1 0 11316 0 1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_16
timestamp 1655484843
transform 1 0 11408 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_17
timestamp 1655484843
transform 1 0 12880 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_18
timestamp 1655484843
transform 1 0 13800 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_19
timestamp 1655484843
transform 1 0 13616 0 1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_20
timestamp 1655484843
transform -1 0 13156 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_21
timestamp 1655484843
transform -1 0 13340 0 -1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_22
timestamp 1655484843
transform 1 0 12328 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_23
timestamp 1655484843
transform 1 0 15088 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_24
timestamp 1655484843
transform 1 0 15916 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_25
timestamp 1655484843
transform 1 0 16376 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_26
timestamp 1655484843
transform 1 0 21896 0 -1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_27
timestamp 1655484843
transform 1 0 21528 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_28
timestamp 1655484843
transform -1 0 22448 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_29
timestamp 1655484843
transform 1 0 22080 0 -1 15504
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_30
timestamp 1655484843
transform 1 0 21620 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_31
timestamp 1655484843
transform -1 0 21988 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_32
timestamp 1655484843
transform 1 0 21896 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_33
timestamp 1655484843
transform 1 0 22080 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_34
timestamp 1655484843
transform -1 0 18308 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_35
timestamp 1655484843
transform 1 0 20700 0 1 6800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_36
timestamp 1655484843
transform -1 0 22448 0 -1 14416
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_37
timestamp 1655484843
transform -1 0 12788 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_38
timestamp 1655484843
transform 1 0 12788 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_39
timestamp 1655484843
transform -1 0 12144 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_40
timestamp 1655484843
transform -1 0 11684 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_41
timestamp 1655484843
transform 1 0 8832 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_42
timestamp 1655484843
transform 1 0 9936 0 -1 10064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_43
timestamp 1655484843
transform 1 0 8924 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_44
timestamp 1655484843
transform -1 0 10304 0 -1 12240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_45
timestamp 1655484843
transform -1 0 10488 0 -1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_46
timestamp 1655484843
transform 1 0 9752 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_47
timestamp 1655484843
transform 1 0 9200 0 -1 16592
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_48
timestamp 1655484843
transform 1 0 10488 0 1 18768
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_49
timestamp 1655484843
transform -1 0 11868 0 1 17680
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_50
timestamp 1655484843
transform -1 0 13248 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_51
timestamp 1655484843
transform -1 0 15364 0 -1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_52
timestamp 1655484843
transform -1 0 16652 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_53
timestamp 1655484843
transform -1 0 19320 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_54
timestamp 1655484843
transform -1 0 19780 0 1 20944
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_55
timestamp 1655484843
transform 1 0 19504 0 -1 22032
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_56
timestamp 1655484843
transform 1 0 6440 0 -1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_57
timestamp 1655484843
transform 1 0 6532 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_58
timestamp 1655484843
transform 1 0 7820 0 1 5712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_59
timestamp 1655484843
transform 1 0 6348 0 1 7888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_60
timestamp 1655484843
transform 1 0 6440 0 1 8976
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_61
timestamp 1655484843
transform 1 0 6624 0 -1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_62
timestamp 1655484843
transform 1 0 6440 0 1 11152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_63
timestamp 1655484843
transform 1 0 7268 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_64
timestamp 1655484843
transform 1 0 6256 0 1 13328
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 13340 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1655484843
transform 1 0 13616 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1655484843
transform 1 0 10028 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1655484843
transform -1 0 12052 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1655484843
transform 1 0 11684 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1655484843
transform 1 0 15824 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1655484843
transform 1 0 18032 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_7
timestamp 1655484843
transform 1 0 6440 0 1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_8
timestamp 1655484843
transform 1 0 10488 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_9
timestamp 1655484843
transform -1 0 7084 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_10
timestamp 1655484843
transform -1 0 7176 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 13984 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 18032 0 1 13328
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1655484843
transform 1 0 17940 0 1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 13892 0 1 7888
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_1
timestamp 1655484843
transform -1 0 18676 0 -1 6800
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_2
timestamp 1655484843
transform 1 0 9200 0 1 6800
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_3
timestamp 1655484843
transform 1 0 18768 0 -1 7888
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_4
timestamp 1655484843
transform 1 0 20056 0 1 12240
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 17848 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_1
timestamp 1655484843
transform 1 0 14536 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 22632 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1655484843
transform 1 0 22632 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1655484843
transform 1 0 22632 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_3
timestamp 1655484843
transform 1 0 22632 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_4
timestamp 1655484843
transform 1 0 22632 0 -1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_5
timestamp 1655484843
transform 1 0 22632 0 -1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_6
timestamp 1655484843
transform 1 0 22632 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_7
timestamp 1655484843
transform 1 0 22632 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_8
timestamp 1655484843
transform 1 0 22632 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_9
timestamp 1655484843
transform 1 0 22632 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_10
timestamp 1655484843
transform 1 0 22632 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_11
timestamp 1655484843
transform 1 0 22632 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_12
timestamp 1655484843
transform 1 0 22632 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_13
timestamp 1655484843
transform 1 0 22632 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_14
timestamp 1655484843
transform 1 0 22632 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_15
timestamp 1655484843
transform 1 0 21344 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_16
timestamp 1655484843
transform 1 0 20056 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_17
timestamp 1655484843
transform 1 0 19688 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_18
timestamp 1655484843
transform 1 0 19228 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_19
timestamp 1655484843
transform 1 0 18952 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_20
timestamp 1655484843
transform 1 0 18492 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_21
timestamp 1655484843
transform 1 0 18216 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_22
timestamp 1655484843
transform 1 0 17664 0 1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_23
timestamp 1655484843
transform 1 0 17480 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_24
timestamp 1655484843
transform 1 0 17480 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_25
timestamp 1655484843
transform 1 0 17480 0 -1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_26
timestamp 1655484843
transform 1 0 17480 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_27
timestamp 1655484843
transform 1 0 17480 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_28
timestamp 1655484843
transform 1 0 16928 0 1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_29
timestamp 1655484843
transform 1 0 16928 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_30
timestamp 1655484843
transform 1 0 16192 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_31
timestamp 1655484843
transform 1 0 16376 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_32
timestamp 1655484843
transform 1 0 15824 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_33
timestamp 1655484843
transform 1 0 14904 0 -1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_34
timestamp 1655484843
transform 1 0 14904 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_35
timestamp 1655484843
transform 1 0 14904 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_36
timestamp 1655484843
transform 1 0 14536 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_37
timestamp 1655484843
transform 1 0 14260 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_38
timestamp 1655484843
transform 1 0 13800 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_39
timestamp 1655484843
transform 1 0 13800 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_40
timestamp 1655484843
transform 1 0 13800 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_41
timestamp 1655484843
transform 1 0 12328 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_42
timestamp 1655484843
transform 1 0 12328 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_43
timestamp 1655484843
transform 1 0 11776 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_44
timestamp 1655484843
transform 1 0 11040 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_45
timestamp 1655484843
transform 1 0 11224 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_46
timestamp 1655484843
transform 1 0 11040 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_47
timestamp 1655484843
transform 1 0 11040 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_48
timestamp 1655484843
transform 1 0 10764 0 -1 19856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_49
timestamp 1655484843
transform 1 0 10672 0 1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_50
timestamp 1655484843
transform 1 0 10672 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_51
timestamp 1655484843
transform 1 0 10304 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_52
timestamp 1655484843
transform 1 0 9752 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_53
timestamp 1655484843
transform 1 0 9752 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_54
timestamp 1655484843
transform 1 0 9384 0 -1 11152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_55
timestamp 1655484843
transform 1 0 9384 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_56
timestamp 1655484843
transform 1 0 8464 0 1 16592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_57
timestamp 1655484843
transform 1 0 8096 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_58
timestamp 1655484843
transform 1 0 8096 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_59
timestamp 1655484843
transform 1 0 8096 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_60
timestamp 1655484843
transform 1 0 7176 0 -1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_61
timestamp 1655484843
transform 1 0 6808 0 -1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_62
timestamp 1655484843
transform 1 0 6808 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_63
timestamp 1655484843
transform 1 0 6624 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_64
timestamp 1655484843
transform 1 0 5888 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_65
timestamp 1655484843
transform 1 0 5888 0 1 14416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 22540 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1655484843
transform 1 0 22172 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1655484843
transform 1 0 21620 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1655484843
transform 1 0 21620 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1655484843
transform 1 0 21528 0 -1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1655484843
transform 1 0 20884 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1655484843
transform 1 0 19688 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1655484843
transform 1 0 19596 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1655484843
transform 1 0 18308 0 1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1655484843
transform 1 0 18308 0 1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_10
timestamp 1655484843
transform 1 0 18308 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_11
timestamp 1655484843
transform 1 0 17756 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_12
timestamp 1655484843
transform 1 0 17480 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_13
timestamp 1655484843
transform 1 0 17664 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_14
timestamp 1655484843
transform 1 0 17020 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_15
timestamp 1655484843
transform 1 0 17020 0 -1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_16
timestamp 1655484843
transform 1 0 17020 0 -1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_17
timestamp 1655484843
transform 1 0 16652 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_18
timestamp 1655484843
transform 1 0 16284 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_19
timestamp 1655484843
transform 1 0 16192 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_20
timestamp 1655484843
transform 1 0 15640 0 1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_21
timestamp 1655484843
transform 1 0 14904 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_22
timestamp 1655484843
transform 1 0 14444 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_23
timestamp 1655484843
transform 1 0 14444 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_24
timestamp 1655484843
transform 1 0 14168 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_25
timestamp 1655484843
transform 1 0 14076 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_26
timestamp 1655484843
transform 1 0 13800 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_27
timestamp 1655484843
transform 1 0 13616 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_28
timestamp 1655484843
transform 1 0 13616 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_29
timestamp 1655484843
transform 1 0 13616 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_30
timestamp 1655484843
transform 1 0 13064 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_31
timestamp 1655484843
transform 1 0 12696 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_32
timestamp 1655484843
transform 1 0 12328 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_33
timestamp 1655484843
transform 1 0 12328 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_34
timestamp 1655484843
transform 1 0 12328 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_35
timestamp 1655484843
transform 1 0 12328 0 -1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_36
timestamp 1655484843
transform 1 0 11868 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_37
timestamp 1655484843
transform 1 0 11684 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_38
timestamp 1655484843
transform 1 0 11316 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_39
timestamp 1655484843
transform 1 0 11040 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_40
timestamp 1655484843
transform 1 0 11040 0 1 11152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_41
timestamp 1655484843
transform 1 0 11132 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_42
timestamp 1655484843
transform 1 0 10580 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_43
timestamp 1655484843
transform 1 0 10580 0 1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_44
timestamp 1655484843
transform 1 0 9752 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_45
timestamp 1655484843
transform 1 0 9844 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_46
timestamp 1655484843
transform 1 0 9292 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_47
timestamp 1655484843
transform 1 0 9292 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_48
timestamp 1655484843
transform 1 0 9292 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_49
timestamp 1655484843
transform 1 0 8832 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_50
timestamp 1655484843
transform 1 0 8740 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_51
timestamp 1655484843
transform 1 0 8464 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_52
timestamp 1655484843
transform 1 0 8464 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_53
timestamp 1655484843
transform 1 0 8464 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_54
timestamp 1655484843
transform 1 0 7728 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_55
timestamp 1655484843
transform 1 0 7360 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_56
timestamp 1655484843
transform 1 0 6716 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_57
timestamp 1655484843
transform 1 0 6624 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_58
timestamp 1655484843
transform 1 0 6256 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_59
timestamp 1655484843
transform 1 0 5888 0 -1 22032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_60
timestamp 1655484843
transform 1 0 5796 0 -1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_61
timestamp 1655484843
transform 1 0 5888 0 1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_62
timestamp 1655484843
transform 1 0 5888 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_63
timestamp 1655484843
transform 1 0 5888 0 1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 21988 0 -1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1655484843
transform 1 0 21988 0 -1 12240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1655484843
transform 1 0 18124 0 1 17680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1655484843
transform 1 0 18124 0 1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1655484843
transform 1 0 18124 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1655484843
transform 1 0 17940 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1655484843
transform 1 0 16836 0 -1 14416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1655484843
transform 1 0 16192 0 1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1655484843
transform 1 0 16284 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1655484843
transform 1 0 14904 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1655484843
transform 1 0 14260 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_11
timestamp 1655484843
transform 1 0 14352 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_12
timestamp 1655484843
transform 1 0 13616 0 1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_13
timestamp 1655484843
transform 1 0 12328 0 -1 17680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_14
timestamp 1655484843
transform 1 0 12512 0 1 7888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_15
timestamp 1655484843
transform 1 0 10396 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_16
timestamp 1655484843
transform 1 0 10396 0 1 12240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_17
timestamp 1655484843
transform 1 0 10396 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_18
timestamp 1655484843
transform 1 0 9752 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_19
timestamp 1655484843
transform 1 0 9844 0 -1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_20
timestamp 1655484843
transform 1 0 9108 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_21
timestamp 1655484843
transform 1 0 8556 0 1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_22
timestamp 1655484843
transform 1 0 8556 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_23
timestamp 1655484843
transform 1 0 8556 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_24
timestamp 1655484843
transform 1 0 8556 0 1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_25
timestamp 1655484843
transform 1 0 8556 0 1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_26
timestamp 1655484843
transform 1 0 8556 0 1 7888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_27
timestamp 1655484843
transform 1 0 8556 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_28
timestamp 1655484843
transform 1 0 7820 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_29
timestamp 1655484843
transform 1 0 7268 0 -1 19856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_30
timestamp 1655484843
transform 1 0 7268 0 -1 14416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_31
timestamp 1655484843
transform 1 0 7176 0 -1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_32
timestamp 1655484843
transform 1 0 7452 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_33
timestamp 1655484843
transform 1 0 6808 0 1 17680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_34
timestamp 1655484843
transform 1 0 5888 0 1 11152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_35
timestamp 1655484843
transform 1 0 5888 0 1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_36
timestamp 1655484843
transform 1 0 5796 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_37
timestamp 1655484843
transform 1 0 5980 0 1 5712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 21804 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1655484843
transform 1 0 20424 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1655484843
transform 1 0 20332 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1655484843
transform 1 0 20332 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1655484843
transform 1 0 19228 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1655484843
transform 1 0 19228 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1655484843
transform 1 0 19228 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1655484843
transform 1 0 18860 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1655484843
transform 1 0 18860 0 1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1655484843
transform 1 0 18860 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1655484843
transform 1 0 18860 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_11
timestamp 1655484843
transform 1 0 18124 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_12
timestamp 1655484843
transform 1 0 17756 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_13
timestamp 1655484843
transform 1 0 17756 0 -1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_14
timestamp 1655484843
transform 1 0 17572 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_15
timestamp 1655484843
transform 1 0 17756 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_16
timestamp 1655484843
transform 1 0 16652 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_17
timestamp 1655484843
transform 1 0 16652 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_18
timestamp 1655484843
transform 1 0 16652 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_19
timestamp 1655484843
transform 1 0 16192 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_20
timestamp 1655484843
transform 1 0 16192 0 1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_21
timestamp 1655484843
transform 1 0 15732 0 -1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_22
timestamp 1655484843
transform 1 0 15364 0 1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_23
timestamp 1655484843
transform 1 0 15180 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_24
timestamp 1655484843
transform 1 0 15180 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_25
timestamp 1655484843
transform 1 0 15180 0 1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_26
timestamp 1655484843
transform 1 0 14996 0 -1 7888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_27
timestamp 1655484843
transform 1 0 14076 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_28
timestamp 1655484843
transform 1 0 14076 0 -1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_29
timestamp 1655484843
transform 1 0 14076 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_30
timestamp 1655484843
transform 1 0 13616 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_31
timestamp 1655484843
transform 1 0 13616 0 1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_32
timestamp 1655484843
transform 1 0 12788 0 1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_33
timestamp 1655484843
transform 1 0 12604 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_34
timestamp 1655484843
transform 1 0 12420 0 -1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_35
timestamp 1655484843
transform 1 0 12604 0 1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_36
timestamp 1655484843
transform 1 0 12604 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_37
timestamp 1655484843
transform 1 0 12604 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_38
timestamp 1655484843
transform 1 0 12052 0 1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_39
timestamp 1655484843
transform 1 0 11500 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_40
timestamp 1655484843
transform 1 0 11040 0 1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_41
timestamp 1655484843
transform 1 0 11040 0 -1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_42
timestamp 1655484843
transform 1 0 11040 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_43
timestamp 1655484843
transform 1 0 11040 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_44
timestamp 1655484843
transform 1 0 9936 0 -1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_45
timestamp 1655484843
transform 1 0 9936 0 -1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_46
timestamp 1655484843
transform 1 0 9752 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_47
timestamp 1655484843
transform 1 0 9844 0 -1 6800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_48
timestamp 1655484843
transform 1 0 8924 0 -1 20944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_49
timestamp 1655484843
transform 1 0 8648 0 1 18768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_50
timestamp 1655484843
transform 1 0 8832 0 1 17680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_51
timestamp 1655484843
transform 1 0 8740 0 1 16592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_52
timestamp 1655484843
transform 1 0 8924 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_53
timestamp 1655484843
transform 1 0 8924 0 -1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_54
timestamp 1655484843
transform 1 0 8924 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_55
timestamp 1655484843
transform 1 0 7360 0 1 12240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_56
timestamp 1655484843
transform 1 0 7360 0 1 10064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_57
timestamp 1655484843
transform 1 0 6072 0 1 19856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_58
timestamp 1655484843
transform 1 0 6164 0 1 15504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_59
timestamp 1655484843
transform 1 0 6164 0 1 14416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_60
timestamp 1655484843
transform 1 0 5796 0 -1 13328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_61
timestamp 1655484843
transform 1 0 5796 0 -1 11152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 21620 0 1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1655484843
transform 1 0 14904 0 1 13328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1655484843
transform 1 0 14904 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1655484843
transform 1 0 8648 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1655484843
transform 1 0 7084 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1655484843
transform 1 0 7084 0 1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1655484843
transform 1 0 7084 0 1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1655484843
transform 1 0 5980 0 1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1655484843
transform 1 0 5980 0 -1 20944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1655484843
transform 1 0 5980 0 -1 19856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1655484843
transform 1 0 5980 0 1 16592
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 12512 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_1
timestamp 1655484843
transform 1 0 18768 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_2
timestamp 1655484843
transform -1 0 11224 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_3
timestamp 1655484843
transform -1 0 18676 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_4
timestamp 1655484843
transform 1 0 18768 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_5
timestamp 1655484843
transform 1 0 18308 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_6
timestamp 1655484843
transform 1 0 20056 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_7
timestamp 1655484843
transform 1 0 18492 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_8
timestamp 1655484843
transform 1 0 18768 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_9
timestamp 1655484843
transform 1 0 18768 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_10
timestamp 1655484843
transform -1 0 21528 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_11
timestamp 1655484843
transform 1 0 18492 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_12
timestamp 1655484843
transform -1 0 21160 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_13
timestamp 1655484843
transform 1 0 18492 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_14
timestamp 1655484843
transform 1 0 18768 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_15
timestamp 1655484843
transform 1 0 16192 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_16
timestamp 1655484843
transform -1 0 18216 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_17
timestamp 1655484843
transform 1 0 15088 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_18
timestamp 1655484843
transform -1 0 14812 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_19
timestamp 1655484843
transform -1 0 18952 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_20
timestamp 1655484843
transform -1 0 17664 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_21
timestamp 1655484843
transform -1 0 18952 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_22
timestamp 1655484843
transform -1 0 17388 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_23
timestamp 1655484843
transform 1 0 14904 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_24
timestamp 1655484843
transform -1 0 17664 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_25
timestamp 1655484843
transform 1 0 13984 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_26
timestamp 1655484843
transform -1 0 16652 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_27
timestamp 1655484843
transform -1 0 16100 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_28
timestamp 1655484843
transform -1 0 18308 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_29
timestamp 1655484843
transform 1 0 16836 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_30
timestamp 1655484843
transform 1 0 13616 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_31
timestamp 1655484843
transform 1 0 12328 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_32
timestamp 1655484843
transform 1 0 15916 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_33
timestamp 1655484843
transform -1 0 18676 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_34
timestamp 1655484843
transform 1 0 15456 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_35
timestamp 1655484843
transform 1 0 13340 0 -1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_36
timestamp 1655484843
transform 1 0 13616 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_37
timestamp 1655484843
transform 1 0 13340 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_38
timestamp 1655484843
transform 1 0 13340 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_39
timestamp 1655484843
transform 1 0 13616 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_40
timestamp 1655484843
transform 1 0 14904 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_41
timestamp 1655484843
transform 1 0 14444 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_42
timestamp 1655484843
transform 1 0 14352 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_43
timestamp 1655484843
transform 1 0 13340 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_44
timestamp 1655484843
transform 1 0 13984 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_45
timestamp 1655484843
transform 1 0 14352 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_46
timestamp 1655484843
transform -1 0 17388 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_47
timestamp 1655484843
transform 1 0 17204 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_48
timestamp 1655484843
transform 1 0 20056 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_49
timestamp 1655484843
transform 1 0 19780 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_50
timestamp 1655484843
transform 1 0 17848 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_51
timestamp 1655484843
transform 1 0 20056 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_52
timestamp 1655484843
transform -1 0 21620 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_53
timestamp 1655484843
transform -1 0 21528 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_54
timestamp 1655484843
transform -1 0 21528 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_55
timestamp 1655484843
transform 1 0 18768 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_56
timestamp 1655484843
transform 1 0 21344 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_57
timestamp 1655484843
transform -1 0 21528 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_58
timestamp 1655484843
transform 1 0 21344 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_59
timestamp 1655484843
transform -1 0 12236 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_60
timestamp 1655484843
transform -1 0 11224 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_61
timestamp 1655484843
transform -1 0 10580 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_62
timestamp 1655484843
transform -1 0 10948 0 1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_63
timestamp 1655484843
transform 1 0 6900 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_64
timestamp 1655484843
transform 1 0 7268 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_65
timestamp 1655484843
transform 1 0 6808 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_66
timestamp 1655484843
transform 1 0 7176 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_67
timestamp 1655484843
transform -1 0 8648 0 -1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_68
timestamp 1655484843
transform 1 0 7360 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_69
timestamp 1655484843
transform 1 0 21344 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_70
timestamp 1655484843
transform 1 0 19228 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_71
timestamp 1655484843
transform 1 0 16192 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_72
timestamp 1655484843
transform 1 0 12328 0 -1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_73
timestamp 1655484843
transform -1 0 12972 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_74
timestamp 1655484843
transform 1 0 12052 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_75
timestamp 1655484843
transform 1 0 12052 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_76
timestamp 1655484843
transform -1 0 13340 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_77
timestamp 1655484843
transform 1 0 12788 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_78
timestamp 1655484843
transform 1 0 12696 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_79
timestamp 1655484843
transform 1 0 12052 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_80
timestamp 1655484843
transform 1 0 10764 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_81
timestamp 1655484843
transform 1 0 12788 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_82
timestamp 1655484843
transform -1 0 15824 0 1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_83
timestamp 1655484843
transform 1 0 16192 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_84
timestamp 1655484843
transform -1 0 20240 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_85
timestamp 1655484843
transform -1 0 23000 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_86
timestamp 1655484843
transform -1 0 22816 0 1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_87
timestamp 1655484843
transform -1 0 22540 0 -1 17680
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_88
timestamp 1655484843
transform -1 0 22816 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_89
timestamp 1655484843
transform -1 0 22540 0 -1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_90
timestamp 1655484843
transform 1 0 21344 0 1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_91
timestamp 1655484843
transform -1 0 22908 0 1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_92
timestamp 1655484843
transform -1 0 22816 0 1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_93
timestamp 1655484843
transform 1 0 18768 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_94
timestamp 1655484843
transform -1 0 22816 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_95
timestamp 1655484843
transform -1 0 22816 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_96
timestamp 1655484843
transform 1 0 20056 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_97
timestamp 1655484843
transform 1 0 19780 0 1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_98
timestamp 1655484843
transform -1 0 19228 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_99
timestamp 1655484843
transform 1 0 15916 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_100
timestamp 1655484843
transform -1 0 15640 0 1 19856
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_101
timestamp 1655484843
transform 1 0 12328 0 -1 20944
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_102
timestamp 1655484843
transform 1 0 10672 0 -1 18768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_103
timestamp 1655484843
transform 1 0 10304 0 -1 16592
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_104
timestamp 1655484843
transform 1 0 9476 0 1 15504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_105
timestamp 1655484843
transform -1 0 12512 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_106
timestamp 1655484843
transform 1 0 7268 0 -1 13328
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_107
timestamp 1655484843
transform 1 0 7452 0 -1 12240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_108
timestamp 1655484843
transform 1 0 9200 0 1 10064
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_109
timestamp 1655484843
transform 1 0 9292 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_110
timestamp 1655484843
transform 1 0 9292 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_111
timestamp 1655484843
transform 1 0 11040 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_112
timestamp 1655484843
transform 1 0 12328 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_113
timestamp 1655484843
transform 1 0 14904 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_114
timestamp 1655484843
transform 1 0 7820 0 -1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_115
timestamp 1655484843
transform 1 0 6900 0 1 14416
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_116
timestamp 1655484843
transform 1 0 6900 0 1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_117
timestamp 1655484843
transform 1 0 7268 0 -1 11152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_118
timestamp 1655484843
transform 1 0 6900 0 1 8976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_119
timestamp 1655484843
transform 1 0 6900 0 1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_120
timestamp 1655484843
transform 1 0 8188 0 -1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_121
timestamp 1655484843
transform 1 0 6900 0 1 6800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  sky130_fd_sc_hd__dfxtp_1_122
timestamp 1655484843
transform 1 0 7176 0 -1 7888
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 21344 0 1 20944
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_1
timestamp 1655484843
transform -1 0 21252 0 1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_2
timestamp 1655484843
transform -1 0 19228 0 -1 19856
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_3
timestamp 1655484843
transform -1 0 16100 0 1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_4
timestamp 1655484843
transform -1 0 14076 0 -1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_5
timestamp 1655484843
transform -1 0 13524 0 1 18768
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_6
timestamp 1655484843
transform 1 0 11868 0 1 17680
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_7
timestamp 1655484843
transform 1 0 11868 0 1 16592
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_8
timestamp 1655484843
transform -1 0 12236 0 -1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_9
timestamp 1655484843
transform 1 0 11132 0 1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_10
timestamp 1655484843
transform 1 0 10580 0 -1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_11
timestamp 1655484843
transform 1 0 10580 0 -1 12240
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_12
timestamp 1655484843
transform 1 0 10396 0 -1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_13
timestamp 1655484843
transform 1 0 10580 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_14
timestamp 1655484843
transform 1 0 10488 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_15
timestamp 1655484843
transform 1 0 20056 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_16
timestamp 1655484843
transform 1 0 20056 0 -1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_17
timestamp 1655484843
transform -1 0 10488 0 1 14416
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_18
timestamp 1655484843
transform 1 0 9200 0 1 13328
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_19
timestamp 1655484843
transform 1 0 8648 0 1 12240
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_20
timestamp 1655484843
transform -1 0 10764 0 1 11152
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_21
timestamp 1655484843
transform -1 0 9384 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_22
timestamp 1655484843
transform -1 0 9660 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_23
timestamp 1655484843
transform 1 0 10580 0 -1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fa_2  sky130_fd_sc_hd__fa_2_24
timestamp 1655484843
transform 1 0 11040 0 1 6800
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 18124 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1655484843
transform 1 0 16192 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1655484843
transform 1 0 12052 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1655484843
transform 1 0 9200 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1655484843
transform 1 0 10304 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1655484843
transform 1 0 8188 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1655484843
transform 1 0 5888 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1655484843
transform 1 0 22908 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1655484843
transform 1 0 18492 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1655484843
transform 1 0 17664 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1655484843
transform 1 0 13340 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1655484843
transform 1 0 12512 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1655484843
transform 1 0 8464 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1655484843
transform 1 0 22908 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1655484843
transform 1 0 7176 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1655484843
transform 1 0 18768 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1655484843
transform 1 0 8188 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1655484843
transform 1 0 6992 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1655484843
transform 1 0 22908 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1655484843
transform 1 0 19596 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1655484843
transform 1 0 18768 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1655484843
transform 1 0 18032 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1655484843
transform 1 0 22908 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1655484843
transform 1 0 20240 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1655484843
transform 1 0 9752 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1655484843
transform 1 0 8648 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1655484843
transform 1 0 22724 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1655484843
transform 1 0 18216 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1655484843
transform 1 0 8188 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1655484843
transform 1 0 5888 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1655484843
transform 1 0 22908 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1655484843
transform 1 0 21528 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1655484843
transform 1 0 22908 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1655484843
transform 1 0 17848 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1655484843
transform 1 0 12328 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1655484843
transform 1 0 13340 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1655484843
transform 1 0 12512 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_37
timestamp 1655484843
transform 1 0 22908 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_38
timestamp 1655484843
transform 1 0 7176 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_39
timestamp 1655484843
transform 1 0 16008 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_40
timestamp 1655484843
transform 1 0 14260 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_41
timestamp 1655484843
transform 1 0 9108 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_42
timestamp 1655484843
transform 1 0 8464 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_43
timestamp 1655484843
transform 1 0 7728 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_44
timestamp 1655484843
transform 1 0 22908 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_45
timestamp 1655484843
transform 1 0 19596 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_46
timestamp 1655484843
transform 1 0 18768 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_47
timestamp 1655484843
transform 1 0 15916 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_48
timestamp 1655484843
transform 1 0 15088 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_49
timestamp 1655484843
transform 1 0 10304 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_50
timestamp 1655484843
transform 1 0 22908 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_51
timestamp 1655484843
transform 1 0 16192 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_52
timestamp 1655484843
transform 1 0 8464 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_53
timestamp 1655484843
transform 1 0 22908 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_54
timestamp 1655484843
transform 1 0 17480 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_55
timestamp 1655484843
transform 1 0 9752 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_56
timestamp 1655484843
transform 1 0 9108 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_57
timestamp 1655484843
transform 1 0 8464 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_58
timestamp 1655484843
transform 1 0 22908 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_59
timestamp 1655484843
transform 1 0 15916 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_60
timestamp 1655484843
transform 1 0 15088 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_61
timestamp 1655484843
transform 1 0 11040 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_62
timestamp 1655484843
transform 1 0 9108 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_63
timestamp 1655484843
transform 1 0 8464 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_64
timestamp 1655484843
transform 1 0 22908 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_65
timestamp 1655484843
transform 1 0 21712 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_66
timestamp 1655484843
transform 1 0 16928 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_67
timestamp 1655484843
transform 1 0 9108 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_68
timestamp 1655484843
transform 1 0 8464 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_69
timestamp 1655484843
transform 1 0 14904 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_70
timestamp 1655484843
transform 1 0 12696 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_71
timestamp 1655484843
transform 1 0 9108 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_72
timestamp 1655484843
transform 1 0 8464 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_73
timestamp 1655484843
transform 1 0 22908 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_74
timestamp 1655484843
transform 1 0 9752 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_75
timestamp 1655484843
transform 1 0 22908 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_76
timestamp 1655484843
transform 1 0 18032 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_77
timestamp 1655484843
transform 1 0 14352 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_78
timestamp 1655484843
transform 1 0 11776 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_79
timestamp 1655484843
transform 1 0 8832 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_80
timestamp 1655484843
transform 1 0 5888 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_81
timestamp 1655484843
transform 1 0 22908 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_82
timestamp 1655484843
transform 1 0 22908 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_83
timestamp 1655484843
transform 1 0 22908 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_84
timestamp 1655484843
transform 1 0 21344 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_85
timestamp 1655484843
transform 1 0 18768 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_86
timestamp 1655484843
transform 1 0 18584 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_87
timestamp 1655484843
transform 1 0 18216 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_88
timestamp 1655484843
transform 1 0 13432 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_89
timestamp 1655484843
transform 1 0 12144 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_90
timestamp 1655484843
transform 1 0 6992 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_91
timestamp 1655484843
transform 1 0 18768 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_92
timestamp 1655484843
transform 1 0 17664 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_93
timestamp 1655484843
transform 1 0 16836 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_94
timestamp 1655484843
transform 1 0 13432 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_95
timestamp 1655484843
transform 1 0 8280 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_96
timestamp 1655484843
transform 1 0 7176 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_97
timestamp 1655484843
transform 1 0 21160 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_98
timestamp 1655484843
transform 1 0 18584 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_99
timestamp 1655484843
transform 1 0 16008 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_100
timestamp 1655484843
transform 1 0 13432 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_101
timestamp 1655484843
transform 1 0 8280 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_102
timestamp 1655484843
transform 1 0 17480 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_103
timestamp 1655484843
transform 1 0 9568 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_104
timestamp 1655484843
transform 1 0 8832 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_105
timestamp 1655484843
transform 1 0 22908 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_106
timestamp 1655484843
transform 1 0 21344 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_107
timestamp 1655484843
transform 1 0 14352 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_108
timestamp 1655484843
transform 1 0 8280 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_109
timestamp 1655484843
transform 1 0 6440 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_110
timestamp 1655484843
transform 1 0 12328 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_111
timestamp 1655484843
transform 1 0 12144 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_112
timestamp 1655484843
transform 1 0 9568 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_113
timestamp 1655484843
transform 1 0 19688 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_114
timestamp 1655484843
transform 1 0 6256 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_115
timestamp 1655484843
transform 1 0 10672 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_116
timestamp 1655484843
transform 1 0 6992 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_117
timestamp 1655484843
transform 1 0 5796 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_118
timestamp 1655484843
transform 1 0 21160 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_119
timestamp 1655484843
transform 1 0 20424 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_120
timestamp 1655484843
transform 1 0 16008 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_121
timestamp 1655484843
transform 1 0 13616 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_122
timestamp 1655484843
transform 1 0 8280 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_123
timestamp 1655484843
transform 1 0 22448 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_124
timestamp 1655484843
transform 1 0 17296 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_125
timestamp 1655484843
transform 1 0 16560 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_126
timestamp 1655484843
transform 1 0 12144 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_127
timestamp 1655484843
transform 1 0 10212 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_128
timestamp 1655484843
transform 1 0 21160 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_129
timestamp 1655484843
transform 1 0 19596 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_130
timestamp 1655484843
transform 1 0 11960 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_131
timestamp 1655484843
transform 1 0 8924 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_132
timestamp 1655484843
transform 1 0 17480 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_133
timestamp 1655484843
transform 1 0 10488 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_134
timestamp 1655484843
transform 1 0 18584 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_135
timestamp 1655484843
transform 1 0 13432 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_136
timestamp 1655484843
transform 1 0 10856 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_137
timestamp 1655484843
transform 1 0 22448 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_138
timestamp 1655484843
transform 1 0 20056 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_139
timestamp 1655484843
transform 1 0 18952 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_140
timestamp 1655484843
transform 1 0 10672 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_141
timestamp 1655484843
transform 1 0 12788 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_142
timestamp 1655484843
transform 1 0 11040 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_143
timestamp 1655484843
transform 1 0 10856 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_144
timestamp 1655484843
transform 1 0 12696 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_145
timestamp 1655484843
transform 1 0 10488 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_146
timestamp 1655484843
transform 1 0 7176 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_147
timestamp 1655484843
transform 1 0 16008 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_148
timestamp 1655484843
transform 1 0 11776 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_149
timestamp 1655484843
transform 1 0 6256 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_150
timestamp 1655484843
transform 1 0 17480 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_151
timestamp 1655484843
transform 1 0 9752 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_152
timestamp 1655484843
transform 1 0 7176 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_153
timestamp 1655484843
transform 1 0 6532 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_154
timestamp 1655484843
transform 1 0 11960 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_155
timestamp 1655484843
transform 1 0 6532 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_156
timestamp 1655484843
transform 1 0 21528 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_157
timestamp 1655484843
transform 1 0 6716 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_158
timestamp 1655484843
transform 1 0 5796 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_159
timestamp 1655484843
transform 1 0 22908 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_160
timestamp 1655484843
transform 1 0 21344 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_161
timestamp 1655484843
transform 1 0 16008 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_162
timestamp 1655484843
transform 1 0 13432 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_163
timestamp 1655484843
transform 1 0 9200 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_164
timestamp 1655484843
transform 1 0 19872 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_165
timestamp 1655484843
transform 1 0 12512 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_166
timestamp 1655484843
transform 1 0 12144 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_167
timestamp 1655484843
transform 1 0 9200 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_168
timestamp 1655484843
transform 1 0 6808 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_169
timestamp 1655484843
transform 1 0 6256 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_170
timestamp 1655484843
transform 1 0 12144 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_171
timestamp 1655484843
transform 1 0 22816 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_172
timestamp 1655484843
transform 1 0 21160 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_173
timestamp 1655484843
transform 1 0 16008 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_174
timestamp 1655484843
transform 1 0 15088 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_175
timestamp 1655484843
transform 1 0 22448 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_176
timestamp 1655484843
transform 1 0 21344 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_177
timestamp 1655484843
transform 1 0 20056 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_178
timestamp 1655484843
transform 1 0 18768 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_179
timestamp 1655484843
transform 1 0 17480 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_180
timestamp 1655484843
transform 1 0 16192 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_181
timestamp 1655484843
transform 1 0 16008 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_182
timestamp 1655484843
transform 1 0 13616 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_183
timestamp 1655484843
transform 1 0 8280 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_184
timestamp 1655484843
transform 1 0 7728 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_185
timestamp 1655484843
transform 1 0 6992 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 13616 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1655484843
transform 1 0 7176 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_2
timestamp 1655484843
transform 1 0 8464 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_3
timestamp 1655484843
transform 1 0 8740 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_4
timestamp 1655484843
transform 1 0 5796 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_5
timestamp 1655484843
transform 1 0 20240 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_6
timestamp 1655484843
transform 1 0 5888 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_7
timestamp 1655484843
transform 1 0 5796 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_8
timestamp 1655484843
transform 1 0 8464 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_9
timestamp 1655484843
transform 1 0 9752 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_10
timestamp 1655484843
transform 1 0 20056 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_11
timestamp 1655484843
transform 1 0 16468 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_12
timestamp 1655484843
transform 1 0 9752 0 -1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_13
timestamp 1655484843
transform 1 0 8740 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_14
timestamp 1655484843
transform 1 0 7176 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_15
timestamp 1655484843
transform 1 0 7176 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_16
timestamp 1655484843
transform 1 0 18676 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_17
timestamp 1655484843
transform 1 0 15916 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_18
timestamp 1655484843
transform 1 0 15456 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_19
timestamp 1655484843
transform 1 0 14904 0 -1 22032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_20
timestamp 1655484843
transform 1 0 17480 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_21
timestamp 1655484843
transform 1 0 16652 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_22
timestamp 1655484843
transform 1 0 14168 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_23
timestamp 1655484843
transform 1 0 13248 0 1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_24
timestamp 1655484843
transform 1 0 15732 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_25
timestamp 1655484843
transform 1 0 14628 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_26
timestamp 1655484843
transform 1 0 14168 0 -1 20944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_27
timestamp 1655484843
transform 1 0 21344 0 1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_28
timestamp 1655484843
transform 1 0 17204 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_29
timestamp 1655484843
transform 1 0 14904 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_30
timestamp 1655484843
transform 1 0 12052 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_31
timestamp 1655484843
transform 1 0 9384 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_32
timestamp 1655484843
transform 1 0 8648 0 -1 19856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_33
timestamp 1655484843
transform 1 0 11040 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_34
timestamp 1655484843
transform 1 0 6256 0 1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_35
timestamp 1655484843
transform 1 0 22356 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_36
timestamp 1655484843
transform 1 0 7176 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_37
timestamp 1655484843
transform 1 0 5796 0 -1 18768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_38
timestamp 1655484843
transform 1 0 22816 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_39
timestamp 1655484843
transform 1 0 16192 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_40
timestamp 1655484843
transform 1 0 8188 0 1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_41
timestamp 1655484843
transform 1 0 14904 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_42
timestamp 1655484843
transform 1 0 9476 0 -1 17680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_43
timestamp 1655484843
transform 1 0 22816 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_44
timestamp 1655484843
transform 1 0 20240 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_45
timestamp 1655484843
transform 1 0 15824 0 1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_46
timestamp 1655484843
transform 1 0 14904 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_47
timestamp 1655484843
transform 1 0 13156 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_48
timestamp 1655484843
transform 1 0 7176 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_49
timestamp 1655484843
transform 1 0 5796 0 -1 16592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_50
timestamp 1655484843
transform 1 0 22816 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_51
timestamp 1655484843
transform 1 0 19412 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_52
timestamp 1655484843
transform 1 0 11500 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_53
timestamp 1655484843
transform 1 0 11040 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_54
timestamp 1655484843
transform 1 0 8740 0 1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_55
timestamp 1655484843
transform 1 0 21896 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_56
timestamp 1655484843
transform 1 0 9752 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_57
timestamp 1655484843
transform 1 0 5796 0 -1 15504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_58
timestamp 1655484843
transform 1 0 22816 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_59
timestamp 1655484843
transform 1 0 15916 0 1 14416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_60
timestamp 1655484843
transform 1 0 22816 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_61
timestamp 1655484843
transform 1 0 13616 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_62
timestamp 1655484843
transform 1 0 13340 0 1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_63
timestamp 1655484843
transform 1 0 15732 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_64
timestamp 1655484843
transform 1 0 14904 0 -1 13328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_65
timestamp 1655484843
transform 1 0 22816 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_66
timestamp 1655484843
transform 1 0 13340 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_67
timestamp 1655484843
transform 1 0 8464 0 1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_68
timestamp 1655484843
transform 1 0 6164 0 -1 12240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_69
timestamp 1655484843
transform 1 0 22816 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_70
timestamp 1655484843
transform 1 0 21068 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_71
timestamp 1655484843
transform 1 0 20240 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_72
timestamp 1655484843
transform 1 0 11868 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_73
timestamp 1655484843
transform 1 0 10764 0 1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_74
timestamp 1655484843
transform 1 0 19780 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_75
timestamp 1655484843
transform 1 0 12052 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_76
timestamp 1655484843
transform 1 0 8740 0 -1 11152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_77
timestamp 1655484843
transform 1 0 22816 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_78
timestamp 1655484843
transform 1 0 11776 0 1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_79
timestamp 1655484843
transform 1 0 19780 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_80
timestamp 1655484843
transform 1 0 10396 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_81
timestamp 1655484843
transform 1 0 9752 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_82
timestamp 1655484843
transform 1 0 6164 0 -1 10064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_83
timestamp 1655484843
transform 1 0 10764 0 1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_84
timestamp 1655484843
transform 1 0 12328 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_85
timestamp 1655484843
transform 1 0 6900 0 -1 8976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_86
timestamp 1655484843
transform 1 0 22816 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_87
timestamp 1655484843
transform 1 0 13340 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_88
timestamp 1655484843
transform 1 0 10764 0 1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_89
timestamp 1655484843
transform 1 0 22356 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_90
timestamp 1655484843
transform 1 0 21712 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_91
timestamp 1655484843
transform 1 0 8648 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_92
timestamp 1655484843
transform 1 0 6900 0 -1 7888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_93
timestamp 1655484843
transform 1 0 17664 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_94
timestamp 1655484843
transform 1 0 6716 0 1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_95
timestamp 1655484843
transform 1 0 21160 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_96
timestamp 1655484843
transform 1 0 6348 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_97
timestamp 1655484843
transform 1 0 5796 0 -1 6800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_98
timestamp 1655484843
transform 1 0 10764 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_99
timestamp 1655484843
transform 1 0 7544 0 1 5712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 15364 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_1
timestamp 1655484843
transform 1 0 13800 0 -1 20944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_2
timestamp 1655484843
transform 1 0 16836 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_3
timestamp 1655484843
transform 1 0 15548 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_4
timestamp 1655484843
transform 1 0 8280 0 -1 19856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_5
timestamp 1655484843
transform 1 0 5888 0 1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_6
timestamp 1655484843
transform 1 0 21528 0 -1 18768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_7
timestamp 1655484843
transform 1 0 7820 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_8
timestamp 1655484843
transform 1 0 5888 0 1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_9
timestamp 1655484843
transform 1 0 21528 0 -1 15504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_10
timestamp 1655484843
transform 1 0 20884 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_11
timestamp 1655484843
transform 1 0 10488 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_12
timestamp 1655484843
transform 1 0 8464 0 1 14416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_13
timestamp 1655484843
transform 1 0 5888 0 1 13328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_14
timestamp 1655484843
transform 1 0 16376 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_15
timestamp 1655484843
transform 1 0 5796 0 -1 12240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_16
timestamp 1655484843
transform 1 0 20884 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_17
timestamp 1655484843
transform 1 0 18308 0 1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_18
timestamp 1655484843
transform 1 0 19412 0 -1 10064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_19
timestamp 1655484843
transform 1 0 20884 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_20
timestamp 1655484843
transform 1 0 18308 0 1 8976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_21
timestamp 1655484843
transform 1 0 20884 0 1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_22
timestamp 1655484843
transform 1 0 6072 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_23
timestamp 1655484843
transform 1 0 18308 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_24
timestamp 1655484843
transform 1 0 15640 0 1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_25
timestamp 1655484843
transform 1 0 7176 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_26
timestamp 1655484843
transform 1 0 7176 0 1 5712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 17480 0 -1 8976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1655484843
transform 1 0 9752 0 1 5712
box -38 -48 774 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 7084 0 -1 15504
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_1
timestamp 1655484843
transform 1 0 5888 0 -1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_2
timestamp 1655484843
transform 1 0 5980 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_3
timestamp 1655484843
transform -1 0 8464 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_4
timestamp 1655484843
transform -1 0 9568 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_5
timestamp 1655484843
transform -1 0 10672 0 1 17680
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_6
timestamp 1655484843
transform -1 0 10488 0 1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_7
timestamp 1655484843
transform 1 0 20056 0 -1 6800
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_8
timestamp 1655484843
transform 1 0 18860 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_9
timestamp 1655484843
transform -1 0 21252 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_10
timestamp 1655484843
transform -1 0 22540 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_11
timestamp 1655484843
transform -1 0 22448 0 -1 6800
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_12
timestamp 1655484843
transform 1 0 21436 0 1 8976
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_13
timestamp 1655484843
transform 1 0 18860 0 -1 18768
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_14
timestamp 1655484843
transform -1 0 22540 0 -1 22032
box -38 -48 1142 592
use sky130_fd_sc_hd__ha_2  sky130_fd_sc_hd__ha_2_15
timestamp 1655484843
transform -1 0 17388 0 1 5712
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 15364 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1655484843
transform 1 0 13064 0 1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1655484843
transform 1 0 8464 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_3
timestamp 1655484843
transform 1 0 11224 0 1 15504
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_4
timestamp 1655484843
transform -1 0 22908 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_5
timestamp 1655484843
transform 1 0 17756 0 1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_6
timestamp 1655484843
transform -1 0 14628 0 -1 20944
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_7
timestamp 1655484843
transform -1 0 6072 0 -1 7888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_8
timestamp 1655484843
transform -1 0 6808 0 -1 13328
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_9
timestamp 1655484843
transform -1 0 6532 0 1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_10
timestamp 1655484843
transform 1 0 7176 0 -1 8976
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 9476 0 -1 17680
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_1
timestamp 1655484843
transform -1 0 12144 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  sky130_fd_sc_hd__nand3_1_2
timestamp 1655484843
transform -1 0 6348 0 -1 6800
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  sky130_fd_sc_hd__nand4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 8924 0 -1 19856
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 13524 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1655484843
transform 1 0 13708 0 1 5712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1655484843
transform -1 0 18584 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1655484843
transform 1 0 15640 0 -1 22032
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1655484843
transform 1 0 11592 0 1 18768
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1655484843
transform -1 0 6624 0 1 12240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_6
timestamp 1655484843
transform -1 0 6164 0 -1 10064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_7
timestamp 1655484843
transform 1 0 7912 0 -1 6800
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  sky130_fd_sc_hd__nor3_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 9200 0 -1 16592
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 20056 0 -1 22032
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_1
timestamp 1655484843
transform 1 0 16928 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_2
timestamp 1655484843
transform 1 0 13616 0 1 20944
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_3
timestamp 1655484843
transform 1 0 11316 0 1 16592
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_4
timestamp 1655484843
transform 1 0 9936 0 -1 15504
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_5
timestamp 1655484843
transform -1 0 7268 0 1 13328
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_6
timestamp 1655484843
transform 1 0 6624 0 1 10064
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_7
timestamp 1655484843
transform 1 0 6348 0 -1 8976
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_8
timestamp 1655484843
transform 1 0 6532 0 -1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  sky130_fd_sc_hd__o21a_1_9
timestamp 1655484843
transform -1 0 6440 0 1 6800
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  sky130_fd_sc_hd__o21ai_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 14076 0 -1 7888
box -38 -48 406 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 16836 0 -1 14416
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_1
timestamp 1655484843
transform 1 0 16468 0 1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_2
timestamp 1655484843
transform -1 0 19872 0 -1 8976
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_3
timestamp 1655484843
transform -1 0 17388 0 -1 7888
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_4
timestamp 1655484843
transform 1 0 13156 0 -1 15504
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_5
timestamp 1655484843
transform -1 0 19412 0 -1 10064
box -38 -48 1694 592
use sky130_fd_sc_hd__sdlclkp_4  sky130_fd_sc_hd__sdlclkp_4_6
timestamp 1655484843
transform 1 0 16376 0 1 17680
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 22540 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1655484843
transform 1 0 21252 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1655484843
transform 1 0 19964 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1655484843
transform 1 0 18676 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1655484843
transform 1 0 17388 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1655484843
transform 1 0 16100 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1655484843
transform 1 0 14812 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1655484843
transform 1 0 13524 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1655484843
transform 1 0 12236 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1655484843
transform 1 0 10948 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1655484843
transform 1 0 9660 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1655484843
transform 1 0 8372 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1655484843
transform 1 0 7084 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1655484843
transform 1 0 5796 0 -1 22032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1655484843
transform 1 0 21252 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1655484843
transform 1 0 18676 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1655484843
transform 1 0 16100 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1655484843
transform 1 0 13524 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1655484843
transform 1 0 10948 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1655484843
transform 1 0 8372 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1655484843
transform 1 0 5796 0 1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1655484843
transform 1 0 22540 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1655484843
transform 1 0 19964 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1655484843
transform 1 0 17388 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1655484843
transform 1 0 14812 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1655484843
transform 1 0 12236 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1655484843
transform 1 0 9660 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1655484843
transform 1 0 7084 0 -1 20944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1655484843
transform 1 0 21252 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1655484843
transform 1 0 18676 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1655484843
transform 1 0 16100 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1655484843
transform 1 0 13524 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1655484843
transform 1 0 10948 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1655484843
transform 1 0 8372 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1655484843
transform 1 0 5796 0 1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1655484843
transform 1 0 22540 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1655484843
transform 1 0 19964 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1655484843
transform 1 0 17388 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1655484843
transform 1 0 14812 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1655484843
transform 1 0 12236 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1655484843
transform 1 0 9660 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1655484843
transform 1 0 7084 0 -1 19856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1655484843
transform 1 0 21252 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1655484843
transform 1 0 18676 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1655484843
transform 1 0 16100 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1655484843
transform 1 0 13524 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1655484843
transform 1 0 10948 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1655484843
transform 1 0 8372 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1655484843
transform 1 0 5796 0 1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1655484843
transform 1 0 22540 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1655484843
transform 1 0 19964 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1655484843
transform 1 0 17388 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1655484843
transform 1 0 14812 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1655484843
transform 1 0 12236 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1655484843
transform 1 0 9660 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1655484843
transform 1 0 7084 0 -1 18768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1655484843
transform 1 0 21252 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1655484843
transform 1 0 18676 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1655484843
transform 1 0 16100 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1655484843
transform 1 0 13524 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1655484843
transform 1 0 10948 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1655484843
transform 1 0 8372 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1655484843
transform 1 0 5796 0 1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1655484843
transform 1 0 22540 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1655484843
transform 1 0 19964 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1655484843
transform 1 0 17388 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1655484843
transform 1 0 14812 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1655484843
transform 1 0 12236 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1655484843
transform 1 0 9660 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1655484843
transform 1 0 7084 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1655484843
transform 1 0 21252 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1655484843
transform 1 0 18676 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1655484843
transform 1 0 16100 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1655484843
transform 1 0 13524 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1655484843
transform 1 0 10948 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1655484843
transform 1 0 8372 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1655484843
transform 1 0 5796 0 1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1655484843
transform 1 0 22540 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1655484843
transform 1 0 19964 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1655484843
transform 1 0 17388 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1655484843
transform 1 0 14812 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1655484843
transform 1 0 12236 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1655484843
transform 1 0 9660 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1655484843
transform 1 0 7084 0 -1 16592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1655484843
transform 1 0 21252 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1655484843
transform 1 0 18676 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1655484843
transform 1 0 16100 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1655484843
transform 1 0 13524 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1655484843
transform 1 0 10948 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1655484843
transform 1 0 8372 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1655484843
transform 1 0 5796 0 1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1655484843
transform 1 0 22540 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1655484843
transform 1 0 19964 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1655484843
transform 1 0 17388 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1655484843
transform 1 0 14812 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1655484843
transform 1 0 12236 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1655484843
transform 1 0 9660 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1655484843
transform 1 0 7084 0 -1 15504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1655484843
transform 1 0 21252 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1655484843
transform 1 0 18676 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1655484843
transform 1 0 16100 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1655484843
transform 1 0 13524 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1655484843
transform 1 0 10948 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1655484843
transform 1 0 8372 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1655484843
transform 1 0 5796 0 1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1655484843
transform 1 0 22540 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1655484843
transform 1 0 19964 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1655484843
transform 1 0 17388 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1655484843
transform 1 0 14812 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1655484843
transform 1 0 12236 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1655484843
transform 1 0 9660 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1655484843
transform 1 0 7084 0 -1 14416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1655484843
transform 1 0 21252 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1655484843
transform 1 0 18676 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1655484843
transform 1 0 16100 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1655484843
transform 1 0 13524 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1655484843
transform 1 0 10948 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1655484843
transform 1 0 8372 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1655484843
transform 1 0 5796 0 1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1655484843
transform 1 0 22540 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1655484843
transform 1 0 19964 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1655484843
transform 1 0 17388 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1655484843
transform 1 0 14812 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1655484843
transform 1 0 12236 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1655484843
transform 1 0 9660 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1655484843
transform 1 0 7084 0 -1 13328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1655484843
transform 1 0 21252 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1655484843
transform 1 0 18676 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1655484843
transform 1 0 16100 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1655484843
transform 1 0 13524 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1655484843
transform 1 0 10948 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1655484843
transform 1 0 8372 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1655484843
transform 1 0 5796 0 1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1655484843
transform 1 0 22540 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1655484843
transform 1 0 19964 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1655484843
transform 1 0 17388 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1655484843
transform 1 0 14812 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1655484843
transform 1 0 12236 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1655484843
transform 1 0 9660 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1655484843
transform 1 0 7084 0 -1 12240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1655484843
transform 1 0 21252 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1655484843
transform 1 0 18676 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1655484843
transform 1 0 16100 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1655484843
transform 1 0 13524 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1655484843
transform 1 0 10948 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1655484843
transform 1 0 8372 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1655484843
transform 1 0 5796 0 1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1655484843
transform 1 0 22540 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1655484843
transform 1 0 19964 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1655484843
transform 1 0 17388 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1655484843
transform 1 0 14812 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1655484843
transform 1 0 12236 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1655484843
transform 1 0 9660 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1655484843
transform 1 0 7084 0 -1 11152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1655484843
transform 1 0 21252 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1655484843
transform 1 0 18676 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1655484843
transform 1 0 16100 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1655484843
transform 1 0 13524 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1655484843
transform 1 0 10948 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1655484843
transform 1 0 8372 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1655484843
transform 1 0 5796 0 1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1655484843
transform 1 0 22540 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1655484843
transform 1 0 19964 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1655484843
transform 1 0 17388 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1655484843
transform 1 0 14812 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1655484843
transform 1 0 12236 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1655484843
transform 1 0 9660 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1655484843
transform 1 0 7084 0 -1 10064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1655484843
transform 1 0 21252 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1655484843
transform 1 0 18676 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1655484843
transform 1 0 16100 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1655484843
transform 1 0 13524 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1655484843
transform 1 0 10948 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1655484843
transform 1 0 8372 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1655484843
transform 1 0 5796 0 1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1655484843
transform 1 0 22540 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1655484843
transform 1 0 19964 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1655484843
transform 1 0 17388 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1655484843
transform 1 0 14812 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1655484843
transform 1 0 12236 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1655484843
transform 1 0 9660 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_181
timestamp 1655484843
transform 1 0 7084 0 -1 8976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1655484843
transform 1 0 21252 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1655484843
transform 1 0 18676 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1655484843
transform 1 0 16100 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1655484843
transform 1 0 13524 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1655484843
transform 1 0 10948 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1655484843
transform 1 0 8372 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1655484843
transform 1 0 5796 0 1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1655484843
transform 1 0 22540 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1655484843
transform 1 0 19964 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1655484843
transform 1 0 17388 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1655484843
transform 1 0 14812 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1655484843
transform 1 0 12236 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1655484843
transform 1 0 9660 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1655484843
transform 1 0 7084 0 -1 7888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_196
timestamp 1655484843
transform 1 0 21252 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_197
timestamp 1655484843
transform 1 0 18676 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_198
timestamp 1655484843
transform 1 0 16100 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_199
timestamp 1655484843
transform 1 0 13524 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_200
timestamp 1655484843
transform 1 0 10948 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_201
timestamp 1655484843
transform 1 0 8372 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_202
timestamp 1655484843
transform 1 0 5796 0 1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_203
timestamp 1655484843
transform 1 0 22540 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_204
timestamp 1655484843
transform 1 0 19964 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_205
timestamp 1655484843
transform 1 0 17388 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_206
timestamp 1655484843
transform 1 0 14812 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_207
timestamp 1655484843
transform 1 0 12236 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_208
timestamp 1655484843
transform 1 0 9660 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_209
timestamp 1655484843
transform 1 0 7084 0 -1 6800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_210
timestamp 1655484843
transform 1 0 22540 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_211
timestamp 1655484843
transform 1 0 21252 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_212
timestamp 1655484843
transform 1 0 19964 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_213
timestamp 1655484843
transform 1 0 18676 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_214
timestamp 1655484843
transform 1 0 17388 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_215
timestamp 1655484843
transform 1 0 16100 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_216
timestamp 1655484843
transform 1 0 14812 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_217
timestamp 1655484843
transform 1 0 13524 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_218
timestamp 1655484843
transform 1 0 12236 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_219
timestamp 1655484843
transform 1 0 10948 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_220
timestamp 1655484843
transform 1 0 9660 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_221
timestamp 1655484843
transform 1 0 8372 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_222
timestamp 1655484843
transform 1 0 7084 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_223
timestamp 1655484843
transform 1 0 5796 0 1 5712
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  sky130_fd_sc_hd__xnor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform -1 0 21252 0 -1 22032
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  sky130_fd_sc_hd__xnor2_1_1
timestamp 1655484843
transform -1 0 6808 0 -1 14416
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655484843
transform 1 0 5980 0 -1 16592
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1655484843
transform 1 0 21896 0 -1 11152
box -38 -48 682 592
<< labels >>
rlabel metal2 s 28736 0 28764 97 4 clk
port 1 nsew
rlabel metal2 s 19168 0 19196 97 4 rst_n
port 2 nsew
rlabel metal2 s 9600 0 9628 97 4 sclk
port 3 nsew
rlabel metal2 s 32 0 60 97 4 cs_n
port 4 nsew
rlabel metal3 s 0 13768 160 13828 4 data_in
port 5 nsew
rlabel metal3 s 28636 104 28796 164 4 data_out[11]
port 6 nsew
rlabel metal3 s 28636 2666 28796 2726 4 data_out[10]
port 7 nsew
rlabel metal3 s 28636 5228 28796 5288 4 data_out[9]
port 8 nsew
rlabel metal3 s 28636 7668 28796 7728 4 data_out[8]
port 9 nsew
rlabel metal3 s 28636 10230 28796 10290 4 data_out[7]
port 10 nsew
rlabel metal3 s 28636 12670 28796 12730 4 data_out[6]
port 11 nsew
rlabel metal3 s 28636 15232 28796 15292 4 data_out[5]
port 12 nsew
rlabel metal3 s 28636 17672 28796 17732 4 data_out[4]
port 13 nsew
rlabel metal3 s 28636 20234 28796 20294 4 data_out[3]
port 14 nsew
rlabel metal3 s 28636 22674 28796 22734 4 data_out[2]
port 15 nsew
rlabel metal3 s 28636 25236 28796 25296 4 data_out[1]
port 16 nsew
rlabel metal3 s 28636 27676 28796 27736 4 data_out[0]
port 17 nsew
rlabel metal2 s 32 27647 60 27744 4 new_data
port 18 nsew
rlabel metal2 s 28736 27647 28764 27744 4 serial_data_out
port 19 nsew
rlabel metal5 s 0 3852 620 4472 4 VSS
port 20 nsew
rlabel metal5 s 0 5092 620 5712 4 VDD
port 21 nsew
<< properties >>
string GDS_END 345230
string GDS_FILE digital_filter_3a.gds
string GDS_START 120
string path 451.950 281.350 456.550 281.350 
<< end >>
