* NGSPICE file created from sc_cmfb.ext - technology: sky130A

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_n416_n136# a_448_n136# 0.02fF
C1 a_n32_n136# a_160_n136# 0.12fF
C2 a_352_n136# a_n508_n136# 0.02fF
C3 w_n646_n356# a_n508_n136# 0.13fF
C4 a_n416_n136# a_n320_n136# 0.33fF
C5 a_n416_n136# a_256_n136# 0.03fF
C6 a_n224_n136# a_n128_n136# 0.33fF
C7 a_352_n136# a_n32_n136# 0.05fF
C8 w_n646_n356# a_n32_n136# 0.05fF
C9 a_448_n136# a_n224_n136# 0.03fF
C10 a_n320_n136# a_n224_n136# 0.33fF
C11 a_n224_n136# a_256_n136# 0.04fF
C12 a_64_n136# a_n128_n136# 0.12fF
C13 a_448_n136# a_64_n136# 0.05fF
C14 a_n512_n234# a_n128_n136# 0.03fF
C15 a_352_n136# a_160_n136# 0.12fF
C16 w_n646_n356# a_160_n136# 0.06fF
C17 a_n320_n136# a_64_n136# 0.05fF
C18 a_64_n136# a_256_n136# 0.12fF
C19 a_n512_n234# a_448_n136# 0.03fF
C20 a_n508_n136# a_n128_n136# 0.05fF
C21 a_n416_n136# a_n224_n136# 0.12fF
C22 w_n646_n356# a_352_n136# 0.08fF
C23 a_n512_n234# a_n320_n136# 0.03fF
C24 a_n512_n234# a_256_n136# 0.03fF
C25 a_448_n136# a_n508_n136# 0.02fF
C26 a_n32_n136# a_n128_n136# 0.33fF
C27 a_n320_n136# a_n508_n136# 0.12fF
C28 a_n508_n136# a_256_n136# 0.02fF
C29 a_448_n136# a_n32_n136# 0.04fF
C30 a_n416_n136# a_64_n136# 0.04fF
C31 a_n32_n136# a_n320_n136# 0.07fF
C32 a_n32_n136# a_256_n136# 0.07fF
C33 a_n416_n136# a_n512_n234# 0.03fF
C34 a_64_n136# a_n224_n136# 0.07fF
C35 a_160_n136# a_n128_n136# 0.07fF
C36 a_n416_n136# a_n508_n136# 0.33fF
C37 a_448_n136# a_160_n136# 0.07fF
C38 a_n512_n234# a_n224_n136# 0.03fF
C39 a_352_n136# a_n128_n136# 0.04fF
C40 w_n646_n356# a_n128_n136# 0.05fF
C41 a_n320_n136# a_160_n136# 0.04fF
C42 a_n416_n136# a_n32_n136# 0.05fF
C43 a_160_n136# a_256_n136# 0.33fF
C44 w_n646_n356# a_448_n136# 0.13fF
C45 a_352_n136# a_448_n136# 0.33fF
C46 a_n508_n136# a_n224_n136# 0.07fF
C47 a_352_n136# a_n320_n136# 0.03fF
C48 w_n646_n356# a_n320_n136# 0.06fF
C49 a_352_n136# a_256_n136# 0.33fF
C50 w_n646_n356# a_256_n136# 0.06fF
C51 a_n512_n234# a_64_n136# 0.03fF
C52 a_n32_n136# a_n224_n136# 0.12fF
C53 a_64_n136# a_n508_n136# 0.03fF
C54 a_n416_n136# a_160_n136# 0.03fF
C55 a_n32_n136# a_64_n136# 0.33fF
C56 a_n512_n234# a_n508_n136# 0.03fF
C57 a_n416_n136# a_352_n136# 0.02fF
C58 w_n646_n356# a_n416_n136# 0.08fF
C59 a_n224_n136# a_160_n136# 0.05fF
C60 a_n512_n234# a_n32_n136# 0.03fF
C61 a_448_n136# a_n128_n136# 0.03fF
C62 a_352_n136# a_n224_n136# 0.03fF
C63 w_n646_n356# a_n224_n136# 0.06fF
C64 a_n320_n136# a_n128_n136# 0.12fF
C65 a_n32_n136# a_n508_n136# 0.04fF
C66 a_256_n136# a_n128_n136# 0.05fF
C67 a_64_n136# a_160_n136# 0.33fF
C68 a_448_n136# a_n320_n136# 0.02fF
C69 a_448_n136# a_256_n136# 0.12fF
C70 a_n320_n136# a_256_n136# 0.03fF
C71 a_n512_n234# a_160_n136# 0.03fF
C72 a_352_n136# a_64_n136# 0.07fF
C73 w_n646_n356# a_64_n136# 0.05fF
C74 a_n508_n136# a_160_n136# 0.03fF
C75 a_n416_n136# a_n128_n136# 0.07fF
C76 a_352_n136# a_n512_n234# 0.03fF
C77 w_n646_n356# a_n512_n234# 1.47fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# a_448_n52# a_n416_n52# a_160_n52#
+ a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149# a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_64_n52# a_n320_n52# 0.02fF
C1 a_352_n52# a_64_n52# 0.03fF
C2 a_n128_n52# a_160_n52# 0.03fF
C3 a_n416_n52# a_256_n52# 0.01fF
C4 a_64_n52# a_n224_n52# 0.03fF
C5 a_256_n52# a_n32_n52# 0.03fF
C6 a_n128_n52# a_n416_n52# 0.03fF
C7 a_n128_n52# a_n32_n52# 0.13fF
C8 a_256_n52# a_64_n52# 0.05fF
C9 a_n128_n52# a_64_n52# 0.05fF
C10 a_352_n52# a_n320_n52# 0.01fF
C11 a_n508_n52# a_448_n52# 0.01fF
C12 a_n320_n52# a_n224_n52# 0.13fF
C13 a_352_n52# a_n224_n52# 0.01fF
C14 a_448_n52# a_n512_n149# 0.03fF
C15 a_256_n52# a_n320_n52# 0.01fF
C16 a_352_n52# a_256_n52# 0.13fF
C17 a_n508_n52# a_n512_n149# 0.03fF
C18 a_n128_n52# a_n320_n52# 0.05fF
C19 a_352_n52# a_n128_n52# 0.02fF
C20 a_256_n52# a_n224_n52# 0.02fF
C21 a_n128_n52# a_n224_n52# 0.13fF
C22 a_448_n52# a_160_n52# 0.03fF
C23 a_n508_n52# a_160_n52# 0.01fF
C24 a_n128_n52# a_256_n52# 0.02fF
C25 a_n416_n52# a_448_n52# 0.01fF
C26 a_n508_n52# a_n416_n52# 0.13fF
C27 a_448_n52# a_n32_n52# 0.02fF
C28 a_n508_n52# a_n32_n52# 0.02fF
C29 a_n512_n149# a_160_n52# 0.03fF
C30 a_448_n52# a_64_n52# 0.02fF
C31 a_n508_n52# a_64_n52# 0.01fF
C32 a_n416_n52# a_n512_n149# 0.03fF
C33 a_n512_n149# a_n32_n52# 0.03fF
C34 a_64_n52# a_n512_n149# 0.03fF
C35 a_n416_n52# a_160_n52# 0.01fF
C36 a_160_n52# a_n32_n52# 0.05fF
C37 a_448_n52# a_n320_n52# 0.01fF
C38 a_352_n52# a_448_n52# 0.13fF
C39 a_n508_n52# a_n320_n52# 0.05fF
C40 a_352_n52# a_n508_n52# 0.01fF
C41 a_64_n52# a_160_n52# 0.13fF
C42 a_n416_n52# a_n32_n52# 0.02fF
C43 a_448_n52# a_n224_n52# 0.01fF
C44 a_n508_n52# a_n224_n52# 0.03fF
C45 a_n416_n52# a_64_n52# 0.02fF
C46 a_64_n52# a_n32_n52# 0.13fF
C47 a_n512_n149# a_n320_n52# 0.03fF
C48 a_352_n52# a_n512_n149# 0.03fF
C49 a_256_n52# a_448_n52# 0.05fF
C50 a_n508_n52# a_256_n52# 0.01fF
C51 a_n128_n52# a_448_n52# 0.01fF
C52 a_n508_n52# a_n128_n52# 0.02fF
C53 a_n512_n149# a_n224_n52# 0.03fF
C54 a_160_n52# a_n320_n52# 0.02fF
C55 a_352_n52# a_160_n52# 0.05fF
C56 a_256_n52# a_n512_n149# 0.03fF
C57 a_n128_n52# a_n512_n149# 0.03fF
C58 a_160_n52# a_n224_n52# 0.02fF
C59 a_n416_n52# a_n320_n52# 0.13fF
C60 a_352_n52# a_n416_n52# 0.01fF
C61 a_n320_n52# a_n32_n52# 0.03fF
C62 a_352_n52# a_n32_n52# 0.02fF
C63 a_n416_n52# a_n224_n52# 0.05fF
C64 a_256_n52# a_160_n52# 0.13fF
C65 a_n224_n52# a_n32_n52# 0.05fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate en en_b VDD in out VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in out in in VSS out in out out en out nmos_tgate
C0 in VDD 0.70fF
C1 en_b en 0.07fF
C2 in en 0.13fF
C3 en_b out 0.01fF
C4 in out 0.77fF
C5 en VDD 0.12fF
C6 out VDD 0.29fF
C7 out en 0.01fF
C8 in en_b 0.15fF
C9 en_b VDD -0.11fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 c1_n530_n480# m3_n630_n580# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb on cm bias_a op cmc p2_b p2 p1_b p1 VDD VSS
Xtransmission_gate_10 p1 p1_b VDD transmission_gate_3/out on VSS transmission_gate
Xtransmission_gate_11 p1 p1_b VDD transmission_gate_4/out op VSS transmission_gate
Xtransmission_gate_0 p1 p1_b VDD cm transmission_gate_7/in VSS transmission_gate
Xtransmission_gate_1 p1 p1_b VDD cm transmission_gate_6/in VSS transmission_gate
Xtransmission_gate_2 p1 p1_b VDD bias_a transmission_gate_8/in VSS transmission_gate
Xtransmission_gate_3 p2 p2_b VDD cm transmission_gate_3/out VSS transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 p2_b VDD cm transmission_gate_4/out VSS transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 p2_b VDD bias_a transmission_gate_9/in VSS transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 p2_b VDD transmission_gate_6/in op VSS transmission_gate
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 p2_b VDD transmission_gate_7/in on VSS transmission_gate
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 p2_b VDD transmission_gate_8/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 p1_b VDD transmission_gate_9/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 transmission_gate_7/in transmission_gate_6/in 0.47fF
C1 p1_b transmission_gate_3/out 0.59fF
C2 transmission_gate_4/out unit_cap_mim_m3m4_30/m3_n630_n580# -0.80fF
C3 transmission_gate_9/in cmc 3.45fF
C4 p2_b transmission_gate_6/in 0.42fF
C5 transmission_gate_3/out unit_cap_mim_m3m4_17/m3_n630_n580# -0.23fF
C6 transmission_gate_6/in unit_cap_mim_m3m4_29/m3_n630_n580# -0.80fF
C7 transmission_gate_9/in cm 0.04fF
C8 transmission_gate_9/in unit_cap_mim_m3m4_16/m3_n630_n580# 0.17fF
C9 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C10 transmission_gate_3/out transmission_gate_7/in 0.30fF
C11 cmc unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C12 p2_b transmission_gate_3/out 0.10fF
C13 p1_b unit_cap_mim_m3m4_18/m3_n630_n580# 0.06fF
C14 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C15 p1 unit_cap_mim_m3m4_29/c1_n530_n480# 0.11fF
C16 op unit_cap_mim_m3m4_30/m3_n630_n580# 0.56fF
C17 transmission_gate_6/in cmc 0.96fF
C18 transmission_gate_9/in on 0.82fF
C19 unit_cap_mim_m3m4_25/c1_n530_n480# p2 0.04fF
C20 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_27/m3_n630_n580# 0.12fF
C21 transmission_gate_6/in cm 0.17fF
C22 transmission_gate_9/in p1 0.70fF
C23 p1_b unit_cap_mim_m3m4_24/m3_n630_n580# 0.06fF
C24 transmission_gate_4/out op 1.12fF
C25 transmission_gate_3/out cmc 0.74fF
C26 transmission_gate_4/out unit_cap_mim_m3m4_31/c1_n530_n480# 0.05fF
C27 unit_cap_mim_m3m4_28/c1_n530_n480# p1_b 0.06fF
C28 transmission_gate_3/out cm 0.17fF
C29 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_8/in 0.17fF
C30 p1_b unit_cap_mim_m3m4_23/m3_n630_n580# 0.05fF
C31 transmission_gate_4/out VDD -0.06fF
C32 unit_cap_mim_m3m4_28/c1_n530_n480# transmission_gate_7/in 0.06fF
C33 unit_cap_mim_m3m4_19/m3_n630_n580# transmission_gate_8/in 0.17fF
C34 on transmission_gate_6/in 0.41fF
C35 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# 0.12fF
C36 cmc unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C37 transmission_gate_9/in unit_cap_mim_m3m4_31/m3_n630_n580# 0.12fF
C38 transmission_gate_6/in p1 0.38fF
C39 op unit_cap_mim_m3m4_31/c1_n530_n480# 0.05fF
C40 transmission_gate_4/out p2 0.15fF
C41 transmission_gate_4/out transmission_gate_8/in 0.27fF
C42 unit_cap_mim_m3m4_27/c1_n530_n480# op 0.01fF
C43 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C44 on transmission_gate_3/out 0.39fF
C45 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C46 transmission_gate_3/out p1 0.72fF
C47 op VDD 0.89fF
C48 unit_cap_mim_m3m4_28/m3_n630_n580# transmission_gate_6/in -0.13fF
C49 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_24/m3_n630_n580# 0.10fF
C50 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C51 transmission_gate_4/out bias_a 0.10fF
C52 transmission_gate_6/in unit_cap_mim_m3m4_27/m3_n630_n580# 0.13fF
C53 op p2 0.16fF
C54 transmission_gate_8/in op 0.40fF
C55 transmission_gate_7/in unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C56 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C57 p2 unit_cap_mim_m3m4_24/c1_n530_n480# 0.04fF
C58 transmission_gate_6/in unit_cap_mim_m3m4_29/c1_n530_n480# -0.37fF
C59 unit_cap_mim_m3m4_18/m3_n630_n580# p1 0.08fF
C60 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_26/c1_n530_n480# -0.35fF
C61 unit_cap_mim_m3m4_27/c1_n530_n480# p2 0.04fF
C62 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580# -0.19fF
C63 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C64 p1_b unit_cap_mim_m3m4_22/m3_n630_n580# 0.05fF
C65 VDD p2 4.16fF
C66 transmission_gate_8/in VDD -0.07fF
C67 p1_b unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C68 transmission_gate_9/in transmission_gate_6/in 0.03fF
C69 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.17fF
C70 transmission_gate_8/in p2 0.63fF
C71 unit_cap_mim_m3m4_24/m3_n630_n580# p1 0.08fF
C72 transmission_gate_8/in unit_cap_mim_m3m4_35/m3_n630_n580# -0.10fF
C73 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C74 transmission_gate_9/in transmission_gate_3/out 1.33fF
C75 unit_cap_mim_m3m4_28/c1_n530_n480# p1 0.11fF
C76 p1_b unit_cap_mim_m3m4_30/m3_n630_n580# 0.01fF
C77 unit_cap_mim_m3m4_20/m3_n630_n580# p1_b 0.05fF
C78 on unit_cap_mim_m3m4_23/m3_n630_n580# 0.47fF
C79 VDD bias_a 0.99fF
C80 unit_cap_mim_m3m4_23/m3_n630_n580# p1 0.06fF
C81 unit_cap_mim_m3m4_19/m3_n630_n580# p1_b 0.06fF
C82 transmission_gate_8/in unit_cap_mim_m3m4_21/c1_n530_n480# -0.41fF
C83 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C84 bias_a p2 0.60fF
C85 transmission_gate_8/in bias_a 0.04fF
C86 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_7/in -0.56fF
C87 transmission_gate_4/out p1_b 0.55fF
C88 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.10fF
C89 transmission_gate_7/in unit_cap_mim_m3m4_20/c1_n530_n480# -0.18fF
C90 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580# -0.33fF
C91 unit_cap_mim_m3m4_26/m3_n630_n580# cmc 0.10fF
C92 unit_cap_mim_m3m4_19/m3_n630_n580# transmission_gate_7/in -0.28fF
C93 cmc unit_cap_mim_m3m4_22/m3_n630_n580# 0.71fF
C94 transmission_gate_3/out transmission_gate_6/in 0.75fF
C95 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C96 transmission_gate_4/out transmission_gate_7/in 0.62fF
C97 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C98 transmission_gate_4/out p2_b 0.05fF
C99 transmission_gate_9/in unit_cap_mim_m3m4_24/m3_n630_n580# 0.23fF
C100 unit_cap_mim_m3m4_22/c1_n530_n480# op 0.07fF
C101 p1_b op 0.28fF
C102 unit_cap_mim_m3m4_23/c1_n530_n480# on 0.19fF
C103 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C104 p1_b unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C105 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C106 transmission_gate_6/in unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C107 p1_b unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C108 transmission_gate_9/in unit_cap_mim_m3m4_23/m3_n630_n580# 0.17fF
C109 op transmission_gate_7/in 2.65fF
C110 transmission_gate_4/out unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C111 p2_b op 0.40fF
C112 op unit_cap_mim_m3m4_29/m3_n630_n580# 0.39fF
C113 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_31/c1_n530_n480# 0.06fF
C114 p1_b VDD 1.01fF
C115 transmission_gate_4/out cmc 0.15fF
C116 unit_cap_mim_m3m4_22/m3_n630_n580# p1 0.06fF
C117 unit_cap_mim_m3m4_26/c1_n530_n480# p2 0.04fF
C118 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580# -0.12fF
C119 on unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C120 unit_cap_mim_m3m4_25/c1_n530_n480# p1 0.11fF
C121 transmission_gate_4/out cm 0.07fF
C122 transmission_gate_4/out unit_cap_mim_m3m4_16/m3_n630_n580# -0.28fF
C123 p1_b p2 5.94fF
C124 transmission_gate_8/in p1_b 0.17fF
C125 p1_b unit_cap_mim_m3m4_35/m3_n630_n580# 0.01fF
C126 unit_cap_mim_m3m4_17/m3_n630_n580# p2 0.04fF
C127 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C128 VDD transmission_gate_7/in -0.16fF
C129 unit_cap_mim_m3m4_28/c1_n530_n480# transmission_gate_6/in 0.05fF
C130 p2_b VDD 1.67fF
C131 unit_cap_mim_m3m4_20/m3_n630_n580# on 0.61fF
C132 transmission_gate_8/in unit_cap_mim_m3m4_21/m3_n630_n580# -1.15fF
C133 transmission_gate_7/in p2 0.60fF
C134 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_27/m3_n630_n580# 0.12fF
C135 transmission_gate_8/in transmission_gate_7/in -0.35fF
C136 unit_cap_mim_m3m4_30/m3_n630_n580# p1 0.06fF
C137 unit_cap_mim_m3m4_20/m3_n630_n580# p1 0.06fF
C138 on unit_cap_mim_m3m4_20/c1_n530_n480# 0.15fF
C139 transmission_gate_4/out unit_cap_mim_m3m4_30/c1_n530_n480# -0.37fF
C140 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C141 p2_b p2 6.58fF
C142 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C143 transmission_gate_8/in p2_b 0.40fF
C144 op cmc -0.30fF
C145 unit_cap_mim_m3m4_33/m3_n630_n580# cmc 0.12fF
C146 transmission_gate_9/in unit_cap_mim_m3m4_25/m3_n630_n580# 0.27fF
C147 unit_cap_mim_m3m4_19/m3_n630_n580# p1 0.08fF
C148 p1_b bias_a 0.52fF
C149 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_19/c1_n530_n480# -0.21fF
C150 transmission_gate_4/out on 3.25fF
C151 transmission_gate_3/out unit_cap_mim_m3m4_23/m3_n630_n580# -0.30fF
C152 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580# -0.19fF
C153 op unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C154 transmission_gate_4/out p1 0.80fF
C155 transmission_gate_7/in bias_a 0.11fF
C156 VDD cmc 1.23fF
C157 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_34/c1_n530_n480# -0.14fF
C158 op unit_cap_mim_m3m4_30/c1_n530_n480# 0.18fF
C159 p2_b bias_a 0.48fF
C160 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580# 0.17fF
C161 transmission_gate_9/in unit_cap_mim_m3m4_22/m3_n630_n580# -0.80fF
C162 VDD cm 1.83fF
C163 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_31/c1_n530_n480# 0.06fF
C164 cmc p2 0.25fF
C165 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580# -0.13fF
C166 transmission_gate_8/in cmc 1.73fF
C167 on op 2.09fF
C168 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C169 cm p2 1.33fF
C170 unit_cap_mim_m3m4_16/m3_n630_n580# p2 0.05fF
C171 transmission_gate_8/in cm 0.03fF
C172 op p1 0.52fF
C173 transmission_gate_4/out unit_cap_mim_m3m4_31/m3_n630_n580# 0.32fF
C174 unit_cap_mim_m3m4_24/c1_n530_n480# p1 0.11fF
C175 unit_cap_mim_m3m4_21/c1_n530_n480# cmc 0.13fF
C176 unit_cap_mim_m3m4_27/c1_n530_n480# p1 0.11fF
C177 on VDD 0.88fF
C178 cm bias_a 1.15fF
C179 unit_cap_mim_m3m4_23/c1_n530_n480# transmission_gate_3/out -0.24fF
C180 p1_b unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C181 VDD p1 1.10fF
C182 unit_cap_mim_m3m4_28/m3_n630_n580# op 0.66fF
C183 on p2 0.24fF
C184 transmission_gate_8/in on 0.56fF
C185 transmission_gate_4/out transmission_gate_9/in -0.11fF
C186 op unit_cap_mim_m3m4_27/m3_n630_n580# 0.48fF
C187 op unit_cap_mim_m3m4_31/m3_n630_n580# 0.03fF
C188 p1_b unit_cap_mim_m3m4_17/m3_n630_n580# 0.06fF
C189 p2 p1 2.82fF
C190 transmission_gate_8/in p1 0.39fF
C191 op unit_cap_mim_m3m4_29/c1_n530_n480# 0.03fF
C192 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_31/c1_n530_n480# -0.25fF
C193 unit_cap_mim_m3m4_35/m3_n630_n580# p1 0.07fF
C194 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580# -0.37fF
C195 p1_b unit_cap_mim_m3m4_21/m3_n630_n580# 0.05fF
C196 p1_b transmission_gate_7/in 0.40fF
C197 unit_cap_mim_m3m4_21/c1_n530_n480# on 0.06fF
C198 p1_b p2_b 2.92fF
C199 p1_b unit_cap_mim_m3m4_29/m3_n630_n580# 0.05fF
C200 transmission_gate_9/in op 0.47fF
C201 transmission_gate_8/in unit_cap_mim_m3m4_28/m3_n630_n580# 0.10fF
C202 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C203 bias_a p1 0.81fF
C204 transmission_gate_4/out transmission_gate_6/in 0.48fF
C205 p2_b transmission_gate_7/in 0.41fF
C206 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480# -0.20fF
C207 p2 unit_cap_mim_m3m4_29/c1_n530_n480# 0.04fF
C208 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C209 transmission_gate_9/in VDD -0.11fF
C210 unit_cap_mim_m3m4_22/c1_n530_n480# cmc 0.13fF
C211 transmission_gate_4/out transmission_gate_3/out 0.38fF
C212 p1_b cmc 0.53fF
C213 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_34/m3_n630_n580# 0.17fF
C214 unit_cap_mim_m3m4_17/m3_n630_n580# cmc 0.17fF
C215 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580# -0.19fF
C216 transmission_gate_9/in p2 0.14fF
C217 p1_b cm 1.15fF
C218 transmission_gate_9/in transmission_gate_8/in 0.93fF
C219 unit_cap_mim_m3m4_16/m3_n630_n580# p1_b 0.06fF
C220 op transmission_gate_6/in 0.61fF
C221 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.12fF
C222 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C223 cmc unit_cap_mim_m3m4_21/m3_n630_n580# 0.69fF
C224 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C225 transmission_gate_7/in cmc 0.11fF
C226 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.12fF
C227 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580# -0.20fF
C228 p2_b cmc 0.12fF
C229 unit_cap_mim_m3m4_27/c1_n530_n480# transmission_gate_6/in -0.13fF
C230 transmission_gate_7/in cm 0.10fF
C231 p2_b cm 1.01fF
C232 op transmission_gate_3/out 0.57fF
C233 VDD transmission_gate_6/in 0.03fF
C234 on unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C235 transmission_gate_9/in bias_a 0.02fF
C236 transmission_gate_8/in unit_cap_mim_m3m4_34/m3_n630_n580# 0.38fF
C237 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_34/m3_n630_n580# 0.17fF
C238 p1_b on 0.45fF
C239 unit_cap_mim_m3m4_26/c1_n530_n480# p1 0.11fF
C240 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580# 0.12fF
C241 transmission_gate_6/in p2 0.61fF
C242 transmission_gate_8/in transmission_gate_6/in -0.41fF
C243 p1_b p1 8.88fF
C244 unit_cap_mim_m3m4_17/m3_n630_n580# p1 0.08fF
C245 transmission_gate_3/out VDD -0.05fF
C246 on transmission_gate_7/in 3.15fF
C247 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_16/c1_n530_n480# -0.21fF
C248 on unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C249 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C250 unit_cap_mim_m3m4_21/m3_n630_n580# p1 0.06fF
C251 p2_b on 0.34fF
C252 transmission_gate_3/out p2 0.15fF
C253 transmission_gate_8/in transmission_gate_3/out 0.16fF
C254 transmission_gate_7/in p1 0.39fF
C255 unit_cap_mim_m3m4_19/c1_n530_n480# transmission_gate_7/in 0.06fF
C256 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C257 p2_b p1 2.16fF
C258 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580# -0.32fF
C259 unit_cap_mim_m3m4_29/m3_n630_n580# p1 0.06fF
C260 transmission_gate_6/in bias_a 0.07fF
C261 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_24/c1_n530_n480# -0.30fF
C262 p1_b unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C263 unit_cap_mim_m3m4_28/c1_n530_n480# op 0.17fF
C264 transmission_gate_3/out bias_a 0.07fF
C265 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.17fF
C266 on cmc -0.58fF
C267 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C268 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C269 transmission_gate_9/in unit_cap_mim_m3m4_22/c1_n530_n480# -0.37fF
C270 cmc p1 0.49fF
C271 transmission_gate_9/in p1_b 0.59fF
C272 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_29/c1_n530_n480# -0.29fF
C273 cm p1 1.50fF
C274 unit_cap_mim_m3m4_16/m3_n630_n580# p1 0.08fF
C275 unit_cap_mim_m3m4_24/m3_n630_n580# p2 0.05fF
C276 transmission_gate_9/in transmission_gate_7/in 0.04fF
C277 transmission_gate_4/out unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C278 unit_cap_mim_m3m4_28/c1_n530_n480# p2 0.04fF
C279 op unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C280 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_33/c1_n530_n480# -0.18fF
C281 transmission_gate_9/in p2_b 0.01fF
C282 cmc unit_cap_mim_m3m4_27/m3_n630_n580# 0.10fF
C283 transmission_gate_4/out unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C284 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580# -0.20fF
C285 p1_b transmission_gate_6/in 0.41fF
C286 on p1 0.49fF
C287 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_20/c1_n530_n480# -0.19fF
C288 unit_cap_mim_m3m4_23/c1_n530_n480# op 0.13fF
C289 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C290 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.39fF
C291 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C292 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.51fF
C293 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C294 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.74fF
C295 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C296 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.51fF
C297 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.51fF
C298 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.82fF
C299 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.60fF
C300 cmc VSS 7.45fF
C301 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.61fF
C302 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.61fF
C303 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C304 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C305 p2 VSS 148.24fF
C306 p2_b VSS 41.62fF
C307 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.84fF
C308 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C309 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.39fF
C310 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C311 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.04fF
C312 transmission_gate_9/in VSS 2.27fF
C313 transmission_gate_4/out VSS -3.31fF
C314 transmission_gate_3/out VSS 2.40fF
C315 transmission_gate_8/in VSS -2.63fF
C316 bias_a VSS 11.61fF
C317 transmission_gate_6/in VSS -13.21fF
C318 transmission_gate_7/in VSS 8.85fF
C319 cm VSS 13.12fF
C320 p1 VSS 111.99fF
C321 op VSS 0.25fF
C322 p1_b VSS 173.74fF
C323 VDD VSS 71.01fF
C324 on VSS -22.35fF
.ends

