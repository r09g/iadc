magic
tech sky130A
timestamp 1654711401
<< error_p >>
rect -765 290 -736 293
rect -686 290 -657 293
rect -607 290 -578 293
rect -528 290 -499 293
rect -449 290 -420 293
rect -370 290 -341 293
rect -291 290 -262 293
rect -212 290 -183 293
rect -133 290 -104 293
rect -54 290 -25 293
rect 25 290 54 293
rect 104 290 133 293
rect 183 290 212 293
rect 262 290 291 293
rect 341 290 370 293
rect 420 290 449 293
rect 499 290 528 293
rect 578 290 607 293
rect 657 290 686 293
rect 736 290 765 293
rect -765 273 -759 290
rect -686 273 -680 290
rect -607 273 -601 290
rect -528 273 -522 290
rect -449 273 -443 290
rect -370 273 -364 290
rect -291 273 -285 290
rect -212 273 -206 290
rect -133 273 -127 290
rect -54 273 -48 290
rect 25 273 31 290
rect 104 273 110 290
rect 183 273 189 290
rect 262 273 268 290
rect 341 273 347 290
rect 420 273 426 290
rect 499 273 505 290
rect 578 273 584 290
rect 657 273 663 290
rect 736 273 742 290
rect -765 270 -736 273
rect -686 270 -657 273
rect -607 270 -578 273
rect -528 270 -499 273
rect -449 270 -420 273
rect -370 270 -341 273
rect -291 270 -262 273
rect -212 270 -183 273
rect -133 270 -104 273
rect -54 270 -25 273
rect 25 270 54 273
rect 104 270 133 273
rect 183 270 212 273
rect 262 270 291 273
rect 341 270 370 273
rect 420 270 449 273
rect 499 270 528 273
rect 578 270 607 273
rect 657 270 686 273
rect 736 270 765 273
rect -765 -273 -736 -270
rect -686 -273 -657 -270
rect -607 -273 -578 -270
rect -528 -273 -499 -270
rect -449 -273 -420 -270
rect -370 -273 -341 -270
rect -291 -273 -262 -270
rect -212 -273 -183 -270
rect -133 -273 -104 -270
rect -54 -273 -25 -270
rect 25 -273 54 -270
rect 104 -273 133 -270
rect 183 -273 212 -270
rect 262 -273 291 -270
rect 341 -273 370 -270
rect 420 -273 449 -270
rect 499 -273 528 -270
rect 578 -273 607 -270
rect 657 -273 686 -270
rect 736 -273 765 -270
rect -765 -290 -759 -273
rect -686 -290 -680 -273
rect -607 -290 -601 -273
rect -528 -290 -522 -273
rect -449 -290 -443 -273
rect -370 -290 -364 -273
rect -291 -290 -285 -273
rect -212 -290 -206 -273
rect -133 -290 -127 -273
rect -54 -290 -48 -273
rect 25 -290 31 -273
rect 104 -290 110 -273
rect 183 -290 189 -273
rect 262 -290 268 -273
rect 341 -290 347 -273
rect 420 -290 426 -273
rect 499 -290 505 -273
rect 578 -290 584 -273
rect 657 -290 663 -273
rect 736 -290 742 -273
rect -765 -293 -736 -290
rect -686 -293 -657 -290
rect -607 -293 -578 -290
rect -528 -293 -499 -290
rect -449 -293 -420 -290
rect -370 -293 -341 -290
rect -291 -293 -262 -290
rect -212 -293 -183 -290
rect -133 -293 -104 -290
rect -54 -293 -25 -290
rect 25 -293 54 -290
rect 104 -293 133 -290
rect 183 -293 212 -290
rect 262 -293 291 -290
rect 341 -293 370 -290
rect 420 -293 449 -290
rect 499 -293 528 -290
rect 578 -293 607 -290
rect 657 -293 686 -290
rect 736 -293 765 -290
<< nwell >>
rect -904 -398 904 398
<< mvpmos >>
rect -775 -250 -725 250
rect -696 -250 -646 250
rect -617 -250 -567 250
rect -538 -250 -488 250
rect -459 -250 -409 250
rect -380 -250 -330 250
rect -301 -250 -251 250
rect -222 -250 -172 250
rect -143 -250 -93 250
rect -64 -250 -14 250
rect 14 -250 64 250
rect 93 -250 143 250
rect 172 -250 222 250
rect 251 -250 301 250
rect 330 -250 380 250
rect 409 -250 459 250
rect 488 -250 538 250
rect 567 -250 617 250
rect 646 -250 696 250
rect 725 -250 775 250
<< mvpdiff >>
rect -804 244 -775 250
rect -804 -244 -798 244
rect -781 -244 -775 244
rect -804 -250 -775 -244
rect -725 244 -696 250
rect -725 -244 -719 244
rect -702 -244 -696 244
rect -725 -250 -696 -244
rect -646 244 -617 250
rect -646 -244 -640 244
rect -623 -244 -617 244
rect -646 -250 -617 -244
rect -567 244 -538 250
rect -567 -244 -561 244
rect -544 -244 -538 244
rect -567 -250 -538 -244
rect -488 244 -459 250
rect -488 -244 -482 244
rect -465 -244 -459 244
rect -488 -250 -459 -244
rect -409 244 -380 250
rect -409 -244 -403 244
rect -386 -244 -380 244
rect -409 -250 -380 -244
rect -330 244 -301 250
rect -330 -244 -324 244
rect -307 -244 -301 244
rect -330 -250 -301 -244
rect -251 244 -222 250
rect -251 -244 -245 244
rect -228 -244 -222 244
rect -251 -250 -222 -244
rect -172 244 -143 250
rect -172 -244 -166 244
rect -149 -244 -143 244
rect -172 -250 -143 -244
rect -93 244 -64 250
rect -93 -244 -87 244
rect -70 -244 -64 244
rect -93 -250 -64 -244
rect -14 244 14 250
rect -14 -244 -8 244
rect 8 -244 14 244
rect -14 -250 14 -244
rect 64 244 93 250
rect 64 -244 70 244
rect 87 -244 93 244
rect 64 -250 93 -244
rect 143 244 172 250
rect 143 -244 149 244
rect 166 -244 172 244
rect 143 -250 172 -244
rect 222 244 251 250
rect 222 -244 228 244
rect 245 -244 251 244
rect 222 -250 251 -244
rect 301 244 330 250
rect 301 -244 307 244
rect 324 -244 330 244
rect 301 -250 330 -244
rect 380 244 409 250
rect 380 -244 386 244
rect 403 -244 409 244
rect 380 -250 409 -244
rect 459 244 488 250
rect 459 -244 465 244
rect 482 -244 488 244
rect 459 -250 488 -244
rect 538 244 567 250
rect 538 -244 544 244
rect 561 -244 567 244
rect 538 -250 567 -244
rect 617 244 646 250
rect 617 -244 623 244
rect 640 -244 646 244
rect 617 -250 646 -244
rect 696 244 725 250
rect 696 -244 702 244
rect 719 -244 725 244
rect 696 -250 725 -244
rect 775 244 804 250
rect 775 -244 781 244
rect 798 -244 804 244
rect 775 -250 804 -244
<< mvpdiffc >>
rect -798 -244 -781 244
rect -719 -244 -702 244
rect -640 -244 -623 244
rect -561 -244 -544 244
rect -482 -244 -465 244
rect -403 -244 -386 244
rect -324 -244 -307 244
rect -245 -244 -228 244
rect -166 -244 -149 244
rect -87 -244 -70 244
rect -8 -244 8 244
rect 70 -244 87 244
rect 149 -244 166 244
rect 228 -244 245 244
rect 307 -244 324 244
rect 386 -244 403 244
rect 465 -244 482 244
rect 544 -244 561 244
rect 623 -244 640 244
rect 702 -244 719 244
rect 781 -244 798 244
<< mvnsubdiff >>
rect -871 359 871 365
rect -871 342 -817 359
rect 817 342 871 359
rect -871 336 871 342
rect -871 311 -842 336
rect -871 -311 -865 311
rect -848 -311 -842 311
rect 842 311 871 336
rect -871 -336 -842 -311
rect 842 -311 848 311
rect 865 -311 871 311
rect 842 -336 871 -311
rect -871 -342 871 -336
rect -871 -359 -817 -342
rect 817 -359 871 -342
rect -871 -365 871 -359
<< mvnsubdiffcont >>
rect -817 342 817 359
rect -865 -311 -848 311
rect 848 -311 865 311
rect -817 -359 817 -342
<< poly >>
rect -775 290 -725 298
rect -775 273 -767 290
rect -733 273 -725 290
rect -775 250 -725 273
rect -696 290 -646 298
rect -696 273 -688 290
rect -654 273 -646 290
rect -696 250 -646 273
rect -617 290 -567 298
rect -617 273 -609 290
rect -575 273 -567 290
rect -617 250 -567 273
rect -538 290 -488 298
rect -538 273 -530 290
rect -496 273 -488 290
rect -538 250 -488 273
rect -459 290 -409 298
rect -459 273 -451 290
rect -417 273 -409 290
rect -459 250 -409 273
rect -380 290 -330 298
rect -380 273 -372 290
rect -338 273 -330 290
rect -380 250 -330 273
rect -301 290 -251 298
rect -301 273 -293 290
rect -259 273 -251 290
rect -301 250 -251 273
rect -222 290 -172 298
rect -222 273 -214 290
rect -180 273 -172 290
rect -222 250 -172 273
rect -143 290 -93 298
rect -143 273 -135 290
rect -101 273 -93 290
rect -143 250 -93 273
rect -64 290 -14 298
rect -64 273 -56 290
rect -22 273 -14 290
rect -64 250 -14 273
rect 14 290 64 298
rect 14 273 22 290
rect 56 273 64 290
rect 14 250 64 273
rect 93 290 143 298
rect 93 273 101 290
rect 135 273 143 290
rect 93 250 143 273
rect 172 290 222 298
rect 172 273 180 290
rect 214 273 222 290
rect 172 250 222 273
rect 251 290 301 298
rect 251 273 259 290
rect 293 273 301 290
rect 251 250 301 273
rect 330 290 380 298
rect 330 273 338 290
rect 372 273 380 290
rect 330 250 380 273
rect 409 290 459 298
rect 409 273 417 290
rect 451 273 459 290
rect 409 250 459 273
rect 488 290 538 298
rect 488 273 496 290
rect 530 273 538 290
rect 488 250 538 273
rect 567 290 617 298
rect 567 273 575 290
rect 609 273 617 290
rect 567 250 617 273
rect 646 290 696 298
rect 646 273 654 290
rect 688 273 696 290
rect 646 250 696 273
rect 725 290 775 298
rect 725 273 733 290
rect 767 273 775 290
rect 725 250 775 273
rect -775 -273 -725 -250
rect -775 -290 -767 -273
rect -733 -290 -725 -273
rect -775 -298 -725 -290
rect -696 -273 -646 -250
rect -696 -290 -688 -273
rect -654 -290 -646 -273
rect -696 -298 -646 -290
rect -617 -273 -567 -250
rect -617 -290 -609 -273
rect -575 -290 -567 -273
rect -617 -298 -567 -290
rect -538 -273 -488 -250
rect -538 -290 -530 -273
rect -496 -290 -488 -273
rect -538 -298 -488 -290
rect -459 -273 -409 -250
rect -459 -290 -451 -273
rect -417 -290 -409 -273
rect -459 -298 -409 -290
rect -380 -273 -330 -250
rect -380 -290 -372 -273
rect -338 -290 -330 -273
rect -380 -298 -330 -290
rect -301 -273 -251 -250
rect -301 -290 -293 -273
rect -259 -290 -251 -273
rect -301 -298 -251 -290
rect -222 -273 -172 -250
rect -222 -290 -214 -273
rect -180 -290 -172 -273
rect -222 -298 -172 -290
rect -143 -273 -93 -250
rect -143 -290 -135 -273
rect -101 -290 -93 -273
rect -143 -298 -93 -290
rect -64 -273 -14 -250
rect -64 -290 -56 -273
rect -22 -290 -14 -273
rect -64 -298 -14 -290
rect 14 -273 64 -250
rect 14 -290 22 -273
rect 56 -290 64 -273
rect 14 -298 64 -290
rect 93 -273 143 -250
rect 93 -290 101 -273
rect 135 -290 143 -273
rect 93 -298 143 -290
rect 172 -273 222 -250
rect 172 -290 180 -273
rect 214 -290 222 -273
rect 172 -298 222 -290
rect 251 -273 301 -250
rect 251 -290 259 -273
rect 293 -290 301 -273
rect 251 -298 301 -290
rect 330 -273 380 -250
rect 330 -290 338 -273
rect 372 -290 380 -273
rect 330 -298 380 -290
rect 409 -273 459 -250
rect 409 -290 417 -273
rect 451 -290 459 -273
rect 409 -298 459 -290
rect 488 -273 538 -250
rect 488 -290 496 -273
rect 530 -290 538 -273
rect 488 -298 538 -290
rect 567 -273 617 -250
rect 567 -290 575 -273
rect 609 -290 617 -273
rect 567 -298 617 -290
rect 646 -273 696 -250
rect 646 -290 654 -273
rect 688 -290 696 -273
rect 646 -298 696 -290
rect 725 -273 775 -250
rect 725 -290 733 -273
rect 767 -290 775 -273
rect 725 -298 775 -290
<< polycont >>
rect -767 273 -733 290
rect -688 273 -654 290
rect -609 273 -575 290
rect -530 273 -496 290
rect -451 273 -417 290
rect -372 273 -338 290
rect -293 273 -259 290
rect -214 273 -180 290
rect -135 273 -101 290
rect -56 273 -22 290
rect 22 273 56 290
rect 101 273 135 290
rect 180 273 214 290
rect 259 273 293 290
rect 338 273 372 290
rect 417 273 451 290
rect 496 273 530 290
rect 575 273 609 290
rect 654 273 688 290
rect 733 273 767 290
rect -767 -290 -733 -273
rect -688 -290 -654 -273
rect -609 -290 -575 -273
rect -530 -290 -496 -273
rect -451 -290 -417 -273
rect -372 -290 -338 -273
rect -293 -290 -259 -273
rect -214 -290 -180 -273
rect -135 -290 -101 -273
rect -56 -290 -22 -273
rect 22 -290 56 -273
rect 101 -290 135 -273
rect 180 -290 214 -273
rect 259 -290 293 -273
rect 338 -290 372 -273
rect 417 -290 451 -273
rect 496 -290 530 -273
rect 575 -290 609 -273
rect 654 -290 688 -273
rect 733 -290 767 -273
<< locali >>
rect -865 342 -817 359
rect 817 342 865 359
rect -865 311 -848 342
rect 848 311 865 342
rect -775 273 -767 290
rect -733 273 -725 290
rect -696 273 -688 290
rect -654 273 -646 290
rect -617 273 -609 290
rect -575 273 -567 290
rect -538 273 -530 290
rect -496 273 -488 290
rect -459 273 -451 290
rect -417 273 -409 290
rect -380 273 -372 290
rect -338 273 -330 290
rect -301 273 -293 290
rect -259 273 -251 290
rect -222 273 -214 290
rect -180 273 -172 290
rect -143 273 -135 290
rect -101 273 -93 290
rect -64 273 -56 290
rect -22 273 -14 290
rect 14 273 22 290
rect 56 273 64 290
rect 93 273 101 290
rect 135 273 143 290
rect 172 273 180 290
rect 214 273 222 290
rect 251 273 259 290
rect 293 273 301 290
rect 330 273 338 290
rect 372 273 380 290
rect 409 273 417 290
rect 451 273 459 290
rect 488 273 496 290
rect 530 273 538 290
rect 567 273 575 290
rect 609 273 617 290
rect 646 273 654 290
rect 688 273 696 290
rect 725 273 733 290
rect 767 273 775 290
rect -798 244 -781 252
rect -798 -252 -781 -244
rect -719 244 -702 252
rect -719 -252 -702 -244
rect -640 244 -623 252
rect -640 -252 -623 -244
rect -561 244 -544 252
rect -561 -252 -544 -244
rect -482 244 -465 252
rect -482 -252 -465 -244
rect -403 244 -386 252
rect -403 -252 -386 -244
rect -324 244 -307 252
rect -324 -252 -307 -244
rect -245 244 -228 252
rect -245 -252 -228 -244
rect -166 244 -149 252
rect -166 -252 -149 -244
rect -87 244 -70 252
rect -87 -252 -70 -244
rect -8 244 8 252
rect -8 -252 8 -244
rect 70 244 87 252
rect 70 -252 87 -244
rect 149 244 166 252
rect 149 -252 166 -244
rect 228 244 245 252
rect 228 -252 245 -244
rect 307 244 324 252
rect 307 -252 324 -244
rect 386 244 403 252
rect 386 -252 403 -244
rect 465 244 482 252
rect 465 -252 482 -244
rect 544 244 561 252
rect 544 -252 561 -244
rect 623 244 640 252
rect 623 -252 640 -244
rect 702 244 719 252
rect 702 -252 719 -244
rect 781 244 798 252
rect 781 -252 798 -244
rect -775 -290 -767 -273
rect -733 -290 -725 -273
rect -696 -290 -688 -273
rect -654 -290 -646 -273
rect -617 -290 -609 -273
rect -575 -290 -567 -273
rect -538 -290 -530 -273
rect -496 -290 -488 -273
rect -459 -290 -451 -273
rect -417 -290 -409 -273
rect -380 -290 -372 -273
rect -338 -290 -330 -273
rect -301 -290 -293 -273
rect -259 -290 -251 -273
rect -222 -290 -214 -273
rect -180 -290 -172 -273
rect -143 -290 -135 -273
rect -101 -290 -93 -273
rect -64 -290 -56 -273
rect -22 -290 -14 -273
rect 14 -290 22 -273
rect 56 -290 64 -273
rect 93 -290 101 -273
rect 135 -290 143 -273
rect 172 -290 180 -273
rect 214 -290 222 -273
rect 251 -290 259 -273
rect 293 -290 301 -273
rect 330 -290 338 -273
rect 372 -290 380 -273
rect 409 -290 417 -273
rect 451 -290 459 -273
rect 488 -290 496 -273
rect 530 -290 538 -273
rect 567 -290 575 -273
rect 609 -290 617 -273
rect 646 -290 654 -273
rect 688 -290 696 -273
rect 725 -290 733 -273
rect 767 -290 775 -273
rect -865 -342 -848 -311
rect 848 -342 865 -311
rect -865 -359 -817 -342
rect 817 -359 865 -342
<< viali >>
rect -759 273 -742 290
rect -680 273 -663 290
rect -601 273 -584 290
rect -522 273 -505 290
rect -443 273 -426 290
rect -364 273 -347 290
rect -285 273 -268 290
rect -206 273 -189 290
rect -127 273 -110 290
rect -48 273 -31 290
rect 31 273 48 290
rect 110 273 127 290
rect 189 273 206 290
rect 268 273 285 290
rect 347 273 364 290
rect 426 273 443 290
rect 505 273 522 290
rect 584 273 601 290
rect 663 273 680 290
rect 742 273 759 290
rect -798 -244 -781 244
rect -719 -244 -702 244
rect -640 -244 -623 244
rect -561 -244 -544 244
rect -482 -244 -465 244
rect -403 -244 -386 244
rect -324 -244 -307 244
rect -245 -244 -228 244
rect -166 -244 -149 244
rect -87 -244 -70 244
rect -8 -244 8 244
rect 70 -244 87 244
rect 149 -244 166 244
rect 228 -244 245 244
rect 307 -244 324 244
rect 386 -244 403 244
rect 465 -244 482 244
rect 544 -244 561 244
rect 623 -244 640 244
rect 702 -244 719 244
rect 781 -244 798 244
rect -759 -290 -742 -273
rect -680 -290 -663 -273
rect -601 -290 -584 -273
rect -522 -290 -505 -273
rect -443 -290 -426 -273
rect -364 -290 -347 -273
rect -285 -290 -268 -273
rect -206 -290 -189 -273
rect -127 -290 -110 -273
rect -48 -290 -31 -273
rect 31 -290 48 -273
rect 110 -290 127 -273
rect 189 -290 206 -273
rect 268 -290 285 -273
rect 347 -290 364 -273
rect 426 -290 443 -273
rect 505 -290 522 -273
rect 584 -290 601 -273
rect 663 -290 680 -273
rect 742 -290 759 -273
<< metal1 >>
rect -765 290 -736 293
rect -765 273 -759 290
rect -742 273 -736 290
rect -765 270 -736 273
rect -686 290 -657 293
rect -686 273 -680 290
rect -663 273 -657 290
rect -686 270 -657 273
rect -607 290 -578 293
rect -607 273 -601 290
rect -584 273 -578 290
rect -607 270 -578 273
rect -528 290 -499 293
rect -528 273 -522 290
rect -505 273 -499 290
rect -528 270 -499 273
rect -449 290 -420 293
rect -449 273 -443 290
rect -426 273 -420 290
rect -449 270 -420 273
rect -370 290 -341 293
rect -370 273 -364 290
rect -347 273 -341 290
rect -370 270 -341 273
rect -291 290 -262 293
rect -291 273 -285 290
rect -268 273 -262 290
rect -291 270 -262 273
rect -212 290 -183 293
rect -212 273 -206 290
rect -189 273 -183 290
rect -212 270 -183 273
rect -133 290 -104 293
rect -133 273 -127 290
rect -110 273 -104 290
rect -133 270 -104 273
rect -54 290 -25 293
rect -54 273 -48 290
rect -31 273 -25 290
rect -54 270 -25 273
rect 25 290 54 293
rect 25 273 31 290
rect 48 273 54 290
rect 25 270 54 273
rect 104 290 133 293
rect 104 273 110 290
rect 127 273 133 290
rect 104 270 133 273
rect 183 290 212 293
rect 183 273 189 290
rect 206 273 212 290
rect 183 270 212 273
rect 262 290 291 293
rect 262 273 268 290
rect 285 273 291 290
rect 262 270 291 273
rect 341 290 370 293
rect 341 273 347 290
rect 364 273 370 290
rect 341 270 370 273
rect 420 290 449 293
rect 420 273 426 290
rect 443 273 449 290
rect 420 270 449 273
rect 499 290 528 293
rect 499 273 505 290
rect 522 273 528 290
rect 499 270 528 273
rect 578 290 607 293
rect 578 273 584 290
rect 601 273 607 290
rect 578 270 607 273
rect 657 290 686 293
rect 657 273 663 290
rect 680 273 686 290
rect 657 270 686 273
rect 736 290 765 293
rect 736 273 742 290
rect 759 273 765 290
rect 736 270 765 273
rect -801 244 -778 250
rect -801 -244 -798 244
rect -781 -244 -778 244
rect -801 -250 -778 -244
rect -722 244 -699 250
rect -722 -244 -719 244
rect -702 -244 -699 244
rect -722 -250 -699 -244
rect -643 244 -620 250
rect -643 -244 -640 244
rect -623 -244 -620 244
rect -643 -250 -620 -244
rect -564 244 -541 250
rect -564 -244 -561 244
rect -544 -244 -541 244
rect -564 -250 -541 -244
rect -485 244 -462 250
rect -485 -244 -482 244
rect -465 -244 -462 244
rect -485 -250 -462 -244
rect -406 244 -383 250
rect -406 -244 -403 244
rect -386 -244 -383 244
rect -406 -250 -383 -244
rect -327 244 -304 250
rect -327 -244 -324 244
rect -307 -244 -304 244
rect -327 -250 -304 -244
rect -248 244 -225 250
rect -248 -244 -245 244
rect -228 -244 -225 244
rect -248 -250 -225 -244
rect -169 244 -146 250
rect -169 -244 -166 244
rect -149 -244 -146 244
rect -169 -250 -146 -244
rect -90 244 -67 250
rect -90 -244 -87 244
rect -70 -244 -67 244
rect -90 -250 -67 -244
rect -11 244 11 250
rect -11 -244 -8 244
rect 8 -244 11 244
rect -11 -250 11 -244
rect 67 244 90 250
rect 67 -244 70 244
rect 87 -244 90 244
rect 67 -250 90 -244
rect 146 244 169 250
rect 146 -244 149 244
rect 166 -244 169 244
rect 146 -250 169 -244
rect 225 244 248 250
rect 225 -244 228 244
rect 245 -244 248 244
rect 225 -250 248 -244
rect 304 244 327 250
rect 304 -244 307 244
rect 324 -244 327 244
rect 304 -250 327 -244
rect 383 244 406 250
rect 383 -244 386 244
rect 403 -244 406 244
rect 383 -250 406 -244
rect 462 244 485 250
rect 462 -244 465 244
rect 482 -244 485 244
rect 462 -250 485 -244
rect 541 244 564 250
rect 541 -244 544 244
rect 561 -244 564 244
rect 541 -250 564 -244
rect 620 244 643 250
rect 620 -244 623 244
rect 640 -244 643 244
rect 620 -250 643 -244
rect 699 244 722 250
rect 699 -244 702 244
rect 719 -244 722 244
rect 699 -250 722 -244
rect 778 244 801 250
rect 778 -244 781 244
rect 798 -244 801 244
rect 778 -250 801 -244
rect -765 -273 -736 -270
rect -765 -290 -759 -273
rect -742 -290 -736 -273
rect -765 -293 -736 -290
rect -686 -273 -657 -270
rect -686 -290 -680 -273
rect -663 -290 -657 -273
rect -686 -293 -657 -290
rect -607 -273 -578 -270
rect -607 -290 -601 -273
rect -584 -290 -578 -273
rect -607 -293 -578 -290
rect -528 -273 -499 -270
rect -528 -290 -522 -273
rect -505 -290 -499 -273
rect -528 -293 -499 -290
rect -449 -273 -420 -270
rect -449 -290 -443 -273
rect -426 -290 -420 -273
rect -449 -293 -420 -290
rect -370 -273 -341 -270
rect -370 -290 -364 -273
rect -347 -290 -341 -273
rect -370 -293 -341 -290
rect -291 -273 -262 -270
rect -291 -290 -285 -273
rect -268 -290 -262 -273
rect -291 -293 -262 -290
rect -212 -273 -183 -270
rect -212 -290 -206 -273
rect -189 -290 -183 -273
rect -212 -293 -183 -290
rect -133 -273 -104 -270
rect -133 -290 -127 -273
rect -110 -290 -104 -273
rect -133 -293 -104 -290
rect -54 -273 -25 -270
rect -54 -290 -48 -273
rect -31 -290 -25 -273
rect -54 -293 -25 -290
rect 25 -273 54 -270
rect 25 -290 31 -273
rect 48 -290 54 -273
rect 25 -293 54 -290
rect 104 -273 133 -270
rect 104 -290 110 -273
rect 127 -290 133 -273
rect 104 -293 133 -290
rect 183 -273 212 -270
rect 183 -290 189 -273
rect 206 -290 212 -273
rect 183 -293 212 -290
rect 262 -273 291 -270
rect 262 -290 268 -273
rect 285 -290 291 -273
rect 262 -293 291 -290
rect 341 -273 370 -270
rect 341 -290 347 -273
rect 364 -290 370 -273
rect 341 -293 370 -290
rect 420 -273 449 -270
rect 420 -290 426 -273
rect 443 -290 449 -273
rect 420 -293 449 -290
rect 499 -273 528 -270
rect 499 -290 505 -273
rect 522 -290 528 -273
rect 499 -293 528 -290
rect 578 -273 607 -270
rect 578 -290 584 -273
rect 601 -290 607 -273
rect 578 -293 607 -290
rect 657 -273 686 -270
rect 657 -290 663 -273
rect 680 -290 686 -273
rect 657 -293 686 -290
rect 736 -273 765 -270
rect 736 -290 742 -273
rect 759 -290 765 -273
rect 736 -293 765 -290
<< properties >>
string FIXED_BBOX -857 -351 857 351
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
