magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< pwell >>
rect -1034 -166 1034 166
<< nmos >>
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
<< ndiff >>
rect -1008 119 -950 140
rect -1008 85 -996 119
rect -962 85 -950 119
rect -1008 51 -950 85
rect -1008 17 -996 51
rect -962 17 -950 51
rect -1008 -17 -950 17
rect -1008 -51 -996 -17
rect -962 -51 -950 -17
rect -1008 -85 -950 -51
rect -1008 -119 -996 -85
rect -962 -119 -950 -85
rect -1008 -140 -950 -119
rect -830 119 -772 140
rect -830 85 -818 119
rect -784 85 -772 119
rect -830 51 -772 85
rect -830 17 -818 51
rect -784 17 -772 51
rect -830 -17 -772 17
rect -830 -51 -818 -17
rect -784 -51 -772 -17
rect -830 -85 -772 -51
rect -830 -119 -818 -85
rect -784 -119 -772 -85
rect -830 -140 -772 -119
rect -652 119 -594 140
rect -652 85 -640 119
rect -606 85 -594 119
rect -652 51 -594 85
rect -652 17 -640 51
rect -606 17 -594 51
rect -652 -17 -594 17
rect -652 -51 -640 -17
rect -606 -51 -594 -17
rect -652 -85 -594 -51
rect -652 -119 -640 -85
rect -606 -119 -594 -85
rect -652 -140 -594 -119
rect -474 119 -416 140
rect -474 85 -462 119
rect -428 85 -416 119
rect -474 51 -416 85
rect -474 17 -462 51
rect -428 17 -416 51
rect -474 -17 -416 17
rect -474 -51 -462 -17
rect -428 -51 -416 -17
rect -474 -85 -416 -51
rect -474 -119 -462 -85
rect -428 -119 -416 -85
rect -474 -140 -416 -119
rect -296 119 -238 140
rect -296 85 -284 119
rect -250 85 -238 119
rect -296 51 -238 85
rect -296 17 -284 51
rect -250 17 -238 51
rect -296 -17 -238 17
rect -296 -51 -284 -17
rect -250 -51 -238 -17
rect -296 -85 -238 -51
rect -296 -119 -284 -85
rect -250 -119 -238 -85
rect -296 -140 -238 -119
rect -118 119 -60 140
rect -118 85 -106 119
rect -72 85 -60 119
rect -118 51 -60 85
rect -118 17 -106 51
rect -72 17 -60 51
rect -118 -17 -60 17
rect -118 -51 -106 -17
rect -72 -51 -60 -17
rect -118 -85 -60 -51
rect -118 -119 -106 -85
rect -72 -119 -60 -85
rect -118 -140 -60 -119
rect 60 119 118 140
rect 60 85 72 119
rect 106 85 118 119
rect 60 51 118 85
rect 60 17 72 51
rect 106 17 118 51
rect 60 -17 118 17
rect 60 -51 72 -17
rect 106 -51 118 -17
rect 60 -85 118 -51
rect 60 -119 72 -85
rect 106 -119 118 -85
rect 60 -140 118 -119
rect 238 119 296 140
rect 238 85 250 119
rect 284 85 296 119
rect 238 51 296 85
rect 238 17 250 51
rect 284 17 296 51
rect 238 -17 296 17
rect 238 -51 250 -17
rect 284 -51 296 -17
rect 238 -85 296 -51
rect 238 -119 250 -85
rect 284 -119 296 -85
rect 238 -140 296 -119
rect 416 119 474 140
rect 416 85 428 119
rect 462 85 474 119
rect 416 51 474 85
rect 416 17 428 51
rect 462 17 474 51
rect 416 -17 474 17
rect 416 -51 428 -17
rect 462 -51 474 -17
rect 416 -85 474 -51
rect 416 -119 428 -85
rect 462 -119 474 -85
rect 416 -140 474 -119
rect 594 119 652 140
rect 594 85 606 119
rect 640 85 652 119
rect 594 51 652 85
rect 594 17 606 51
rect 640 17 652 51
rect 594 -17 652 17
rect 594 -51 606 -17
rect 640 -51 652 -17
rect 594 -85 652 -51
rect 594 -119 606 -85
rect 640 -119 652 -85
rect 594 -140 652 -119
rect 772 119 830 140
rect 772 85 784 119
rect 818 85 830 119
rect 772 51 830 85
rect 772 17 784 51
rect 818 17 830 51
rect 772 -17 830 17
rect 772 -51 784 -17
rect 818 -51 830 -17
rect 772 -85 830 -51
rect 772 -119 784 -85
rect 818 -119 830 -85
rect 772 -140 830 -119
rect 950 119 1008 140
rect 950 85 962 119
rect 996 85 1008 119
rect 950 51 1008 85
rect 950 17 962 51
rect 996 17 1008 51
rect 950 -17 1008 17
rect 950 -51 962 -17
rect 996 -51 1008 -17
rect 950 -85 1008 -51
rect 950 -119 962 -85
rect 996 -119 1008 -85
rect 950 -140 1008 -119
<< ndiffc >>
rect -996 85 -962 119
rect -996 17 -962 51
rect -996 -51 -962 -17
rect -996 -119 -962 -85
rect -818 85 -784 119
rect -818 17 -784 51
rect -818 -51 -784 -17
rect -818 -119 -784 -85
rect -640 85 -606 119
rect -640 17 -606 51
rect -640 -51 -606 -17
rect -640 -119 -606 -85
rect -462 85 -428 119
rect -462 17 -428 51
rect -462 -51 -428 -17
rect -462 -119 -428 -85
rect -284 85 -250 119
rect -284 17 -250 51
rect -284 -51 -250 -17
rect -284 -119 -250 -85
rect -106 85 -72 119
rect -106 17 -72 51
rect -106 -51 -72 -17
rect -106 -119 -72 -85
rect 72 85 106 119
rect 72 17 106 51
rect 72 -51 106 -17
rect 72 -119 106 -85
rect 250 85 284 119
rect 250 17 284 51
rect 250 -51 284 -17
rect 250 -119 284 -85
rect 428 85 462 119
rect 428 17 462 51
rect 428 -51 462 -17
rect 428 -119 462 -85
rect 606 85 640 119
rect 606 17 640 51
rect 606 -51 640 -17
rect 606 -119 640 -85
rect 784 85 818 119
rect 784 17 818 51
rect 784 -51 818 -17
rect 784 -119 818 -85
rect 962 85 996 119
rect 962 17 996 51
rect 962 -51 996 -17
rect 962 -119 996 -85
<< poly >>
rect -928 212 -852 228
rect -928 194 -907 212
rect -950 178 -907 194
rect -873 194 -852 212
rect -750 212 -674 228
rect -750 194 -729 212
rect -873 178 -830 194
rect -950 140 -830 178
rect -772 178 -729 194
rect -695 194 -674 212
rect -572 212 -496 228
rect -572 194 -551 212
rect -695 178 -652 194
rect -772 140 -652 178
rect -594 178 -551 194
rect -517 194 -496 212
rect -394 212 -318 228
rect -394 194 -373 212
rect -517 178 -474 194
rect -594 140 -474 178
rect -416 178 -373 194
rect -339 194 -318 212
rect -216 212 -140 228
rect -216 194 -195 212
rect -339 178 -296 194
rect -416 140 -296 178
rect -238 178 -195 194
rect -161 194 -140 212
rect -38 212 38 228
rect -38 194 -17 212
rect -161 178 -118 194
rect -238 140 -118 178
rect -60 178 -17 194
rect 17 194 38 212
rect 140 212 216 228
rect 140 194 161 212
rect 17 178 60 194
rect -60 140 60 178
rect 118 178 161 194
rect 195 194 216 212
rect 318 212 394 228
rect 318 194 339 212
rect 195 178 238 194
rect 118 140 238 178
rect 296 178 339 194
rect 373 194 394 212
rect 496 212 572 228
rect 496 194 517 212
rect 373 178 416 194
rect 296 140 416 178
rect 474 178 517 194
rect 551 194 572 212
rect 674 212 750 228
rect 674 194 695 212
rect 551 178 594 194
rect 474 140 594 178
rect 652 178 695 194
rect 729 194 750 212
rect 852 212 928 228
rect 852 194 873 212
rect 729 178 772 194
rect 652 140 772 178
rect 830 178 873 194
rect 907 194 928 212
rect 907 178 950 194
rect 830 140 950 178
rect -950 -178 -830 -140
rect -950 -194 -907 -178
rect -928 -212 -907 -194
rect -873 -194 -830 -178
rect -772 -178 -652 -140
rect -772 -194 -729 -178
rect -873 -212 -852 -194
rect -928 -228 -852 -212
rect -750 -212 -729 -194
rect -695 -194 -652 -178
rect -594 -178 -474 -140
rect -594 -194 -551 -178
rect -695 -212 -674 -194
rect -750 -228 -674 -212
rect -572 -212 -551 -194
rect -517 -194 -474 -178
rect -416 -178 -296 -140
rect -416 -194 -373 -178
rect -517 -212 -496 -194
rect -572 -228 -496 -212
rect -394 -212 -373 -194
rect -339 -194 -296 -178
rect -238 -178 -118 -140
rect -238 -194 -195 -178
rect -339 -212 -318 -194
rect -394 -228 -318 -212
rect -216 -212 -195 -194
rect -161 -194 -118 -178
rect -60 -178 60 -140
rect -60 -194 -17 -178
rect -161 -212 -140 -194
rect -216 -228 -140 -212
rect -38 -212 -17 -194
rect 17 -194 60 -178
rect 118 -178 238 -140
rect 118 -194 161 -178
rect 17 -212 38 -194
rect -38 -228 38 -212
rect 140 -212 161 -194
rect 195 -194 238 -178
rect 296 -178 416 -140
rect 296 -194 339 -178
rect 195 -212 216 -194
rect 140 -228 216 -212
rect 318 -212 339 -194
rect 373 -194 416 -178
rect 474 -178 594 -140
rect 474 -194 517 -178
rect 373 -212 394 -194
rect 318 -228 394 -212
rect 496 -212 517 -194
rect 551 -194 594 -178
rect 652 -178 772 -140
rect 652 -194 695 -178
rect 551 -212 572 -194
rect 496 -228 572 -212
rect 674 -212 695 -194
rect 729 -194 772 -178
rect 830 -178 950 -140
rect 830 -194 873 -178
rect 729 -212 750 -194
rect 674 -228 750 -212
rect 852 -212 873 -194
rect 907 -194 950 -178
rect 907 -212 928 -194
rect 852 -228 928 -212
<< polycont >>
rect -907 178 -873 212
rect -729 178 -695 212
rect -551 178 -517 212
rect -373 178 -339 212
rect -195 178 -161 212
rect -17 178 17 212
rect 161 178 195 212
rect 339 178 373 212
rect 517 178 551 212
rect 695 178 729 212
rect 873 178 907 212
rect -907 -212 -873 -178
rect -729 -212 -695 -178
rect -551 -212 -517 -178
rect -373 -212 -339 -178
rect -195 -212 -161 -178
rect -17 -212 17 -178
rect 161 -212 195 -178
rect 339 -212 373 -178
rect 517 -212 551 -178
rect 695 -212 729 -178
rect 873 -212 907 -178
<< locali >>
rect -928 178 -907 212
rect -873 178 -852 212
rect -750 178 -729 212
rect -695 178 -674 212
rect -572 178 -551 212
rect -517 178 -496 212
rect -394 178 -373 212
rect -339 178 -318 212
rect -216 178 -195 212
rect -161 178 -140 212
rect -38 178 -17 212
rect 17 178 38 212
rect 140 178 161 212
rect 195 178 216 212
rect 318 178 339 212
rect 373 178 394 212
rect 496 178 517 212
rect 551 178 572 212
rect 674 178 695 212
rect 729 178 750 212
rect 852 178 873 212
rect 907 178 928 212
rect -996 125 -962 144
rect -996 53 -962 85
rect -996 -17 -962 17
rect -996 -85 -962 -53
rect -996 -144 -962 -125
rect -818 125 -784 144
rect -818 53 -784 85
rect -818 -17 -784 17
rect -818 -85 -784 -53
rect -818 -144 -784 -125
rect -640 125 -606 144
rect -640 53 -606 85
rect -640 -17 -606 17
rect -640 -85 -606 -53
rect -640 -144 -606 -125
rect -462 125 -428 144
rect -462 53 -428 85
rect -462 -17 -428 17
rect -462 -85 -428 -53
rect -462 -144 -428 -125
rect -284 125 -250 144
rect -284 53 -250 85
rect -284 -17 -250 17
rect -284 -85 -250 -53
rect -284 -144 -250 -125
rect -106 125 -72 144
rect -106 53 -72 85
rect -106 -17 -72 17
rect -106 -85 -72 -53
rect -106 -144 -72 -125
rect 72 125 106 144
rect 72 53 106 85
rect 72 -17 106 17
rect 72 -85 106 -53
rect 72 -144 106 -125
rect 250 125 284 144
rect 250 53 284 85
rect 250 -17 284 17
rect 250 -85 284 -53
rect 250 -144 284 -125
rect 428 125 462 144
rect 428 53 462 85
rect 428 -17 462 17
rect 428 -85 462 -53
rect 428 -144 462 -125
rect 606 125 640 144
rect 606 53 640 85
rect 606 -17 640 17
rect 606 -85 640 -53
rect 606 -144 640 -125
rect 784 125 818 144
rect 784 53 818 85
rect 784 -17 818 17
rect 784 -85 818 -53
rect 784 -144 818 -125
rect 962 125 996 144
rect 962 53 996 85
rect 962 -17 996 17
rect 962 -85 996 -53
rect 962 -144 996 -125
rect -928 -212 -907 -178
rect -873 -212 -852 -178
rect -750 -212 -729 -178
rect -695 -212 -674 -178
rect -572 -212 -551 -178
rect -517 -212 -496 -178
rect -394 -212 -373 -178
rect -339 -212 -318 -178
rect -216 -212 -195 -178
rect -161 -212 -140 -178
rect -38 -212 -17 -178
rect 17 -212 38 -178
rect 140 -212 161 -178
rect 195 -212 216 -178
rect 318 -212 339 -178
rect 373 -212 394 -178
rect 496 -212 517 -178
rect 551 -212 572 -178
rect 674 -212 695 -178
rect 729 -212 750 -178
rect 852 -212 873 -178
rect 907 -212 928 -178
<< viali >>
rect -907 178 -873 212
rect -729 178 -695 212
rect -551 178 -517 212
rect -373 178 -339 212
rect -195 178 -161 212
rect -17 178 17 212
rect 161 178 195 212
rect 339 178 373 212
rect 517 178 551 212
rect 695 178 729 212
rect 873 178 907 212
rect -996 119 -962 125
rect -996 91 -962 119
rect -996 51 -962 53
rect -996 19 -962 51
rect -996 -51 -962 -19
rect -996 -53 -962 -51
rect -996 -119 -962 -91
rect -996 -125 -962 -119
rect -818 119 -784 125
rect -818 91 -784 119
rect -818 51 -784 53
rect -818 19 -784 51
rect -818 -51 -784 -19
rect -818 -53 -784 -51
rect -818 -119 -784 -91
rect -818 -125 -784 -119
rect -640 119 -606 125
rect -640 91 -606 119
rect -640 51 -606 53
rect -640 19 -606 51
rect -640 -51 -606 -19
rect -640 -53 -606 -51
rect -640 -119 -606 -91
rect -640 -125 -606 -119
rect -462 119 -428 125
rect -462 91 -428 119
rect -462 51 -428 53
rect -462 19 -428 51
rect -462 -51 -428 -19
rect -462 -53 -428 -51
rect -462 -119 -428 -91
rect -462 -125 -428 -119
rect -284 119 -250 125
rect -284 91 -250 119
rect -284 51 -250 53
rect -284 19 -250 51
rect -284 -51 -250 -19
rect -284 -53 -250 -51
rect -284 -119 -250 -91
rect -284 -125 -250 -119
rect -106 119 -72 125
rect -106 91 -72 119
rect -106 51 -72 53
rect -106 19 -72 51
rect -106 -51 -72 -19
rect -106 -53 -72 -51
rect -106 -119 -72 -91
rect -106 -125 -72 -119
rect 72 119 106 125
rect 72 91 106 119
rect 72 51 106 53
rect 72 19 106 51
rect 72 -51 106 -19
rect 72 -53 106 -51
rect 72 -119 106 -91
rect 72 -125 106 -119
rect 250 119 284 125
rect 250 91 284 119
rect 250 51 284 53
rect 250 19 284 51
rect 250 -51 284 -19
rect 250 -53 284 -51
rect 250 -119 284 -91
rect 250 -125 284 -119
rect 428 119 462 125
rect 428 91 462 119
rect 428 51 462 53
rect 428 19 462 51
rect 428 -51 462 -19
rect 428 -53 462 -51
rect 428 -119 462 -91
rect 428 -125 462 -119
rect 606 119 640 125
rect 606 91 640 119
rect 606 51 640 53
rect 606 19 640 51
rect 606 -51 640 -19
rect 606 -53 640 -51
rect 606 -119 640 -91
rect 606 -125 640 -119
rect 784 119 818 125
rect 784 91 818 119
rect 784 51 818 53
rect 784 19 818 51
rect 784 -51 818 -19
rect 784 -53 818 -51
rect 784 -119 818 -91
rect 784 -125 818 -119
rect 962 119 996 125
rect 962 91 996 119
rect 962 51 996 53
rect 962 19 996 51
rect 962 -51 996 -19
rect 962 -53 996 -51
rect 962 -119 996 -91
rect 962 -125 996 -119
rect -907 -212 -873 -178
rect -729 -212 -695 -178
rect -551 -212 -517 -178
rect -373 -212 -339 -178
rect -195 -212 -161 -178
rect -17 -212 17 -178
rect 161 -212 195 -178
rect 339 -212 373 -178
rect 517 -212 551 -178
rect 695 -212 729 -178
rect 873 -212 907 -178
<< metal1 >>
rect -928 212 -852 228
rect -928 178 -907 212
rect -873 178 -852 212
rect -928 172 -852 178
rect -750 212 -674 228
rect -750 178 -729 212
rect -695 178 -674 212
rect -750 172 -674 178
rect -572 212 -496 228
rect -572 178 -551 212
rect -517 178 -496 212
rect -572 172 -496 178
rect -394 212 -318 228
rect -394 178 -373 212
rect -339 178 -318 212
rect -394 172 -318 178
rect -216 212 -140 228
rect -216 178 -195 212
rect -161 178 -140 212
rect -216 172 -140 178
rect -38 212 38 228
rect -38 178 -17 212
rect 17 178 38 212
rect -38 172 38 178
rect 140 212 216 228
rect 140 178 161 212
rect 195 178 216 212
rect 140 172 216 178
rect 318 212 394 228
rect 318 178 339 212
rect 373 178 394 212
rect 318 172 394 178
rect 496 212 572 228
rect 496 178 517 212
rect 551 178 572 212
rect 496 172 572 178
rect 674 212 750 228
rect 674 178 695 212
rect 729 178 750 212
rect 674 172 750 178
rect 852 212 928 228
rect 852 178 873 212
rect 907 178 928 212
rect 852 172 928 178
rect -1002 125 -956 140
rect -1002 91 -996 125
rect -962 91 -956 125
rect -1002 53 -956 91
rect -1002 19 -996 53
rect -962 19 -956 53
rect -1002 -19 -956 19
rect -1002 -53 -996 -19
rect -962 -53 -956 -19
rect -1002 -91 -956 -53
rect -1002 -125 -996 -91
rect -962 -125 -956 -91
rect -1002 -140 -956 -125
rect -824 125 -778 140
rect -824 91 -818 125
rect -784 91 -778 125
rect -824 53 -778 91
rect -824 19 -818 53
rect -784 19 -778 53
rect -824 -19 -778 19
rect -824 -53 -818 -19
rect -784 -53 -778 -19
rect -824 -91 -778 -53
rect -824 -125 -818 -91
rect -784 -125 -778 -91
rect -824 -140 -778 -125
rect -646 125 -600 140
rect -646 91 -640 125
rect -606 91 -600 125
rect -646 53 -600 91
rect -646 19 -640 53
rect -606 19 -600 53
rect -646 -19 -600 19
rect -646 -53 -640 -19
rect -606 -53 -600 -19
rect -646 -91 -600 -53
rect -646 -125 -640 -91
rect -606 -125 -600 -91
rect -646 -140 -600 -125
rect -468 125 -422 140
rect -468 91 -462 125
rect -428 91 -422 125
rect -468 53 -422 91
rect -468 19 -462 53
rect -428 19 -422 53
rect -468 -19 -422 19
rect -468 -53 -462 -19
rect -428 -53 -422 -19
rect -468 -91 -422 -53
rect -468 -125 -462 -91
rect -428 -125 -422 -91
rect -468 -140 -422 -125
rect -290 125 -244 140
rect -290 91 -284 125
rect -250 91 -244 125
rect -290 53 -244 91
rect -290 19 -284 53
rect -250 19 -244 53
rect -290 -19 -244 19
rect -290 -53 -284 -19
rect -250 -53 -244 -19
rect -290 -91 -244 -53
rect -290 -125 -284 -91
rect -250 -125 -244 -91
rect -290 -140 -244 -125
rect -112 125 -66 140
rect -112 91 -106 125
rect -72 91 -66 125
rect -112 53 -66 91
rect -112 19 -106 53
rect -72 19 -66 53
rect -112 -19 -66 19
rect -112 -53 -106 -19
rect -72 -53 -66 -19
rect -112 -91 -66 -53
rect -112 -125 -106 -91
rect -72 -125 -66 -91
rect -112 -140 -66 -125
rect 66 125 112 140
rect 66 91 72 125
rect 106 91 112 125
rect 66 53 112 91
rect 66 19 72 53
rect 106 19 112 53
rect 66 -19 112 19
rect 66 -53 72 -19
rect 106 -53 112 -19
rect 66 -91 112 -53
rect 66 -125 72 -91
rect 106 -125 112 -91
rect 66 -140 112 -125
rect 244 125 290 140
rect 244 91 250 125
rect 284 91 290 125
rect 244 53 290 91
rect 244 19 250 53
rect 284 19 290 53
rect 244 -19 290 19
rect 244 -53 250 -19
rect 284 -53 290 -19
rect 244 -91 290 -53
rect 244 -125 250 -91
rect 284 -125 290 -91
rect 244 -140 290 -125
rect 422 125 468 140
rect 422 91 428 125
rect 462 91 468 125
rect 422 53 468 91
rect 422 19 428 53
rect 462 19 468 53
rect 422 -19 468 19
rect 422 -53 428 -19
rect 462 -53 468 -19
rect 422 -91 468 -53
rect 422 -125 428 -91
rect 462 -125 468 -91
rect 422 -140 468 -125
rect 600 125 646 140
rect 600 91 606 125
rect 640 91 646 125
rect 600 53 646 91
rect 600 19 606 53
rect 640 19 646 53
rect 600 -19 646 19
rect 600 -53 606 -19
rect 640 -53 646 -19
rect 600 -91 646 -53
rect 600 -125 606 -91
rect 640 -125 646 -91
rect 600 -140 646 -125
rect 778 125 824 140
rect 778 91 784 125
rect 818 91 824 125
rect 778 53 824 91
rect 778 19 784 53
rect 818 19 824 53
rect 778 -19 824 19
rect 778 -53 784 -19
rect 818 -53 824 -19
rect 778 -91 824 -53
rect 778 -125 784 -91
rect 818 -125 824 -91
rect 778 -140 824 -125
rect 956 125 1002 140
rect 956 91 962 125
rect 996 91 1002 125
rect 956 53 1002 91
rect 956 19 962 53
rect 996 19 1002 53
rect 956 -19 1002 19
rect 956 -53 962 -19
rect 996 -53 1002 -19
rect 956 -91 1002 -53
rect 956 -125 962 -91
rect 996 -125 1002 -91
rect 956 -140 1002 -125
rect -928 -178 -852 -172
rect -928 -212 -907 -178
rect -873 -212 -852 -178
rect -928 -228 -852 -212
rect -750 -178 -674 -172
rect -750 -212 -729 -178
rect -695 -212 -674 -178
rect -750 -228 -674 -212
rect -572 -178 -496 -172
rect -572 -212 -551 -178
rect -517 -212 -496 -178
rect -572 -228 -496 -212
rect -394 -178 -318 -172
rect -394 -212 -373 -178
rect -339 -212 -318 -178
rect -394 -228 -318 -212
rect -216 -178 -140 -172
rect -216 -212 -195 -178
rect -161 -212 -140 -178
rect -216 -228 -140 -212
rect -38 -178 38 -172
rect -38 -212 -17 -178
rect 17 -212 38 -178
rect -38 -228 38 -212
rect 140 -178 216 -172
rect 140 -212 161 -178
rect 195 -212 216 -178
rect 140 -228 216 -212
rect 318 -178 394 -172
rect 318 -212 339 -178
rect 373 -212 394 -178
rect 318 -228 394 -212
rect 496 -178 572 -172
rect 496 -212 517 -178
rect 551 -212 572 -178
rect 496 -228 572 -212
rect 674 -178 750 -172
rect 674 -212 695 -178
rect 729 -212 750 -178
rect 674 -228 750 -212
rect 852 -178 928 -172
rect 852 -212 873 -178
rect 907 -212 928 -178
rect 852 -228 928 -212
<< end >>
