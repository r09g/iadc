magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< pwell >>
rect -3615 -166 3615 166
<< nmos >>
rect -3531 -140 -3411 140
rect -3353 -140 -3233 140
rect -3175 -140 -3055 140
rect -2997 -140 -2877 140
rect -2819 -140 -2699 140
rect -2641 -140 -2521 140
rect -2463 -140 -2343 140
rect -2285 -140 -2165 140
rect -2107 -140 -1987 140
rect -1929 -140 -1809 140
rect -1751 -140 -1631 140
rect -1573 -140 -1453 140
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
rect 1453 -140 1573 140
rect 1631 -140 1751 140
rect 1809 -140 1929 140
rect 1987 -140 2107 140
rect 2165 -140 2285 140
rect 2343 -140 2463 140
rect 2521 -140 2641 140
rect 2699 -140 2819 140
rect 2877 -140 2997 140
rect 3055 -140 3175 140
rect 3233 -140 3353 140
rect 3411 -140 3531 140
<< ndiff >>
rect -3589 119 -3531 140
rect -3589 85 -3577 119
rect -3543 85 -3531 119
rect -3589 51 -3531 85
rect -3589 17 -3577 51
rect -3543 17 -3531 51
rect -3589 -17 -3531 17
rect -3589 -51 -3577 -17
rect -3543 -51 -3531 -17
rect -3589 -85 -3531 -51
rect -3589 -119 -3577 -85
rect -3543 -119 -3531 -85
rect -3589 -140 -3531 -119
rect -3411 119 -3353 140
rect -3411 85 -3399 119
rect -3365 85 -3353 119
rect -3411 51 -3353 85
rect -3411 17 -3399 51
rect -3365 17 -3353 51
rect -3411 -17 -3353 17
rect -3411 -51 -3399 -17
rect -3365 -51 -3353 -17
rect -3411 -85 -3353 -51
rect -3411 -119 -3399 -85
rect -3365 -119 -3353 -85
rect -3411 -140 -3353 -119
rect -3233 119 -3175 140
rect -3233 85 -3221 119
rect -3187 85 -3175 119
rect -3233 51 -3175 85
rect -3233 17 -3221 51
rect -3187 17 -3175 51
rect -3233 -17 -3175 17
rect -3233 -51 -3221 -17
rect -3187 -51 -3175 -17
rect -3233 -85 -3175 -51
rect -3233 -119 -3221 -85
rect -3187 -119 -3175 -85
rect -3233 -140 -3175 -119
rect -3055 119 -2997 140
rect -3055 85 -3043 119
rect -3009 85 -2997 119
rect -3055 51 -2997 85
rect -3055 17 -3043 51
rect -3009 17 -2997 51
rect -3055 -17 -2997 17
rect -3055 -51 -3043 -17
rect -3009 -51 -2997 -17
rect -3055 -85 -2997 -51
rect -3055 -119 -3043 -85
rect -3009 -119 -2997 -85
rect -3055 -140 -2997 -119
rect -2877 119 -2819 140
rect -2877 85 -2865 119
rect -2831 85 -2819 119
rect -2877 51 -2819 85
rect -2877 17 -2865 51
rect -2831 17 -2819 51
rect -2877 -17 -2819 17
rect -2877 -51 -2865 -17
rect -2831 -51 -2819 -17
rect -2877 -85 -2819 -51
rect -2877 -119 -2865 -85
rect -2831 -119 -2819 -85
rect -2877 -140 -2819 -119
rect -2699 119 -2641 140
rect -2699 85 -2687 119
rect -2653 85 -2641 119
rect -2699 51 -2641 85
rect -2699 17 -2687 51
rect -2653 17 -2641 51
rect -2699 -17 -2641 17
rect -2699 -51 -2687 -17
rect -2653 -51 -2641 -17
rect -2699 -85 -2641 -51
rect -2699 -119 -2687 -85
rect -2653 -119 -2641 -85
rect -2699 -140 -2641 -119
rect -2521 119 -2463 140
rect -2521 85 -2509 119
rect -2475 85 -2463 119
rect -2521 51 -2463 85
rect -2521 17 -2509 51
rect -2475 17 -2463 51
rect -2521 -17 -2463 17
rect -2521 -51 -2509 -17
rect -2475 -51 -2463 -17
rect -2521 -85 -2463 -51
rect -2521 -119 -2509 -85
rect -2475 -119 -2463 -85
rect -2521 -140 -2463 -119
rect -2343 119 -2285 140
rect -2343 85 -2331 119
rect -2297 85 -2285 119
rect -2343 51 -2285 85
rect -2343 17 -2331 51
rect -2297 17 -2285 51
rect -2343 -17 -2285 17
rect -2343 -51 -2331 -17
rect -2297 -51 -2285 -17
rect -2343 -85 -2285 -51
rect -2343 -119 -2331 -85
rect -2297 -119 -2285 -85
rect -2343 -140 -2285 -119
rect -2165 119 -2107 140
rect -2165 85 -2153 119
rect -2119 85 -2107 119
rect -2165 51 -2107 85
rect -2165 17 -2153 51
rect -2119 17 -2107 51
rect -2165 -17 -2107 17
rect -2165 -51 -2153 -17
rect -2119 -51 -2107 -17
rect -2165 -85 -2107 -51
rect -2165 -119 -2153 -85
rect -2119 -119 -2107 -85
rect -2165 -140 -2107 -119
rect -1987 119 -1929 140
rect -1987 85 -1975 119
rect -1941 85 -1929 119
rect -1987 51 -1929 85
rect -1987 17 -1975 51
rect -1941 17 -1929 51
rect -1987 -17 -1929 17
rect -1987 -51 -1975 -17
rect -1941 -51 -1929 -17
rect -1987 -85 -1929 -51
rect -1987 -119 -1975 -85
rect -1941 -119 -1929 -85
rect -1987 -140 -1929 -119
rect -1809 119 -1751 140
rect -1809 85 -1797 119
rect -1763 85 -1751 119
rect -1809 51 -1751 85
rect -1809 17 -1797 51
rect -1763 17 -1751 51
rect -1809 -17 -1751 17
rect -1809 -51 -1797 -17
rect -1763 -51 -1751 -17
rect -1809 -85 -1751 -51
rect -1809 -119 -1797 -85
rect -1763 -119 -1751 -85
rect -1809 -140 -1751 -119
rect -1631 119 -1573 140
rect -1631 85 -1619 119
rect -1585 85 -1573 119
rect -1631 51 -1573 85
rect -1631 17 -1619 51
rect -1585 17 -1573 51
rect -1631 -17 -1573 17
rect -1631 -51 -1619 -17
rect -1585 -51 -1573 -17
rect -1631 -85 -1573 -51
rect -1631 -119 -1619 -85
rect -1585 -119 -1573 -85
rect -1631 -140 -1573 -119
rect -1453 119 -1395 140
rect -1453 85 -1441 119
rect -1407 85 -1395 119
rect -1453 51 -1395 85
rect -1453 17 -1441 51
rect -1407 17 -1395 51
rect -1453 -17 -1395 17
rect -1453 -51 -1441 -17
rect -1407 -51 -1395 -17
rect -1453 -85 -1395 -51
rect -1453 -119 -1441 -85
rect -1407 -119 -1395 -85
rect -1453 -140 -1395 -119
rect -1275 119 -1217 140
rect -1275 85 -1263 119
rect -1229 85 -1217 119
rect -1275 51 -1217 85
rect -1275 17 -1263 51
rect -1229 17 -1217 51
rect -1275 -17 -1217 17
rect -1275 -51 -1263 -17
rect -1229 -51 -1217 -17
rect -1275 -85 -1217 -51
rect -1275 -119 -1263 -85
rect -1229 -119 -1217 -85
rect -1275 -140 -1217 -119
rect -1097 119 -1039 140
rect -1097 85 -1085 119
rect -1051 85 -1039 119
rect -1097 51 -1039 85
rect -1097 17 -1085 51
rect -1051 17 -1039 51
rect -1097 -17 -1039 17
rect -1097 -51 -1085 -17
rect -1051 -51 -1039 -17
rect -1097 -85 -1039 -51
rect -1097 -119 -1085 -85
rect -1051 -119 -1039 -85
rect -1097 -140 -1039 -119
rect -919 119 -861 140
rect -919 85 -907 119
rect -873 85 -861 119
rect -919 51 -861 85
rect -919 17 -907 51
rect -873 17 -861 51
rect -919 -17 -861 17
rect -919 -51 -907 -17
rect -873 -51 -861 -17
rect -919 -85 -861 -51
rect -919 -119 -907 -85
rect -873 -119 -861 -85
rect -919 -140 -861 -119
rect -741 119 -683 140
rect -741 85 -729 119
rect -695 85 -683 119
rect -741 51 -683 85
rect -741 17 -729 51
rect -695 17 -683 51
rect -741 -17 -683 17
rect -741 -51 -729 -17
rect -695 -51 -683 -17
rect -741 -85 -683 -51
rect -741 -119 -729 -85
rect -695 -119 -683 -85
rect -741 -140 -683 -119
rect -563 119 -505 140
rect -563 85 -551 119
rect -517 85 -505 119
rect -563 51 -505 85
rect -563 17 -551 51
rect -517 17 -505 51
rect -563 -17 -505 17
rect -563 -51 -551 -17
rect -517 -51 -505 -17
rect -563 -85 -505 -51
rect -563 -119 -551 -85
rect -517 -119 -505 -85
rect -563 -140 -505 -119
rect -385 119 -327 140
rect -385 85 -373 119
rect -339 85 -327 119
rect -385 51 -327 85
rect -385 17 -373 51
rect -339 17 -327 51
rect -385 -17 -327 17
rect -385 -51 -373 -17
rect -339 -51 -327 -17
rect -385 -85 -327 -51
rect -385 -119 -373 -85
rect -339 -119 -327 -85
rect -385 -140 -327 -119
rect -207 119 -149 140
rect -207 85 -195 119
rect -161 85 -149 119
rect -207 51 -149 85
rect -207 17 -195 51
rect -161 17 -149 51
rect -207 -17 -149 17
rect -207 -51 -195 -17
rect -161 -51 -149 -17
rect -207 -85 -149 -51
rect -207 -119 -195 -85
rect -161 -119 -149 -85
rect -207 -140 -149 -119
rect -29 119 29 140
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -140 29 -119
rect 149 119 207 140
rect 149 85 161 119
rect 195 85 207 119
rect 149 51 207 85
rect 149 17 161 51
rect 195 17 207 51
rect 149 -17 207 17
rect 149 -51 161 -17
rect 195 -51 207 -17
rect 149 -85 207 -51
rect 149 -119 161 -85
rect 195 -119 207 -85
rect 149 -140 207 -119
rect 327 119 385 140
rect 327 85 339 119
rect 373 85 385 119
rect 327 51 385 85
rect 327 17 339 51
rect 373 17 385 51
rect 327 -17 385 17
rect 327 -51 339 -17
rect 373 -51 385 -17
rect 327 -85 385 -51
rect 327 -119 339 -85
rect 373 -119 385 -85
rect 327 -140 385 -119
rect 505 119 563 140
rect 505 85 517 119
rect 551 85 563 119
rect 505 51 563 85
rect 505 17 517 51
rect 551 17 563 51
rect 505 -17 563 17
rect 505 -51 517 -17
rect 551 -51 563 -17
rect 505 -85 563 -51
rect 505 -119 517 -85
rect 551 -119 563 -85
rect 505 -140 563 -119
rect 683 119 741 140
rect 683 85 695 119
rect 729 85 741 119
rect 683 51 741 85
rect 683 17 695 51
rect 729 17 741 51
rect 683 -17 741 17
rect 683 -51 695 -17
rect 729 -51 741 -17
rect 683 -85 741 -51
rect 683 -119 695 -85
rect 729 -119 741 -85
rect 683 -140 741 -119
rect 861 119 919 140
rect 861 85 873 119
rect 907 85 919 119
rect 861 51 919 85
rect 861 17 873 51
rect 907 17 919 51
rect 861 -17 919 17
rect 861 -51 873 -17
rect 907 -51 919 -17
rect 861 -85 919 -51
rect 861 -119 873 -85
rect 907 -119 919 -85
rect 861 -140 919 -119
rect 1039 119 1097 140
rect 1039 85 1051 119
rect 1085 85 1097 119
rect 1039 51 1097 85
rect 1039 17 1051 51
rect 1085 17 1097 51
rect 1039 -17 1097 17
rect 1039 -51 1051 -17
rect 1085 -51 1097 -17
rect 1039 -85 1097 -51
rect 1039 -119 1051 -85
rect 1085 -119 1097 -85
rect 1039 -140 1097 -119
rect 1217 119 1275 140
rect 1217 85 1229 119
rect 1263 85 1275 119
rect 1217 51 1275 85
rect 1217 17 1229 51
rect 1263 17 1275 51
rect 1217 -17 1275 17
rect 1217 -51 1229 -17
rect 1263 -51 1275 -17
rect 1217 -85 1275 -51
rect 1217 -119 1229 -85
rect 1263 -119 1275 -85
rect 1217 -140 1275 -119
rect 1395 119 1453 140
rect 1395 85 1407 119
rect 1441 85 1453 119
rect 1395 51 1453 85
rect 1395 17 1407 51
rect 1441 17 1453 51
rect 1395 -17 1453 17
rect 1395 -51 1407 -17
rect 1441 -51 1453 -17
rect 1395 -85 1453 -51
rect 1395 -119 1407 -85
rect 1441 -119 1453 -85
rect 1395 -140 1453 -119
rect 1573 119 1631 140
rect 1573 85 1585 119
rect 1619 85 1631 119
rect 1573 51 1631 85
rect 1573 17 1585 51
rect 1619 17 1631 51
rect 1573 -17 1631 17
rect 1573 -51 1585 -17
rect 1619 -51 1631 -17
rect 1573 -85 1631 -51
rect 1573 -119 1585 -85
rect 1619 -119 1631 -85
rect 1573 -140 1631 -119
rect 1751 119 1809 140
rect 1751 85 1763 119
rect 1797 85 1809 119
rect 1751 51 1809 85
rect 1751 17 1763 51
rect 1797 17 1809 51
rect 1751 -17 1809 17
rect 1751 -51 1763 -17
rect 1797 -51 1809 -17
rect 1751 -85 1809 -51
rect 1751 -119 1763 -85
rect 1797 -119 1809 -85
rect 1751 -140 1809 -119
rect 1929 119 1987 140
rect 1929 85 1941 119
rect 1975 85 1987 119
rect 1929 51 1987 85
rect 1929 17 1941 51
rect 1975 17 1987 51
rect 1929 -17 1987 17
rect 1929 -51 1941 -17
rect 1975 -51 1987 -17
rect 1929 -85 1987 -51
rect 1929 -119 1941 -85
rect 1975 -119 1987 -85
rect 1929 -140 1987 -119
rect 2107 119 2165 140
rect 2107 85 2119 119
rect 2153 85 2165 119
rect 2107 51 2165 85
rect 2107 17 2119 51
rect 2153 17 2165 51
rect 2107 -17 2165 17
rect 2107 -51 2119 -17
rect 2153 -51 2165 -17
rect 2107 -85 2165 -51
rect 2107 -119 2119 -85
rect 2153 -119 2165 -85
rect 2107 -140 2165 -119
rect 2285 119 2343 140
rect 2285 85 2297 119
rect 2331 85 2343 119
rect 2285 51 2343 85
rect 2285 17 2297 51
rect 2331 17 2343 51
rect 2285 -17 2343 17
rect 2285 -51 2297 -17
rect 2331 -51 2343 -17
rect 2285 -85 2343 -51
rect 2285 -119 2297 -85
rect 2331 -119 2343 -85
rect 2285 -140 2343 -119
rect 2463 119 2521 140
rect 2463 85 2475 119
rect 2509 85 2521 119
rect 2463 51 2521 85
rect 2463 17 2475 51
rect 2509 17 2521 51
rect 2463 -17 2521 17
rect 2463 -51 2475 -17
rect 2509 -51 2521 -17
rect 2463 -85 2521 -51
rect 2463 -119 2475 -85
rect 2509 -119 2521 -85
rect 2463 -140 2521 -119
rect 2641 119 2699 140
rect 2641 85 2653 119
rect 2687 85 2699 119
rect 2641 51 2699 85
rect 2641 17 2653 51
rect 2687 17 2699 51
rect 2641 -17 2699 17
rect 2641 -51 2653 -17
rect 2687 -51 2699 -17
rect 2641 -85 2699 -51
rect 2641 -119 2653 -85
rect 2687 -119 2699 -85
rect 2641 -140 2699 -119
rect 2819 119 2877 140
rect 2819 85 2831 119
rect 2865 85 2877 119
rect 2819 51 2877 85
rect 2819 17 2831 51
rect 2865 17 2877 51
rect 2819 -17 2877 17
rect 2819 -51 2831 -17
rect 2865 -51 2877 -17
rect 2819 -85 2877 -51
rect 2819 -119 2831 -85
rect 2865 -119 2877 -85
rect 2819 -140 2877 -119
rect 2997 119 3055 140
rect 2997 85 3009 119
rect 3043 85 3055 119
rect 2997 51 3055 85
rect 2997 17 3009 51
rect 3043 17 3055 51
rect 2997 -17 3055 17
rect 2997 -51 3009 -17
rect 3043 -51 3055 -17
rect 2997 -85 3055 -51
rect 2997 -119 3009 -85
rect 3043 -119 3055 -85
rect 2997 -140 3055 -119
rect 3175 119 3233 140
rect 3175 85 3187 119
rect 3221 85 3233 119
rect 3175 51 3233 85
rect 3175 17 3187 51
rect 3221 17 3233 51
rect 3175 -17 3233 17
rect 3175 -51 3187 -17
rect 3221 -51 3233 -17
rect 3175 -85 3233 -51
rect 3175 -119 3187 -85
rect 3221 -119 3233 -85
rect 3175 -140 3233 -119
rect 3353 119 3411 140
rect 3353 85 3365 119
rect 3399 85 3411 119
rect 3353 51 3411 85
rect 3353 17 3365 51
rect 3399 17 3411 51
rect 3353 -17 3411 17
rect 3353 -51 3365 -17
rect 3399 -51 3411 -17
rect 3353 -85 3411 -51
rect 3353 -119 3365 -85
rect 3399 -119 3411 -85
rect 3353 -140 3411 -119
rect 3531 119 3589 140
rect 3531 85 3543 119
rect 3577 85 3589 119
rect 3531 51 3589 85
rect 3531 17 3543 51
rect 3577 17 3589 51
rect 3531 -17 3589 17
rect 3531 -51 3543 -17
rect 3577 -51 3589 -17
rect 3531 -85 3589 -51
rect 3531 -119 3543 -85
rect 3577 -119 3589 -85
rect 3531 -140 3589 -119
<< ndiffc >>
rect -3577 85 -3543 119
rect -3577 17 -3543 51
rect -3577 -51 -3543 -17
rect -3577 -119 -3543 -85
rect -3399 85 -3365 119
rect -3399 17 -3365 51
rect -3399 -51 -3365 -17
rect -3399 -119 -3365 -85
rect -3221 85 -3187 119
rect -3221 17 -3187 51
rect -3221 -51 -3187 -17
rect -3221 -119 -3187 -85
rect -3043 85 -3009 119
rect -3043 17 -3009 51
rect -3043 -51 -3009 -17
rect -3043 -119 -3009 -85
rect -2865 85 -2831 119
rect -2865 17 -2831 51
rect -2865 -51 -2831 -17
rect -2865 -119 -2831 -85
rect -2687 85 -2653 119
rect -2687 17 -2653 51
rect -2687 -51 -2653 -17
rect -2687 -119 -2653 -85
rect -2509 85 -2475 119
rect -2509 17 -2475 51
rect -2509 -51 -2475 -17
rect -2509 -119 -2475 -85
rect -2331 85 -2297 119
rect -2331 17 -2297 51
rect -2331 -51 -2297 -17
rect -2331 -119 -2297 -85
rect -2153 85 -2119 119
rect -2153 17 -2119 51
rect -2153 -51 -2119 -17
rect -2153 -119 -2119 -85
rect -1975 85 -1941 119
rect -1975 17 -1941 51
rect -1975 -51 -1941 -17
rect -1975 -119 -1941 -85
rect -1797 85 -1763 119
rect -1797 17 -1763 51
rect -1797 -51 -1763 -17
rect -1797 -119 -1763 -85
rect -1619 85 -1585 119
rect -1619 17 -1585 51
rect -1619 -51 -1585 -17
rect -1619 -119 -1585 -85
rect -1441 85 -1407 119
rect -1441 17 -1407 51
rect -1441 -51 -1407 -17
rect -1441 -119 -1407 -85
rect -1263 85 -1229 119
rect -1263 17 -1229 51
rect -1263 -51 -1229 -17
rect -1263 -119 -1229 -85
rect -1085 85 -1051 119
rect -1085 17 -1051 51
rect -1085 -51 -1051 -17
rect -1085 -119 -1051 -85
rect -907 85 -873 119
rect -907 17 -873 51
rect -907 -51 -873 -17
rect -907 -119 -873 -85
rect -729 85 -695 119
rect -729 17 -695 51
rect -729 -51 -695 -17
rect -729 -119 -695 -85
rect -551 85 -517 119
rect -551 17 -517 51
rect -551 -51 -517 -17
rect -551 -119 -517 -85
rect -373 85 -339 119
rect -373 17 -339 51
rect -373 -51 -339 -17
rect -373 -119 -339 -85
rect -195 85 -161 119
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect 161 -119 195 -85
rect 339 85 373 119
rect 339 17 373 51
rect 339 -51 373 -17
rect 339 -119 373 -85
rect 517 85 551 119
rect 517 17 551 51
rect 517 -51 551 -17
rect 517 -119 551 -85
rect 695 85 729 119
rect 695 17 729 51
rect 695 -51 729 -17
rect 695 -119 729 -85
rect 873 85 907 119
rect 873 17 907 51
rect 873 -51 907 -17
rect 873 -119 907 -85
rect 1051 85 1085 119
rect 1051 17 1085 51
rect 1051 -51 1085 -17
rect 1051 -119 1085 -85
rect 1229 85 1263 119
rect 1229 17 1263 51
rect 1229 -51 1263 -17
rect 1229 -119 1263 -85
rect 1407 85 1441 119
rect 1407 17 1441 51
rect 1407 -51 1441 -17
rect 1407 -119 1441 -85
rect 1585 85 1619 119
rect 1585 17 1619 51
rect 1585 -51 1619 -17
rect 1585 -119 1619 -85
rect 1763 85 1797 119
rect 1763 17 1797 51
rect 1763 -51 1797 -17
rect 1763 -119 1797 -85
rect 1941 85 1975 119
rect 1941 17 1975 51
rect 1941 -51 1975 -17
rect 1941 -119 1975 -85
rect 2119 85 2153 119
rect 2119 17 2153 51
rect 2119 -51 2153 -17
rect 2119 -119 2153 -85
rect 2297 85 2331 119
rect 2297 17 2331 51
rect 2297 -51 2331 -17
rect 2297 -119 2331 -85
rect 2475 85 2509 119
rect 2475 17 2509 51
rect 2475 -51 2509 -17
rect 2475 -119 2509 -85
rect 2653 85 2687 119
rect 2653 17 2687 51
rect 2653 -51 2687 -17
rect 2653 -119 2687 -85
rect 2831 85 2865 119
rect 2831 17 2865 51
rect 2831 -51 2865 -17
rect 2831 -119 2865 -85
rect 3009 85 3043 119
rect 3009 17 3043 51
rect 3009 -51 3043 -17
rect 3009 -119 3043 -85
rect 3187 85 3221 119
rect 3187 17 3221 51
rect 3187 -51 3221 -17
rect 3187 -119 3221 -85
rect 3365 85 3399 119
rect 3365 17 3399 51
rect 3365 -51 3399 -17
rect 3365 -119 3399 -85
rect 3543 85 3577 119
rect 3543 17 3577 51
rect 3543 -51 3577 -17
rect 3543 -119 3577 -85
<< poly >>
rect -3509 212 -3433 228
rect -3509 194 -3488 212
rect -3531 178 -3488 194
rect -3454 194 -3433 212
rect -3331 212 -3255 228
rect -3331 194 -3310 212
rect -3454 178 -3411 194
rect -3531 140 -3411 178
rect -3353 178 -3310 194
rect -3276 194 -3255 212
rect -3153 212 -3077 228
rect -3153 194 -3132 212
rect -3276 178 -3233 194
rect -3353 140 -3233 178
rect -3175 178 -3132 194
rect -3098 194 -3077 212
rect -2975 212 -2899 228
rect -2975 194 -2954 212
rect -3098 178 -3055 194
rect -3175 140 -3055 178
rect -2997 178 -2954 194
rect -2920 194 -2899 212
rect -2797 212 -2721 228
rect -2797 194 -2776 212
rect -2920 178 -2877 194
rect -2997 140 -2877 178
rect -2819 178 -2776 194
rect -2742 194 -2721 212
rect -2619 212 -2543 228
rect -2619 194 -2598 212
rect -2742 178 -2699 194
rect -2819 140 -2699 178
rect -2641 178 -2598 194
rect -2564 194 -2543 212
rect -2441 212 -2365 228
rect -2441 194 -2420 212
rect -2564 178 -2521 194
rect -2641 140 -2521 178
rect -2463 178 -2420 194
rect -2386 194 -2365 212
rect -2263 212 -2187 228
rect -2263 194 -2242 212
rect -2386 178 -2343 194
rect -2463 140 -2343 178
rect -2285 178 -2242 194
rect -2208 194 -2187 212
rect -2085 212 -2009 228
rect -2085 194 -2064 212
rect -2208 178 -2165 194
rect -2285 140 -2165 178
rect -2107 178 -2064 194
rect -2030 194 -2009 212
rect -1907 212 -1831 228
rect -1907 194 -1886 212
rect -2030 178 -1987 194
rect -2107 140 -1987 178
rect -1929 178 -1886 194
rect -1852 194 -1831 212
rect -1729 212 -1653 228
rect -1729 194 -1708 212
rect -1852 178 -1809 194
rect -1929 140 -1809 178
rect -1751 178 -1708 194
rect -1674 194 -1653 212
rect -1551 212 -1475 228
rect -1551 194 -1530 212
rect -1674 178 -1631 194
rect -1751 140 -1631 178
rect -1573 178 -1530 194
rect -1496 194 -1475 212
rect -1373 212 -1297 228
rect -1373 194 -1352 212
rect -1496 178 -1453 194
rect -1573 140 -1453 178
rect -1395 178 -1352 194
rect -1318 194 -1297 212
rect -1195 212 -1119 228
rect -1195 194 -1174 212
rect -1318 178 -1275 194
rect -1395 140 -1275 178
rect -1217 178 -1174 194
rect -1140 194 -1119 212
rect -1017 212 -941 228
rect -1017 194 -996 212
rect -1140 178 -1097 194
rect -1217 140 -1097 178
rect -1039 178 -996 194
rect -962 194 -941 212
rect -839 212 -763 228
rect -839 194 -818 212
rect -962 178 -919 194
rect -1039 140 -919 178
rect -861 178 -818 194
rect -784 194 -763 212
rect -661 212 -585 228
rect -661 194 -640 212
rect -784 178 -741 194
rect -861 140 -741 178
rect -683 178 -640 194
rect -606 194 -585 212
rect -483 212 -407 228
rect -483 194 -462 212
rect -606 178 -563 194
rect -683 140 -563 178
rect -505 178 -462 194
rect -428 194 -407 212
rect -305 212 -229 228
rect -305 194 -284 212
rect -428 178 -385 194
rect -505 140 -385 178
rect -327 178 -284 194
rect -250 194 -229 212
rect -127 212 -51 228
rect -127 194 -106 212
rect -250 178 -207 194
rect -327 140 -207 178
rect -149 178 -106 194
rect -72 194 -51 212
rect 51 212 127 228
rect 51 194 72 212
rect -72 178 -29 194
rect -149 140 -29 178
rect 29 178 72 194
rect 106 194 127 212
rect 229 212 305 228
rect 229 194 250 212
rect 106 178 149 194
rect 29 140 149 178
rect 207 178 250 194
rect 284 194 305 212
rect 407 212 483 228
rect 407 194 428 212
rect 284 178 327 194
rect 207 140 327 178
rect 385 178 428 194
rect 462 194 483 212
rect 585 212 661 228
rect 585 194 606 212
rect 462 178 505 194
rect 385 140 505 178
rect 563 178 606 194
rect 640 194 661 212
rect 763 212 839 228
rect 763 194 784 212
rect 640 178 683 194
rect 563 140 683 178
rect 741 178 784 194
rect 818 194 839 212
rect 941 212 1017 228
rect 941 194 962 212
rect 818 178 861 194
rect 741 140 861 178
rect 919 178 962 194
rect 996 194 1017 212
rect 1119 212 1195 228
rect 1119 194 1140 212
rect 996 178 1039 194
rect 919 140 1039 178
rect 1097 178 1140 194
rect 1174 194 1195 212
rect 1297 212 1373 228
rect 1297 194 1318 212
rect 1174 178 1217 194
rect 1097 140 1217 178
rect 1275 178 1318 194
rect 1352 194 1373 212
rect 1475 212 1551 228
rect 1475 194 1496 212
rect 1352 178 1395 194
rect 1275 140 1395 178
rect 1453 178 1496 194
rect 1530 194 1551 212
rect 1653 212 1729 228
rect 1653 194 1674 212
rect 1530 178 1573 194
rect 1453 140 1573 178
rect 1631 178 1674 194
rect 1708 194 1729 212
rect 1831 212 1907 228
rect 1831 194 1852 212
rect 1708 178 1751 194
rect 1631 140 1751 178
rect 1809 178 1852 194
rect 1886 194 1907 212
rect 2009 212 2085 228
rect 2009 194 2030 212
rect 1886 178 1929 194
rect 1809 140 1929 178
rect 1987 178 2030 194
rect 2064 194 2085 212
rect 2187 212 2263 228
rect 2187 194 2208 212
rect 2064 178 2107 194
rect 1987 140 2107 178
rect 2165 178 2208 194
rect 2242 194 2263 212
rect 2365 212 2441 228
rect 2365 194 2386 212
rect 2242 178 2285 194
rect 2165 140 2285 178
rect 2343 178 2386 194
rect 2420 194 2441 212
rect 2543 212 2619 228
rect 2543 194 2564 212
rect 2420 178 2463 194
rect 2343 140 2463 178
rect 2521 178 2564 194
rect 2598 194 2619 212
rect 2721 212 2797 228
rect 2721 194 2742 212
rect 2598 178 2641 194
rect 2521 140 2641 178
rect 2699 178 2742 194
rect 2776 194 2797 212
rect 2899 212 2975 228
rect 2899 194 2920 212
rect 2776 178 2819 194
rect 2699 140 2819 178
rect 2877 178 2920 194
rect 2954 194 2975 212
rect 3077 212 3153 228
rect 3077 194 3098 212
rect 2954 178 2997 194
rect 2877 140 2997 178
rect 3055 178 3098 194
rect 3132 194 3153 212
rect 3255 212 3331 228
rect 3255 194 3276 212
rect 3132 178 3175 194
rect 3055 140 3175 178
rect 3233 178 3276 194
rect 3310 194 3331 212
rect 3433 212 3509 228
rect 3433 194 3454 212
rect 3310 178 3353 194
rect 3233 140 3353 178
rect 3411 178 3454 194
rect 3488 194 3509 212
rect 3488 178 3531 194
rect 3411 140 3531 178
rect -3531 -178 -3411 -140
rect -3531 -194 -3488 -178
rect -3509 -212 -3488 -194
rect -3454 -194 -3411 -178
rect -3353 -178 -3233 -140
rect -3353 -194 -3310 -178
rect -3454 -212 -3433 -194
rect -3509 -228 -3433 -212
rect -3331 -212 -3310 -194
rect -3276 -194 -3233 -178
rect -3175 -178 -3055 -140
rect -3175 -194 -3132 -178
rect -3276 -212 -3255 -194
rect -3331 -228 -3255 -212
rect -3153 -212 -3132 -194
rect -3098 -194 -3055 -178
rect -2997 -178 -2877 -140
rect -2997 -194 -2954 -178
rect -3098 -212 -3077 -194
rect -3153 -228 -3077 -212
rect -2975 -212 -2954 -194
rect -2920 -194 -2877 -178
rect -2819 -178 -2699 -140
rect -2819 -194 -2776 -178
rect -2920 -212 -2899 -194
rect -2975 -228 -2899 -212
rect -2797 -212 -2776 -194
rect -2742 -194 -2699 -178
rect -2641 -178 -2521 -140
rect -2641 -194 -2598 -178
rect -2742 -212 -2721 -194
rect -2797 -228 -2721 -212
rect -2619 -212 -2598 -194
rect -2564 -194 -2521 -178
rect -2463 -178 -2343 -140
rect -2463 -194 -2420 -178
rect -2564 -212 -2543 -194
rect -2619 -228 -2543 -212
rect -2441 -212 -2420 -194
rect -2386 -194 -2343 -178
rect -2285 -178 -2165 -140
rect -2285 -194 -2242 -178
rect -2386 -212 -2365 -194
rect -2441 -228 -2365 -212
rect -2263 -212 -2242 -194
rect -2208 -194 -2165 -178
rect -2107 -178 -1987 -140
rect -2107 -194 -2064 -178
rect -2208 -212 -2187 -194
rect -2263 -228 -2187 -212
rect -2085 -212 -2064 -194
rect -2030 -194 -1987 -178
rect -1929 -178 -1809 -140
rect -1929 -194 -1886 -178
rect -2030 -212 -2009 -194
rect -2085 -228 -2009 -212
rect -1907 -212 -1886 -194
rect -1852 -194 -1809 -178
rect -1751 -178 -1631 -140
rect -1751 -194 -1708 -178
rect -1852 -212 -1831 -194
rect -1907 -228 -1831 -212
rect -1729 -212 -1708 -194
rect -1674 -194 -1631 -178
rect -1573 -178 -1453 -140
rect -1573 -194 -1530 -178
rect -1674 -212 -1653 -194
rect -1729 -228 -1653 -212
rect -1551 -212 -1530 -194
rect -1496 -194 -1453 -178
rect -1395 -178 -1275 -140
rect -1395 -194 -1352 -178
rect -1496 -212 -1475 -194
rect -1551 -228 -1475 -212
rect -1373 -212 -1352 -194
rect -1318 -194 -1275 -178
rect -1217 -178 -1097 -140
rect -1217 -194 -1174 -178
rect -1318 -212 -1297 -194
rect -1373 -228 -1297 -212
rect -1195 -212 -1174 -194
rect -1140 -194 -1097 -178
rect -1039 -178 -919 -140
rect -1039 -194 -996 -178
rect -1140 -212 -1119 -194
rect -1195 -228 -1119 -212
rect -1017 -212 -996 -194
rect -962 -194 -919 -178
rect -861 -178 -741 -140
rect -861 -194 -818 -178
rect -962 -212 -941 -194
rect -1017 -228 -941 -212
rect -839 -212 -818 -194
rect -784 -194 -741 -178
rect -683 -178 -563 -140
rect -683 -194 -640 -178
rect -784 -212 -763 -194
rect -839 -228 -763 -212
rect -661 -212 -640 -194
rect -606 -194 -563 -178
rect -505 -178 -385 -140
rect -505 -194 -462 -178
rect -606 -212 -585 -194
rect -661 -228 -585 -212
rect -483 -212 -462 -194
rect -428 -194 -385 -178
rect -327 -178 -207 -140
rect -327 -194 -284 -178
rect -428 -212 -407 -194
rect -483 -228 -407 -212
rect -305 -212 -284 -194
rect -250 -194 -207 -178
rect -149 -178 -29 -140
rect -149 -194 -106 -178
rect -250 -212 -229 -194
rect -305 -228 -229 -212
rect -127 -212 -106 -194
rect -72 -194 -29 -178
rect 29 -178 149 -140
rect 29 -194 72 -178
rect -72 -212 -51 -194
rect -127 -228 -51 -212
rect 51 -212 72 -194
rect 106 -194 149 -178
rect 207 -178 327 -140
rect 207 -194 250 -178
rect 106 -212 127 -194
rect 51 -228 127 -212
rect 229 -212 250 -194
rect 284 -194 327 -178
rect 385 -178 505 -140
rect 385 -194 428 -178
rect 284 -212 305 -194
rect 229 -228 305 -212
rect 407 -212 428 -194
rect 462 -194 505 -178
rect 563 -178 683 -140
rect 563 -194 606 -178
rect 462 -212 483 -194
rect 407 -228 483 -212
rect 585 -212 606 -194
rect 640 -194 683 -178
rect 741 -178 861 -140
rect 741 -194 784 -178
rect 640 -212 661 -194
rect 585 -228 661 -212
rect 763 -212 784 -194
rect 818 -194 861 -178
rect 919 -178 1039 -140
rect 919 -194 962 -178
rect 818 -212 839 -194
rect 763 -228 839 -212
rect 941 -212 962 -194
rect 996 -194 1039 -178
rect 1097 -178 1217 -140
rect 1097 -194 1140 -178
rect 996 -212 1017 -194
rect 941 -228 1017 -212
rect 1119 -212 1140 -194
rect 1174 -194 1217 -178
rect 1275 -178 1395 -140
rect 1275 -194 1318 -178
rect 1174 -212 1195 -194
rect 1119 -228 1195 -212
rect 1297 -212 1318 -194
rect 1352 -194 1395 -178
rect 1453 -178 1573 -140
rect 1453 -194 1496 -178
rect 1352 -212 1373 -194
rect 1297 -228 1373 -212
rect 1475 -212 1496 -194
rect 1530 -194 1573 -178
rect 1631 -178 1751 -140
rect 1631 -194 1674 -178
rect 1530 -212 1551 -194
rect 1475 -228 1551 -212
rect 1653 -212 1674 -194
rect 1708 -194 1751 -178
rect 1809 -178 1929 -140
rect 1809 -194 1852 -178
rect 1708 -212 1729 -194
rect 1653 -228 1729 -212
rect 1831 -212 1852 -194
rect 1886 -194 1929 -178
rect 1987 -178 2107 -140
rect 1987 -194 2030 -178
rect 1886 -212 1907 -194
rect 1831 -228 1907 -212
rect 2009 -212 2030 -194
rect 2064 -194 2107 -178
rect 2165 -178 2285 -140
rect 2165 -194 2208 -178
rect 2064 -212 2085 -194
rect 2009 -228 2085 -212
rect 2187 -212 2208 -194
rect 2242 -194 2285 -178
rect 2343 -178 2463 -140
rect 2343 -194 2386 -178
rect 2242 -212 2263 -194
rect 2187 -228 2263 -212
rect 2365 -212 2386 -194
rect 2420 -194 2463 -178
rect 2521 -178 2641 -140
rect 2521 -194 2564 -178
rect 2420 -212 2441 -194
rect 2365 -228 2441 -212
rect 2543 -212 2564 -194
rect 2598 -194 2641 -178
rect 2699 -178 2819 -140
rect 2699 -194 2742 -178
rect 2598 -212 2619 -194
rect 2543 -228 2619 -212
rect 2721 -212 2742 -194
rect 2776 -194 2819 -178
rect 2877 -178 2997 -140
rect 2877 -194 2920 -178
rect 2776 -212 2797 -194
rect 2721 -228 2797 -212
rect 2899 -212 2920 -194
rect 2954 -194 2997 -178
rect 3055 -178 3175 -140
rect 3055 -194 3098 -178
rect 2954 -212 2975 -194
rect 2899 -228 2975 -212
rect 3077 -212 3098 -194
rect 3132 -194 3175 -178
rect 3233 -178 3353 -140
rect 3233 -194 3276 -178
rect 3132 -212 3153 -194
rect 3077 -228 3153 -212
rect 3255 -212 3276 -194
rect 3310 -194 3353 -178
rect 3411 -178 3531 -140
rect 3411 -194 3454 -178
rect 3310 -212 3331 -194
rect 3255 -228 3331 -212
rect 3433 -212 3454 -194
rect 3488 -194 3531 -178
rect 3488 -212 3509 -194
rect 3433 -228 3509 -212
<< polycont >>
rect -3488 178 -3454 212
rect -3310 178 -3276 212
rect -3132 178 -3098 212
rect -2954 178 -2920 212
rect -2776 178 -2742 212
rect -2598 178 -2564 212
rect -2420 178 -2386 212
rect -2242 178 -2208 212
rect -2064 178 -2030 212
rect -1886 178 -1852 212
rect -1708 178 -1674 212
rect -1530 178 -1496 212
rect -1352 178 -1318 212
rect -1174 178 -1140 212
rect -996 178 -962 212
rect -818 178 -784 212
rect -640 178 -606 212
rect -462 178 -428 212
rect -284 178 -250 212
rect -106 178 -72 212
rect 72 178 106 212
rect 250 178 284 212
rect 428 178 462 212
rect 606 178 640 212
rect 784 178 818 212
rect 962 178 996 212
rect 1140 178 1174 212
rect 1318 178 1352 212
rect 1496 178 1530 212
rect 1674 178 1708 212
rect 1852 178 1886 212
rect 2030 178 2064 212
rect 2208 178 2242 212
rect 2386 178 2420 212
rect 2564 178 2598 212
rect 2742 178 2776 212
rect 2920 178 2954 212
rect 3098 178 3132 212
rect 3276 178 3310 212
rect 3454 178 3488 212
rect -3488 -212 -3454 -178
rect -3310 -212 -3276 -178
rect -3132 -212 -3098 -178
rect -2954 -212 -2920 -178
rect -2776 -212 -2742 -178
rect -2598 -212 -2564 -178
rect -2420 -212 -2386 -178
rect -2242 -212 -2208 -178
rect -2064 -212 -2030 -178
rect -1886 -212 -1852 -178
rect -1708 -212 -1674 -178
rect -1530 -212 -1496 -178
rect -1352 -212 -1318 -178
rect -1174 -212 -1140 -178
rect -996 -212 -962 -178
rect -818 -212 -784 -178
rect -640 -212 -606 -178
rect -462 -212 -428 -178
rect -284 -212 -250 -178
rect -106 -212 -72 -178
rect 72 -212 106 -178
rect 250 -212 284 -178
rect 428 -212 462 -178
rect 606 -212 640 -178
rect 784 -212 818 -178
rect 962 -212 996 -178
rect 1140 -212 1174 -178
rect 1318 -212 1352 -178
rect 1496 -212 1530 -178
rect 1674 -212 1708 -178
rect 1852 -212 1886 -178
rect 2030 -212 2064 -178
rect 2208 -212 2242 -178
rect 2386 -212 2420 -178
rect 2564 -212 2598 -178
rect 2742 -212 2776 -178
rect 2920 -212 2954 -178
rect 3098 -212 3132 -178
rect 3276 -212 3310 -178
rect 3454 -212 3488 -178
<< locali >>
rect -3509 178 -3488 212
rect -3454 178 -3433 212
rect -3331 178 -3310 212
rect -3276 178 -3255 212
rect -3153 178 -3132 212
rect -3098 178 -3077 212
rect -2975 178 -2954 212
rect -2920 178 -2899 212
rect -2797 178 -2776 212
rect -2742 178 -2721 212
rect -2619 178 -2598 212
rect -2564 178 -2543 212
rect -2441 178 -2420 212
rect -2386 178 -2365 212
rect -2263 178 -2242 212
rect -2208 178 -2187 212
rect -2085 178 -2064 212
rect -2030 178 -2009 212
rect -1907 178 -1886 212
rect -1852 178 -1831 212
rect -1729 178 -1708 212
rect -1674 178 -1653 212
rect -1551 178 -1530 212
rect -1496 178 -1475 212
rect -1373 178 -1352 212
rect -1318 178 -1297 212
rect -1195 178 -1174 212
rect -1140 178 -1119 212
rect -1017 178 -996 212
rect -962 178 -941 212
rect -839 178 -818 212
rect -784 178 -763 212
rect -661 178 -640 212
rect -606 178 -585 212
rect -483 178 -462 212
rect -428 178 -407 212
rect -305 178 -284 212
rect -250 178 -229 212
rect -127 178 -106 212
rect -72 178 -51 212
rect 51 178 72 212
rect 106 178 127 212
rect 229 178 250 212
rect 284 178 305 212
rect 407 178 428 212
rect 462 178 483 212
rect 585 178 606 212
rect 640 178 661 212
rect 763 178 784 212
rect 818 178 839 212
rect 941 178 962 212
rect 996 178 1017 212
rect 1119 178 1140 212
rect 1174 178 1195 212
rect 1297 178 1318 212
rect 1352 178 1373 212
rect 1475 178 1496 212
rect 1530 178 1551 212
rect 1653 178 1674 212
rect 1708 178 1729 212
rect 1831 178 1852 212
rect 1886 178 1907 212
rect 2009 178 2030 212
rect 2064 178 2085 212
rect 2187 178 2208 212
rect 2242 178 2263 212
rect 2365 178 2386 212
rect 2420 178 2441 212
rect 2543 178 2564 212
rect 2598 178 2619 212
rect 2721 178 2742 212
rect 2776 178 2797 212
rect 2899 178 2920 212
rect 2954 178 2975 212
rect 3077 178 3098 212
rect 3132 178 3153 212
rect 3255 178 3276 212
rect 3310 178 3331 212
rect 3433 178 3454 212
rect 3488 178 3509 212
rect -3577 125 -3543 144
rect -3577 53 -3543 85
rect -3577 -17 -3543 17
rect -3577 -85 -3543 -53
rect -3577 -144 -3543 -125
rect -3399 125 -3365 144
rect -3399 53 -3365 85
rect -3399 -17 -3365 17
rect -3399 -85 -3365 -53
rect -3399 -144 -3365 -125
rect -3221 125 -3187 144
rect -3221 53 -3187 85
rect -3221 -17 -3187 17
rect -3221 -85 -3187 -53
rect -3221 -144 -3187 -125
rect -3043 125 -3009 144
rect -3043 53 -3009 85
rect -3043 -17 -3009 17
rect -3043 -85 -3009 -53
rect -3043 -144 -3009 -125
rect -2865 125 -2831 144
rect -2865 53 -2831 85
rect -2865 -17 -2831 17
rect -2865 -85 -2831 -53
rect -2865 -144 -2831 -125
rect -2687 125 -2653 144
rect -2687 53 -2653 85
rect -2687 -17 -2653 17
rect -2687 -85 -2653 -53
rect -2687 -144 -2653 -125
rect -2509 125 -2475 144
rect -2509 53 -2475 85
rect -2509 -17 -2475 17
rect -2509 -85 -2475 -53
rect -2509 -144 -2475 -125
rect -2331 125 -2297 144
rect -2331 53 -2297 85
rect -2331 -17 -2297 17
rect -2331 -85 -2297 -53
rect -2331 -144 -2297 -125
rect -2153 125 -2119 144
rect -2153 53 -2119 85
rect -2153 -17 -2119 17
rect -2153 -85 -2119 -53
rect -2153 -144 -2119 -125
rect -1975 125 -1941 144
rect -1975 53 -1941 85
rect -1975 -17 -1941 17
rect -1975 -85 -1941 -53
rect -1975 -144 -1941 -125
rect -1797 125 -1763 144
rect -1797 53 -1763 85
rect -1797 -17 -1763 17
rect -1797 -85 -1763 -53
rect -1797 -144 -1763 -125
rect -1619 125 -1585 144
rect -1619 53 -1585 85
rect -1619 -17 -1585 17
rect -1619 -85 -1585 -53
rect -1619 -144 -1585 -125
rect -1441 125 -1407 144
rect -1441 53 -1407 85
rect -1441 -17 -1407 17
rect -1441 -85 -1407 -53
rect -1441 -144 -1407 -125
rect -1263 125 -1229 144
rect -1263 53 -1229 85
rect -1263 -17 -1229 17
rect -1263 -85 -1229 -53
rect -1263 -144 -1229 -125
rect -1085 125 -1051 144
rect -1085 53 -1051 85
rect -1085 -17 -1051 17
rect -1085 -85 -1051 -53
rect -1085 -144 -1051 -125
rect -907 125 -873 144
rect -907 53 -873 85
rect -907 -17 -873 17
rect -907 -85 -873 -53
rect -907 -144 -873 -125
rect -729 125 -695 144
rect -729 53 -695 85
rect -729 -17 -695 17
rect -729 -85 -695 -53
rect -729 -144 -695 -125
rect -551 125 -517 144
rect -551 53 -517 85
rect -551 -17 -517 17
rect -551 -85 -517 -53
rect -551 -144 -517 -125
rect -373 125 -339 144
rect -373 53 -339 85
rect -373 -17 -339 17
rect -373 -85 -339 -53
rect -373 -144 -339 -125
rect -195 125 -161 144
rect -195 53 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -53
rect -195 -144 -161 -125
rect -17 125 17 144
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -144 17 -125
rect 161 125 195 144
rect 161 53 195 85
rect 161 -17 195 17
rect 161 -85 195 -53
rect 161 -144 195 -125
rect 339 125 373 144
rect 339 53 373 85
rect 339 -17 373 17
rect 339 -85 373 -53
rect 339 -144 373 -125
rect 517 125 551 144
rect 517 53 551 85
rect 517 -17 551 17
rect 517 -85 551 -53
rect 517 -144 551 -125
rect 695 125 729 144
rect 695 53 729 85
rect 695 -17 729 17
rect 695 -85 729 -53
rect 695 -144 729 -125
rect 873 125 907 144
rect 873 53 907 85
rect 873 -17 907 17
rect 873 -85 907 -53
rect 873 -144 907 -125
rect 1051 125 1085 144
rect 1051 53 1085 85
rect 1051 -17 1085 17
rect 1051 -85 1085 -53
rect 1051 -144 1085 -125
rect 1229 125 1263 144
rect 1229 53 1263 85
rect 1229 -17 1263 17
rect 1229 -85 1263 -53
rect 1229 -144 1263 -125
rect 1407 125 1441 144
rect 1407 53 1441 85
rect 1407 -17 1441 17
rect 1407 -85 1441 -53
rect 1407 -144 1441 -125
rect 1585 125 1619 144
rect 1585 53 1619 85
rect 1585 -17 1619 17
rect 1585 -85 1619 -53
rect 1585 -144 1619 -125
rect 1763 125 1797 144
rect 1763 53 1797 85
rect 1763 -17 1797 17
rect 1763 -85 1797 -53
rect 1763 -144 1797 -125
rect 1941 125 1975 144
rect 1941 53 1975 85
rect 1941 -17 1975 17
rect 1941 -85 1975 -53
rect 1941 -144 1975 -125
rect 2119 125 2153 144
rect 2119 53 2153 85
rect 2119 -17 2153 17
rect 2119 -85 2153 -53
rect 2119 -144 2153 -125
rect 2297 125 2331 144
rect 2297 53 2331 85
rect 2297 -17 2331 17
rect 2297 -85 2331 -53
rect 2297 -144 2331 -125
rect 2475 125 2509 144
rect 2475 53 2509 85
rect 2475 -17 2509 17
rect 2475 -85 2509 -53
rect 2475 -144 2509 -125
rect 2653 125 2687 144
rect 2653 53 2687 85
rect 2653 -17 2687 17
rect 2653 -85 2687 -53
rect 2653 -144 2687 -125
rect 2831 125 2865 144
rect 2831 53 2865 85
rect 2831 -17 2865 17
rect 2831 -85 2865 -53
rect 2831 -144 2865 -125
rect 3009 125 3043 144
rect 3009 53 3043 85
rect 3009 -17 3043 17
rect 3009 -85 3043 -53
rect 3009 -144 3043 -125
rect 3187 125 3221 144
rect 3187 53 3221 85
rect 3187 -17 3221 17
rect 3187 -85 3221 -53
rect 3187 -144 3221 -125
rect 3365 125 3399 144
rect 3365 53 3399 85
rect 3365 -17 3399 17
rect 3365 -85 3399 -53
rect 3365 -144 3399 -125
rect 3543 125 3577 144
rect 3543 53 3577 85
rect 3543 -17 3577 17
rect 3543 -85 3577 -53
rect 3543 -144 3577 -125
rect -3509 -212 -3488 -178
rect -3454 -212 -3433 -178
rect -3331 -212 -3310 -178
rect -3276 -212 -3255 -178
rect -3153 -212 -3132 -178
rect -3098 -212 -3077 -178
rect -2975 -212 -2954 -178
rect -2920 -212 -2899 -178
rect -2797 -212 -2776 -178
rect -2742 -212 -2721 -178
rect -2619 -212 -2598 -178
rect -2564 -212 -2543 -178
rect -2441 -212 -2420 -178
rect -2386 -212 -2365 -178
rect -2263 -212 -2242 -178
rect -2208 -212 -2187 -178
rect -2085 -212 -2064 -178
rect -2030 -212 -2009 -178
rect -1907 -212 -1886 -178
rect -1852 -212 -1831 -178
rect -1729 -212 -1708 -178
rect -1674 -212 -1653 -178
rect -1551 -212 -1530 -178
rect -1496 -212 -1475 -178
rect -1373 -212 -1352 -178
rect -1318 -212 -1297 -178
rect -1195 -212 -1174 -178
rect -1140 -212 -1119 -178
rect -1017 -212 -996 -178
rect -962 -212 -941 -178
rect -839 -212 -818 -178
rect -784 -212 -763 -178
rect -661 -212 -640 -178
rect -606 -212 -585 -178
rect -483 -212 -462 -178
rect -428 -212 -407 -178
rect -305 -212 -284 -178
rect -250 -212 -229 -178
rect -127 -212 -106 -178
rect -72 -212 -51 -178
rect 51 -212 72 -178
rect 106 -212 127 -178
rect 229 -212 250 -178
rect 284 -212 305 -178
rect 407 -212 428 -178
rect 462 -212 483 -178
rect 585 -212 606 -178
rect 640 -212 661 -178
rect 763 -212 784 -178
rect 818 -212 839 -178
rect 941 -212 962 -178
rect 996 -212 1017 -178
rect 1119 -212 1140 -178
rect 1174 -212 1195 -178
rect 1297 -212 1318 -178
rect 1352 -212 1373 -178
rect 1475 -212 1496 -178
rect 1530 -212 1551 -178
rect 1653 -212 1674 -178
rect 1708 -212 1729 -178
rect 1831 -212 1852 -178
rect 1886 -212 1907 -178
rect 2009 -212 2030 -178
rect 2064 -212 2085 -178
rect 2187 -212 2208 -178
rect 2242 -212 2263 -178
rect 2365 -212 2386 -178
rect 2420 -212 2441 -178
rect 2543 -212 2564 -178
rect 2598 -212 2619 -178
rect 2721 -212 2742 -178
rect 2776 -212 2797 -178
rect 2899 -212 2920 -178
rect 2954 -212 2975 -178
rect 3077 -212 3098 -178
rect 3132 -212 3153 -178
rect 3255 -212 3276 -178
rect 3310 -212 3331 -178
rect 3433 -212 3454 -178
rect 3488 -212 3509 -178
<< viali >>
rect -3488 178 -3454 212
rect -3310 178 -3276 212
rect -3132 178 -3098 212
rect -2954 178 -2920 212
rect -2776 178 -2742 212
rect -2598 178 -2564 212
rect -2420 178 -2386 212
rect -2242 178 -2208 212
rect -2064 178 -2030 212
rect -1886 178 -1852 212
rect -1708 178 -1674 212
rect -1530 178 -1496 212
rect -1352 178 -1318 212
rect -1174 178 -1140 212
rect -996 178 -962 212
rect -818 178 -784 212
rect -640 178 -606 212
rect -462 178 -428 212
rect -284 178 -250 212
rect -106 178 -72 212
rect 72 178 106 212
rect 250 178 284 212
rect 428 178 462 212
rect 606 178 640 212
rect 784 178 818 212
rect 962 178 996 212
rect 1140 178 1174 212
rect 1318 178 1352 212
rect 1496 178 1530 212
rect 1674 178 1708 212
rect 1852 178 1886 212
rect 2030 178 2064 212
rect 2208 178 2242 212
rect 2386 178 2420 212
rect 2564 178 2598 212
rect 2742 178 2776 212
rect 2920 178 2954 212
rect 3098 178 3132 212
rect 3276 178 3310 212
rect 3454 178 3488 212
rect -3577 119 -3543 125
rect -3577 91 -3543 119
rect -3577 51 -3543 53
rect -3577 19 -3543 51
rect -3577 -51 -3543 -19
rect -3577 -53 -3543 -51
rect -3577 -119 -3543 -91
rect -3577 -125 -3543 -119
rect -3399 119 -3365 125
rect -3399 91 -3365 119
rect -3399 51 -3365 53
rect -3399 19 -3365 51
rect -3399 -51 -3365 -19
rect -3399 -53 -3365 -51
rect -3399 -119 -3365 -91
rect -3399 -125 -3365 -119
rect -3221 119 -3187 125
rect -3221 91 -3187 119
rect -3221 51 -3187 53
rect -3221 19 -3187 51
rect -3221 -51 -3187 -19
rect -3221 -53 -3187 -51
rect -3221 -119 -3187 -91
rect -3221 -125 -3187 -119
rect -3043 119 -3009 125
rect -3043 91 -3009 119
rect -3043 51 -3009 53
rect -3043 19 -3009 51
rect -3043 -51 -3009 -19
rect -3043 -53 -3009 -51
rect -3043 -119 -3009 -91
rect -3043 -125 -3009 -119
rect -2865 119 -2831 125
rect -2865 91 -2831 119
rect -2865 51 -2831 53
rect -2865 19 -2831 51
rect -2865 -51 -2831 -19
rect -2865 -53 -2831 -51
rect -2865 -119 -2831 -91
rect -2865 -125 -2831 -119
rect -2687 119 -2653 125
rect -2687 91 -2653 119
rect -2687 51 -2653 53
rect -2687 19 -2653 51
rect -2687 -51 -2653 -19
rect -2687 -53 -2653 -51
rect -2687 -119 -2653 -91
rect -2687 -125 -2653 -119
rect -2509 119 -2475 125
rect -2509 91 -2475 119
rect -2509 51 -2475 53
rect -2509 19 -2475 51
rect -2509 -51 -2475 -19
rect -2509 -53 -2475 -51
rect -2509 -119 -2475 -91
rect -2509 -125 -2475 -119
rect -2331 119 -2297 125
rect -2331 91 -2297 119
rect -2331 51 -2297 53
rect -2331 19 -2297 51
rect -2331 -51 -2297 -19
rect -2331 -53 -2297 -51
rect -2331 -119 -2297 -91
rect -2331 -125 -2297 -119
rect -2153 119 -2119 125
rect -2153 91 -2119 119
rect -2153 51 -2119 53
rect -2153 19 -2119 51
rect -2153 -51 -2119 -19
rect -2153 -53 -2119 -51
rect -2153 -119 -2119 -91
rect -2153 -125 -2119 -119
rect -1975 119 -1941 125
rect -1975 91 -1941 119
rect -1975 51 -1941 53
rect -1975 19 -1941 51
rect -1975 -51 -1941 -19
rect -1975 -53 -1941 -51
rect -1975 -119 -1941 -91
rect -1975 -125 -1941 -119
rect -1797 119 -1763 125
rect -1797 91 -1763 119
rect -1797 51 -1763 53
rect -1797 19 -1763 51
rect -1797 -51 -1763 -19
rect -1797 -53 -1763 -51
rect -1797 -119 -1763 -91
rect -1797 -125 -1763 -119
rect -1619 119 -1585 125
rect -1619 91 -1585 119
rect -1619 51 -1585 53
rect -1619 19 -1585 51
rect -1619 -51 -1585 -19
rect -1619 -53 -1585 -51
rect -1619 -119 -1585 -91
rect -1619 -125 -1585 -119
rect -1441 119 -1407 125
rect -1441 91 -1407 119
rect -1441 51 -1407 53
rect -1441 19 -1407 51
rect -1441 -51 -1407 -19
rect -1441 -53 -1407 -51
rect -1441 -119 -1407 -91
rect -1441 -125 -1407 -119
rect -1263 119 -1229 125
rect -1263 91 -1229 119
rect -1263 51 -1229 53
rect -1263 19 -1229 51
rect -1263 -51 -1229 -19
rect -1263 -53 -1229 -51
rect -1263 -119 -1229 -91
rect -1263 -125 -1229 -119
rect -1085 119 -1051 125
rect -1085 91 -1051 119
rect -1085 51 -1051 53
rect -1085 19 -1051 51
rect -1085 -51 -1051 -19
rect -1085 -53 -1051 -51
rect -1085 -119 -1051 -91
rect -1085 -125 -1051 -119
rect -907 119 -873 125
rect -907 91 -873 119
rect -907 51 -873 53
rect -907 19 -873 51
rect -907 -51 -873 -19
rect -907 -53 -873 -51
rect -907 -119 -873 -91
rect -907 -125 -873 -119
rect -729 119 -695 125
rect -729 91 -695 119
rect -729 51 -695 53
rect -729 19 -695 51
rect -729 -51 -695 -19
rect -729 -53 -695 -51
rect -729 -119 -695 -91
rect -729 -125 -695 -119
rect -551 119 -517 125
rect -551 91 -517 119
rect -551 51 -517 53
rect -551 19 -517 51
rect -551 -51 -517 -19
rect -551 -53 -517 -51
rect -551 -119 -517 -91
rect -551 -125 -517 -119
rect -373 119 -339 125
rect -373 91 -339 119
rect -373 51 -339 53
rect -373 19 -339 51
rect -373 -51 -339 -19
rect -373 -53 -339 -51
rect -373 -119 -339 -91
rect -373 -125 -339 -119
rect -195 119 -161 125
rect -195 91 -161 119
rect -195 51 -161 53
rect -195 19 -161 51
rect -195 -51 -161 -19
rect -195 -53 -161 -51
rect -195 -119 -161 -91
rect -195 -125 -161 -119
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect 161 119 195 125
rect 161 91 195 119
rect 161 51 195 53
rect 161 19 195 51
rect 161 -51 195 -19
rect 161 -53 195 -51
rect 161 -119 195 -91
rect 161 -125 195 -119
rect 339 119 373 125
rect 339 91 373 119
rect 339 51 373 53
rect 339 19 373 51
rect 339 -51 373 -19
rect 339 -53 373 -51
rect 339 -119 373 -91
rect 339 -125 373 -119
rect 517 119 551 125
rect 517 91 551 119
rect 517 51 551 53
rect 517 19 551 51
rect 517 -51 551 -19
rect 517 -53 551 -51
rect 517 -119 551 -91
rect 517 -125 551 -119
rect 695 119 729 125
rect 695 91 729 119
rect 695 51 729 53
rect 695 19 729 51
rect 695 -51 729 -19
rect 695 -53 729 -51
rect 695 -119 729 -91
rect 695 -125 729 -119
rect 873 119 907 125
rect 873 91 907 119
rect 873 51 907 53
rect 873 19 907 51
rect 873 -51 907 -19
rect 873 -53 907 -51
rect 873 -119 907 -91
rect 873 -125 907 -119
rect 1051 119 1085 125
rect 1051 91 1085 119
rect 1051 51 1085 53
rect 1051 19 1085 51
rect 1051 -51 1085 -19
rect 1051 -53 1085 -51
rect 1051 -119 1085 -91
rect 1051 -125 1085 -119
rect 1229 119 1263 125
rect 1229 91 1263 119
rect 1229 51 1263 53
rect 1229 19 1263 51
rect 1229 -51 1263 -19
rect 1229 -53 1263 -51
rect 1229 -119 1263 -91
rect 1229 -125 1263 -119
rect 1407 119 1441 125
rect 1407 91 1441 119
rect 1407 51 1441 53
rect 1407 19 1441 51
rect 1407 -51 1441 -19
rect 1407 -53 1441 -51
rect 1407 -119 1441 -91
rect 1407 -125 1441 -119
rect 1585 119 1619 125
rect 1585 91 1619 119
rect 1585 51 1619 53
rect 1585 19 1619 51
rect 1585 -51 1619 -19
rect 1585 -53 1619 -51
rect 1585 -119 1619 -91
rect 1585 -125 1619 -119
rect 1763 119 1797 125
rect 1763 91 1797 119
rect 1763 51 1797 53
rect 1763 19 1797 51
rect 1763 -51 1797 -19
rect 1763 -53 1797 -51
rect 1763 -119 1797 -91
rect 1763 -125 1797 -119
rect 1941 119 1975 125
rect 1941 91 1975 119
rect 1941 51 1975 53
rect 1941 19 1975 51
rect 1941 -51 1975 -19
rect 1941 -53 1975 -51
rect 1941 -119 1975 -91
rect 1941 -125 1975 -119
rect 2119 119 2153 125
rect 2119 91 2153 119
rect 2119 51 2153 53
rect 2119 19 2153 51
rect 2119 -51 2153 -19
rect 2119 -53 2153 -51
rect 2119 -119 2153 -91
rect 2119 -125 2153 -119
rect 2297 119 2331 125
rect 2297 91 2331 119
rect 2297 51 2331 53
rect 2297 19 2331 51
rect 2297 -51 2331 -19
rect 2297 -53 2331 -51
rect 2297 -119 2331 -91
rect 2297 -125 2331 -119
rect 2475 119 2509 125
rect 2475 91 2509 119
rect 2475 51 2509 53
rect 2475 19 2509 51
rect 2475 -51 2509 -19
rect 2475 -53 2509 -51
rect 2475 -119 2509 -91
rect 2475 -125 2509 -119
rect 2653 119 2687 125
rect 2653 91 2687 119
rect 2653 51 2687 53
rect 2653 19 2687 51
rect 2653 -51 2687 -19
rect 2653 -53 2687 -51
rect 2653 -119 2687 -91
rect 2653 -125 2687 -119
rect 2831 119 2865 125
rect 2831 91 2865 119
rect 2831 51 2865 53
rect 2831 19 2865 51
rect 2831 -51 2865 -19
rect 2831 -53 2865 -51
rect 2831 -119 2865 -91
rect 2831 -125 2865 -119
rect 3009 119 3043 125
rect 3009 91 3043 119
rect 3009 51 3043 53
rect 3009 19 3043 51
rect 3009 -51 3043 -19
rect 3009 -53 3043 -51
rect 3009 -119 3043 -91
rect 3009 -125 3043 -119
rect 3187 119 3221 125
rect 3187 91 3221 119
rect 3187 51 3221 53
rect 3187 19 3221 51
rect 3187 -51 3221 -19
rect 3187 -53 3221 -51
rect 3187 -119 3221 -91
rect 3187 -125 3221 -119
rect 3365 119 3399 125
rect 3365 91 3399 119
rect 3365 51 3399 53
rect 3365 19 3399 51
rect 3365 -51 3399 -19
rect 3365 -53 3399 -51
rect 3365 -119 3399 -91
rect 3365 -125 3399 -119
rect 3543 119 3577 125
rect 3543 91 3577 119
rect 3543 51 3577 53
rect 3543 19 3577 51
rect 3543 -51 3577 -19
rect 3543 -53 3577 -51
rect 3543 -119 3577 -91
rect 3543 -125 3577 -119
rect -3488 -212 -3454 -178
rect -3310 -212 -3276 -178
rect -3132 -212 -3098 -178
rect -2954 -212 -2920 -178
rect -2776 -212 -2742 -178
rect -2598 -212 -2564 -178
rect -2420 -212 -2386 -178
rect -2242 -212 -2208 -178
rect -2064 -212 -2030 -178
rect -1886 -212 -1852 -178
rect -1708 -212 -1674 -178
rect -1530 -212 -1496 -178
rect -1352 -212 -1318 -178
rect -1174 -212 -1140 -178
rect -996 -212 -962 -178
rect -818 -212 -784 -178
rect -640 -212 -606 -178
rect -462 -212 -428 -178
rect -284 -212 -250 -178
rect -106 -212 -72 -178
rect 72 -212 106 -178
rect 250 -212 284 -178
rect 428 -212 462 -178
rect 606 -212 640 -178
rect 784 -212 818 -178
rect 962 -212 996 -178
rect 1140 -212 1174 -178
rect 1318 -212 1352 -178
rect 1496 -212 1530 -178
rect 1674 -212 1708 -178
rect 1852 -212 1886 -178
rect 2030 -212 2064 -178
rect 2208 -212 2242 -178
rect 2386 -212 2420 -178
rect 2564 -212 2598 -178
rect 2742 -212 2776 -178
rect 2920 -212 2954 -178
rect 3098 -212 3132 -178
rect 3276 -212 3310 -178
rect 3454 -212 3488 -178
<< metal1 >>
rect -3509 212 -3433 228
rect -3509 178 -3488 212
rect -3454 178 -3433 212
rect -3509 172 -3433 178
rect -3331 212 -3255 228
rect -3331 178 -3310 212
rect -3276 178 -3255 212
rect -3331 172 -3255 178
rect -3153 212 -3077 228
rect -3153 178 -3132 212
rect -3098 178 -3077 212
rect -3153 172 -3077 178
rect -2975 212 -2899 228
rect -2975 178 -2954 212
rect -2920 178 -2899 212
rect -2975 172 -2899 178
rect -2797 212 -2721 228
rect -2797 178 -2776 212
rect -2742 178 -2721 212
rect -2797 172 -2721 178
rect -2619 212 -2543 228
rect -2619 178 -2598 212
rect -2564 178 -2543 212
rect -2619 172 -2543 178
rect -2441 212 -2365 228
rect -2441 178 -2420 212
rect -2386 178 -2365 212
rect -2441 172 -2365 178
rect -2263 212 -2187 228
rect -2263 178 -2242 212
rect -2208 178 -2187 212
rect -2263 172 -2187 178
rect -2085 212 -2009 228
rect -2085 178 -2064 212
rect -2030 178 -2009 212
rect -2085 172 -2009 178
rect -1907 212 -1831 228
rect -1907 178 -1886 212
rect -1852 178 -1831 212
rect -1907 172 -1831 178
rect -1729 212 -1653 228
rect -1729 178 -1708 212
rect -1674 178 -1653 212
rect -1729 172 -1653 178
rect -1551 212 -1475 228
rect -1551 178 -1530 212
rect -1496 178 -1475 212
rect -1551 172 -1475 178
rect -1373 212 -1297 228
rect -1373 178 -1352 212
rect -1318 178 -1297 212
rect -1373 172 -1297 178
rect -1195 212 -1119 228
rect -1195 178 -1174 212
rect -1140 178 -1119 212
rect -1195 172 -1119 178
rect -1017 212 -941 228
rect -1017 178 -996 212
rect -962 178 -941 212
rect -1017 172 -941 178
rect -839 212 -763 228
rect -839 178 -818 212
rect -784 178 -763 212
rect -839 172 -763 178
rect -661 212 -585 228
rect -661 178 -640 212
rect -606 178 -585 212
rect -661 172 -585 178
rect -483 212 -407 228
rect -483 178 -462 212
rect -428 178 -407 212
rect -483 172 -407 178
rect -305 212 -229 228
rect -305 178 -284 212
rect -250 178 -229 212
rect -305 172 -229 178
rect -127 212 -51 228
rect -127 178 -106 212
rect -72 178 -51 212
rect -127 172 -51 178
rect 51 212 127 228
rect 51 178 72 212
rect 106 178 127 212
rect 51 172 127 178
rect 229 212 305 228
rect 229 178 250 212
rect 284 178 305 212
rect 229 172 305 178
rect 407 212 483 228
rect 407 178 428 212
rect 462 178 483 212
rect 407 172 483 178
rect 585 212 661 228
rect 585 178 606 212
rect 640 178 661 212
rect 585 172 661 178
rect 763 212 839 228
rect 763 178 784 212
rect 818 178 839 212
rect 763 172 839 178
rect 941 212 1017 228
rect 941 178 962 212
rect 996 178 1017 212
rect 941 172 1017 178
rect 1119 212 1195 228
rect 1119 178 1140 212
rect 1174 178 1195 212
rect 1119 172 1195 178
rect 1297 212 1373 228
rect 1297 178 1318 212
rect 1352 178 1373 212
rect 1297 172 1373 178
rect 1475 212 1551 228
rect 1475 178 1496 212
rect 1530 178 1551 212
rect 1475 172 1551 178
rect 1653 212 1729 228
rect 1653 178 1674 212
rect 1708 178 1729 212
rect 1653 172 1729 178
rect 1831 212 1907 228
rect 1831 178 1852 212
rect 1886 178 1907 212
rect 1831 172 1907 178
rect 2009 212 2085 228
rect 2009 178 2030 212
rect 2064 178 2085 212
rect 2009 172 2085 178
rect 2187 212 2263 228
rect 2187 178 2208 212
rect 2242 178 2263 212
rect 2187 172 2263 178
rect 2365 212 2441 228
rect 2365 178 2386 212
rect 2420 178 2441 212
rect 2365 172 2441 178
rect 2543 212 2619 228
rect 2543 178 2564 212
rect 2598 178 2619 212
rect 2543 172 2619 178
rect 2721 212 2797 228
rect 2721 178 2742 212
rect 2776 178 2797 212
rect 2721 172 2797 178
rect 2899 212 2975 228
rect 2899 178 2920 212
rect 2954 178 2975 212
rect 2899 172 2975 178
rect 3077 212 3153 228
rect 3077 178 3098 212
rect 3132 178 3153 212
rect 3077 172 3153 178
rect 3255 212 3331 228
rect 3255 178 3276 212
rect 3310 178 3331 212
rect 3255 172 3331 178
rect 3433 212 3509 228
rect 3433 178 3454 212
rect 3488 178 3509 212
rect 3433 172 3509 178
rect -3583 125 -3537 140
rect -3583 91 -3577 125
rect -3543 91 -3537 125
rect -3583 53 -3537 91
rect -3583 19 -3577 53
rect -3543 19 -3537 53
rect -3583 -19 -3537 19
rect -3583 -53 -3577 -19
rect -3543 -53 -3537 -19
rect -3583 -91 -3537 -53
rect -3583 -125 -3577 -91
rect -3543 -125 -3537 -91
rect -3583 -140 -3537 -125
rect -3405 125 -3359 140
rect -3405 91 -3399 125
rect -3365 91 -3359 125
rect -3405 53 -3359 91
rect -3405 19 -3399 53
rect -3365 19 -3359 53
rect -3405 -19 -3359 19
rect -3405 -53 -3399 -19
rect -3365 -53 -3359 -19
rect -3405 -91 -3359 -53
rect -3405 -125 -3399 -91
rect -3365 -125 -3359 -91
rect -3405 -140 -3359 -125
rect -3227 125 -3181 140
rect -3227 91 -3221 125
rect -3187 91 -3181 125
rect -3227 53 -3181 91
rect -3227 19 -3221 53
rect -3187 19 -3181 53
rect -3227 -19 -3181 19
rect -3227 -53 -3221 -19
rect -3187 -53 -3181 -19
rect -3227 -91 -3181 -53
rect -3227 -125 -3221 -91
rect -3187 -125 -3181 -91
rect -3227 -140 -3181 -125
rect -3049 125 -3003 140
rect -3049 91 -3043 125
rect -3009 91 -3003 125
rect -3049 53 -3003 91
rect -3049 19 -3043 53
rect -3009 19 -3003 53
rect -3049 -19 -3003 19
rect -3049 -53 -3043 -19
rect -3009 -53 -3003 -19
rect -3049 -91 -3003 -53
rect -3049 -125 -3043 -91
rect -3009 -125 -3003 -91
rect -3049 -140 -3003 -125
rect -2871 125 -2825 140
rect -2871 91 -2865 125
rect -2831 91 -2825 125
rect -2871 53 -2825 91
rect -2871 19 -2865 53
rect -2831 19 -2825 53
rect -2871 -19 -2825 19
rect -2871 -53 -2865 -19
rect -2831 -53 -2825 -19
rect -2871 -91 -2825 -53
rect -2871 -125 -2865 -91
rect -2831 -125 -2825 -91
rect -2871 -140 -2825 -125
rect -2693 125 -2647 140
rect -2693 91 -2687 125
rect -2653 91 -2647 125
rect -2693 53 -2647 91
rect -2693 19 -2687 53
rect -2653 19 -2647 53
rect -2693 -19 -2647 19
rect -2693 -53 -2687 -19
rect -2653 -53 -2647 -19
rect -2693 -91 -2647 -53
rect -2693 -125 -2687 -91
rect -2653 -125 -2647 -91
rect -2693 -140 -2647 -125
rect -2515 125 -2469 140
rect -2515 91 -2509 125
rect -2475 91 -2469 125
rect -2515 53 -2469 91
rect -2515 19 -2509 53
rect -2475 19 -2469 53
rect -2515 -19 -2469 19
rect -2515 -53 -2509 -19
rect -2475 -53 -2469 -19
rect -2515 -91 -2469 -53
rect -2515 -125 -2509 -91
rect -2475 -125 -2469 -91
rect -2515 -140 -2469 -125
rect -2337 125 -2291 140
rect -2337 91 -2331 125
rect -2297 91 -2291 125
rect -2337 53 -2291 91
rect -2337 19 -2331 53
rect -2297 19 -2291 53
rect -2337 -19 -2291 19
rect -2337 -53 -2331 -19
rect -2297 -53 -2291 -19
rect -2337 -91 -2291 -53
rect -2337 -125 -2331 -91
rect -2297 -125 -2291 -91
rect -2337 -140 -2291 -125
rect -2159 125 -2113 140
rect -2159 91 -2153 125
rect -2119 91 -2113 125
rect -2159 53 -2113 91
rect -2159 19 -2153 53
rect -2119 19 -2113 53
rect -2159 -19 -2113 19
rect -2159 -53 -2153 -19
rect -2119 -53 -2113 -19
rect -2159 -91 -2113 -53
rect -2159 -125 -2153 -91
rect -2119 -125 -2113 -91
rect -2159 -140 -2113 -125
rect -1981 125 -1935 140
rect -1981 91 -1975 125
rect -1941 91 -1935 125
rect -1981 53 -1935 91
rect -1981 19 -1975 53
rect -1941 19 -1935 53
rect -1981 -19 -1935 19
rect -1981 -53 -1975 -19
rect -1941 -53 -1935 -19
rect -1981 -91 -1935 -53
rect -1981 -125 -1975 -91
rect -1941 -125 -1935 -91
rect -1981 -140 -1935 -125
rect -1803 125 -1757 140
rect -1803 91 -1797 125
rect -1763 91 -1757 125
rect -1803 53 -1757 91
rect -1803 19 -1797 53
rect -1763 19 -1757 53
rect -1803 -19 -1757 19
rect -1803 -53 -1797 -19
rect -1763 -53 -1757 -19
rect -1803 -91 -1757 -53
rect -1803 -125 -1797 -91
rect -1763 -125 -1757 -91
rect -1803 -140 -1757 -125
rect -1625 125 -1579 140
rect -1625 91 -1619 125
rect -1585 91 -1579 125
rect -1625 53 -1579 91
rect -1625 19 -1619 53
rect -1585 19 -1579 53
rect -1625 -19 -1579 19
rect -1625 -53 -1619 -19
rect -1585 -53 -1579 -19
rect -1625 -91 -1579 -53
rect -1625 -125 -1619 -91
rect -1585 -125 -1579 -91
rect -1625 -140 -1579 -125
rect -1447 125 -1401 140
rect -1447 91 -1441 125
rect -1407 91 -1401 125
rect -1447 53 -1401 91
rect -1447 19 -1441 53
rect -1407 19 -1401 53
rect -1447 -19 -1401 19
rect -1447 -53 -1441 -19
rect -1407 -53 -1401 -19
rect -1447 -91 -1401 -53
rect -1447 -125 -1441 -91
rect -1407 -125 -1401 -91
rect -1447 -140 -1401 -125
rect -1269 125 -1223 140
rect -1269 91 -1263 125
rect -1229 91 -1223 125
rect -1269 53 -1223 91
rect -1269 19 -1263 53
rect -1229 19 -1223 53
rect -1269 -19 -1223 19
rect -1269 -53 -1263 -19
rect -1229 -53 -1223 -19
rect -1269 -91 -1223 -53
rect -1269 -125 -1263 -91
rect -1229 -125 -1223 -91
rect -1269 -140 -1223 -125
rect -1091 125 -1045 140
rect -1091 91 -1085 125
rect -1051 91 -1045 125
rect -1091 53 -1045 91
rect -1091 19 -1085 53
rect -1051 19 -1045 53
rect -1091 -19 -1045 19
rect -1091 -53 -1085 -19
rect -1051 -53 -1045 -19
rect -1091 -91 -1045 -53
rect -1091 -125 -1085 -91
rect -1051 -125 -1045 -91
rect -1091 -140 -1045 -125
rect -913 125 -867 140
rect -913 91 -907 125
rect -873 91 -867 125
rect -913 53 -867 91
rect -913 19 -907 53
rect -873 19 -867 53
rect -913 -19 -867 19
rect -913 -53 -907 -19
rect -873 -53 -867 -19
rect -913 -91 -867 -53
rect -913 -125 -907 -91
rect -873 -125 -867 -91
rect -913 -140 -867 -125
rect -735 125 -689 140
rect -735 91 -729 125
rect -695 91 -689 125
rect -735 53 -689 91
rect -735 19 -729 53
rect -695 19 -689 53
rect -735 -19 -689 19
rect -735 -53 -729 -19
rect -695 -53 -689 -19
rect -735 -91 -689 -53
rect -735 -125 -729 -91
rect -695 -125 -689 -91
rect -735 -140 -689 -125
rect -557 125 -511 140
rect -557 91 -551 125
rect -517 91 -511 125
rect -557 53 -511 91
rect -557 19 -551 53
rect -517 19 -511 53
rect -557 -19 -511 19
rect -557 -53 -551 -19
rect -517 -53 -511 -19
rect -557 -91 -511 -53
rect -557 -125 -551 -91
rect -517 -125 -511 -91
rect -557 -140 -511 -125
rect -379 125 -333 140
rect -379 91 -373 125
rect -339 91 -333 125
rect -379 53 -333 91
rect -379 19 -373 53
rect -339 19 -333 53
rect -379 -19 -333 19
rect -379 -53 -373 -19
rect -339 -53 -333 -19
rect -379 -91 -333 -53
rect -379 -125 -373 -91
rect -339 -125 -333 -91
rect -379 -140 -333 -125
rect -201 125 -155 140
rect -201 91 -195 125
rect -161 91 -155 125
rect -201 53 -155 91
rect -201 19 -195 53
rect -161 19 -155 53
rect -201 -19 -155 19
rect -201 -53 -195 -19
rect -161 -53 -155 -19
rect -201 -91 -155 -53
rect -201 -125 -195 -91
rect -161 -125 -155 -91
rect -201 -140 -155 -125
rect -23 125 23 140
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -140 23 -125
rect 155 125 201 140
rect 155 91 161 125
rect 195 91 201 125
rect 155 53 201 91
rect 155 19 161 53
rect 195 19 201 53
rect 155 -19 201 19
rect 155 -53 161 -19
rect 195 -53 201 -19
rect 155 -91 201 -53
rect 155 -125 161 -91
rect 195 -125 201 -91
rect 155 -140 201 -125
rect 333 125 379 140
rect 333 91 339 125
rect 373 91 379 125
rect 333 53 379 91
rect 333 19 339 53
rect 373 19 379 53
rect 333 -19 379 19
rect 333 -53 339 -19
rect 373 -53 379 -19
rect 333 -91 379 -53
rect 333 -125 339 -91
rect 373 -125 379 -91
rect 333 -140 379 -125
rect 511 125 557 140
rect 511 91 517 125
rect 551 91 557 125
rect 511 53 557 91
rect 511 19 517 53
rect 551 19 557 53
rect 511 -19 557 19
rect 511 -53 517 -19
rect 551 -53 557 -19
rect 511 -91 557 -53
rect 511 -125 517 -91
rect 551 -125 557 -91
rect 511 -140 557 -125
rect 689 125 735 140
rect 689 91 695 125
rect 729 91 735 125
rect 689 53 735 91
rect 689 19 695 53
rect 729 19 735 53
rect 689 -19 735 19
rect 689 -53 695 -19
rect 729 -53 735 -19
rect 689 -91 735 -53
rect 689 -125 695 -91
rect 729 -125 735 -91
rect 689 -140 735 -125
rect 867 125 913 140
rect 867 91 873 125
rect 907 91 913 125
rect 867 53 913 91
rect 867 19 873 53
rect 907 19 913 53
rect 867 -19 913 19
rect 867 -53 873 -19
rect 907 -53 913 -19
rect 867 -91 913 -53
rect 867 -125 873 -91
rect 907 -125 913 -91
rect 867 -140 913 -125
rect 1045 125 1091 140
rect 1045 91 1051 125
rect 1085 91 1091 125
rect 1045 53 1091 91
rect 1045 19 1051 53
rect 1085 19 1091 53
rect 1045 -19 1091 19
rect 1045 -53 1051 -19
rect 1085 -53 1091 -19
rect 1045 -91 1091 -53
rect 1045 -125 1051 -91
rect 1085 -125 1091 -91
rect 1045 -140 1091 -125
rect 1223 125 1269 140
rect 1223 91 1229 125
rect 1263 91 1269 125
rect 1223 53 1269 91
rect 1223 19 1229 53
rect 1263 19 1269 53
rect 1223 -19 1269 19
rect 1223 -53 1229 -19
rect 1263 -53 1269 -19
rect 1223 -91 1269 -53
rect 1223 -125 1229 -91
rect 1263 -125 1269 -91
rect 1223 -140 1269 -125
rect 1401 125 1447 140
rect 1401 91 1407 125
rect 1441 91 1447 125
rect 1401 53 1447 91
rect 1401 19 1407 53
rect 1441 19 1447 53
rect 1401 -19 1447 19
rect 1401 -53 1407 -19
rect 1441 -53 1447 -19
rect 1401 -91 1447 -53
rect 1401 -125 1407 -91
rect 1441 -125 1447 -91
rect 1401 -140 1447 -125
rect 1579 125 1625 140
rect 1579 91 1585 125
rect 1619 91 1625 125
rect 1579 53 1625 91
rect 1579 19 1585 53
rect 1619 19 1625 53
rect 1579 -19 1625 19
rect 1579 -53 1585 -19
rect 1619 -53 1625 -19
rect 1579 -91 1625 -53
rect 1579 -125 1585 -91
rect 1619 -125 1625 -91
rect 1579 -140 1625 -125
rect 1757 125 1803 140
rect 1757 91 1763 125
rect 1797 91 1803 125
rect 1757 53 1803 91
rect 1757 19 1763 53
rect 1797 19 1803 53
rect 1757 -19 1803 19
rect 1757 -53 1763 -19
rect 1797 -53 1803 -19
rect 1757 -91 1803 -53
rect 1757 -125 1763 -91
rect 1797 -125 1803 -91
rect 1757 -140 1803 -125
rect 1935 125 1981 140
rect 1935 91 1941 125
rect 1975 91 1981 125
rect 1935 53 1981 91
rect 1935 19 1941 53
rect 1975 19 1981 53
rect 1935 -19 1981 19
rect 1935 -53 1941 -19
rect 1975 -53 1981 -19
rect 1935 -91 1981 -53
rect 1935 -125 1941 -91
rect 1975 -125 1981 -91
rect 1935 -140 1981 -125
rect 2113 125 2159 140
rect 2113 91 2119 125
rect 2153 91 2159 125
rect 2113 53 2159 91
rect 2113 19 2119 53
rect 2153 19 2159 53
rect 2113 -19 2159 19
rect 2113 -53 2119 -19
rect 2153 -53 2159 -19
rect 2113 -91 2159 -53
rect 2113 -125 2119 -91
rect 2153 -125 2159 -91
rect 2113 -140 2159 -125
rect 2291 125 2337 140
rect 2291 91 2297 125
rect 2331 91 2337 125
rect 2291 53 2337 91
rect 2291 19 2297 53
rect 2331 19 2337 53
rect 2291 -19 2337 19
rect 2291 -53 2297 -19
rect 2331 -53 2337 -19
rect 2291 -91 2337 -53
rect 2291 -125 2297 -91
rect 2331 -125 2337 -91
rect 2291 -140 2337 -125
rect 2469 125 2515 140
rect 2469 91 2475 125
rect 2509 91 2515 125
rect 2469 53 2515 91
rect 2469 19 2475 53
rect 2509 19 2515 53
rect 2469 -19 2515 19
rect 2469 -53 2475 -19
rect 2509 -53 2515 -19
rect 2469 -91 2515 -53
rect 2469 -125 2475 -91
rect 2509 -125 2515 -91
rect 2469 -140 2515 -125
rect 2647 125 2693 140
rect 2647 91 2653 125
rect 2687 91 2693 125
rect 2647 53 2693 91
rect 2647 19 2653 53
rect 2687 19 2693 53
rect 2647 -19 2693 19
rect 2647 -53 2653 -19
rect 2687 -53 2693 -19
rect 2647 -91 2693 -53
rect 2647 -125 2653 -91
rect 2687 -125 2693 -91
rect 2647 -140 2693 -125
rect 2825 125 2871 140
rect 2825 91 2831 125
rect 2865 91 2871 125
rect 2825 53 2871 91
rect 2825 19 2831 53
rect 2865 19 2871 53
rect 2825 -19 2871 19
rect 2825 -53 2831 -19
rect 2865 -53 2871 -19
rect 2825 -91 2871 -53
rect 2825 -125 2831 -91
rect 2865 -125 2871 -91
rect 2825 -140 2871 -125
rect 3003 125 3049 140
rect 3003 91 3009 125
rect 3043 91 3049 125
rect 3003 53 3049 91
rect 3003 19 3009 53
rect 3043 19 3049 53
rect 3003 -19 3049 19
rect 3003 -53 3009 -19
rect 3043 -53 3049 -19
rect 3003 -91 3049 -53
rect 3003 -125 3009 -91
rect 3043 -125 3049 -91
rect 3003 -140 3049 -125
rect 3181 125 3227 140
rect 3181 91 3187 125
rect 3221 91 3227 125
rect 3181 53 3227 91
rect 3181 19 3187 53
rect 3221 19 3227 53
rect 3181 -19 3227 19
rect 3181 -53 3187 -19
rect 3221 -53 3227 -19
rect 3181 -91 3227 -53
rect 3181 -125 3187 -91
rect 3221 -125 3227 -91
rect 3181 -140 3227 -125
rect 3359 125 3405 140
rect 3359 91 3365 125
rect 3399 91 3405 125
rect 3359 53 3405 91
rect 3359 19 3365 53
rect 3399 19 3405 53
rect 3359 -19 3405 19
rect 3359 -53 3365 -19
rect 3399 -53 3405 -19
rect 3359 -91 3405 -53
rect 3359 -125 3365 -91
rect 3399 -125 3405 -91
rect 3359 -140 3405 -125
rect 3537 125 3583 140
rect 3537 91 3543 125
rect 3577 91 3583 125
rect 3537 53 3583 91
rect 3537 19 3543 53
rect 3577 19 3583 53
rect 3537 -19 3583 19
rect 3537 -53 3543 -19
rect 3577 -53 3583 -19
rect 3537 -91 3583 -53
rect 3537 -125 3543 -91
rect 3577 -125 3583 -91
rect 3537 -140 3583 -125
rect -3509 -178 -3433 -172
rect -3509 -212 -3488 -178
rect -3454 -212 -3433 -178
rect -3509 -228 -3433 -212
rect -3331 -178 -3255 -172
rect -3331 -212 -3310 -178
rect -3276 -212 -3255 -178
rect -3331 -228 -3255 -212
rect -3153 -178 -3077 -172
rect -3153 -212 -3132 -178
rect -3098 -212 -3077 -178
rect -3153 -228 -3077 -212
rect -2975 -178 -2899 -172
rect -2975 -212 -2954 -178
rect -2920 -212 -2899 -178
rect -2975 -228 -2899 -212
rect -2797 -178 -2721 -172
rect -2797 -212 -2776 -178
rect -2742 -212 -2721 -178
rect -2797 -228 -2721 -212
rect -2619 -178 -2543 -172
rect -2619 -212 -2598 -178
rect -2564 -212 -2543 -178
rect -2619 -228 -2543 -212
rect -2441 -178 -2365 -172
rect -2441 -212 -2420 -178
rect -2386 -212 -2365 -178
rect -2441 -228 -2365 -212
rect -2263 -178 -2187 -172
rect -2263 -212 -2242 -178
rect -2208 -212 -2187 -178
rect -2263 -228 -2187 -212
rect -2085 -178 -2009 -172
rect -2085 -212 -2064 -178
rect -2030 -212 -2009 -178
rect -2085 -228 -2009 -212
rect -1907 -178 -1831 -172
rect -1907 -212 -1886 -178
rect -1852 -212 -1831 -178
rect -1907 -228 -1831 -212
rect -1729 -178 -1653 -172
rect -1729 -212 -1708 -178
rect -1674 -212 -1653 -178
rect -1729 -228 -1653 -212
rect -1551 -178 -1475 -172
rect -1551 -212 -1530 -178
rect -1496 -212 -1475 -178
rect -1551 -228 -1475 -212
rect -1373 -178 -1297 -172
rect -1373 -212 -1352 -178
rect -1318 -212 -1297 -178
rect -1373 -228 -1297 -212
rect -1195 -178 -1119 -172
rect -1195 -212 -1174 -178
rect -1140 -212 -1119 -178
rect -1195 -228 -1119 -212
rect -1017 -178 -941 -172
rect -1017 -212 -996 -178
rect -962 -212 -941 -178
rect -1017 -228 -941 -212
rect -839 -178 -763 -172
rect -839 -212 -818 -178
rect -784 -212 -763 -178
rect -839 -228 -763 -212
rect -661 -178 -585 -172
rect -661 -212 -640 -178
rect -606 -212 -585 -178
rect -661 -228 -585 -212
rect -483 -178 -407 -172
rect -483 -212 -462 -178
rect -428 -212 -407 -178
rect -483 -228 -407 -212
rect -305 -178 -229 -172
rect -305 -212 -284 -178
rect -250 -212 -229 -178
rect -305 -228 -229 -212
rect -127 -178 -51 -172
rect -127 -212 -106 -178
rect -72 -212 -51 -178
rect -127 -228 -51 -212
rect 51 -178 127 -172
rect 51 -212 72 -178
rect 106 -212 127 -178
rect 51 -228 127 -212
rect 229 -178 305 -172
rect 229 -212 250 -178
rect 284 -212 305 -178
rect 229 -228 305 -212
rect 407 -178 483 -172
rect 407 -212 428 -178
rect 462 -212 483 -178
rect 407 -228 483 -212
rect 585 -178 661 -172
rect 585 -212 606 -178
rect 640 -212 661 -178
rect 585 -228 661 -212
rect 763 -178 839 -172
rect 763 -212 784 -178
rect 818 -212 839 -178
rect 763 -228 839 -212
rect 941 -178 1017 -172
rect 941 -212 962 -178
rect 996 -212 1017 -178
rect 941 -228 1017 -212
rect 1119 -178 1195 -172
rect 1119 -212 1140 -178
rect 1174 -212 1195 -178
rect 1119 -228 1195 -212
rect 1297 -178 1373 -172
rect 1297 -212 1318 -178
rect 1352 -212 1373 -178
rect 1297 -228 1373 -212
rect 1475 -178 1551 -172
rect 1475 -212 1496 -178
rect 1530 -212 1551 -178
rect 1475 -228 1551 -212
rect 1653 -178 1729 -172
rect 1653 -212 1674 -178
rect 1708 -212 1729 -178
rect 1653 -228 1729 -212
rect 1831 -178 1907 -172
rect 1831 -212 1852 -178
rect 1886 -212 1907 -178
rect 1831 -228 1907 -212
rect 2009 -178 2085 -172
rect 2009 -212 2030 -178
rect 2064 -212 2085 -178
rect 2009 -228 2085 -212
rect 2187 -178 2263 -172
rect 2187 -212 2208 -178
rect 2242 -212 2263 -178
rect 2187 -228 2263 -212
rect 2365 -178 2441 -172
rect 2365 -212 2386 -178
rect 2420 -212 2441 -178
rect 2365 -228 2441 -212
rect 2543 -178 2619 -172
rect 2543 -212 2564 -178
rect 2598 -212 2619 -178
rect 2543 -228 2619 -212
rect 2721 -178 2797 -172
rect 2721 -212 2742 -178
rect 2776 -212 2797 -178
rect 2721 -228 2797 -212
rect 2899 -178 2975 -172
rect 2899 -212 2920 -178
rect 2954 -212 2975 -178
rect 2899 -228 2975 -212
rect 3077 -178 3153 -172
rect 3077 -212 3098 -178
rect 3132 -212 3153 -178
rect 3077 -228 3153 -212
rect 3255 -178 3331 -172
rect 3255 -212 3276 -178
rect 3310 -212 3331 -178
rect 3255 -228 3331 -212
rect 3433 -178 3509 -172
rect 3433 -212 3454 -178
rect 3488 -212 3509 -178
rect 3433 -228 3509 -212
<< end >>
