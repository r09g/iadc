magic
tech sky130A
magscale 1 2
timestamp 1653030110
<< nmos >>
rect -3086 -140 -2966 140
rect -2908 -140 -2788 140
rect -2730 -140 -2610 140
rect -2552 -140 -2432 140
rect -2374 -140 -2254 140
rect -2196 -140 -2076 140
rect -2018 -140 -1898 140
rect -1840 -140 -1720 140
rect -1662 -140 -1542 140
rect -1484 -140 -1364 140
rect -1306 -140 -1186 140
rect -1128 -140 -1008 140
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
rect 1008 -140 1128 140
rect 1186 -140 1306 140
rect 1364 -140 1484 140
rect 1542 -140 1662 140
rect 1720 -140 1840 140
rect 1898 -140 2018 140
rect 2076 -140 2196 140
rect 2254 -140 2374 140
rect 2432 -140 2552 140
rect 2610 -140 2730 140
rect 2788 -140 2908 140
rect 2966 -140 3086 140
<< ndiff >>
rect -3144 128 -3086 140
rect -3144 -128 -3132 128
rect -3098 -128 -3086 128
rect -3144 -140 -3086 -128
rect -2966 128 -2908 140
rect -2966 -128 -2954 128
rect -2920 -128 -2908 128
rect -2966 -140 -2908 -128
rect -2788 128 -2730 140
rect -2788 -128 -2776 128
rect -2742 -128 -2730 128
rect -2788 -140 -2730 -128
rect -2610 128 -2552 140
rect -2610 -128 -2598 128
rect -2564 -128 -2552 128
rect -2610 -140 -2552 -128
rect -2432 128 -2374 140
rect -2432 -128 -2420 128
rect -2386 -128 -2374 128
rect -2432 -140 -2374 -128
rect -2254 128 -2196 140
rect -2254 -128 -2242 128
rect -2208 -128 -2196 128
rect -2254 -140 -2196 -128
rect -2076 128 -2018 140
rect -2076 -128 -2064 128
rect -2030 -128 -2018 128
rect -2076 -140 -2018 -128
rect -1898 128 -1840 140
rect -1898 -128 -1886 128
rect -1852 -128 -1840 128
rect -1898 -140 -1840 -128
rect -1720 128 -1662 140
rect -1720 -128 -1708 128
rect -1674 -128 -1662 128
rect -1720 -140 -1662 -128
rect -1542 128 -1484 140
rect -1542 -128 -1530 128
rect -1496 -128 -1484 128
rect -1542 -140 -1484 -128
rect -1364 128 -1306 140
rect -1364 -128 -1352 128
rect -1318 -128 -1306 128
rect -1364 -140 -1306 -128
rect -1186 128 -1128 140
rect -1186 -128 -1174 128
rect -1140 -128 -1128 128
rect -1186 -140 -1128 -128
rect -1008 128 -950 140
rect -1008 -128 -996 128
rect -962 -128 -950 128
rect -1008 -140 -950 -128
rect -830 128 -772 140
rect -830 -128 -818 128
rect -784 -128 -772 128
rect -830 -140 -772 -128
rect -652 128 -594 140
rect -652 -128 -640 128
rect -606 -128 -594 128
rect -652 -140 -594 -128
rect -474 128 -416 140
rect -474 -128 -462 128
rect -428 -128 -416 128
rect -474 -140 -416 -128
rect -296 128 -238 140
rect -296 -128 -284 128
rect -250 -128 -238 128
rect -296 -140 -238 -128
rect -118 128 -60 140
rect -118 -128 -106 128
rect -72 -128 -60 128
rect -118 -140 -60 -128
rect 60 128 118 140
rect 60 -128 72 128
rect 106 -128 118 128
rect 60 -140 118 -128
rect 238 128 296 140
rect 238 -128 250 128
rect 284 -128 296 128
rect 238 -140 296 -128
rect 416 128 474 140
rect 416 -128 428 128
rect 462 -128 474 128
rect 416 -140 474 -128
rect 594 128 652 140
rect 594 -128 606 128
rect 640 -128 652 128
rect 594 -140 652 -128
rect 772 128 830 140
rect 772 -128 784 128
rect 818 -128 830 128
rect 772 -140 830 -128
rect 950 128 1008 140
rect 950 -128 962 128
rect 996 -128 1008 128
rect 950 -140 1008 -128
rect 1128 128 1186 140
rect 1128 -128 1140 128
rect 1174 -128 1186 128
rect 1128 -140 1186 -128
rect 1306 128 1364 140
rect 1306 -128 1318 128
rect 1352 -128 1364 128
rect 1306 -140 1364 -128
rect 1484 128 1542 140
rect 1484 -128 1496 128
rect 1530 -128 1542 128
rect 1484 -140 1542 -128
rect 1662 128 1720 140
rect 1662 -128 1674 128
rect 1708 -128 1720 128
rect 1662 -140 1720 -128
rect 1840 128 1898 140
rect 1840 -128 1852 128
rect 1886 -128 1898 128
rect 1840 -140 1898 -128
rect 2018 128 2076 140
rect 2018 -128 2030 128
rect 2064 -128 2076 128
rect 2018 -140 2076 -128
rect 2196 128 2254 140
rect 2196 -128 2208 128
rect 2242 -128 2254 128
rect 2196 -140 2254 -128
rect 2374 128 2432 140
rect 2374 -128 2386 128
rect 2420 -128 2432 128
rect 2374 -140 2432 -128
rect 2552 128 2610 140
rect 2552 -128 2564 128
rect 2598 -128 2610 128
rect 2552 -140 2610 -128
rect 2730 128 2788 140
rect 2730 -128 2742 128
rect 2776 -128 2788 128
rect 2730 -140 2788 -128
rect 2908 128 2966 140
rect 2908 -128 2920 128
rect 2954 -128 2966 128
rect 2908 -140 2966 -128
rect 3086 128 3144 140
rect 3086 -128 3098 128
rect 3132 -128 3144 128
rect 3086 -140 3144 -128
<< ndiffc >>
rect -3132 -128 -3098 128
rect -2954 -128 -2920 128
rect -2776 -128 -2742 128
rect -2598 -128 -2564 128
rect -2420 -128 -2386 128
rect -2242 -128 -2208 128
rect -2064 -128 -2030 128
rect -1886 -128 -1852 128
rect -1708 -128 -1674 128
rect -1530 -128 -1496 128
rect -1352 -128 -1318 128
rect -1174 -128 -1140 128
rect -996 -128 -962 128
rect -818 -128 -784 128
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect 784 -128 818 128
rect 962 -128 996 128
rect 1140 -128 1174 128
rect 1318 -128 1352 128
rect 1496 -128 1530 128
rect 1674 -128 1708 128
rect 1852 -128 1886 128
rect 2030 -128 2064 128
rect 2208 -128 2242 128
rect 2386 -128 2420 128
rect 2564 -128 2598 128
rect 2742 -128 2776 128
rect 2920 -128 2954 128
rect 3098 -128 3132 128
<< poly >>
rect -3064 212 -2988 228
rect -3064 195 -3048 212
rect -3086 178 -3048 195
rect -3004 195 -2988 212
rect -2886 212 -2810 228
rect -2886 195 -2870 212
rect -3004 178 -2966 195
rect -3086 140 -2966 178
rect -2908 178 -2870 195
rect -2826 195 -2810 212
rect -2708 212 -2632 228
rect -2708 195 -2692 212
rect -2826 178 -2788 195
rect -2908 140 -2788 178
rect -2730 178 -2692 195
rect -2648 195 -2632 212
rect -2530 212 -2454 228
rect -2530 195 -2514 212
rect -2648 178 -2610 195
rect -2730 140 -2610 178
rect -2552 178 -2514 195
rect -2470 195 -2454 212
rect -2352 212 -2276 228
rect -2352 195 -2336 212
rect -2470 178 -2432 195
rect -2552 140 -2432 178
rect -2374 178 -2336 195
rect -2292 195 -2276 212
rect -2174 212 -2098 228
rect -2174 195 -2158 212
rect -2292 178 -2254 195
rect -2374 140 -2254 178
rect -2196 178 -2158 195
rect -2114 195 -2098 212
rect -1996 212 -1920 228
rect -1996 195 -1980 212
rect -2114 178 -2076 195
rect -2196 140 -2076 178
rect -2018 178 -1980 195
rect -1936 195 -1920 212
rect -1818 212 -1742 228
rect -1818 195 -1802 212
rect -1936 178 -1898 195
rect -2018 140 -1898 178
rect -1840 178 -1802 195
rect -1758 195 -1742 212
rect -1640 212 -1564 228
rect -1640 195 -1624 212
rect -1758 178 -1720 195
rect -1840 140 -1720 178
rect -1662 178 -1624 195
rect -1580 195 -1564 212
rect -1462 212 -1386 228
rect -1462 195 -1446 212
rect -1580 178 -1542 195
rect -1662 140 -1542 178
rect -1484 178 -1446 195
rect -1402 195 -1386 212
rect -1284 212 -1208 228
rect -1284 195 -1268 212
rect -1402 178 -1364 195
rect -1484 140 -1364 178
rect -1306 178 -1268 195
rect -1224 195 -1208 212
rect -1106 212 -1030 228
rect -1106 195 -1090 212
rect -1224 178 -1186 195
rect -1306 140 -1186 178
rect -1128 178 -1090 195
rect -1046 195 -1030 212
rect -928 212 -852 228
rect -928 195 -912 212
rect -1046 178 -1008 195
rect -1128 140 -1008 178
rect -950 178 -912 195
rect -868 195 -852 212
rect -750 212 -674 228
rect -750 195 -734 212
rect -868 178 -830 195
rect -950 140 -830 178
rect -772 178 -734 195
rect -690 195 -674 212
rect -572 212 -496 228
rect -572 195 -556 212
rect -690 178 -652 195
rect -772 140 -652 178
rect -594 178 -556 195
rect -512 195 -496 212
rect -394 212 -318 228
rect -394 195 -378 212
rect -512 178 -474 195
rect -594 140 -474 178
rect -416 178 -378 195
rect -334 195 -318 212
rect -216 212 -140 228
rect -216 195 -200 212
rect -334 178 -296 195
rect -416 140 -296 178
rect -238 178 -200 195
rect -156 195 -140 212
rect -38 212 38 228
rect -38 195 -22 212
rect -156 178 -118 195
rect -238 140 -118 178
rect -60 178 -22 195
rect 22 195 38 212
rect 140 212 216 228
rect 140 195 156 212
rect 22 178 60 195
rect -60 140 60 178
rect 118 178 156 195
rect 200 195 216 212
rect 318 212 394 228
rect 318 195 334 212
rect 200 178 238 195
rect 118 140 238 178
rect 296 178 334 195
rect 378 195 394 212
rect 496 212 572 228
rect 496 195 512 212
rect 378 178 416 195
rect 296 140 416 178
rect 474 178 512 195
rect 556 195 572 212
rect 674 212 750 228
rect 674 195 690 212
rect 556 178 594 195
rect 474 140 594 178
rect 652 178 690 195
rect 734 195 750 212
rect 852 212 928 228
rect 852 195 868 212
rect 734 178 772 195
rect 652 140 772 178
rect 830 178 868 195
rect 912 195 928 212
rect 1030 212 1106 228
rect 1030 195 1046 212
rect 912 178 950 195
rect 830 140 950 178
rect 1008 178 1046 195
rect 1090 195 1106 212
rect 1208 212 1284 228
rect 1208 195 1224 212
rect 1090 178 1128 195
rect 1008 140 1128 178
rect 1186 178 1224 195
rect 1268 195 1284 212
rect 1386 212 1462 228
rect 1386 195 1402 212
rect 1268 178 1306 195
rect 1186 140 1306 178
rect 1364 178 1402 195
rect 1446 195 1462 212
rect 1564 212 1640 228
rect 1564 195 1580 212
rect 1446 178 1484 195
rect 1364 140 1484 178
rect 1542 178 1580 195
rect 1624 195 1640 212
rect 1742 212 1818 228
rect 1742 195 1758 212
rect 1624 178 1662 195
rect 1542 140 1662 178
rect 1720 178 1758 195
rect 1802 195 1818 212
rect 1920 212 1996 228
rect 1920 195 1936 212
rect 1802 178 1840 195
rect 1720 140 1840 178
rect 1898 178 1936 195
rect 1980 195 1996 212
rect 2098 212 2174 228
rect 2098 195 2114 212
rect 1980 178 2018 195
rect 1898 140 2018 178
rect 2076 178 2114 195
rect 2158 195 2174 212
rect 2276 212 2352 228
rect 2276 195 2292 212
rect 2158 178 2196 195
rect 2076 140 2196 178
rect 2254 178 2292 195
rect 2336 195 2352 212
rect 2454 212 2530 228
rect 2454 195 2470 212
rect 2336 178 2374 195
rect 2254 140 2374 178
rect 2432 178 2470 195
rect 2514 195 2530 212
rect 2632 212 2708 228
rect 2632 195 2648 212
rect 2514 178 2552 195
rect 2432 140 2552 178
rect 2610 178 2648 195
rect 2692 195 2708 212
rect 2810 212 2886 228
rect 2810 195 2826 212
rect 2692 178 2730 195
rect 2610 140 2730 178
rect 2788 178 2826 195
rect 2870 195 2886 212
rect 2988 212 3064 228
rect 2988 195 3004 212
rect 2870 178 2908 195
rect 2788 140 2908 178
rect 2966 178 3004 195
rect 3048 195 3064 212
rect 3048 178 3086 195
rect 2966 140 3086 178
rect -3086 -178 -2966 -140
rect -3086 -195 -3048 -178
rect -3064 -212 -3048 -195
rect -3004 -195 -2966 -178
rect -2908 -178 -2788 -140
rect -2908 -195 -2870 -178
rect -3004 -212 -2988 -195
rect -3064 -228 -2988 -212
rect -2886 -212 -2870 -195
rect -2826 -195 -2788 -178
rect -2730 -178 -2610 -140
rect -2730 -195 -2692 -178
rect -2826 -212 -2810 -195
rect -2886 -228 -2810 -212
rect -2708 -212 -2692 -195
rect -2648 -195 -2610 -178
rect -2552 -178 -2432 -140
rect -2552 -195 -2514 -178
rect -2648 -212 -2632 -195
rect -2708 -228 -2632 -212
rect -2530 -212 -2514 -195
rect -2470 -195 -2432 -178
rect -2374 -178 -2254 -140
rect -2374 -195 -2336 -178
rect -2470 -212 -2454 -195
rect -2530 -228 -2454 -212
rect -2352 -212 -2336 -195
rect -2292 -195 -2254 -178
rect -2196 -178 -2076 -140
rect -2196 -195 -2158 -178
rect -2292 -212 -2276 -195
rect -2352 -228 -2276 -212
rect -2174 -212 -2158 -195
rect -2114 -195 -2076 -178
rect -2018 -178 -1898 -140
rect -2018 -195 -1980 -178
rect -2114 -212 -2098 -195
rect -2174 -228 -2098 -212
rect -1996 -212 -1980 -195
rect -1936 -195 -1898 -178
rect -1840 -178 -1720 -140
rect -1840 -195 -1802 -178
rect -1936 -212 -1920 -195
rect -1996 -228 -1920 -212
rect -1818 -212 -1802 -195
rect -1758 -195 -1720 -178
rect -1662 -178 -1542 -140
rect -1662 -195 -1624 -178
rect -1758 -212 -1742 -195
rect -1818 -228 -1742 -212
rect -1640 -212 -1624 -195
rect -1580 -195 -1542 -178
rect -1484 -178 -1364 -140
rect -1484 -195 -1446 -178
rect -1580 -212 -1564 -195
rect -1640 -228 -1564 -212
rect -1462 -212 -1446 -195
rect -1402 -195 -1364 -178
rect -1306 -178 -1186 -140
rect -1306 -195 -1268 -178
rect -1402 -212 -1386 -195
rect -1462 -228 -1386 -212
rect -1284 -212 -1268 -195
rect -1224 -195 -1186 -178
rect -1128 -178 -1008 -140
rect -1128 -195 -1090 -178
rect -1224 -212 -1208 -195
rect -1284 -228 -1208 -212
rect -1106 -212 -1090 -195
rect -1046 -195 -1008 -178
rect -950 -178 -830 -140
rect -950 -195 -912 -178
rect -1046 -212 -1030 -195
rect -1106 -228 -1030 -212
rect -928 -212 -912 -195
rect -868 -195 -830 -178
rect -772 -178 -652 -140
rect -772 -195 -734 -178
rect -868 -212 -852 -195
rect -928 -228 -852 -212
rect -750 -212 -734 -195
rect -690 -195 -652 -178
rect -594 -178 -474 -140
rect -594 -195 -556 -178
rect -690 -212 -674 -195
rect -750 -228 -674 -212
rect -572 -212 -556 -195
rect -512 -195 -474 -178
rect -416 -178 -296 -140
rect -416 -195 -378 -178
rect -512 -212 -496 -195
rect -572 -228 -496 -212
rect -394 -212 -378 -195
rect -334 -195 -296 -178
rect -238 -178 -118 -140
rect -238 -195 -200 -178
rect -334 -212 -318 -195
rect -394 -228 -318 -212
rect -216 -212 -200 -195
rect -156 -195 -118 -178
rect -60 -178 60 -140
rect -60 -195 -22 -178
rect -156 -212 -140 -195
rect -216 -228 -140 -212
rect -38 -212 -22 -195
rect 22 -195 60 -178
rect 118 -178 238 -140
rect 118 -195 156 -178
rect 22 -212 38 -195
rect -38 -228 38 -212
rect 140 -212 156 -195
rect 200 -195 238 -178
rect 296 -178 416 -140
rect 296 -195 334 -178
rect 200 -212 216 -195
rect 140 -228 216 -212
rect 318 -212 334 -195
rect 378 -195 416 -178
rect 474 -178 594 -140
rect 474 -195 512 -178
rect 378 -212 394 -195
rect 318 -228 394 -212
rect 496 -212 512 -195
rect 556 -195 594 -178
rect 652 -178 772 -140
rect 652 -195 690 -178
rect 556 -212 572 -195
rect 496 -228 572 -212
rect 674 -212 690 -195
rect 734 -195 772 -178
rect 830 -178 950 -140
rect 830 -195 868 -178
rect 734 -212 750 -195
rect 674 -228 750 -212
rect 852 -212 868 -195
rect 912 -195 950 -178
rect 1008 -178 1128 -140
rect 1008 -195 1046 -178
rect 912 -212 928 -195
rect 852 -228 928 -212
rect 1030 -212 1046 -195
rect 1090 -195 1128 -178
rect 1186 -178 1306 -140
rect 1186 -195 1224 -178
rect 1090 -212 1106 -195
rect 1030 -228 1106 -212
rect 1208 -212 1224 -195
rect 1268 -195 1306 -178
rect 1364 -178 1484 -140
rect 1364 -195 1402 -178
rect 1268 -212 1284 -195
rect 1208 -228 1284 -212
rect 1386 -212 1402 -195
rect 1446 -195 1484 -178
rect 1542 -178 1662 -140
rect 1542 -195 1580 -178
rect 1446 -212 1462 -195
rect 1386 -228 1462 -212
rect 1564 -212 1580 -195
rect 1624 -195 1662 -178
rect 1720 -178 1840 -140
rect 1720 -195 1758 -178
rect 1624 -212 1640 -195
rect 1564 -228 1640 -212
rect 1742 -212 1758 -195
rect 1802 -195 1840 -178
rect 1898 -178 2018 -140
rect 1898 -195 1936 -178
rect 1802 -212 1818 -195
rect 1742 -228 1818 -212
rect 1920 -212 1936 -195
rect 1980 -195 2018 -178
rect 2076 -178 2196 -140
rect 2076 -195 2114 -178
rect 1980 -212 1996 -195
rect 1920 -228 1996 -212
rect 2098 -212 2114 -195
rect 2158 -195 2196 -178
rect 2254 -178 2374 -140
rect 2254 -195 2292 -178
rect 2158 -212 2174 -195
rect 2098 -228 2174 -212
rect 2276 -212 2292 -195
rect 2336 -195 2374 -178
rect 2432 -178 2552 -140
rect 2432 -195 2470 -178
rect 2336 -212 2352 -195
rect 2276 -228 2352 -212
rect 2454 -212 2470 -195
rect 2514 -195 2552 -178
rect 2610 -178 2730 -140
rect 2610 -195 2648 -178
rect 2514 -212 2530 -195
rect 2454 -228 2530 -212
rect 2632 -212 2648 -195
rect 2692 -195 2730 -178
rect 2788 -178 2908 -140
rect 2788 -195 2826 -178
rect 2692 -212 2708 -195
rect 2632 -228 2708 -212
rect 2810 -212 2826 -195
rect 2870 -195 2908 -178
rect 2966 -178 3086 -140
rect 2966 -195 3004 -178
rect 2870 -212 2886 -195
rect 2810 -228 2886 -212
rect 2988 -212 3004 -195
rect 3048 -195 3086 -178
rect 3048 -212 3064 -195
rect 2988 -228 3064 -212
<< polycont >>
rect -3048 178 -3004 212
rect -2870 178 -2826 212
rect -2692 178 -2648 212
rect -2514 178 -2470 212
rect -2336 178 -2292 212
rect -2158 178 -2114 212
rect -1980 178 -1936 212
rect -1802 178 -1758 212
rect -1624 178 -1580 212
rect -1446 178 -1402 212
rect -1268 178 -1224 212
rect -1090 178 -1046 212
rect -912 178 -868 212
rect -734 178 -690 212
rect -556 178 -512 212
rect -378 178 -334 212
rect -200 178 -156 212
rect -22 178 22 212
rect 156 178 200 212
rect 334 178 378 212
rect 512 178 556 212
rect 690 178 734 212
rect 868 178 912 212
rect 1046 178 1090 212
rect 1224 178 1268 212
rect 1402 178 1446 212
rect 1580 178 1624 212
rect 1758 178 1802 212
rect 1936 178 1980 212
rect 2114 178 2158 212
rect 2292 178 2336 212
rect 2470 178 2514 212
rect 2648 178 2692 212
rect 2826 178 2870 212
rect 3004 178 3048 212
rect -3048 -212 -3004 -178
rect -2870 -212 -2826 -178
rect -2692 -212 -2648 -178
rect -2514 -212 -2470 -178
rect -2336 -212 -2292 -178
rect -2158 -212 -2114 -178
rect -1980 -212 -1936 -178
rect -1802 -212 -1758 -178
rect -1624 -212 -1580 -178
rect -1446 -212 -1402 -178
rect -1268 -212 -1224 -178
rect -1090 -212 -1046 -178
rect -912 -212 -868 -178
rect -734 -212 -690 -178
rect -556 -212 -512 -178
rect -378 -212 -334 -178
rect -200 -212 -156 -178
rect -22 -212 22 -178
rect 156 -212 200 -178
rect 334 -212 378 -178
rect 512 -212 556 -178
rect 690 -212 734 -178
rect 868 -212 912 -178
rect 1046 -212 1090 -178
rect 1224 -212 1268 -178
rect 1402 -212 1446 -178
rect 1580 -212 1624 -178
rect 1758 -212 1802 -178
rect 1936 -212 1980 -178
rect 2114 -212 2158 -178
rect 2292 -212 2336 -178
rect 2470 -212 2514 -178
rect 2648 -212 2692 -178
rect 2826 -212 2870 -178
rect 3004 -212 3048 -178
<< locali >>
rect -3064 178 -3048 212
rect -3004 178 -2988 212
rect -2886 178 -2870 212
rect -2826 178 -2810 212
rect -2708 178 -2692 212
rect -2648 178 -2632 212
rect -2530 178 -2514 212
rect -2470 178 -2454 212
rect -2352 178 -2336 212
rect -2292 178 -2276 212
rect -2174 178 -2158 212
rect -2114 178 -2098 212
rect -1996 178 -1980 212
rect -1936 178 -1920 212
rect -1818 178 -1802 212
rect -1758 178 -1742 212
rect -1640 178 -1624 212
rect -1580 178 -1564 212
rect -1462 178 -1446 212
rect -1402 178 -1386 212
rect -1284 178 -1268 212
rect -1224 178 -1208 212
rect -1106 178 -1090 212
rect -1046 178 -1030 212
rect -928 178 -912 212
rect -868 178 -852 212
rect -750 178 -734 212
rect -690 178 -674 212
rect -572 178 -556 212
rect -512 178 -496 212
rect -394 178 -378 212
rect -334 178 -318 212
rect -216 178 -200 212
rect -156 178 -140 212
rect -38 178 -22 212
rect 22 178 38 212
rect 140 178 156 212
rect 200 178 216 212
rect 318 178 334 212
rect 378 178 394 212
rect 496 178 512 212
rect 556 178 572 212
rect 674 178 690 212
rect 734 178 750 212
rect 852 178 868 212
rect 912 178 928 212
rect 1030 178 1046 212
rect 1090 178 1106 212
rect 1208 178 1224 212
rect 1268 178 1284 212
rect 1386 178 1402 212
rect 1446 178 1462 212
rect 1564 178 1580 212
rect 1624 178 1640 212
rect 1742 178 1758 212
rect 1802 178 1818 212
rect 1920 178 1936 212
rect 1980 178 1996 212
rect 2098 178 2114 212
rect 2158 178 2174 212
rect 2276 178 2292 212
rect 2336 178 2352 212
rect 2454 178 2470 212
rect 2514 178 2530 212
rect 2632 178 2648 212
rect 2692 178 2708 212
rect 2810 178 2826 212
rect 2870 178 2886 212
rect 2988 178 3004 212
rect 3048 178 3064 212
rect -3132 128 -3098 144
rect -3132 -144 -3098 -128
rect -2954 128 -2920 144
rect -2954 -144 -2920 -128
rect -2776 128 -2742 144
rect -2776 -144 -2742 -128
rect -2598 128 -2564 144
rect -2598 -144 -2564 -128
rect -2420 128 -2386 144
rect -2420 -144 -2386 -128
rect -2242 128 -2208 144
rect -2242 -144 -2208 -128
rect -2064 128 -2030 144
rect -2064 -144 -2030 -128
rect -1886 128 -1852 144
rect -1886 -144 -1852 -128
rect -1708 128 -1674 144
rect -1708 -144 -1674 -128
rect -1530 128 -1496 144
rect -1530 -144 -1496 -128
rect -1352 128 -1318 144
rect -1352 -144 -1318 -128
rect -1174 128 -1140 144
rect -1174 -144 -1140 -128
rect -996 128 -962 144
rect -996 -144 -962 -128
rect -818 128 -784 144
rect -818 -144 -784 -128
rect -640 128 -606 144
rect -640 -144 -606 -128
rect -462 128 -428 144
rect -462 -144 -428 -128
rect -284 128 -250 144
rect -284 -144 -250 -128
rect -106 128 -72 144
rect -106 -144 -72 -128
rect 72 128 106 144
rect 72 -144 106 -128
rect 250 128 284 144
rect 250 -144 284 -128
rect 428 128 462 144
rect 428 -144 462 -128
rect 606 128 640 144
rect 606 -144 640 -128
rect 784 128 818 144
rect 784 -144 818 -128
rect 962 128 996 144
rect 962 -144 996 -128
rect 1140 128 1174 144
rect 1140 -144 1174 -128
rect 1318 128 1352 144
rect 1318 -144 1352 -128
rect 1496 128 1530 144
rect 1496 -144 1530 -128
rect 1674 128 1708 144
rect 1674 -144 1708 -128
rect 1852 128 1886 144
rect 1852 -144 1886 -128
rect 2030 128 2064 144
rect 2030 -144 2064 -128
rect 2208 128 2242 144
rect 2208 -144 2242 -128
rect 2386 128 2420 144
rect 2386 -144 2420 -128
rect 2564 128 2598 144
rect 2564 -144 2598 -128
rect 2742 128 2776 144
rect 2742 -144 2776 -128
rect 2920 128 2954 144
rect 2920 -144 2954 -128
rect 3098 128 3132 144
rect 3098 -144 3132 -128
rect -3064 -212 -3048 -178
rect -3004 -212 -2988 -178
rect -2886 -212 -2870 -178
rect -2826 -212 -2810 -178
rect -2708 -212 -2692 -178
rect -2648 -212 -2632 -178
rect -2530 -212 -2514 -178
rect -2470 -212 -2454 -178
rect -2352 -212 -2336 -178
rect -2292 -212 -2276 -178
rect -2174 -212 -2158 -178
rect -2114 -212 -2098 -178
rect -1996 -212 -1980 -178
rect -1936 -212 -1920 -178
rect -1818 -212 -1802 -178
rect -1758 -212 -1742 -178
rect -1640 -212 -1624 -178
rect -1580 -212 -1564 -178
rect -1462 -212 -1446 -178
rect -1402 -212 -1386 -178
rect -1284 -212 -1268 -178
rect -1224 -212 -1208 -178
rect -1106 -212 -1090 -178
rect -1046 -212 -1030 -178
rect -928 -212 -912 -178
rect -868 -212 -852 -178
rect -750 -212 -734 -178
rect -690 -212 -674 -178
rect -572 -212 -556 -178
rect -512 -212 -496 -178
rect -394 -212 -378 -178
rect -334 -212 -318 -178
rect -216 -212 -200 -178
rect -156 -212 -140 -178
rect -38 -212 -22 -178
rect 22 -212 38 -178
rect 140 -212 156 -178
rect 200 -212 216 -178
rect 318 -212 334 -178
rect 378 -212 394 -178
rect 496 -212 512 -178
rect 556 -212 572 -178
rect 674 -212 690 -178
rect 734 -212 750 -178
rect 852 -212 868 -178
rect 912 -212 928 -178
rect 1030 -212 1046 -178
rect 1090 -212 1106 -178
rect 1208 -212 1224 -178
rect 1268 -212 1284 -178
rect 1386 -212 1402 -178
rect 1446 -212 1462 -178
rect 1564 -212 1580 -178
rect 1624 -212 1640 -178
rect 1742 -212 1758 -178
rect 1802 -212 1818 -178
rect 1920 -212 1936 -178
rect 1980 -212 1996 -178
rect 2098 -212 2114 -178
rect 2158 -212 2174 -178
rect 2276 -212 2292 -178
rect 2336 -212 2352 -178
rect 2454 -212 2470 -178
rect 2514 -212 2530 -178
rect 2632 -212 2648 -178
rect 2692 -212 2708 -178
rect 2810 -212 2826 -178
rect 2870 -212 2886 -178
rect 2988 -212 3004 -178
rect 3048 -212 3064 -178
<< viali >>
rect -3048 178 -3004 212
rect -2870 178 -2826 212
rect -2692 178 -2648 212
rect -2514 178 -2470 212
rect -2336 178 -2292 212
rect -2158 178 -2114 212
rect -1980 178 -1936 212
rect -1802 178 -1758 212
rect -1624 178 -1580 212
rect -1446 178 -1402 212
rect -1268 178 -1224 212
rect -1090 178 -1046 212
rect -912 178 -868 212
rect -734 178 -690 212
rect -556 178 -512 212
rect -378 178 -334 212
rect -200 178 -156 212
rect -22 178 22 212
rect 156 178 200 212
rect 334 178 378 212
rect 512 178 556 212
rect 690 178 734 212
rect 868 178 912 212
rect 1046 178 1090 212
rect 1224 178 1268 212
rect 1402 178 1446 212
rect 1580 178 1624 212
rect 1758 178 1802 212
rect 1936 178 1980 212
rect 2114 178 2158 212
rect 2292 178 2336 212
rect 2470 178 2514 212
rect 2648 178 2692 212
rect 2826 178 2870 212
rect 3004 178 3048 212
rect -3132 -128 -3098 128
rect -2954 -128 -2920 128
rect -2776 -128 -2742 128
rect -2598 -128 -2564 128
rect -2420 -128 -2386 128
rect -2242 -128 -2208 128
rect -2064 -128 -2030 128
rect -1886 -128 -1852 128
rect -1708 -128 -1674 128
rect -1530 -128 -1496 128
rect -1352 -128 -1318 128
rect -1174 -128 -1140 128
rect -996 -128 -962 128
rect -818 -128 -784 128
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect 784 -128 818 128
rect 962 -128 996 128
rect 1140 -128 1174 128
rect 1318 -128 1352 128
rect 1496 -128 1530 128
rect 1674 -128 1708 128
rect 1852 -128 1886 128
rect 2030 -128 2064 128
rect 2208 -128 2242 128
rect 2386 -128 2420 128
rect 2564 -128 2598 128
rect 2742 -128 2776 128
rect 2920 -128 2954 128
rect 3098 -128 3132 128
rect -3048 -212 -3004 -178
rect -2870 -212 -2826 -178
rect -2692 -212 -2648 -178
rect -2514 -212 -2470 -178
rect -2336 -212 -2292 -178
rect -2158 -212 -2114 -178
rect -1980 -212 -1936 -178
rect -1802 -212 -1758 -178
rect -1624 -212 -1580 -178
rect -1446 -212 -1402 -178
rect -1268 -212 -1224 -178
rect -1090 -212 -1046 -178
rect -912 -212 -868 -178
rect -734 -212 -690 -178
rect -556 -212 -512 -178
rect -378 -212 -334 -178
rect -200 -212 -156 -178
rect -22 -212 22 -178
rect 156 -212 200 -178
rect 334 -212 378 -178
rect 512 -212 556 -178
rect 690 -212 734 -178
rect 868 -212 912 -178
rect 1046 -212 1090 -178
rect 1224 -212 1268 -178
rect 1402 -212 1446 -178
rect 1580 -212 1624 -178
rect 1758 -212 1802 -178
rect 1936 -212 1980 -178
rect 2114 -212 2158 -178
rect 2292 -212 2336 -178
rect 2470 -212 2514 -178
rect 2648 -212 2692 -178
rect 2826 -212 2870 -178
rect 3004 -212 3048 -178
<< metal1 >>
rect -3064 212 -2988 228
rect -3064 178 -3048 212
rect -3004 178 -2988 212
rect -3064 172 -2988 178
rect -2886 212 -2810 228
rect -2886 178 -2870 212
rect -2826 178 -2810 212
rect -2886 172 -2810 178
rect -2708 212 -2632 228
rect -2708 178 -2692 212
rect -2648 178 -2632 212
rect -2708 172 -2632 178
rect -2530 212 -2454 228
rect -2530 178 -2514 212
rect -2470 178 -2454 212
rect -2530 172 -2454 178
rect -2352 212 -2276 228
rect -2352 178 -2336 212
rect -2292 178 -2276 212
rect -2352 172 -2276 178
rect -2174 212 -2098 228
rect -2174 178 -2158 212
rect -2114 178 -2098 212
rect -2174 172 -2098 178
rect -1996 212 -1920 228
rect -1996 178 -1980 212
rect -1936 178 -1920 212
rect -1996 172 -1920 178
rect -1818 212 -1742 228
rect -1818 178 -1802 212
rect -1758 178 -1742 212
rect -1818 172 -1742 178
rect -1640 212 -1564 228
rect -1640 178 -1624 212
rect -1580 178 -1564 212
rect -1640 172 -1564 178
rect -1462 212 -1386 228
rect -1462 178 -1446 212
rect -1402 178 -1386 212
rect -1462 172 -1386 178
rect -1284 212 -1208 228
rect -1284 178 -1268 212
rect -1224 178 -1208 212
rect -1284 172 -1208 178
rect -1106 212 -1030 228
rect -1106 178 -1090 212
rect -1046 178 -1030 212
rect -1106 172 -1030 178
rect -928 212 -852 228
rect -928 178 -912 212
rect -868 178 -852 212
rect -928 172 -852 178
rect -750 212 -674 228
rect -750 178 -734 212
rect -690 178 -674 212
rect -750 172 -674 178
rect -572 212 -496 228
rect -572 178 -556 212
rect -512 178 -496 212
rect -572 172 -496 178
rect -394 212 -318 228
rect -394 178 -378 212
rect -334 178 -318 212
rect -394 172 -318 178
rect -216 212 -140 228
rect -216 178 -200 212
rect -156 178 -140 212
rect -216 172 -140 178
rect -38 212 38 228
rect -38 178 -22 212
rect 22 178 38 212
rect -38 172 38 178
rect 140 212 216 228
rect 140 178 156 212
rect 200 178 216 212
rect 140 172 216 178
rect 318 212 394 228
rect 318 178 334 212
rect 378 178 394 212
rect 318 172 394 178
rect 496 212 572 228
rect 496 178 512 212
rect 556 178 572 212
rect 496 172 572 178
rect 674 212 750 228
rect 674 178 690 212
rect 734 178 750 212
rect 674 172 750 178
rect 852 212 928 228
rect 852 178 868 212
rect 912 178 928 212
rect 852 172 928 178
rect 1030 212 1106 228
rect 1030 178 1046 212
rect 1090 178 1106 212
rect 1030 172 1106 178
rect 1208 212 1284 228
rect 1208 178 1224 212
rect 1268 178 1284 212
rect 1208 172 1284 178
rect 1386 212 1462 228
rect 1386 178 1402 212
rect 1446 178 1462 212
rect 1386 172 1462 178
rect 1564 212 1640 228
rect 1564 178 1580 212
rect 1624 178 1640 212
rect 1564 172 1640 178
rect 1742 212 1818 228
rect 1742 178 1758 212
rect 1802 178 1818 212
rect 1742 172 1818 178
rect 1920 212 1996 228
rect 1920 178 1936 212
rect 1980 178 1996 212
rect 1920 172 1996 178
rect 2098 212 2174 228
rect 2098 178 2114 212
rect 2158 178 2174 212
rect 2098 172 2174 178
rect 2276 212 2352 228
rect 2276 178 2292 212
rect 2336 178 2352 212
rect 2276 172 2352 178
rect 2454 212 2530 228
rect 2454 178 2470 212
rect 2514 178 2530 212
rect 2454 172 2530 178
rect 2632 212 2708 228
rect 2632 178 2648 212
rect 2692 178 2708 212
rect 2632 172 2708 178
rect 2810 212 2886 228
rect 2810 178 2826 212
rect 2870 178 2886 212
rect 2810 172 2886 178
rect 2988 212 3064 228
rect 2988 178 3004 212
rect 3048 178 3064 212
rect 2988 172 3064 178
rect -3138 128 -3092 140
rect -3138 -128 -3132 128
rect -3098 -128 -3092 128
rect -3138 -140 -3092 -128
rect -2960 128 -2914 140
rect -2960 -128 -2954 128
rect -2920 -128 -2914 128
rect -2960 -140 -2914 -128
rect -2782 128 -2736 140
rect -2782 -128 -2776 128
rect -2742 -128 -2736 128
rect -2782 -140 -2736 -128
rect -2604 128 -2558 140
rect -2604 -128 -2598 128
rect -2564 -128 -2558 128
rect -2604 -140 -2558 -128
rect -2426 128 -2380 140
rect -2426 -128 -2420 128
rect -2386 -128 -2380 128
rect -2426 -140 -2380 -128
rect -2248 128 -2202 140
rect -2248 -128 -2242 128
rect -2208 -128 -2202 128
rect -2248 -140 -2202 -128
rect -2070 128 -2024 140
rect -2070 -128 -2064 128
rect -2030 -128 -2024 128
rect -2070 -140 -2024 -128
rect -1892 128 -1846 140
rect -1892 -128 -1886 128
rect -1852 -128 -1846 128
rect -1892 -140 -1846 -128
rect -1714 128 -1668 140
rect -1714 -128 -1708 128
rect -1674 -128 -1668 128
rect -1714 -140 -1668 -128
rect -1536 128 -1490 140
rect -1536 -128 -1530 128
rect -1496 -128 -1490 128
rect -1536 -140 -1490 -128
rect -1358 128 -1312 140
rect -1358 -128 -1352 128
rect -1318 -128 -1312 128
rect -1358 -140 -1312 -128
rect -1180 128 -1134 140
rect -1180 -128 -1174 128
rect -1140 -128 -1134 128
rect -1180 -140 -1134 -128
rect -1002 128 -956 140
rect -1002 -128 -996 128
rect -962 -128 -956 128
rect -1002 -140 -956 -128
rect -824 128 -778 140
rect -824 -128 -818 128
rect -784 -128 -778 128
rect -824 -140 -778 -128
rect -646 128 -600 140
rect -646 -128 -640 128
rect -606 -128 -600 128
rect -646 -140 -600 -128
rect -468 128 -422 140
rect -468 -128 -462 128
rect -428 -128 -422 128
rect -468 -140 -422 -128
rect -290 128 -244 140
rect -290 -128 -284 128
rect -250 -128 -244 128
rect -290 -140 -244 -128
rect -112 128 -66 140
rect -112 -128 -106 128
rect -72 -128 -66 128
rect -112 -140 -66 -128
rect 66 128 112 140
rect 66 -128 72 128
rect 106 -128 112 128
rect 66 -140 112 -128
rect 244 128 290 140
rect 244 -128 250 128
rect 284 -128 290 128
rect 244 -140 290 -128
rect 422 128 468 140
rect 422 -128 428 128
rect 462 -128 468 128
rect 422 -140 468 -128
rect 600 128 646 140
rect 600 -128 606 128
rect 640 -128 646 128
rect 600 -140 646 -128
rect 778 128 824 140
rect 778 -128 784 128
rect 818 -128 824 128
rect 778 -140 824 -128
rect 956 128 1002 140
rect 956 -128 962 128
rect 996 -128 1002 128
rect 956 -140 1002 -128
rect 1134 128 1180 140
rect 1134 -128 1140 128
rect 1174 -128 1180 128
rect 1134 -140 1180 -128
rect 1312 128 1358 140
rect 1312 -128 1318 128
rect 1352 -128 1358 128
rect 1312 -140 1358 -128
rect 1490 128 1536 140
rect 1490 -128 1496 128
rect 1530 -128 1536 128
rect 1490 -140 1536 -128
rect 1668 128 1714 140
rect 1668 -128 1674 128
rect 1708 -128 1714 128
rect 1668 -140 1714 -128
rect 1846 128 1892 140
rect 1846 -128 1852 128
rect 1886 -128 1892 128
rect 1846 -140 1892 -128
rect 2024 128 2070 140
rect 2024 -128 2030 128
rect 2064 -128 2070 128
rect 2024 -140 2070 -128
rect 2202 128 2248 140
rect 2202 -128 2208 128
rect 2242 -128 2248 128
rect 2202 -140 2248 -128
rect 2380 128 2426 140
rect 2380 -128 2386 128
rect 2420 -128 2426 128
rect 2380 -140 2426 -128
rect 2558 128 2604 140
rect 2558 -128 2564 128
rect 2598 -128 2604 128
rect 2558 -140 2604 -128
rect 2736 128 2782 140
rect 2736 -128 2742 128
rect 2776 -128 2782 128
rect 2736 -140 2782 -128
rect 2914 128 2960 140
rect 2914 -128 2920 128
rect 2954 -128 2960 128
rect 2914 -140 2960 -128
rect 3092 128 3138 140
rect 3092 -128 3098 128
rect 3132 -128 3138 128
rect 3092 -140 3138 -128
rect -3064 -178 -2988 -172
rect -3064 -212 -3048 -178
rect -3004 -212 -2988 -178
rect -3064 -228 -2988 -212
rect -2886 -178 -2810 -172
rect -2886 -212 -2870 -178
rect -2826 -212 -2810 -178
rect -2886 -228 -2810 -212
rect -2708 -178 -2632 -172
rect -2708 -212 -2692 -178
rect -2648 -212 -2632 -178
rect -2708 -228 -2632 -212
rect -2530 -178 -2454 -172
rect -2530 -212 -2514 -178
rect -2470 -212 -2454 -178
rect -2530 -228 -2454 -212
rect -2352 -178 -2276 -172
rect -2352 -212 -2336 -178
rect -2292 -212 -2276 -178
rect -2352 -228 -2276 -212
rect -2174 -178 -2098 -172
rect -2174 -212 -2158 -178
rect -2114 -212 -2098 -178
rect -2174 -228 -2098 -212
rect -1996 -178 -1920 -172
rect -1996 -212 -1980 -178
rect -1936 -212 -1920 -178
rect -1996 -228 -1920 -212
rect -1818 -178 -1742 -172
rect -1818 -212 -1802 -178
rect -1758 -212 -1742 -178
rect -1818 -228 -1742 -212
rect -1640 -178 -1564 -172
rect -1640 -212 -1624 -178
rect -1580 -212 -1564 -178
rect -1640 -228 -1564 -212
rect -1462 -178 -1386 -172
rect -1462 -212 -1446 -178
rect -1402 -212 -1386 -178
rect -1462 -228 -1386 -212
rect -1284 -178 -1208 -172
rect -1284 -212 -1268 -178
rect -1224 -212 -1208 -178
rect -1284 -228 -1208 -212
rect -1106 -178 -1030 -172
rect -1106 -212 -1090 -178
rect -1046 -212 -1030 -178
rect -1106 -228 -1030 -212
rect -928 -178 -852 -172
rect -928 -212 -912 -178
rect -868 -212 -852 -178
rect -928 -228 -852 -212
rect -750 -178 -674 -172
rect -750 -212 -734 -178
rect -690 -212 -674 -178
rect -750 -228 -674 -212
rect -572 -178 -496 -172
rect -572 -212 -556 -178
rect -512 -212 -496 -178
rect -572 -228 -496 -212
rect -394 -178 -318 -172
rect -394 -212 -378 -178
rect -334 -212 -318 -178
rect -394 -228 -318 -212
rect -216 -178 -140 -172
rect -216 -212 -200 -178
rect -156 -212 -140 -178
rect -216 -228 -140 -212
rect -38 -178 38 -172
rect -38 -212 -22 -178
rect 22 -212 38 -178
rect -38 -228 38 -212
rect 140 -178 216 -172
rect 140 -212 156 -178
rect 200 -212 216 -178
rect 140 -228 216 -212
rect 318 -178 394 -172
rect 318 -212 334 -178
rect 378 -212 394 -178
rect 318 -228 394 -212
rect 496 -178 572 -172
rect 496 -212 512 -178
rect 556 -212 572 -178
rect 496 -228 572 -212
rect 674 -178 750 -172
rect 674 -212 690 -178
rect 734 -212 750 -178
rect 674 -228 750 -212
rect 852 -178 928 -172
rect 852 -212 868 -178
rect 912 -212 928 -178
rect 852 -228 928 -212
rect 1030 -178 1106 -172
rect 1030 -212 1046 -178
rect 1090 -212 1106 -178
rect 1030 -228 1106 -212
rect 1208 -178 1284 -172
rect 1208 -212 1224 -178
rect 1268 -212 1284 -178
rect 1208 -228 1284 -212
rect 1386 -178 1462 -172
rect 1386 -212 1402 -178
rect 1446 -212 1462 -178
rect 1386 -228 1462 -212
rect 1564 -178 1640 -172
rect 1564 -212 1580 -178
rect 1624 -212 1640 -178
rect 1564 -228 1640 -212
rect 1742 -178 1818 -172
rect 1742 -212 1758 -178
rect 1802 -212 1818 -178
rect 1742 -228 1818 -212
rect 1920 -178 1996 -172
rect 1920 -212 1936 -178
rect 1980 -212 1996 -178
rect 1920 -228 1996 -212
rect 2098 -178 2174 -172
rect 2098 -212 2114 -178
rect 2158 -212 2174 -178
rect 2098 -228 2174 -212
rect 2276 -178 2352 -172
rect 2276 -212 2292 -178
rect 2336 -212 2352 -178
rect 2276 -228 2352 -212
rect 2454 -178 2530 -172
rect 2454 -212 2470 -178
rect 2514 -212 2530 -178
rect 2454 -228 2530 -212
rect 2632 -178 2708 -172
rect 2632 -212 2648 -178
rect 2692 -212 2708 -178
rect 2632 -228 2708 -212
rect 2810 -178 2886 -172
rect 2810 -212 2826 -178
rect 2870 -212 2886 -178
rect 2810 -228 2886 -212
rect 2988 -178 3064 -172
rect 2988 -212 3004 -178
rect 3048 -212 3064 -178
rect 2988 -228 3064 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 35 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
