magic
tech sky130A
magscale 1 2
timestamp 1654713294
<< locali >>
rect 6609 19960 6865 20216
rect -61 8576 5805 8582
rect -61 8332 5555 8576
rect 5799 8332 5805 8576
rect -61 8326 5805 8332
rect 23491 8569 23747 8575
rect -61 18 195 8326
rect 23491 8325 23497 8569
rect 23741 8325 23747 8569
rect 7193 6918 7449 7996
rect 11584 6968 11840 7996
rect 16315 6980 16571 7996
rect 21581 6945 21837 8022
rect 23491 280 23747 8325
rect 21894 24 23747 280
<< viali >>
rect 8715 8761 8971 9017
rect 19650 8749 19906 9005
rect 5555 8332 5799 8576
rect 23497 8325 23741 8569
<< metal1 >>
rect 6805 14170 6815 14689
rect 6910 14170 6920 14689
rect 5451 13073 5457 13485
rect 5869 13073 5875 13485
rect 6338 11514 6348 11637
rect 6458 11514 6468 11637
rect 6329 11102 6335 11514
rect 6747 11102 6753 11514
rect 21875 11225 21885 11732
rect 21996 11539 22006 11732
rect 21997 11429 22006 11539
rect 21996 11225 22006 11429
rect 6338 11097 6348 11102
rect 6458 11097 6468 11102
rect 22389 9295 22399 9835
rect 22509 9295 22519 9835
rect 8703 9017 8983 9023
rect 8703 8761 8715 9017
rect 8971 8761 8983 9017
rect 8703 8755 8983 8761
rect 19638 9005 19918 9011
rect 8715 8582 8971 8755
rect 19638 8749 19650 9005
rect 19906 8749 19918 9005
rect 19638 8743 19918 8749
rect 5543 8576 8971 8582
rect 5543 8332 5555 8576
rect 5799 8332 8971 8576
rect 5543 8326 8971 8332
rect 19650 8575 19906 8743
rect 19650 8569 23753 8575
rect 19650 8325 23497 8569
rect 23741 8325 23753 8569
rect 19650 8319 23753 8325
rect 2937 4263 2993 5118
rect 4720 4263 4776 5118
rect 9761 4008 17630 4125
rect 647 3692 657 3802
rect 767 3692 777 3802
rect 21251 1092 22312 1220
<< via1 >>
rect 6815 14170 6910 14689
rect 5457 13073 5869 13485
rect 6348 11514 6458 11637
rect 6335 11102 6747 11514
rect 21885 11539 21996 11732
rect 21885 11429 21997 11539
rect 21885 11225 21996 11429
rect 6348 11097 6458 11102
rect 22399 9295 22509 9835
rect 657 3692 767 3802
<< metal2 >>
rect 6815 14689 6910 14699
rect 613 14302 6815 14508
rect 613 3802 819 14302
rect 6910 14302 6912 14508
rect 6815 14160 6910 14170
rect 5457 13485 5869 13491
rect 5457 10415 5869 13073
rect 21885 11732 21996 11742
rect 6335 11649 6747 11670
rect 6331 11637 6747 11649
rect 6331 11514 6348 11637
rect 6458 11514 6747 11637
rect 23475 11592 23656 11602
rect 6331 11443 6335 11514
rect 6334 11102 6335 11105
rect 21881 11429 21885 11539
rect 21997 11429 23475 11539
rect 23475 11363 23656 11373
rect 21885 11215 21996 11225
rect 6334 11097 6348 11102
rect 6458 11097 6747 11102
rect 6334 10899 6747 11097
rect 5457 4656 5870 10415
rect 5457 4254 5462 4656
rect 5864 4455 5870 4656
rect 5457 4249 5664 4254
rect 5462 4245 5870 4249
rect 5664 4210 5870 4245
rect 613 3692 657 3802
rect 767 3692 819 3802
rect 613 3682 819 3692
rect 6335 3586 6747 10899
rect 22387 9835 22593 9877
rect 22387 9295 22399 9835
rect 22509 9295 22593 9835
rect 19353 4834 19411 5532
rect 20331 5141 20462 5841
rect 8757 4454 8881 4464
rect 8757 4239 8881 4249
rect 11452 3588 11558 3598
rect 6331 3184 6340 3586
rect 6742 3184 6751 3586
rect 11558 3379 11561 3388
rect 6335 3179 6747 3184
rect 11558 3270 11561 3279
rect 11452 3172 11558 3182
rect 17433 3017 17535 3018
rect 17432 3008 17542 3017
rect 17432 3007 17433 3008
rect 17535 3007 17542 3008
rect 17432 2887 17433 2897
rect 17535 2887 17542 2897
rect 22387 3004 22593 9295
rect 17433 2793 17535 2803
rect 22387 2788 22593 2798
<< via2 >>
rect 23475 11373 23656 11592
rect 5462 4455 5864 4656
rect 5462 4254 5870 4455
rect 5664 4249 5870 4254
rect 8757 4249 8881 4454
rect 6340 3184 6742 3586
rect 11452 3379 11558 3588
rect 11452 3279 11561 3379
rect 11452 3182 11558 3279
rect 17433 3007 17535 3008
rect 17432 2897 17542 3007
rect 17433 2803 17535 2897
rect 22387 2798 22593 3004
<< metal3 >>
rect 23462 11592 23668 11618
rect 23462 11373 23475 11592
rect 23656 11373 23668 11592
rect 5457 4656 8891 4661
rect 5457 4254 5462 4656
rect 5864 4455 8891 4656
rect 5870 4454 8891 4455
rect 5457 4249 5664 4254
rect 5870 4249 8757 4454
rect 8881 4249 8891 4454
rect 5654 4244 5880 4249
rect 8747 4244 8891 4249
rect 23462 3833 23668 11373
rect 13209 3627 23668 3833
rect 11442 3591 11568 3593
rect 6335 3588 11579 3591
rect 6335 3586 11452 3588
rect 6335 3394 6340 3586
rect 6333 3210 6340 3394
rect 6335 3184 6340 3210
rect 6742 3184 11452 3586
rect 11558 3379 11579 3588
rect 11561 3279 11579 3379
rect 6335 3182 11452 3184
rect 11558 3182 11579 3279
rect 6335 3179 11579 3182
rect 11442 3177 11568 3179
rect 13209 2681 13415 3627
rect 17423 3012 17545 3013
rect 17422 3008 17552 3012
rect 17422 3007 17433 3008
rect 17535 3007 17552 3008
rect 17422 2897 17432 3007
rect 17542 3006 17552 3007
rect 22377 3006 22603 3009
rect 17542 3004 22603 3006
rect 17542 2897 22387 3004
rect 17422 2892 17433 2897
rect 17423 2803 17433 2892
rect 17535 2803 22387 2897
rect 17423 2800 22387 2803
rect 17423 2798 17545 2800
rect 22377 2798 22387 2800
rect 22593 2798 22603 3004
rect 22377 2793 22603 2798
rect -170 2475 13415 2681
<< metal4 >>
rect 7353 20556 21191 20620
rect 7272 20156 7581 20220
rect 7272 19756 7872 19820
rect 7272 19356 8182 19420
use ota_v2_without_cmfb  ota_v2_without_cmfb_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/ota_v2
timestamp 1654712441
transform -1 0 21026 0 1 335
box -1045 -334 21142 6713
use sc_cmfb  sc_cmfb_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout_v2/sc_cmfb
timestamp 1654713294
transform 1 0 11071 0 1 10659
box -5376 -2919 11546 9969
<< labels >>
flabel metal1 2965 4960 2965 4960 1 FreeSans 800 0 0 0 in
port 2 n
flabel metal1 4751 4964 4751 4964 1 FreeSans 800 0 0 0 ip
port 1 n
flabel metal4 7524 20588 7524 20588 1 FreeSans 800 0 0 0 p2_b
port 6 n
flabel metal4 7520 20183 7520 20183 1 FreeSans 800 0 0 0 p2
port 5 n
flabel metal4 7522 19788 7522 19788 1 FreeSans 800 0 0 0 p1_b
port 4 n
flabel metal4 7522 19380 7522 19380 1 FreeSans 800 0 0 0 p1
port 3 n
flabel metal2 5790 8141 5790 8141 1 FreeSans 800 0 0 0 op
port 7 n
flabel metal2 6403 8150 6403 8150 1 FreeSans 800 0 0 0 on
port 8 n
flabel metal1 22248 1153 22248 1153 1 FreeSans 800 0 0 0 i_bias
port 9 n
flabel metal3 -153 2588 -153 2588 1 FreeSans 800 0 0 0 cm
port 10 n
flabel locali 6730 20089 6730 20089 1 FreeSans 800 0 0 0 VDD
port 16 n power bidirectional
flabel locali 11 93 11 93 1 FreeSans 800 0 0 0 VSS
port 17 n power bidirectional
flabel metal2 22492 5814 22492 5814 1 FreeSans 800 0 0 0 bias_a
port 11 n
flabel metal2 19379 5290 19379 5290 1 FreeSans 800 0 0 0 bias_c
port 13 n
flabel metal2 20397 5292 20397 5292 1 FreeSans 800 0 0 0 bias_b
port 12 n
flabel metal2 708 5110 708 5110 1 FreeSans 800 0 0 0 cmc
port 15 n
flabel metal1 16024 4072 16024 4072 1 FreeSans 800 0 0 0 bias_d
port 14 n
<< end >>
