magic
tech sky130A
magscale 1 2
timestamp 1654899744
<< metal2 >>
rect 372200 516868 372209 516928
rect 372269 516912 372278 516928
rect 373663 516912 373691 522678
rect 402367 519092 402395 520676
rect 424601 519108 424661 519117
rect 402367 519064 424601 519092
rect 424601 519039 424661 519048
rect 372269 516884 373691 516912
rect 372269 516868 372278 516884
rect 373663 504711 373691 507736
rect 383231 504757 383259 507813
rect 373647 504702 373707 504711
rect 383206 504697 383215 504757
rect 383275 504697 383284 504757
rect 392799 504716 392827 507951
rect 392774 504656 392783 504716
rect 392843 504656 392852 504716
rect 373647 504633 373707 504642
rect 481589 44783 481598 44895
rect 481710 44783 481719 44895
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 44783
rect 485135 44774 485144 44886
rect 485256 44774 485265 44886
rect 482771 16673 482780 16785
rect 482892 16673 482901 16785
rect 482780 -800 482892 16673
rect 483962 -800 484074 480
rect 485144 -800 485256 44774
rect 488681 44762 488690 44874
rect 488802 44762 488811 44874
rect 486317 16718 486326 16830
rect 486438 16718 486447 16830
rect 486326 -800 486438 16718
rect 487508 -800 487620 480
rect 488690 -800 488802 44762
rect 489872 16753 489984 16762
rect 489872 -800 489984 16641
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 372209 516868 372269 516928
rect 424601 519048 424661 519108
rect 373647 504642 373707 504702
rect 383215 504697 383275 504757
rect 392783 504656 392843 504716
rect 481598 44783 481710 44895
rect 485144 44774 485256 44886
rect 482780 16673 482892 16785
rect 488690 44762 488802 44874
rect 486326 16718 486438 16830
rect 489872 16641 489984 16753
<< metal3 >>
rect 16194 702737 21194 704800
rect 15877 695646 21331 702737
rect 68194 702547 73194 704800
rect 120194 702701 125194 704800
rect 49727 695646 55181 695653
rect 15877 690192 55181 695646
rect 558 685242 41326 685356
rect -800 680242 41326 685242
rect 558 679902 41326 680242
rect 5371 648752 8383 648776
rect 805 648642 8383 648752
rect -800 643842 8383 648642
rect 805 643688 8383 643842
rect 13471 643688 13477 648776
rect 805 643686 5945 643688
rect 5371 638726 8391 638742
rect 805 638642 8391 638726
rect -800 633842 8391 638642
rect 805 633670 8391 633842
rect 13463 633670 13469 638742
rect 805 633660 5945 633670
rect 35872 617459 41326 679902
rect 49727 657865 55181 690192
rect 68098 673045 73321 702547
rect 119810 690196 125221 702701
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702955 418394 704800
rect 465394 703014 470394 704800
rect 413191 690689 418453 702955
rect 119810 684785 260348 690196
rect 68098 667822 227958 673045
rect 49727 652411 203813 657865
rect 198359 646060 203813 652411
rect 222735 646060 227958 667822
rect 254937 646060 260348 684785
rect 285478 685427 418453 690689
rect 465252 702300 470394 703014
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 703689 571594 704800
rect 285478 646060 290740 685427
rect 465252 675437 470365 702300
rect 566410 693330 571704 703689
rect 308691 670324 470365 675437
rect 501739 688036 571704 693330
rect 308691 646060 313804 670324
rect 501739 655869 507033 688036
rect 571542 682984 582953 683337
rect 571542 677984 584800 682984
rect 571542 677569 582953 677984
rect 571542 665727 577310 677569
rect 342062 650575 507033 655869
rect 530161 659959 577310 665727
rect 342062 646060 347356 650575
rect 199510 623965 200510 646060
rect 224356 628106 225356 646060
rect 257844 640529 258844 646060
rect 238371 639529 258844 640529
rect 224356 627106 232299 628106
rect 199510 622965 217854 623965
rect 35872 615141 171201 617459
rect 35872 614141 210863 615141
rect 35872 612005 171201 614141
rect 209863 588028 210863 614141
rect 216854 588501 217854 622965
rect 231299 588737 232299 627106
rect 238371 587555 239371 639529
rect 287552 633507 288552 646060
rect 248373 632507 288552 633507
rect 248373 588028 249373 632507
rect 310957 628466 311957 646060
rect 259248 627466 311957 628466
rect 259248 587083 260248 627466
rect 344265 622344 345265 646060
rect 267558 621344 345265 622344
rect 267558 587733 268558 621344
rect 530161 618189 535929 659959
rect 570812 639592 570818 644694
rect 575920 644684 580012 644694
rect 575920 644584 583353 644684
rect 575920 639784 584800 644584
rect 575920 639592 583353 639784
rect 578927 639578 583353 639592
rect 579387 634674 583813 634748
rect 570867 629638 570873 634674
rect 575909 634584 583813 634674
rect 575909 629784 584800 634584
rect 575909 629642 583813 629784
rect 575909 629638 580012 629642
rect 356710 616223 535929 618189
rect 276898 615223 535929 616223
rect 276898 587124 277898 615223
rect 356710 612421 535929 615223
rect 286354 602558 487607 603558
rect 488607 602558 488613 603558
rect 286354 587425 287354 602558
rect 288354 596090 482433 597090
rect 483433 596090 483439 597090
rect 288354 587536 289354 596090
rect 290346 589077 477776 590077
rect 478776 589077 478782 590077
rect 565585 589584 565697 589590
rect 565697 589472 584800 589584
rect 565585 589466 565697 589472
rect 290346 589012 291354 589077
rect 290346 586827 291346 589012
rect 577012 588290 584800 588402
rect 510491 587292 576060 587293
rect 510486 586294 510492 587292
rect 511490 586958 576060 587292
rect 577012 586958 577124 588290
rect 583473 587108 584800 587220
rect 511490 586846 577124 586958
rect 511490 586294 576060 586846
rect 510491 586293 576060 586294
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 156592 580061 158820 580222
rect 156592 578063 156708 580061
rect 158706 578063 158820 580061
rect 156592 576250 158820 578063
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 145434 525406 171100 576250
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 425730 535389 425794 535395
rect 402219 535327 425730 535387
rect 425730 535319 425794 535325
rect 423449 532949 423513 532955
rect 402264 532887 423449 532947
rect 423449 532879 423513 532885
rect 355561 532597 356561 532603
rect 338673 531597 355561 532597
rect 356561 531597 366475 532597
rect 355561 531591 356561 531597
rect 365475 522025 366475 531597
rect 421586 530387 421650 530393
rect 402219 530325 421586 530385
rect 421586 530317 421650 530323
rect 419511 527947 419575 527953
rect 402230 527885 419511 527945
rect 419511 527877 419575 527883
rect 417539 525383 417545 525385
rect 402078 525323 417545 525383
rect 417539 525321 417545 525323
rect 417609 525321 417615 525385
rect 415539 522943 415545 522945
rect 401983 522883 415545 522943
rect 415539 522881 415545 522883
rect 415609 522881 415615 522945
rect 365475 522007 368109 522025
rect 365475 521479 372498 522007
rect 365475 521419 373965 521479
rect 365475 521025 372498 521419
rect 367231 521007 372498 521025
rect 413516 520383 413580 520389
rect 401504 520321 413516 520381
rect 413516 520313 413580 520319
rect 510491 519692 511491 519698
rect 424147 519108 510491 519692
rect 424147 519048 424601 519108
rect 424661 519048 510491 519108
rect 424147 518692 510491 519048
rect 510491 518686 511491 518692
rect 411487 517943 411551 517949
rect 402002 517881 411487 517941
rect 411487 517873 411551 517879
rect 365528 517349 366528 517355
rect 366528 516928 372498 517349
rect 366528 516868 372209 516928
rect 372269 516868 372498 516928
rect 366528 516349 372498 516868
rect 365528 516343 366528 516349
rect 409483 515381 409547 515387
rect 402220 515319 409483 515379
rect 409483 515311 409547 515317
rect 407542 512941 407606 512947
rect 402309 512879 407542 512939
rect 407542 512871 407606 512877
rect -800 511530 480 511642
rect -800 510348 480 510460
rect 405502 510379 405566 510385
rect 401843 510317 405502 510377
rect 405502 510309 405566 510315
rect -800 509166 480 509278
rect 83456 509247 84454 509252
rect 13939 509246 84455 509247
rect 12230 508887 12340 508892
rect 13939 508887 83456 509246
rect 12229 508886 83456 508887
rect 12229 508776 12230 508886
rect 12340 508776 83456 508886
rect 12229 508775 83456 508776
rect 12230 508770 12340 508775
rect 13939 508248 83456 508775
rect 84454 508248 84455 509246
rect 13939 508247 84455 508248
rect 83456 508242 84454 508247
rect -800 507984 480 508096
rect 403541 507817 403605 507823
rect 387908 507753 387914 507817
rect 387978 507815 387984 507817
rect 387978 507755 388477 507815
rect 402339 507755 403541 507815
rect 387978 507753 387984 507755
rect 403541 507747 403605 507753
rect 12229 506914 12341 506920
rect -800 506802 12229 506914
rect 12229 506796 12341 506802
rect -800 505620 25370 505732
rect 25482 505620 25488 505732
rect 373560 504707 373808 504793
rect 373560 504637 373642 504707
rect 373712 504637 373808 504707
rect 383174 504762 383339 504801
rect 383174 504757 383216 504762
rect 383174 504697 383215 504757
rect 383174 504692 383216 504697
rect 383280 504692 383339 504762
rect 383174 504647 383339 504692
rect 373560 504536 373808 504637
rect 387425 504447 388425 504968
rect 392669 504721 392960 504847
rect 392669 504716 392784 504721
rect 392669 504656 392783 504716
rect 392669 504651 392784 504656
rect 392848 504651 392960 504721
rect 392669 504545 392960 504651
rect 559955 500162 560067 500168
rect 559949 500052 559955 500162
rect 560067 500050 584800 500162
rect 559955 500044 560067 500050
rect 583520 498868 584800 498980
rect 549985 498323 578145 498324
rect 549980 497325 549986 498323
rect 550984 497798 578145 498323
rect 550984 497686 584800 497798
rect 550984 497325 578145 497686
rect 549985 497324 578145 497325
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 549985 480109 550985 480115
rect 382734 480108 549985 480109
rect 382729 479110 382735 480108
rect 383733 479110 549985 480108
rect 382734 479109 549985 479110
rect 549985 479103 550985 479109
rect 373156 476016 374154 476021
rect 373155 476015 549890 476016
rect 373155 475017 373156 476015
rect 374154 475017 549890 476015
rect 373155 475016 549890 475017
rect 550890 475016 550896 476016
rect 373156 475011 374154 475016
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect 78270 465202 79268 465207
rect 15018 465201 79269 465202
rect -800 464762 480 464874
rect 15018 464769 78270 465201
rect 13362 464768 78270 464769
rect 13357 464658 13363 464768
rect 13473 464658 78270 464768
rect 13362 464657 78270 464658
rect 15018 464203 78270 464657
rect 79268 464203 79269 465201
rect 15018 464202 79269 464203
rect 78270 464197 79268 464202
rect 13362 463692 13474 463698
rect -800 463580 13362 463692
rect 13362 463574 13474 463580
rect 25407 462510 25519 462516
rect -800 462398 25407 462510
rect 25407 462392 25519 462398
rect 240180 457761 241180 459480
rect 240180 456755 241180 456761
rect 250981 457761 251981 459175
rect 250981 456755 251981 456761
rect 560008 455740 560120 455746
rect 560120 455628 584800 455740
rect 560008 455622 560120 455628
rect 583520 454446 584800 454558
rect 549890 453859 578427 453860
rect 549885 452861 549891 453859
rect 550889 453376 578427 453859
rect 550889 453264 584800 453376
rect 550889 452861 578427 453264
rect 549890 452860 578427 452861
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 392312 426639 393310 426644
rect 243838 426633 324048 426639
rect 240180 426632 324048 426633
rect 240175 425634 240181 426632
rect 241179 425639 324048 426632
rect 325048 426638 393311 426639
rect 325048 425640 392312 426638
rect 393310 425640 393311 426638
rect 325048 425639 393311 425640
rect 241179 425634 245025 425639
rect 392312 425634 393310 425639
rect 240180 425633 245025 425634
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 250982 421100 251980 421105
rect 336048 421100 337048 421106
rect 250981 421099 336048 421100
rect 72633 420888 73631 420893
rect 15289 420887 73632 420888
rect 15289 420470 72633 420887
rect -800 420358 72633 420470
rect 15289 419889 72633 420358
rect 73631 419889 73632 420887
rect 250981 420101 250982 421099
rect 251980 420101 336048 421099
rect 250981 420100 336048 420101
rect 337048 420100 387407 421100
rect 388407 420100 388413 421100
rect 250982 420095 251980 420100
rect 336048 420094 337048 420100
rect 15289 419888 73632 419889
rect 72633 419883 73631 419888
rect 25438 419288 25550 419294
rect -800 419176 25438 419288
rect 25438 419170 25550 419176
rect 560017 411318 560129 411324
rect 560129 411206 584800 411318
rect 560017 411200 560129 411206
rect 583520 410024 584800 410136
rect 549018 409466 550016 409471
rect 549017 409465 579376 409466
rect 549017 408467 549018 409465
rect 550016 408954 579376 409465
rect 550016 408842 584800 408954
rect 550016 408467 579376 408842
rect 549017 408466 579376 408467
rect 549018 408461 550016 408466
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 336049 387271 337047 387276
rect 548986 387271 550037 387302
rect 336048 387270 549017 387271
rect 336048 386272 336049 387270
rect 337047 386272 549017 387270
rect 336048 386271 549017 386272
rect 550017 386271 550037 387271
rect 336049 386266 337047 386271
rect 548986 386232 550037 386271
rect -800 381864 480 381976
rect 324048 381237 548896 381238
rect -800 380682 480 380794
rect 324043 380239 324049 381237
rect 325047 380239 548896 381237
rect 324048 380238 548896 380239
rect 549896 380238 550017 381238
rect -800 379500 480 379612
rect 65787 378990 66785 378995
rect 14217 378989 66786 378990
rect 12758 378524 12868 378529
rect 14217 378524 65787 378989
rect 12757 378523 65787 378524
rect -800 378318 480 378430
rect 12757 378413 12758 378523
rect 12868 378413 65787 378523
rect 12757 378412 65787 378413
rect 12758 378407 12868 378412
rect 14217 377991 65787 378412
rect 66785 377991 66786 378989
rect 14217 377990 66786 377991
rect 65787 377985 66785 377990
rect 12757 377248 12869 377254
rect -800 377136 12757 377248
rect 12757 377130 12869 377136
rect -800 375954 25430 376066
rect 25542 375954 25548 376066
rect 560038 364896 560150 364902
rect 560150 364784 584800 364896
rect 560038 364778 560150 364784
rect 583520 363602 584800 363714
rect 548897 363047 549895 363052
rect 548896 363046 578945 363047
rect 548896 362048 548897 363046
rect 549895 362532 578945 363046
rect 549895 362420 584800 362532
rect 549895 362048 578945 362420
rect 548896 362047 578945 362048
rect 548897 362042 549895 362047
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect 14352 335076 59670 335077
rect 14352 334684 58671 335076
rect 13037 334683 58671 334684
rect 13032 334573 13038 334683
rect 13148 334573 58671 334683
rect 13037 334572 58671 334573
rect 14352 334078 58671 334572
rect 59669 334078 59675 335076
rect 14352 334077 59670 334078
rect 13037 334026 13149 334032
rect -800 333914 13037 334026
rect 13037 333908 13149 333914
rect 25372 332844 25484 332850
rect -800 332732 25372 332844
rect 25484 332734 25490 332844
rect 25372 332726 25484 332732
rect 565606 319674 565718 319680
rect 565718 319562 584800 319674
rect 565606 319556 565718 319562
rect 578500 318380 584800 318492
rect 365529 317851 366527 317856
rect 365528 317850 576625 317851
rect 365528 316852 365529 317850
rect 366527 317496 576625 317850
rect 578500 317496 578612 318380
rect 366527 317384 578612 317496
rect 366527 316852 576625 317384
rect 583520 317198 584800 317310
rect 365528 316851 576625 316852
rect 365529 316846 366527 316851
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 355562 296500 356560 296505
rect 549082 296500 550082 296506
rect 355561 296499 549082 296500
rect -800 295420 480 295532
rect 355561 295501 355562 296499
rect 356560 295501 549082 296499
rect 355561 295500 549082 295501
rect 355562 295495 356560 295500
rect 549082 295494 550082 295500
rect -800 294238 480 294350
rect -800 293056 480 293168
rect 49270 292102 50268 292107
rect 14352 292101 50269 292102
rect -800 291874 480 291986
rect 13045 291699 13155 291704
rect 14352 291699 49270 292101
rect 13044 291698 49270 291699
rect 13044 291588 13045 291698
rect 13155 291588 49270 291698
rect 13044 291587 49270 291588
rect 13045 291582 13155 291587
rect 14352 291103 49270 291587
rect 50268 291103 50269 292101
rect 14352 291102 50269 291103
rect 49270 291097 50268 291102
rect 13044 290804 13156 290810
rect -800 290692 13044 290804
rect 13044 290686 13156 290692
rect 25372 289622 25484 289628
rect -800 289510 25372 289622
rect 25372 289504 25484 289510
rect 565650 275140 565656 275252
rect 565768 275140 584800 275252
rect 549072 274464 550093 274475
rect 549072 274463 580774 274464
rect 549072 273465 549083 274463
rect 550081 274070 580774 274463
rect 550081 273958 584800 274070
rect 550081 273465 580774 273958
rect 549072 273464 580774 273465
rect 549072 273450 550093 273464
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 83449 268390 83455 269390
rect 84455 268390 425035 269390
rect 426035 268390 426041 269390
rect 583520 269230 584800 269342
rect 78269 267390 79269 267396
rect 79269 266390 423042 267390
rect 424042 266390 424048 267390
rect 78269 266384 79269 266390
rect 72626 264390 72632 265390
rect 73632 264390 421075 265390
rect 422075 264390 422081 265390
rect 65786 263390 66786 263396
rect 66786 262390 419082 263390
rect 420082 262390 420088 263390
rect 65786 262384 66786 262390
rect 58670 261390 59670 261396
rect 59670 260390 417049 261390
rect 418049 260390 418055 261390
rect 58670 260384 59670 260390
rect 49263 258390 49269 259390
rect 50269 258390 415074 259390
rect 416074 258390 416080 259390
rect 49269 257390 50269 257396
rect 50269 256390 413046 257390
rect 414046 256390 414052 257390
rect 49269 256384 50269 256390
rect 58938 255390 59938 255396
rect 59938 254390 411018 255390
rect 412018 254390 412024 255390
rect 58938 254384 59938 254390
rect 65894 253390 66894 253396
rect -800 252398 480 252510
rect 66894 252390 409097 253390
rect 410097 252390 410103 253390
rect 65894 252384 66894 252390
rect 72906 251390 73906 251396
rect -800 251216 480 251328
rect 73906 250390 407015 251390
rect 408015 250390 408021 251390
rect 72906 250384 73906 250390
rect -800 250034 480 250146
rect 78414 249390 79414 249396
rect -800 248852 480 248964
rect 79414 248390 405094 249390
rect 406094 248390 406100 249390
rect 78414 248384 79414 248390
rect 14889 248052 50269 248053
rect 14889 247782 49270 248052
rect -800 247670 49270 247782
rect 14889 247054 49270 247670
rect 50268 247054 50274 248052
rect 83668 247390 84668 247396
rect 403025 247390 404061 247405
rect 14889 247053 50269 247054
rect 25415 246600 25527 246606
rect -800 246488 25415 246600
rect 25415 246482 25527 246488
rect 84668 247389 404061 247390
rect 84668 246391 403046 247389
rect 404044 246391 404061 247389
rect 84668 246390 404061 246391
rect 83668 246384 84668 246390
rect 403025 246376 404061 246390
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 570495 191330 570501 196290
rect 575461 196288 580012 196290
rect 575461 196230 583067 196288
rect 575461 191430 584800 196230
rect 575461 191330 583067 191430
rect 578955 191312 583067 191330
rect 570408 181252 570414 186370
rect 575532 186368 580012 186370
rect 575532 186230 583645 186368
rect 575532 181430 584800 186230
rect 575532 181256 583643 181430
rect 575532 181252 580012 181256
rect 990 177688 13066 177860
rect -800 172888 13066 177688
rect 990 172742 13066 172888
rect 18184 172742 18190 177860
rect 808 167688 13374 167862
rect -800 162888 13374 167688
rect 808 162744 13374 162888
rect 18492 162744 18498 167862
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect 58939 120855 59937 120860
rect 14112 120854 59938 120855
rect 14112 120160 58939 120854
rect -800 120048 58939 120160
rect 14112 119856 58939 120048
rect 59937 119856 59938 120854
rect 14112 119855 59938 119856
rect 58939 119850 59937 119855
rect 25403 118978 25515 118984
rect -800 118866 25403 118978
rect 25403 118860 25515 118866
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 14112 79051 66894 79052
rect 12334 78528 12444 78533
rect 14112 78528 65895 79051
rect 12333 78527 65895 78528
rect 12333 78417 12334 78527
rect 12444 78417 65895 78527
rect 12333 78416 65895 78417
rect 12334 78411 12444 78416
rect -800 78008 480 78120
rect 14112 78053 65895 78416
rect 66893 78053 66899 79051
rect 14112 78052 66894 78053
rect 12333 76938 12445 76944
rect -800 76826 12333 76938
rect 12333 76820 12445 76826
rect 25414 75756 25526 75762
rect -800 75644 25414 75756
rect 25414 75638 25526 75644
rect 72894 66137 73915 66152
rect 15445 66136 73915 66137
rect 12619 65629 12729 65634
rect 15445 65629 72907 66136
rect 12618 65628 72907 65629
rect 12618 65518 12619 65628
rect 12729 65518 72907 65628
rect 12618 65517 72907 65518
rect 12619 65512 12729 65517
rect 15445 65138 72907 65517
rect 73905 65138 73915 66136
rect 15445 65137 73915 65138
rect 72894 65128 73915 65137
rect 78386 62396 79436 62431
rect 15445 62395 79436 62396
rect 14459 62017 14569 62022
rect 15445 62017 78415 62395
rect 14458 62016 78415 62017
rect 14458 61906 14459 62016
rect 14569 61906 78415 62016
rect 14458 61905 78415 61906
rect 14459 61900 14569 61905
rect 15445 61397 78415 61905
rect 79413 61397 79436 62395
rect 15445 61396 79436 61397
rect 78386 61367 79436 61396
rect 83660 59107 84676 59115
rect 15445 59106 84676 59107
rect 15445 58593 83669 59106
rect 15445 58483 16146 58593
rect 16256 58483 83669 58593
rect 15445 58108 83669 58483
rect 84667 58108 84676 59106
rect 15445 58107 84676 58108
rect 83660 58099 84676 58107
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 478104 44895 478216 44901
rect 481593 44895 481715 44900
rect 478216 44783 481598 44895
rect 481710 44783 481715 44895
rect 478104 44777 478216 44783
rect 481593 44778 481715 44783
rect 482769 44886 482881 44892
rect 485139 44886 485261 44891
rect 482881 44774 485144 44886
rect 485256 44774 485261 44886
rect 482769 44768 482881 44774
rect 485139 44769 485261 44774
rect 488005 44874 488117 44880
rect 488685 44874 488807 44879
rect 488117 44762 488690 44874
rect 488802 44762 488807 44874
rect 488005 44756 488117 44762
rect 488685 44757 488807 44762
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect 12618 33716 12730 33722
rect -800 33604 12618 33716
rect 12618 33598 12730 33604
rect -800 32422 25408 32534
rect 25520 32422 25526 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 25446 18906 25558 18912
rect 21662 18905 25446 18906
rect 21657 18795 21663 18905
rect 21773 18795 25446 18905
rect 21662 18794 25446 18795
rect 25446 18788 25558 18794
rect 583520 18092 584800 18204
rect 25438 18068 25550 18074
rect 22608 18067 25438 18068
rect 22603 17957 22609 18067
rect 22719 17957 25438 18067
rect 22608 17956 25438 17957
rect 25438 17950 25550 17956
rect 24982 17174 25982 17180
rect 565200 17174 566198 17179
rect -800 16910 480 17022
rect 25982 17173 566199 17174
rect 25982 16830 565200 17173
rect 25982 16785 486326 16830
rect 25982 16673 482780 16785
rect 482892 16718 486326 16785
rect 486438 16753 565200 16830
rect 486438 16718 489872 16753
rect 482892 16673 489872 16718
rect 25982 16641 489872 16673
rect 489984 16641 565200 16753
rect 25982 16175 565200 16641
rect 566198 16175 566199 17173
rect 583520 16910 584800 17022
rect 25982 16174 566199 16175
rect 24982 16168 25982 16174
rect 565200 16169 566198 16174
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect 14458 12294 14570 12300
rect -800 12182 14458 12294
rect 583520 12182 584800 12294
rect 14458 12176 14570 12182
rect 21662 11112 21774 11118
rect -800 11000 21662 11112
rect 583520 11000 584800 11112
rect 21662 10994 21774 11000
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect 16145 7566 16257 7572
rect -800 7454 16145 7566
rect 583520 7454 584800 7566
rect 16145 7448 16257 7454
rect 22608 6384 22720 6390
rect -800 6272 22608 6384
rect 583520 6272 584800 6384
rect 22608 6266 22720 6272
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 8383 643688 13471 648776
rect 8391 633670 13463 638742
rect 570818 639592 575920 644694
rect 570873 629638 575909 634674
rect 487607 602558 488607 603558
rect 482433 596090 483433 597090
rect 477776 589077 478776 590077
rect 565585 589472 565697 589584
rect 510492 586294 511490 587292
rect 156708 578063 158706 580061
rect 425730 535325 425794 535389
rect 423449 532885 423513 532949
rect 355561 531597 356561 532597
rect 421586 530323 421650 530387
rect 419511 527883 419575 527947
rect 417545 525321 417609 525385
rect 415545 522881 415609 522945
rect 413516 520319 413580 520383
rect 510491 518692 511491 519692
rect 411487 517879 411551 517943
rect 365528 516349 366528 517349
rect 409483 515317 409547 515381
rect 407542 512877 407606 512941
rect 405502 510315 405566 510379
rect 12230 508776 12340 508886
rect 83456 508248 84454 509246
rect 387914 507753 387978 507817
rect 403541 507753 403605 507817
rect 12229 506802 12341 506914
rect 25370 505620 25482 505732
rect 373642 504702 373712 504707
rect 373642 504642 373647 504702
rect 373647 504642 373707 504702
rect 373707 504642 373712 504702
rect 373642 504637 373712 504642
rect 383216 504757 383280 504762
rect 383216 504697 383275 504757
rect 383275 504697 383280 504757
rect 383216 504692 383280 504697
rect 392784 504716 392848 504721
rect 392784 504656 392843 504716
rect 392843 504656 392848 504716
rect 392784 504651 392848 504656
rect 559955 500050 560067 500162
rect 549986 497325 550984 498323
rect 382735 479110 383733 480108
rect 549985 479109 550985 480109
rect 373156 475017 374154 476015
rect 549890 475016 550890 476016
rect 13363 464658 13473 464768
rect 78270 464203 79268 465201
rect 13362 463580 13474 463692
rect 25407 462398 25519 462510
rect 240180 456761 241180 457761
rect 250981 456761 251981 457761
rect 560008 455628 560120 455740
rect 549891 452861 550889 453859
rect 240181 425634 241179 426632
rect 324048 425639 325048 426639
rect 392312 425640 393310 426638
rect 72633 419889 73631 420887
rect 250982 420101 251980 421099
rect 336048 420100 337048 421100
rect 387407 420100 388407 421100
rect 25438 419176 25550 419288
rect 560017 411206 560129 411318
rect 549018 408467 550016 409465
rect 336049 386272 337047 387270
rect 549017 386271 550017 387271
rect 324049 380239 325047 381237
rect 548896 380238 549896 381238
rect 12758 378413 12868 378523
rect 65787 377991 66785 378989
rect 12757 377136 12869 377248
rect 25430 375954 25542 376066
rect 560038 364784 560150 364896
rect 548897 362048 549895 363046
rect 13038 334573 13148 334683
rect 58671 334078 59669 335076
rect 13037 333914 13149 334026
rect 25372 332732 25484 332844
rect 565606 319562 565718 319674
rect 365529 316852 366527 317850
rect 355562 295501 356560 296499
rect 549082 295500 550082 296500
rect 13045 291588 13155 291698
rect 49270 291103 50268 292101
rect 13044 290692 13156 290804
rect 25372 289510 25484 289622
rect 565656 275140 565768 275252
rect 549083 273465 550081 274463
rect 83455 268390 84455 269390
rect 425035 268390 426035 269390
rect 78269 266390 79269 267390
rect 423042 266390 424042 267390
rect 72632 264390 73632 265390
rect 421075 264390 422075 265390
rect 65786 262390 66786 263390
rect 419082 262390 420082 263390
rect 58670 260390 59670 261390
rect 417049 260390 418049 261390
rect 49269 258390 50269 259390
rect 415074 258390 416074 259390
rect 49269 256390 50269 257390
rect 413046 256390 414046 257390
rect 58938 254390 59938 255390
rect 411018 254390 412018 255390
rect 65894 252390 66894 253390
rect 409097 252390 410097 253390
rect 72906 250390 73906 251390
rect 407015 250390 408015 251390
rect 78414 248390 79414 249390
rect 405094 248390 406094 249390
rect 49270 247054 50268 248052
rect 25415 246488 25527 246600
rect 83668 246390 84668 247390
rect 403046 246391 404044 247389
rect 570501 191330 575461 196290
rect 570414 181252 575532 186370
rect 13066 172742 18184 177860
rect 13374 162744 18492 167862
rect 58939 119856 59937 120854
rect 25403 118866 25515 118978
rect 12334 78417 12444 78527
rect 65895 78053 66893 79051
rect 12333 76826 12445 76938
rect 25414 75644 25526 75756
rect 12619 65518 12729 65628
rect 72907 65138 73905 66136
rect 14459 61906 14569 62016
rect 78415 61397 79413 62395
rect 16146 58483 16256 58593
rect 83669 58108 84667 59106
rect 478104 44783 478216 44895
rect 482769 44774 482881 44886
rect 488005 44762 488117 44874
rect 12618 33604 12730 33716
rect 25408 32422 25520 32534
rect 21663 18795 21773 18905
rect 25446 18794 25558 18906
rect 22609 17957 22719 18067
rect 25438 17956 25550 18068
rect 24982 16174 25982 17174
rect 565200 16175 566198 17173
rect 14458 12182 14570 12294
rect 21662 11000 21774 11112
rect 16145 7454 16257 7566
rect 22608 6272 22720 6384
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 131021 648752 136109 649974
rect 131021 643712 131219 648752
rect 131021 638718 136109 643712
rect 131021 633694 131043 638718
rect 136067 633694 136109 638718
rect 118328 580341 123446 614371
rect 131021 584235 136109 633694
rect 559614 644687 560614 645250
rect 559614 639595 559620 644687
rect 559614 634721 560614 639595
rect 560609 629629 560614 634721
rect 437075 605496 442175 629601
rect 378807 584076 379427 584275
rect 437075 584137 442163 605496
rect 396631 584080 397251 584136
rect 118328 577835 118354 580341
rect 123274 577835 123446 580341
rect 12229 508886 12341 508887
rect 12229 508776 12230 508886
rect 12340 508776 12341 508886
rect 12229 506915 12341 508776
rect 12228 506914 12342 506915
rect 12228 506802 12229 506914
rect 12341 506802 12342 506914
rect 12228 506801 12342 506802
rect 24982 505732 25982 520014
rect 24982 505620 25370 505732
rect 25482 505620 25982 505732
rect 13362 464768 13474 464769
rect 13362 464658 13363 464768
rect 13473 464658 13474 464768
rect 13362 463693 13474 464658
rect 13361 463692 13475 463693
rect 13361 463580 13362 463692
rect 13474 463580 13475 463692
rect 13361 463579 13475 463580
rect 24982 462510 25982 505620
rect 83455 509246 84455 509247
rect 83455 508248 83456 509246
rect 84454 508248 84455 509246
rect 24982 462398 25407 462510
rect 25519 462398 25982 462510
rect 24982 419288 25982 462398
rect 78269 465201 79269 465202
rect 78269 464203 78270 465201
rect 79268 464203 79269 465201
rect 24982 419176 25438 419288
rect 25550 419176 25982 419288
rect 12757 378523 12869 378524
rect 12757 378413 12758 378523
rect 12868 378413 12869 378523
rect 12757 377249 12869 378413
rect 12756 377248 12870 377249
rect 12756 377136 12757 377248
rect 12869 377136 12870 377248
rect 12756 377135 12870 377136
rect 24982 376066 25982 419176
rect 72632 420887 73632 420888
rect 72632 419889 72633 420887
rect 73631 419889 73632 420887
rect 24982 375954 25430 376066
rect 25542 375954 25982 376066
rect 13037 334683 13149 334684
rect 13037 334573 13038 334683
rect 13148 334573 13149 334683
rect 13037 334027 13149 334573
rect 13036 334026 13150 334027
rect 13036 333914 13037 334026
rect 13149 333914 13150 334026
rect 13036 333913 13150 333914
rect 24982 332844 25982 375954
rect 65786 378989 66786 378990
rect 65786 377991 65787 378989
rect 66785 377991 66786 378989
rect 24982 332732 25372 332844
rect 25484 332732 25982 332844
rect 13044 291698 13156 291699
rect 13044 291588 13045 291698
rect 13155 291588 13156 291698
rect 13044 290805 13156 291588
rect 13043 290804 13157 290805
rect 13043 290692 13044 290804
rect 13156 290692 13157 290804
rect 13043 290691 13157 290692
rect 24982 289622 25982 332732
rect 58670 335076 59670 335345
rect 58670 334078 58671 335076
rect 59669 334078 59670 335076
rect 24982 289510 25372 289622
rect 25484 289510 25982 289622
rect 24982 246600 25982 289510
rect 49269 292101 50269 292102
rect 49269 291103 49270 292101
rect 50268 291103 50269 292101
rect 49269 259391 50269 291103
rect 58670 261391 59670 334078
rect 65786 263391 66786 377991
rect 72632 265391 73632 419889
rect 78269 267391 79269 464203
rect 83455 269391 84455 508248
rect 118328 467391 123446 577835
rect 131021 548284 136109 581875
rect 156666 580061 158779 580122
rect 156666 578063 156708 580061
rect 158706 578063 158779 580061
rect 156666 577968 158779 578063
rect 131021 543196 148197 548284
rect 83454 269390 84456 269391
rect 83454 268390 83455 269390
rect 84455 268390 84456 269390
rect 83454 268389 84456 268390
rect 78268 267390 79270 267391
rect 78268 266390 78269 267390
rect 79269 266390 79270 267390
rect 78268 266389 79270 266390
rect 72631 265390 73633 265391
rect 72631 264390 72632 265390
rect 73632 264390 73633 265390
rect 72631 264389 73633 264390
rect 65785 263390 66787 263391
rect 65785 262390 65786 263390
rect 66786 262390 66787 263390
rect 65785 262389 66787 262390
rect 58669 261390 59671 261391
rect 58669 260390 58670 261390
rect 59670 260390 59671 261390
rect 58669 260389 59671 260390
rect 49268 259390 50270 259391
rect 49268 258390 49269 259390
rect 50269 258390 50270 259390
rect 49268 258389 50270 258390
rect 49268 257390 50270 257391
rect 49268 256390 49269 257390
rect 50269 256390 50270 257390
rect 49268 256389 50270 256390
rect 49269 248052 50269 256389
rect 58937 255390 59939 255391
rect 58937 254390 58938 255390
rect 59938 254390 59939 255390
rect 58937 254389 59939 254390
rect 49269 247054 49270 248052
rect 50268 247054 50269 248052
rect 49269 247053 50269 247054
rect 24982 246488 25415 246600
rect 25527 246488 25982 246600
rect 24982 177806 25982 246488
rect 24982 167760 25982 172855
rect 24982 162809 25000 167760
rect 24982 118978 25982 162809
rect 58938 120854 59938 254389
rect 65893 253390 66895 253391
rect 65893 252390 65894 253390
rect 66894 252390 66895 253390
rect 65893 252389 66895 252390
rect 58938 119856 58939 120854
rect 59937 119856 59938 120854
rect 58938 119855 59938 119856
rect 24982 118866 25403 118978
rect 25515 118866 25982 118978
rect 12333 78527 12445 78528
rect 12333 78417 12334 78527
rect 12444 78417 12445 78527
rect 12333 76939 12445 78417
rect 12332 76938 12446 76939
rect 12332 76826 12333 76938
rect 12445 76826 12446 76938
rect 12332 76825 12446 76826
rect 24982 75756 25982 118866
rect 65894 79051 66894 252389
rect 72905 251390 73907 251391
rect 72905 250390 72906 251390
rect 73906 250390 73907 251390
rect 72905 250389 73907 250390
rect 65894 78053 65895 79051
rect 66893 78053 66894 79051
rect 65894 78052 66894 78053
rect 24982 75644 25414 75756
rect 25526 75644 25982 75756
rect 12618 65628 12730 65629
rect 12618 65518 12619 65628
rect 12729 65518 12730 65628
rect 12618 33717 12730 65518
rect 14458 62016 14570 62017
rect 14458 61906 14459 62016
rect 14569 61906 14570 62016
rect 12617 33716 12731 33717
rect 12617 33604 12618 33716
rect 12730 33604 12731 33716
rect 12617 33603 12731 33604
rect 14458 12295 14570 61906
rect 16145 58593 16257 58594
rect 16145 58483 16146 58593
rect 16256 58483 16257 58593
rect 14457 12294 14571 12295
rect 14457 12182 14458 12294
rect 14570 12182 14571 12294
rect 14457 12181 14571 12182
rect 16145 7567 16257 58483
rect 24982 32534 25982 75644
rect 72906 66152 73906 250389
rect 78413 249390 79415 249391
rect 78413 248390 78414 249390
rect 79414 248390 79415 249390
rect 78413 248389 79415 248390
rect 72894 66136 73915 66152
rect 72894 65138 72907 66136
rect 73905 65138 73915 66136
rect 72894 65128 73915 65138
rect 72906 65038 73906 65128
rect 78414 62431 79414 248389
rect 83667 247390 84669 247391
rect 83667 246390 83668 247390
rect 84668 246390 84669 247390
rect 83667 246389 84669 246390
rect 78386 62395 79436 62431
rect 78386 61397 78415 62395
rect 79413 61397 79436 62395
rect 78386 61367 79436 61397
rect 78414 61319 79414 61367
rect 83668 59115 84668 246389
rect 118328 177836 123446 465128
rect 131021 463295 136109 543196
rect 377567 534554 378187 578103
rect 378807 534486 379427 582061
rect 396631 534614 397251 582065
rect 397871 580068 398491 580202
rect 437075 578606 442163 581960
rect 449668 580116 454786 612029
rect 487606 603558 488608 603559
rect 487606 602558 487607 603558
rect 488607 602558 488608 603558
rect 487606 602557 488608 602558
rect 482432 597090 483434 597091
rect 482432 596090 482433 597090
rect 483433 596090 483434 597090
rect 482432 596089 483434 596090
rect 477775 590077 478777 590078
rect 477775 589077 477776 590077
rect 478776 589077 478777 590077
rect 477775 589076 478777 589077
rect 397871 534943 398491 578053
rect 425729 535389 425795 535390
rect 425729 535325 425730 535389
rect 425794 535325 425795 535389
rect 425729 535324 425795 535325
rect 425732 533985 425792 535324
rect 423448 532949 423514 532950
rect 423448 532885 423449 532949
rect 423513 532885 423514 532949
rect 423448 532884 423514 532885
rect 355560 532597 356562 532598
rect 355560 531597 355561 532597
rect 356561 531597 356562 532597
rect 355560 531596 356562 531597
rect 136035 461032 136109 463295
rect 131021 201242 136109 461032
rect 240179 457761 241181 457762
rect 240179 456761 240180 457761
rect 241180 456761 241181 457761
rect 240179 456760 241181 456761
rect 250980 457761 251982 457762
rect 250980 456761 250981 457761
rect 251981 456761 251982 457761
rect 250980 456760 251982 456761
rect 240180 426632 241180 456760
rect 240180 425634 240181 426632
rect 241179 425634 241180 426632
rect 240180 425633 241180 425634
rect 250981 421099 251981 456760
rect 324047 426639 325049 426640
rect 324047 425639 324048 426639
rect 325048 425639 325049 426639
rect 324047 425638 325049 425639
rect 250981 420101 250982 421099
rect 251980 420101 251981 421099
rect 250981 420100 251981 420101
rect 324048 381237 325048 425638
rect 336047 421100 337049 421101
rect 336047 420100 336048 421100
rect 337048 420100 337049 421100
rect 336047 420099 337049 420100
rect 336048 387270 337048 420099
rect 336048 386272 336049 387270
rect 337047 386272 337048 387270
rect 336048 386271 337048 386272
rect 324048 380239 324049 381237
rect 325047 380239 325048 381237
rect 324048 380238 325048 380239
rect 355561 296499 356561 531596
rect 423451 531548 423511 532884
rect 421585 530387 421651 530388
rect 421585 530323 421586 530387
rect 421650 530323 421651 530387
rect 421585 530322 421651 530323
rect 421588 528704 421648 530322
rect 419510 527947 419576 527948
rect 419510 527883 419511 527947
rect 419575 527883 419576 527947
rect 419510 527882 419576 527883
rect 419513 526413 419573 527882
rect 417544 525385 417610 525386
rect 417544 525321 417545 525385
rect 417609 525321 417610 525385
rect 417544 525320 417610 525321
rect 417547 523744 417607 525320
rect 415544 522945 415610 522946
rect 415544 522881 415545 522945
rect 415609 522881 415610 522945
rect 415544 522880 415610 522881
rect 415547 521278 415607 522880
rect 413515 520383 413581 520384
rect 413515 520319 413516 520383
rect 413580 520319 413581 520383
rect 413515 520318 413581 520319
rect 413518 518914 413578 520318
rect 411486 517943 411552 517944
rect 411486 517879 411487 517943
rect 411551 517879 411552 517943
rect 411486 517878 411552 517879
rect 365527 517349 366529 517350
rect 365527 516349 365528 517349
rect 366528 516349 366529 517349
rect 365527 516348 366529 516349
rect 365528 317850 366528 516348
rect 411489 516312 411549 517878
rect 409482 515381 409548 515382
rect 409482 515317 409483 515381
rect 409547 515317 409548 515381
rect 409482 515316 409548 515317
rect 409485 513846 409545 515316
rect 407541 512941 407607 512942
rect 407541 512877 407542 512941
rect 407606 512877 407607 512941
rect 407541 512876 407607 512877
rect 407544 511313 407604 512876
rect 405501 510379 405567 510380
rect 405501 510315 405502 510379
rect 405566 510315 405567 510379
rect 405501 510314 405567 510315
rect 405504 508779 405564 510314
rect 373152 504829 374155 504968
rect 373155 504707 374155 504829
rect 373155 504637 373642 504707
rect 373712 504637 374155 504707
rect 373155 476015 374155 504637
rect 373155 475017 373156 476015
rect 374154 475017 374155 476015
rect 373155 475016 374155 475017
rect 377567 467291 378187 508101
rect 377567 465237 378187 465285
rect 378807 463289 379427 508379
rect 387913 507817 387979 507818
rect 387913 507753 387914 507817
rect 387978 507753 387979 507817
rect 387913 507752 387979 507753
rect 382734 504762 383734 505017
rect 387916 504968 387976 507752
rect 382734 504692 383216 504762
rect 383280 504692 383734 504762
rect 382734 480108 383734 504692
rect 387425 486995 388425 504968
rect 392312 504721 393312 504968
rect 392312 504651 392784 504721
rect 392848 504651 393312 504721
rect 392312 504631 393312 504651
rect 382734 479110 382735 480108
rect 383733 479110 383734 480108
rect 382734 479109 383734 479110
rect 387407 485497 388425 486995
rect 392311 504474 393312 504631
rect 387407 421101 388407 485497
rect 392311 426638 393311 504474
rect 396631 463277 397251 507704
rect 397871 467290 398491 507962
rect 403540 507817 403606 507818
rect 403540 507753 403541 507817
rect 403605 507753 403606 507817
rect 403540 507752 403606 507753
rect 403543 506068 403603 507752
rect 392311 425640 392312 426638
rect 393310 425640 393311 426638
rect 392311 425639 393311 425640
rect 387406 421100 388408 421101
rect 387406 420100 387407 421100
rect 388407 420100 388408 421100
rect 387406 420099 388408 420100
rect 365528 316852 365529 317850
rect 366527 316852 366528 317850
rect 365528 316851 366528 316852
rect 355561 295501 355562 296499
rect 356560 295501 356561 296499
rect 355561 295500 356561 295501
rect 403045 247405 404045 506068
rect 405045 249391 406045 508779
rect 407045 251391 408045 511313
rect 409045 253391 410045 513846
rect 411045 255391 412045 516312
rect 413045 257391 414045 518914
rect 415045 259391 416045 521278
rect 417045 261391 418045 523744
rect 419045 263391 420045 526413
rect 421045 265391 422045 528704
rect 423045 267391 424045 531548
rect 425045 269391 426045 533985
rect 437075 530351 442175 578606
rect 442149 529681 442175 530351
rect 437075 513406 442175 529681
rect 449668 531568 454786 577998
rect 449668 530898 449712 531568
rect 437075 512736 437103 513406
rect 437075 463376 442175 512736
rect 449668 512175 454786 530898
rect 449668 511505 449671 512175
rect 454772 511505 454786 512175
rect 449668 467421 454786 511505
rect 449668 465158 449674 467421
rect 425034 269390 426045 269391
rect 425034 268390 425035 269390
rect 426035 268390 426045 269390
rect 425034 268389 426045 268390
rect 425045 268228 426045 268389
rect 423041 267390 424045 267391
rect 423041 266390 423042 267390
rect 424042 266390 424045 267390
rect 423041 266389 424045 266390
rect 423045 266279 424045 266389
rect 421045 265390 422076 265391
rect 421045 264390 421075 265390
rect 422075 264390 422076 265390
rect 421045 264389 422076 264390
rect 421045 264274 422045 264389
rect 419045 263390 420083 263391
rect 419045 262390 419082 263390
rect 420082 262390 420083 263390
rect 419045 262389 420083 262390
rect 419045 262214 420045 262389
rect 417045 261390 418050 261391
rect 417045 260390 417049 261390
rect 418049 260390 418050 261390
rect 417045 260389 418050 260390
rect 417045 260265 418045 260389
rect 415045 259390 416075 259391
rect 415045 258390 415074 259390
rect 416074 258390 416075 259390
rect 415045 258389 416075 258390
rect 415045 258205 416045 258389
rect 413045 257390 414047 257391
rect 413045 256390 413046 257390
rect 414046 256390 414047 257390
rect 413045 256389 414047 256390
rect 413045 256256 414045 256389
rect 411017 255390 412045 255391
rect 411017 254390 411018 255390
rect 412018 254390 412045 255390
rect 411017 254389 412045 254390
rect 411045 254252 412045 254389
rect 409045 253390 410098 253391
rect 409045 252390 409097 253390
rect 410097 252390 410098 253390
rect 409045 252389 410098 252390
rect 409045 252247 410045 252389
rect 407014 251390 408045 251391
rect 407014 250390 407015 251390
rect 408015 250390 408045 251390
rect 407014 250389 408045 250390
rect 407045 250197 408045 250389
rect 405045 249390 406095 249391
rect 405045 248390 405094 249390
rect 406094 248390 406095 249390
rect 405045 248389 406095 248390
rect 405045 248355 406045 248389
rect 403025 247389 404061 247405
rect 403025 246391 403046 247389
rect 404044 246391 404061 247389
rect 403025 246376 404061 246391
rect 437075 195272 442175 461113
rect 449668 196266 454786 465158
rect 454435 191354 454786 196266
rect 449668 186346 454786 191354
rect 454514 181276 454786 186346
rect 123398 172766 123446 177836
rect 118328 167838 123446 172766
rect 123264 162768 123446 167838
rect 449668 177836 454786 181276
rect 449668 172766 449876 177836
rect 449668 167838 454786 172766
rect 449668 162995 449738 167838
rect 118328 160061 123446 162768
rect 83660 59106 84676 59115
rect 83660 58108 83669 59106
rect 84667 58108 84676 59106
rect 83660 58099 84676 58108
rect 477776 54057 478776 589076
rect 482433 54057 483433 596089
rect 487607 54057 488607 602557
rect 510491 587292 511491 587293
rect 510491 586294 510492 587292
rect 511490 586294 511491 587292
rect 510491 519693 511491 586294
rect 510490 519692 511492 519693
rect 510490 518692 510491 519692
rect 511491 518692 511492 519692
rect 510490 518691 511492 518692
rect 559614 500162 560614 629629
rect 559614 500050 559955 500162
rect 560067 500050 560614 500162
rect 549985 498323 550985 498324
rect 549985 497325 549986 498323
rect 550984 497325 550985 498323
rect 549985 480110 550985 497325
rect 549984 480109 550986 480110
rect 549984 479109 549985 480109
rect 550985 479109 550986 480109
rect 549984 479108 550986 479109
rect 549889 476016 550891 476017
rect 549889 475016 549890 476016
rect 550890 475016 550891 476016
rect 549889 475015 550891 475016
rect 549890 453859 550890 475015
rect 549890 452861 549891 453859
rect 550889 452861 550890 453859
rect 549890 452860 550890 452861
rect 559614 455740 560614 500050
rect 559614 455628 560008 455740
rect 560120 455628 560614 455740
rect 559614 411318 560614 455628
rect 559614 411206 560017 411318
rect 560129 411206 560614 411318
rect 549017 409465 550017 409466
rect 549017 408467 549018 409465
rect 550016 408467 550017 409465
rect 549017 387302 550017 408467
rect 548986 387271 550037 387302
rect 548986 386271 549017 387271
rect 550017 386271 550037 387271
rect 548986 386232 550037 386271
rect 548895 381238 549897 381239
rect 548895 380238 548896 381238
rect 549896 380238 549897 381238
rect 548895 380237 549897 380238
rect 548896 363046 549896 380237
rect 548896 362048 548897 363046
rect 549895 362048 549896 363046
rect 548896 362047 549896 362048
rect 559614 364896 560614 411206
rect 559614 364784 560038 364896
rect 560150 364784 560614 364896
rect 559614 352599 560614 364784
rect 565199 589584 566199 604185
rect 565199 589472 565585 589584
rect 565697 589472 566199 589584
rect 565199 319674 566199 589472
rect 565199 319562 565606 319674
rect 565718 319562 566199 319674
rect 549081 296500 550083 296501
rect 549081 295500 549082 296500
rect 550082 295500 550083 296500
rect 549081 295499 550083 295500
rect 549082 274475 550082 295499
rect 565199 275252 566199 319562
rect 565199 275140 565656 275252
rect 565768 275140 566199 275252
rect 549072 274463 550093 274475
rect 549072 273465 549083 274463
rect 550081 273465 550093 274463
rect 549072 273450 550093 273465
rect 549082 273312 550082 273450
rect 565199 196299 566199 275140
rect 566194 191348 566199 196299
rect 565199 186266 566199 191348
rect 575460 196290 575462 196291
rect 575461 191330 575462 196290
rect 575460 191329 575462 191330
rect 565199 181315 565206 186266
rect 478104 44896 478216 54057
rect 478103 44895 478217 44896
rect 478103 44783 478104 44895
rect 478216 44783 478217 44895
rect 482769 44887 482881 54057
rect 478103 44782 478217 44783
rect 482768 44886 482882 44887
rect 482768 44774 482769 44886
rect 482881 44774 482882 44886
rect 488005 44875 488117 54057
rect 482768 44773 482882 44774
rect 488004 44874 488118 44875
rect 488004 44762 488005 44874
rect 488117 44762 488118 44874
rect 488004 44761 488118 44762
rect 24982 32422 25408 32534
rect 25520 32422 25982 32534
rect 24982 18906 25982 32422
rect 21662 18905 21774 18906
rect 21662 18795 21663 18905
rect 21773 18795 21774 18905
rect 21662 11113 21774 18795
rect 24982 18794 25446 18906
rect 25558 18794 25982 18906
rect 24982 18068 25982 18794
rect 22608 18067 22720 18068
rect 22608 17957 22609 18067
rect 22719 17957 22720 18067
rect 21661 11112 21775 11113
rect 21661 11000 21662 11112
rect 21774 11000 21775 11112
rect 21661 10999 21775 11000
rect 16144 7566 16258 7567
rect 16144 7454 16145 7566
rect 16257 7454 16258 7566
rect 16144 7453 16258 7454
rect 22608 6385 22720 17957
rect 24982 17956 25438 18068
rect 25550 17956 25982 18068
rect 24982 17175 25982 17956
rect 24981 17174 25983 17175
rect 24981 16174 24982 17174
rect 25982 16174 25983 17174
rect 565199 17173 566199 181315
rect 565199 16175 565200 17173
rect 566198 16175 566199 17173
rect 565199 16174 566199 16175
rect 24981 16173 25983 16174
rect 22607 6384 22721 6385
rect 22607 6272 22608 6384
rect 22720 6272 22721 6384
rect 22607 6271 22721 6272
<< via4 >>
rect 8382 648776 13472 648777
rect 8382 643688 8383 648776
rect 8383 643688 13471 648776
rect 13471 643688 13472 648776
rect 8382 643687 13472 643688
rect 131219 643712 136259 648752
rect 8390 638742 13464 638743
rect 8390 633670 8391 638742
rect 8391 633670 13463 638742
rect 13463 633670 13464 638742
rect 8390 633669 13464 633670
rect 131043 633694 136067 638718
rect 437023 629601 442234 648802
rect 570817 644694 575921 644695
rect 559620 639595 560618 644687
rect 570817 639592 570818 644694
rect 570818 639592 575920 644694
rect 575920 639592 575921 644694
rect 570817 639591 575921 639592
rect 559611 629629 560609 634721
rect 570872 634674 575910 634675
rect 570872 629638 570873 634674
rect 570873 629638 575909 634674
rect 575909 629638 575910 634674
rect 570872 629637 575910 629638
rect 130984 581875 136121 584235
rect 378792 582061 379469 584076
rect 396584 582065 397261 584080
rect 118354 577835 123274 580341
rect 156731 578086 158683 580038
rect 377445 578103 378296 580049
rect 118302 465128 123454 467391
rect 13065 177860 18185 177861
rect 13065 172742 13066 177860
rect 13066 172742 18184 177860
rect 18184 172742 18185 177860
rect 24981 172855 25988 177806
rect 13065 172741 18185 172742
rect 13373 167862 18493 167863
rect 13373 162744 13374 167862
rect 13374 162744 18492 167862
rect 18492 162744 18493 167862
rect 13373 162743 18493 162744
rect 25000 162809 26007 167760
rect 437037 581960 442172 584137
rect 397858 578053 398535 580068
rect 130883 461032 136035 463295
rect 377512 465285 378229 467291
rect 378782 461283 379499 463289
rect 397854 465284 398571 467290
rect 396581 461271 397298 463277
rect 449647 577998 454787 580116
rect 437048 529681 442149 530351
rect 449712 530898 454813 531568
rect 437103 512736 442204 513406
rect 449671 511505 454772 512175
rect 449674 465158 454826 467421
rect 437058 461113 442210 463376
rect 449523 191354 454435 196266
rect 449444 181276 454514 186346
rect 118328 172766 123398 177836
rect 118194 162768 123264 167838
rect 449876 172766 454946 177836
rect 449738 162768 454808 167838
rect 565187 191348 566194 196299
rect 570500 196290 575460 196291
rect 570500 191330 570501 196290
rect 570501 191330 575460 196290
rect 570500 191329 575460 191330
rect 570413 186370 575533 186371
rect 565206 181315 566213 186266
rect 570413 181252 570414 186370
rect 570414 181252 575532 186370
rect 575532 181252 575533 186370
rect 570413 181251 575533 181252
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 436999 648802 442258 648826
rect 8358 648777 13496 648801
rect 8358 643687 8382 648777
rect 13472 648776 13496 648777
rect 436999 648776 437023 648802
rect 13472 648752 437023 648776
rect 13472 643712 131219 648752
rect 136259 643712 437023 648752
rect 13472 643688 437023 643712
rect 13472 643687 13496 643688
rect 8358 643663 13496 643687
rect 8366 638743 13488 638767
rect 8366 633669 8390 638743
rect 13464 638742 13488 638743
rect 436999 638742 437023 643688
rect 13464 638718 437023 638742
rect 13464 633694 131043 638718
rect 136067 633694 437023 638718
rect 13464 633670 437023 633694
rect 13464 633669 13488 633670
rect 8366 633645 13488 633669
rect 436999 629601 437023 633670
rect 442234 644694 442258 648802
rect 559596 644694 560642 644711
rect 570793 644695 575945 644719
rect 570793 644694 570817 644695
rect 442234 644687 570817 644694
rect 442234 639595 559620 644687
rect 560618 639595 570817 644687
rect 442234 639592 570817 639595
rect 442234 634674 442258 639592
rect 559596 639571 560642 639592
rect 570793 639591 570817 639592
rect 575921 639591 575945 644695
rect 570793 639567 575945 639591
rect 559587 634721 560633 634745
rect 559587 634674 559611 634721
rect 442234 629638 559611 634674
rect 442234 629601 442258 629638
rect 559587 629629 559611 629638
rect 560609 634674 560633 634721
rect 570848 634675 575934 634699
rect 570848 634674 570872 634675
rect 560609 629638 570872 634674
rect 560609 629629 560633 629638
rect 559587 629605 560633 629629
rect 570848 629637 570872 629638
rect 575910 629637 575934 634675
rect 570848 629613 575934 629637
rect 436999 629577 442258 629601
rect 130960 584235 136145 584259
rect 130960 581875 130984 584235
rect 136121 584062 136145 584235
rect 437013 584137 442196 584161
rect 378768 584076 379493 584100
rect 378768 584062 378792 584076
rect 136121 582062 181559 584062
rect 338673 582062 378792 584062
rect 136121 581875 136145 582062
rect 378768 582061 378792 582062
rect 379469 584062 379493 584076
rect 396560 584080 397285 584104
rect 396560 584062 396584 584080
rect 379469 582065 396584 584062
rect 397261 584062 397285 584080
rect 437013 584062 437037 584137
rect 397261 582065 437037 584062
rect 379469 582062 437037 582065
rect 379469 582061 379493 582062
rect 378768 582037 379493 582061
rect 396560 582041 397285 582062
rect 437013 581960 437037 582062
rect 442172 581960 442196 584137
rect 437013 581936 442196 581960
rect 130960 581851 136145 581875
rect 118330 580341 123298 580365
rect 118330 577835 118354 580341
rect 123274 580062 123298 580341
rect 449623 580116 454811 580140
rect 377421 580062 378320 580073
rect 397834 580068 398559 580092
rect 397834 580062 397858 580068
rect 123274 580038 179747 580062
rect 123274 578086 156731 580038
rect 158683 578086 179747 580038
rect 123274 578062 179747 578086
rect 338673 580049 397858 580062
rect 338673 578103 377445 580049
rect 378296 578103 397858 580049
rect 338673 578062 397858 578103
rect 123274 577835 123298 578062
rect 397834 578053 397858 578062
rect 398535 580062 398559 580068
rect 449623 580062 449647 580116
rect 398535 578062 449647 580062
rect 398535 578053 398559 578062
rect 397834 578029 398559 578053
rect 449623 577998 449647 578062
rect 454787 580062 454811 580116
rect 454787 578062 454847 580062
rect 454787 577998 454811 578062
rect 449623 577974 454811 577998
rect 118330 577811 123298 577835
rect 449688 531568 454837 531592
rect 449688 531548 449712 531568
rect 401948 530928 449712 531548
rect 449688 530898 449712 530928
rect 454813 530898 454837 531568
rect 449688 530874 454837 530898
rect 437024 530351 442173 530375
rect 437024 530308 437048 530351
rect 401922 529688 437048 530308
rect 437024 529681 437048 529688
rect 442149 529681 442173 530351
rect 437024 529657 442173 529681
rect 437079 513406 442228 513430
rect 437079 513368 437103 513406
rect 402069 512748 437103 513368
rect 437079 512736 437103 512748
rect 442204 512736 442228 513406
rect 437079 512712 442228 512736
rect 449647 512175 454796 512199
rect 449647 512128 449671 512175
rect 401970 511508 449671 512128
rect 449647 511505 449671 511508
rect 454772 511505 454796 512175
rect 449647 511481 454796 511505
rect 449650 467421 454850 467445
rect 118278 467391 123478 467415
rect 118278 467280 118302 467391
rect 118170 465280 118302 467280
rect 118278 465128 118302 465280
rect 123454 467280 123478 467391
rect 377488 467291 378253 467315
rect 377488 467280 377512 467291
rect 123454 465280 180364 467280
rect 338673 465285 377512 467280
rect 378229 467280 378253 467291
rect 397830 467290 398595 467314
rect 397830 467280 397854 467290
rect 378229 465285 397854 467280
rect 338673 465284 397854 465285
rect 398571 467280 398595 467290
rect 449650 467280 449674 467421
rect 398571 465284 449674 467280
rect 338673 465280 449674 465284
rect 123454 465128 123478 465280
rect 377488 465261 378253 465280
rect 397830 465260 398595 465280
rect 449650 465158 449674 465280
rect 454826 465158 454850 467421
rect 449650 465134 454850 465158
rect 118278 465104 123478 465128
rect 437034 463376 442234 463400
rect 130859 463295 136059 463319
rect 130859 463280 130883 463295
rect 130434 461280 130883 463280
rect 130859 461032 130883 461280
rect 136035 463280 136059 463295
rect 378758 463289 379523 463313
rect 378758 463280 378782 463289
rect 136035 461280 180216 463280
rect 338673 461283 378782 463280
rect 379499 463280 379523 463289
rect 396557 463280 397322 463301
rect 437034 463280 437058 463376
rect 379499 463277 437058 463280
rect 379499 461283 396581 463277
rect 338673 461280 396581 461283
rect 136035 461032 136059 461280
rect 378758 461259 379523 461280
rect 396557 461271 396581 461280
rect 397298 461280 437058 463277
rect 397298 461271 397322 461280
rect 396557 461247 397322 461271
rect 437034 461113 437058 461280
rect 442210 463280 442234 463376
rect 442210 461280 442485 463280
rect 442210 461113 442234 461280
rect 437034 461089 442234 461113
rect 130859 461008 136059 461032
rect 565163 196299 566218 196323
rect 565163 196290 565187 196299
rect 449499 196266 565187 196290
rect 449499 191354 449523 196266
rect 454435 191354 565187 196266
rect 449499 191348 565187 191354
rect 566194 196290 566218 196299
rect 570476 196291 575484 196315
rect 570476 196290 570500 196291
rect 566194 191348 570500 196290
rect 449499 191330 570500 191348
rect 565163 191324 566218 191330
rect 570476 191329 570500 191330
rect 575460 191329 575484 196291
rect 570476 191305 575484 191329
rect 570389 186371 575557 186395
rect 570389 186370 570413 186371
rect 449420 186346 570413 186370
rect 449420 181276 449444 186346
rect 454514 186266 570413 186346
rect 454514 181315 565206 186266
rect 566213 181315 570413 186266
rect 454514 181276 570413 181315
rect 449420 181252 570413 181276
rect 570389 181251 570413 181252
rect 575533 181251 575557 186371
rect 570389 181227 575557 181251
rect 13041 177861 18209 177885
rect 13041 172741 13065 177861
rect 18185 177860 18209 177861
rect 18185 177836 454970 177860
rect 18185 177806 118328 177836
rect 18185 172855 24981 177806
rect 25988 172855 118328 177806
rect 18185 172766 118328 172855
rect 123398 172766 449876 177836
rect 454946 172766 454970 177836
rect 18185 172742 454970 172766
rect 18185 172741 18209 172742
rect 13041 172717 18209 172741
rect 13349 167863 18517 167887
rect 13349 162743 13373 167863
rect 18493 167862 18517 167863
rect 18493 167838 454832 167862
rect 18493 167760 118194 167838
rect 18493 162809 25000 167760
rect 26007 162809 118194 167760
rect 18493 162768 118194 162809
rect 123264 162768 449738 167838
rect 454808 162768 454832 167838
rect 18493 162744 454832 162768
rect 18493 162743 18517 162744
rect 13349 162719 18517 162743
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use analog_top  analog_top_0
timestamp 1654899744
transform 1 0 173490 0 1 497666
box 4703 -40917 166970 91353
use digital_filter  digital_filter_0
timestamp 1654899744
transform 1 0 373631 0 1 507651
box 0 0 28796 27744
use sky130_fd_pr__cap_mim_m3_1_PXTAZD  sky130_fd_pr__cap_mim_m3_1_PXTAZD_0
timestamp 1654898484
transform 1 0 158372 0 1 550806
box -12624 -25192 12624 25192
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
<< end >>
