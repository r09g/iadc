magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< pwell >>
rect -646 260 647 261
rect -647 -261 647 260
<< nmos >>
rect -447 -51 -417 51
rect -351 -51 -321 51
rect -255 -51 -225 51
rect -159 -51 -129 51
rect -63 -51 -33 51
rect 33 -51 63 51
rect 129 -51 159 51
rect 225 -51 255 51
rect 321 -51 351 51
rect 417 -51 447 51
<< ndiff >>
rect -509 39 -447 51
rect -509 -39 -497 39
rect -463 -39 -447 39
rect -509 -51 -447 -39
rect -417 39 -351 51
rect -417 -39 -401 39
rect -367 -39 -351 39
rect -417 -51 -351 -39
rect -321 39 -255 51
rect -321 -39 -305 39
rect -271 -39 -255 39
rect -321 -51 -255 -39
rect -225 39 -159 51
rect -225 -39 -209 39
rect -175 -39 -159 39
rect -225 -51 -159 -39
rect -129 39 -63 51
rect -129 -39 -113 39
rect -79 -39 -63 39
rect -129 -51 -63 -39
rect -33 39 33 51
rect -33 -39 -17 39
rect 17 -39 33 39
rect -33 -51 33 -39
rect 63 39 129 51
rect 63 -39 79 39
rect 113 -39 129 39
rect 63 -51 129 -39
rect 159 39 225 51
rect 159 -39 175 39
rect 209 -39 225 39
rect 159 -51 225 -39
rect 255 39 321 51
rect 255 -39 271 39
rect 305 -39 321 39
rect 255 -51 321 -39
rect 351 39 417 51
rect 351 -39 367 39
rect 401 -39 417 39
rect 351 -51 417 -39
rect 447 39 509 51
rect 447 -39 463 39
rect 497 -39 509 39
rect 447 -51 509 -39
<< ndiffc >>
rect -497 -39 -463 39
rect -401 -39 -367 39
rect -305 -39 -271 39
rect -209 -39 -175 39
rect -113 -39 -79 39
rect -17 -39 17 39
rect 79 -39 113 39
rect 175 -39 209 39
rect 271 -39 305 39
rect 367 -39 401 39
rect 463 -39 497 39
<< psubdiff >>
rect -611 191 -515 225
rect 515 191 611 225
rect -611 129 -577 191
rect 577 129 611 191
rect -611 -191 -577 -129
rect 577 -191 611 -129
rect -611 -225 -515 -191
rect 515 -225 611 -191
<< psubdiffcont >>
rect -515 191 515 225
rect -611 -129 -577 129
rect 577 -129 611 129
rect -515 -225 515 -191
<< poly >>
rect -483 123 -417 139
rect -483 89 -467 123
rect -433 89 -417 123
rect -483 73 -417 89
rect -447 51 -417 73
rect -351 123 351 139
rect -351 89 -287 123
rect -253 89 -113 123
rect -79 89 79 123
rect 113 89 271 123
rect 305 89 351 123
rect -351 73 351 89
rect -351 51 -321 73
rect -255 51 -225 73
rect -159 51 -129 73
rect -63 51 -33 73
rect 33 51 63 73
rect 129 51 159 73
rect 225 51 255 73
rect 321 51 351 73
rect 417 123 483 139
rect 417 89 433 123
rect 467 89 483 123
rect 417 73 483 89
rect 417 51 447 73
rect -447 -73 -417 -51
rect -483 -89 -417 -73
rect -351 -77 -321 -51
rect -255 -77 -225 -51
rect -159 -77 -129 -51
rect -63 -77 -33 -51
rect 33 -77 63 -51
rect 129 -77 159 -51
rect 225 -77 255 -51
rect 321 -77 351 -51
rect 417 -73 447 -51
rect -483 -123 -467 -89
rect -433 -123 -417 -89
rect -483 -139 -417 -123
rect 417 -89 483 -73
rect 417 -123 433 -89
rect 467 -123 483 -89
rect 417 -139 483 -123
<< polycont >>
rect -467 89 -433 123
rect -287 89 -253 123
rect -113 89 -79 123
rect 79 89 113 123
rect 271 89 305 123
rect 433 89 467 123
rect -467 -123 -433 -89
rect 433 -123 467 -89
<< locali >>
rect -611 191 -515 225
rect 515 191 611 225
rect -611 129 -577 191
rect -611 -191 -577 -129
rect -497 123 -463 191
rect 463 123 497 191
rect -497 89 -467 123
rect -433 89 -417 123
rect -303 89 -287 123
rect -253 89 -237 123
rect -129 89 -113 123
rect -79 89 -63 123
rect 63 89 79 123
rect 113 89 129 123
rect 255 89 271 123
rect 305 89 321 123
rect 417 89 433 123
rect 467 89 497 123
rect -497 39 -463 89
rect -497 -89 -463 -39
rect -401 39 -367 55
rect -401 -55 -367 -39
rect -305 39 -271 55
rect -497 -123 -467 -89
rect -433 -123 -417 -89
rect -497 -191 -463 -123
rect -305 -191 -271 -39
rect -209 39 -175 55
rect -209 -55 -175 -39
rect -113 39 -79 55
rect -113 -191 -79 -39
rect -17 39 17 55
rect -17 -55 17 -39
rect 79 39 113 55
rect 79 -191 113 -39
rect 175 39 209 55
rect 175 -55 209 -39
rect 271 39 305 55
rect 271 -191 305 -39
rect 367 39 401 55
rect 367 -55 401 -39
rect 463 39 497 89
rect 463 -89 497 -39
rect 417 -123 433 -89
rect 467 -123 497 -89
rect 463 -191 497 -123
rect 577 129 611 191
rect 577 -191 611 -129
rect -611 -225 -515 -191
rect 515 -225 611 -191
<< viali >>
rect -287 89 -253 123
rect -113 89 -79 123
rect 79 89 113 123
rect 271 89 305 123
rect -401 -17 -367 17
rect -209 -17 -175 17
rect -17 -17 17 17
rect 175 -17 209 17
rect 367 -17 401 17
<< metal1 >>
rect -299 123 -241 129
rect -125 123 -67 129
rect 67 123 125 129
rect 259 123 317 129
rect -351 89 -287 123
rect -253 89 -113 123
rect -79 89 79 123
rect 113 89 271 123
rect 305 89 351 123
rect -299 83 -241 89
rect -125 83 -67 89
rect 67 83 125 89
rect 259 83 317 89
rect -413 17 -355 23
rect -221 17 -163 23
rect -29 17 29 23
rect 163 17 221 23
rect 355 17 413 23
rect -413 -17 -401 17
rect -367 -17 -209 17
rect -175 -17 -17 17
rect 17 -17 175 17
rect 209 -17 367 17
rect 401 -17 413 17
rect -413 -23 -355 -17
rect -221 -23 -163 -17
rect -29 -23 29 -17
rect 163 -23 221 -17
rect 355 -23 413 -17
<< properties >>
string FIXED_BBOX -594 -206 594 206
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
