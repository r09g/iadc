magic
tech sky130A
magscale 1 2
timestamp 1654572275
<< error_s >>
rect 257 359 315 365
rect 677 359 735 365
rect 1097 359 1155 365
rect 1517 359 1575 365
rect 1937 359 1995 365
rect 2357 359 2415 365
rect 2777 359 2835 365
rect 3197 359 3255 365
rect 3617 359 3675 365
rect 4037 359 4095 365
rect 4457 359 4515 365
rect 4877 359 4935 365
rect 5297 359 5355 365
rect 5717 359 5775 365
rect 6137 359 6195 365
rect 6557 359 6615 365
rect 6977 359 7035 365
rect 7397 359 7455 365
rect 7817 359 7875 365
rect 8237 359 8295 365
rect 257 325 269 359
rect 677 325 689 359
rect 1097 325 1109 359
rect 1517 325 1529 359
rect 1937 325 1949 359
rect 2357 325 2369 359
rect 2777 325 2789 359
rect 3197 325 3209 359
rect 3617 325 3629 359
rect 4037 325 4049 359
rect 4457 325 4469 359
rect 4877 325 4889 359
rect 5297 325 5309 359
rect 5717 325 5729 359
rect 6137 325 6149 359
rect 6557 325 6569 359
rect 6977 325 6989 359
rect 7397 325 7409 359
rect 7817 325 7829 359
rect 8237 325 8249 359
rect 257 319 315 325
rect 677 319 735 325
rect 1097 319 1155 325
rect 1517 319 1575 325
rect 1937 319 1995 325
rect 2357 319 2415 325
rect 2777 319 2835 325
rect 3197 319 3255 325
rect 3617 319 3675 325
rect 4037 319 4095 325
rect 4457 319 4515 325
rect 4877 319 4935 325
rect 5297 319 5355 325
rect 5717 319 5775 325
rect 6137 319 6195 325
rect 6557 319 6615 325
rect 6977 319 7035 325
rect 7397 319 7455 325
rect 7817 319 7875 325
rect 8237 319 8295 325
rect 467 49 525 55
rect 887 49 945 55
rect 1307 49 1365 55
rect 1727 49 1785 55
rect 2147 49 2205 55
rect 2567 49 2625 55
rect 2987 49 3045 55
rect 3407 49 3465 55
rect 3827 49 3885 55
rect 4247 49 4305 55
rect 4667 49 4725 55
rect 5087 49 5145 55
rect 5507 49 5565 55
rect 5927 49 5985 55
rect 6347 49 6405 55
rect 6767 49 6825 55
rect 7187 49 7245 55
rect 7607 49 7665 55
rect 8027 49 8085 55
rect 8447 49 8505 55
rect 467 15 479 49
rect 887 15 899 49
rect 1307 15 1319 49
rect 1727 15 1739 49
rect 2147 15 2159 49
rect 2567 15 2579 49
rect 2987 15 2999 49
rect 3407 15 3419 49
rect 3827 15 3839 49
rect 4247 15 4259 49
rect 4667 15 4679 49
rect 5087 15 5099 49
rect 5507 15 5519 49
rect 5927 15 5939 49
rect 6347 15 6359 49
rect 6767 15 6779 49
rect 7187 15 7199 49
rect 7607 15 7619 49
rect 8027 15 8039 49
rect 8447 15 8459 49
rect 467 9 525 15
rect 887 9 945 15
rect 1307 9 1365 15
rect 1727 9 1785 15
rect 2147 9 2205 15
rect 2567 9 2625 15
rect 2987 9 3045 15
rect 3407 9 3465 15
rect 3827 9 3885 15
rect 4247 9 4305 15
rect 4667 9 4725 15
rect 5087 9 5145 15
rect 5507 9 5565 15
rect 5927 9 5985 15
rect 6347 9 6405 15
rect 6767 9 6825 15
rect 7187 9 7245 15
rect 7607 9 7665 15
rect 8027 9 8085 15
rect 8447 9 8505 15
rect 257 -81 315 -75
rect 677 -81 735 -75
rect 1097 -81 1155 -75
rect 1517 -81 1575 -75
rect 1937 -81 1995 -75
rect 2357 -81 2415 -75
rect 2777 -81 2835 -75
rect 3197 -81 3255 -75
rect 3617 -81 3675 -75
rect 4037 -81 4095 -75
rect 4457 -81 4515 -75
rect 4877 -81 4935 -75
rect 5297 -81 5355 -75
rect 5717 -81 5775 -75
rect 6137 -81 6195 -75
rect 6557 -81 6615 -75
rect 6977 -81 7035 -75
rect 7397 -81 7455 -75
rect 7817 -81 7875 -75
rect 8237 -81 8295 -75
rect 257 -115 269 -81
rect 677 -115 689 -81
rect 1097 -115 1109 -81
rect 1517 -115 1529 -81
rect 1937 -115 1949 -81
rect 2357 -115 2369 -81
rect 2777 -115 2789 -81
rect 3197 -115 3209 -81
rect 3617 -115 3629 -81
rect 4037 -115 4049 -81
rect 4457 -115 4469 -81
rect 4877 -115 4889 -81
rect 5297 -115 5309 -81
rect 5717 -115 5729 -81
rect 6137 -115 6149 -81
rect 6557 -115 6569 -81
rect 6977 -115 6989 -81
rect 7397 -115 7409 -81
rect 7817 -115 7829 -81
rect 8237 -115 8249 -81
rect 257 -121 315 -115
rect 677 -121 735 -115
rect 1097 -121 1155 -115
rect 1517 -121 1575 -115
rect 1937 -121 1995 -115
rect 2357 -121 2415 -115
rect 2777 -121 2835 -115
rect 3197 -121 3255 -115
rect 3617 -121 3675 -115
rect 4037 -121 4095 -115
rect 4457 -121 4515 -115
rect 4877 -121 4935 -115
rect 5297 -121 5355 -115
rect 5717 -121 5775 -115
rect 6137 -121 6195 -115
rect 6557 -121 6615 -115
rect 6977 -121 7035 -115
rect 7397 -121 7455 -115
rect 7817 -121 7875 -115
rect 8237 -121 8295 -115
rect 467 -391 525 -385
rect 887 -391 945 -385
rect 1307 -391 1365 -385
rect 1727 -391 1785 -385
rect 2147 -391 2205 -385
rect 2567 -391 2625 -385
rect 2987 -391 3045 -385
rect 3407 -391 3465 -385
rect 3827 -391 3885 -385
rect 4247 -391 4305 -385
rect 4667 -391 4725 -385
rect 5087 -391 5145 -385
rect 5507 -391 5565 -385
rect 5927 -391 5985 -385
rect 6347 -391 6405 -385
rect 6767 -391 6825 -385
rect 7187 -391 7245 -385
rect 7607 -391 7665 -385
rect 8027 -391 8085 -385
rect 8447 -391 8505 -385
rect 467 -425 479 -391
rect 887 -425 899 -391
rect 1307 -425 1319 -391
rect 1727 -425 1739 -391
rect 2147 -425 2159 -391
rect 2567 -425 2579 -391
rect 2987 -425 2999 -391
rect 3407 -425 3419 -391
rect 3827 -425 3839 -391
rect 4247 -425 4259 -391
rect 4667 -425 4679 -391
rect 5087 -425 5099 -391
rect 5507 -425 5519 -391
rect 5927 -425 5939 -391
rect 6347 -425 6359 -391
rect 6767 -425 6779 -391
rect 7187 -425 7199 -391
rect 7607 -425 7619 -391
rect 8027 -425 8039 -391
rect 8447 -425 8459 -391
rect 467 -431 525 -425
rect 887 -431 945 -425
rect 1307 -431 1365 -425
rect 1727 -431 1785 -425
rect 2147 -431 2205 -425
rect 2567 -431 2625 -425
rect 2987 -431 3045 -425
rect 3407 -431 3465 -425
rect 3827 -431 3885 -425
rect 4247 -431 4305 -425
rect 4667 -431 4725 -425
rect 5087 -431 5145 -425
rect 5507 -431 5565 -425
rect 5927 -431 5985 -425
rect 6347 -431 6405 -425
rect 6767 -431 6825 -425
rect 7187 -431 7245 -425
rect 7607 -431 7665 -425
rect 8027 -431 8085 -425
rect 8447 -431 8505 -425
rect 257 -521 315 -515
rect 677 -521 735 -515
rect 1097 -521 1155 -515
rect 1517 -521 1575 -515
rect 1937 -521 1995 -515
rect 2357 -521 2415 -515
rect 2777 -521 2835 -515
rect 3197 -521 3255 -515
rect 3617 -521 3675 -515
rect 4037 -521 4095 -515
rect 4457 -521 4515 -515
rect 4877 -521 4935 -515
rect 5297 -521 5355 -515
rect 5717 -521 5775 -515
rect 6137 -521 6195 -515
rect 6557 -521 6615 -515
rect 6977 -521 7035 -515
rect 7397 -521 7455 -515
rect 7817 -521 7875 -515
rect 8237 -521 8295 -515
rect 257 -555 269 -521
rect 677 -555 689 -521
rect 1097 -555 1109 -521
rect 1517 -555 1529 -521
rect 1937 -555 1949 -521
rect 2357 -555 2369 -521
rect 2777 -555 2789 -521
rect 3197 -555 3209 -521
rect 3617 -555 3629 -521
rect 4037 -555 4049 -521
rect 4457 -555 4469 -521
rect 4877 -555 4889 -521
rect 5297 -555 5309 -521
rect 5717 -555 5729 -521
rect 6137 -555 6149 -521
rect 6557 -555 6569 -521
rect 6977 -555 6989 -521
rect 7397 -555 7409 -521
rect 7817 -555 7829 -521
rect 8237 -555 8249 -521
rect 257 -561 315 -555
rect 677 -561 735 -555
rect 1097 -561 1155 -555
rect 1517 -561 1575 -555
rect 1937 -561 1995 -555
rect 2357 -561 2415 -555
rect 2777 -561 2835 -555
rect 3197 -561 3255 -555
rect 3617 -561 3675 -555
rect 4037 -561 4095 -555
rect 4457 -561 4515 -555
rect 4877 -561 4935 -555
rect 5297 -561 5355 -555
rect 5717 -561 5775 -555
rect 6137 -561 6195 -555
rect 6557 -561 6615 -555
rect 6977 -561 7035 -555
rect 7397 -561 7455 -555
rect 7817 -561 7875 -555
rect 8237 -561 8295 -555
rect 467 -831 525 -825
rect 887 -831 945 -825
rect 1307 -831 1365 -825
rect 1727 -831 1785 -825
rect 2147 -831 2205 -825
rect 2567 -831 2625 -825
rect 2987 -831 3045 -825
rect 3407 -831 3465 -825
rect 3827 -831 3885 -825
rect 4247 -831 4305 -825
rect 4667 -831 4725 -825
rect 5087 -831 5145 -825
rect 5507 -831 5565 -825
rect 5927 -831 5985 -825
rect 6347 -831 6405 -825
rect 6767 -831 6825 -825
rect 7187 -831 7245 -825
rect 7607 -831 7665 -825
rect 8027 -831 8085 -825
rect 8447 -831 8505 -825
rect 467 -865 479 -831
rect 887 -865 899 -831
rect 1307 -865 1319 -831
rect 1727 -865 1739 -831
rect 2147 -865 2159 -831
rect 2567 -865 2579 -831
rect 2987 -865 2999 -831
rect 3407 -865 3419 -831
rect 3827 -865 3839 -831
rect 4247 -865 4259 -831
rect 4667 -865 4679 -831
rect 5087 -865 5099 -831
rect 5507 -865 5519 -831
rect 5927 -865 5939 -831
rect 6347 -865 6359 -831
rect 6767 -865 6779 -831
rect 7187 -865 7199 -831
rect 7607 -865 7619 -831
rect 8027 -865 8039 -831
rect 8447 -865 8459 -831
rect 467 -871 525 -865
rect 887 -871 945 -865
rect 1307 -871 1365 -865
rect 1727 -871 1785 -865
rect 2147 -871 2205 -865
rect 2567 -871 2625 -865
rect 2987 -871 3045 -865
rect 3407 -871 3465 -865
rect 3827 -871 3885 -865
rect 4247 -871 4305 -865
rect 4667 -871 4725 -865
rect 5087 -871 5145 -865
rect 5507 -871 5565 -865
rect 5927 -871 5985 -865
rect 6347 -871 6405 -865
rect 6767 -871 6825 -865
rect 7187 -871 7245 -865
rect 7607 -871 7665 -865
rect 8027 -871 8085 -865
rect 8447 -871 8505 -865
rect 257 -961 315 -955
rect 677 -961 735 -955
rect 1097 -961 1155 -955
rect 1517 -961 1575 -955
rect 1937 -961 1995 -955
rect 2357 -961 2415 -955
rect 2777 -961 2835 -955
rect 3197 -961 3255 -955
rect 3617 -961 3675 -955
rect 4037 -961 4095 -955
rect 4457 -961 4515 -955
rect 4877 -961 4935 -955
rect 5297 -961 5355 -955
rect 5717 -961 5775 -955
rect 6137 -961 6195 -955
rect 6557 -961 6615 -955
rect 6977 -961 7035 -955
rect 7397 -961 7455 -955
rect 7817 -961 7875 -955
rect 8237 -961 8295 -955
rect 257 -995 269 -961
rect 677 -995 689 -961
rect 1097 -995 1109 -961
rect 1517 -995 1529 -961
rect 1937 -995 1949 -961
rect 2357 -995 2369 -961
rect 2777 -995 2789 -961
rect 3197 -995 3209 -961
rect 3617 -995 3629 -961
rect 4037 -995 4049 -961
rect 4457 -995 4469 -961
rect 4877 -995 4889 -961
rect 5297 -995 5309 -961
rect 5717 -995 5729 -961
rect 6137 -995 6149 -961
rect 6557 -995 6569 -961
rect 6977 -995 6989 -961
rect 7397 -995 7409 -961
rect 7817 -995 7829 -961
rect 8237 -995 8249 -961
rect 257 -1001 315 -995
rect 677 -1001 735 -995
rect 1097 -1001 1155 -995
rect 1517 -1001 1575 -995
rect 1937 -1001 1995 -995
rect 2357 -1001 2415 -995
rect 2777 -1001 2835 -995
rect 3197 -1001 3255 -995
rect 3617 -1001 3675 -995
rect 4037 -1001 4095 -995
rect 4457 -1001 4515 -995
rect 4877 -1001 4935 -995
rect 5297 -1001 5355 -995
rect 5717 -1001 5775 -995
rect 6137 -1001 6195 -995
rect 6557 -1001 6615 -995
rect 6977 -1001 7035 -995
rect 7397 -1001 7455 -995
rect 7817 -1001 7875 -995
rect 8237 -1001 8295 -995
rect 467 -1271 525 -1265
rect 887 -1271 945 -1265
rect 1307 -1271 1365 -1265
rect 1727 -1271 1785 -1265
rect 2147 -1271 2205 -1265
rect 2567 -1271 2625 -1265
rect 2987 -1271 3045 -1265
rect 3407 -1271 3465 -1265
rect 3827 -1271 3885 -1265
rect 4247 -1271 4305 -1265
rect 4667 -1271 4725 -1265
rect 5087 -1271 5145 -1265
rect 5507 -1271 5565 -1265
rect 5927 -1271 5985 -1265
rect 6347 -1271 6405 -1265
rect 6767 -1271 6825 -1265
rect 7187 -1271 7245 -1265
rect 7607 -1271 7665 -1265
rect 8027 -1271 8085 -1265
rect 8447 -1271 8505 -1265
rect 467 -1305 479 -1271
rect 887 -1305 899 -1271
rect 1307 -1305 1319 -1271
rect 1727 -1305 1739 -1271
rect 2147 -1305 2159 -1271
rect 2567 -1305 2579 -1271
rect 2987 -1305 2999 -1271
rect 3407 -1305 3419 -1271
rect 3827 -1305 3839 -1271
rect 4247 -1305 4259 -1271
rect 4667 -1305 4679 -1271
rect 5087 -1305 5099 -1271
rect 5507 -1305 5519 -1271
rect 5927 -1305 5939 -1271
rect 6347 -1305 6359 -1271
rect 6767 -1305 6779 -1271
rect 7187 -1305 7199 -1271
rect 7607 -1305 7619 -1271
rect 8027 -1305 8039 -1271
rect 8447 -1305 8459 -1271
rect 467 -1311 525 -1305
rect 887 -1311 945 -1305
rect 1307 -1311 1365 -1305
rect 1727 -1311 1785 -1305
rect 2147 -1311 2205 -1305
rect 2567 -1311 2625 -1305
rect 2987 -1311 3045 -1305
rect 3407 -1311 3465 -1305
rect 3827 -1311 3885 -1305
rect 4247 -1311 4305 -1305
rect 4667 -1311 4725 -1305
rect 5087 -1311 5145 -1305
rect 5507 -1311 5565 -1305
rect 5927 -1311 5985 -1305
rect 6347 -1311 6405 -1305
rect 6767 -1311 6825 -1305
rect 7187 -1311 7245 -1305
rect 7607 -1311 7665 -1305
rect 8027 -1311 8085 -1305
rect 8447 -1311 8505 -1305
rect 257 -1401 315 -1395
rect 677 -1401 735 -1395
rect 1097 -1401 1155 -1395
rect 1517 -1401 1575 -1395
rect 1937 -1401 1995 -1395
rect 2357 -1401 2415 -1395
rect 2777 -1401 2835 -1395
rect 3197 -1401 3255 -1395
rect 3617 -1401 3675 -1395
rect 4037 -1401 4095 -1395
rect 4457 -1401 4515 -1395
rect 4877 -1401 4935 -1395
rect 5297 -1401 5355 -1395
rect 5717 -1401 5775 -1395
rect 6137 -1401 6195 -1395
rect 6557 -1401 6615 -1395
rect 6977 -1401 7035 -1395
rect 7397 -1401 7455 -1395
rect 7817 -1401 7875 -1395
rect 8237 -1401 8295 -1395
rect 257 -1435 269 -1401
rect 677 -1435 689 -1401
rect 1097 -1435 1109 -1401
rect 1517 -1435 1529 -1401
rect 1937 -1435 1949 -1401
rect 2357 -1435 2369 -1401
rect 2777 -1435 2789 -1401
rect 3197 -1435 3209 -1401
rect 3617 -1435 3629 -1401
rect 4037 -1435 4049 -1401
rect 4457 -1435 4469 -1401
rect 4877 -1435 4889 -1401
rect 5297 -1435 5309 -1401
rect 5717 -1435 5729 -1401
rect 6137 -1435 6149 -1401
rect 6557 -1435 6569 -1401
rect 6977 -1435 6989 -1401
rect 7397 -1435 7409 -1401
rect 7817 -1435 7829 -1401
rect 8237 -1435 8249 -1401
rect 257 -1441 315 -1435
rect 677 -1441 735 -1435
rect 1097 -1441 1155 -1435
rect 1517 -1441 1575 -1435
rect 1937 -1441 1995 -1435
rect 2357 -1441 2415 -1435
rect 2777 -1441 2835 -1435
rect 3197 -1441 3255 -1435
rect 3617 -1441 3675 -1435
rect 4037 -1441 4095 -1435
rect 4457 -1441 4515 -1435
rect 4877 -1441 4935 -1435
rect 5297 -1441 5355 -1435
rect 5717 -1441 5775 -1435
rect 6137 -1441 6195 -1435
rect 6557 -1441 6615 -1435
rect 6977 -1441 7035 -1435
rect 7397 -1441 7455 -1435
rect 7817 -1441 7875 -1435
rect 8237 -1441 8295 -1435
rect 467 -1711 525 -1705
rect 887 -1711 945 -1705
rect 1307 -1711 1365 -1705
rect 1727 -1711 1785 -1705
rect 2147 -1711 2205 -1705
rect 2567 -1711 2625 -1705
rect 2987 -1711 3045 -1705
rect 3407 -1711 3465 -1705
rect 3827 -1711 3885 -1705
rect 4247 -1711 4305 -1705
rect 4667 -1711 4725 -1705
rect 5087 -1711 5145 -1705
rect 5507 -1711 5565 -1705
rect 5927 -1711 5985 -1705
rect 6347 -1711 6405 -1705
rect 6767 -1711 6825 -1705
rect 7187 -1711 7245 -1705
rect 7607 -1711 7665 -1705
rect 8027 -1711 8085 -1705
rect 8447 -1711 8505 -1705
rect 467 -1745 479 -1711
rect 887 -1745 899 -1711
rect 1307 -1745 1319 -1711
rect 1727 -1745 1739 -1711
rect 2147 -1745 2159 -1711
rect 2567 -1745 2579 -1711
rect 2987 -1745 2999 -1711
rect 3407 -1745 3419 -1711
rect 3827 -1745 3839 -1711
rect 4247 -1745 4259 -1711
rect 4667 -1745 4679 -1711
rect 5087 -1745 5099 -1711
rect 5507 -1745 5519 -1711
rect 5927 -1745 5939 -1711
rect 6347 -1745 6359 -1711
rect 6767 -1745 6779 -1711
rect 7187 -1745 7199 -1711
rect 7607 -1745 7619 -1711
rect 8027 -1745 8039 -1711
rect 8447 -1745 8459 -1711
rect 467 -1751 525 -1745
rect 887 -1751 945 -1745
rect 1307 -1751 1365 -1745
rect 1727 -1751 1785 -1745
rect 2147 -1751 2205 -1745
rect 2567 -1751 2625 -1745
rect 2987 -1751 3045 -1745
rect 3407 -1751 3465 -1745
rect 3827 -1751 3885 -1745
rect 4247 -1751 4305 -1745
rect 4667 -1751 4725 -1745
rect 5087 -1751 5145 -1745
rect 5507 -1751 5565 -1745
rect 5927 -1751 5985 -1745
rect 6347 -1751 6405 -1745
rect 6767 -1751 6825 -1745
rect 7187 -1751 7245 -1745
rect 7607 -1751 7665 -1745
rect 8027 -1751 8085 -1745
rect 8447 -1751 8505 -1745
rect 257 -1841 315 -1835
rect 677 -1841 735 -1835
rect 1097 -1841 1155 -1835
rect 1517 -1841 1575 -1835
rect 1937 -1841 1995 -1835
rect 2357 -1841 2415 -1835
rect 2777 -1841 2835 -1835
rect 3197 -1841 3255 -1835
rect 3617 -1841 3675 -1835
rect 4037 -1841 4095 -1835
rect 4457 -1841 4515 -1835
rect 4877 -1841 4935 -1835
rect 5297 -1841 5355 -1835
rect 5717 -1841 5775 -1835
rect 6137 -1841 6195 -1835
rect 6557 -1841 6615 -1835
rect 6977 -1841 7035 -1835
rect 7397 -1841 7455 -1835
rect 7817 -1841 7875 -1835
rect 8237 -1841 8295 -1835
rect 257 -1875 269 -1841
rect 677 -1875 689 -1841
rect 1097 -1875 1109 -1841
rect 1517 -1875 1529 -1841
rect 1937 -1875 1949 -1841
rect 2357 -1875 2369 -1841
rect 2777 -1875 2789 -1841
rect 3197 -1875 3209 -1841
rect 3617 -1875 3629 -1841
rect 4037 -1875 4049 -1841
rect 4457 -1875 4469 -1841
rect 4877 -1875 4889 -1841
rect 5297 -1875 5309 -1841
rect 5717 -1875 5729 -1841
rect 6137 -1875 6149 -1841
rect 6557 -1875 6569 -1841
rect 6977 -1875 6989 -1841
rect 7397 -1875 7409 -1841
rect 7817 -1875 7829 -1841
rect 8237 -1875 8249 -1841
rect 257 -1881 315 -1875
rect 677 -1881 735 -1875
rect 1097 -1881 1155 -1875
rect 1517 -1881 1575 -1875
rect 1937 -1881 1995 -1875
rect 2357 -1881 2415 -1875
rect 2777 -1881 2835 -1875
rect 3197 -1881 3255 -1875
rect 3617 -1881 3675 -1875
rect 4037 -1881 4095 -1875
rect 4457 -1881 4515 -1875
rect 4877 -1881 4935 -1875
rect 5297 -1881 5355 -1875
rect 5717 -1881 5775 -1875
rect 6137 -1881 6195 -1875
rect 6557 -1881 6615 -1875
rect 6977 -1881 7035 -1875
rect 7397 -1881 7455 -1875
rect 7817 -1881 7875 -1875
rect 8237 -1881 8295 -1875
rect 467 -2151 525 -2145
rect 887 -2151 945 -2145
rect 1307 -2151 1365 -2145
rect 1727 -2151 1785 -2145
rect 2147 -2151 2205 -2145
rect 2567 -2151 2625 -2145
rect 2987 -2151 3045 -2145
rect 3407 -2151 3465 -2145
rect 3827 -2151 3885 -2145
rect 4247 -2151 4305 -2145
rect 4667 -2151 4725 -2145
rect 5087 -2151 5145 -2145
rect 5507 -2151 5565 -2145
rect 5927 -2151 5985 -2145
rect 6347 -2151 6405 -2145
rect 6767 -2151 6825 -2145
rect 7187 -2151 7245 -2145
rect 7607 -2151 7665 -2145
rect 8027 -2151 8085 -2145
rect 8447 -2151 8505 -2145
rect 467 -2185 479 -2151
rect 887 -2185 899 -2151
rect 1307 -2185 1319 -2151
rect 1727 -2185 1739 -2151
rect 2147 -2185 2159 -2151
rect 2567 -2185 2579 -2151
rect 2987 -2185 2999 -2151
rect 3407 -2185 3419 -2151
rect 3827 -2185 3839 -2151
rect 4247 -2185 4259 -2151
rect 4667 -2185 4679 -2151
rect 5087 -2185 5099 -2151
rect 5507 -2185 5519 -2151
rect 5927 -2185 5939 -2151
rect 6347 -2185 6359 -2151
rect 6767 -2185 6779 -2151
rect 7187 -2185 7199 -2151
rect 7607 -2185 7619 -2151
rect 8027 -2185 8039 -2151
rect 8447 -2185 8459 -2151
rect 467 -2191 525 -2185
rect 887 -2191 945 -2185
rect 1307 -2191 1365 -2185
rect 1727 -2191 1785 -2185
rect 2147 -2191 2205 -2185
rect 2567 -2191 2625 -2185
rect 2987 -2191 3045 -2185
rect 3407 -2191 3465 -2185
rect 3827 -2191 3885 -2185
rect 4247 -2191 4305 -2185
rect 4667 -2191 4725 -2185
rect 5087 -2191 5145 -2185
rect 5507 -2191 5565 -2185
rect 5927 -2191 5985 -2185
rect 6347 -2191 6405 -2185
rect 6767 -2191 6825 -2185
rect 7187 -2191 7245 -2185
rect 7607 -2191 7665 -2185
rect 8027 -2191 8085 -2185
rect 8447 -2191 8505 -2185
rect 257 -2281 315 -2275
rect 677 -2281 735 -2275
rect 1097 -2281 1155 -2275
rect 1517 -2281 1575 -2275
rect 1937 -2281 1995 -2275
rect 2357 -2281 2415 -2275
rect 2777 -2281 2835 -2275
rect 3197 -2281 3255 -2275
rect 3617 -2281 3675 -2275
rect 4037 -2281 4095 -2275
rect 4457 -2281 4515 -2275
rect 4877 -2281 4935 -2275
rect 5297 -2281 5355 -2275
rect 5717 -2281 5775 -2275
rect 6137 -2281 6195 -2275
rect 6557 -2281 6615 -2275
rect 6977 -2281 7035 -2275
rect 7397 -2281 7455 -2275
rect 7817 -2281 7875 -2275
rect 8237 -2281 8295 -2275
rect 257 -2315 269 -2281
rect 677 -2315 689 -2281
rect 1097 -2315 1109 -2281
rect 1517 -2315 1529 -2281
rect 1937 -2315 1949 -2281
rect 2357 -2315 2369 -2281
rect 2777 -2315 2789 -2281
rect 3197 -2315 3209 -2281
rect 3617 -2315 3629 -2281
rect 4037 -2315 4049 -2281
rect 4457 -2315 4469 -2281
rect 4877 -2315 4889 -2281
rect 5297 -2315 5309 -2281
rect 5717 -2315 5729 -2281
rect 6137 -2315 6149 -2281
rect 6557 -2315 6569 -2281
rect 6977 -2315 6989 -2281
rect 7397 -2315 7409 -2281
rect 7817 -2315 7829 -2281
rect 8237 -2315 8249 -2281
rect 257 -2321 315 -2315
rect 677 -2321 735 -2315
rect 1097 -2321 1155 -2315
rect 1517 -2321 1575 -2315
rect 1937 -2321 1995 -2315
rect 2357 -2321 2415 -2315
rect 2777 -2321 2835 -2315
rect 3197 -2321 3255 -2315
rect 3617 -2321 3675 -2315
rect 4037 -2321 4095 -2315
rect 4457 -2321 4515 -2315
rect 4877 -2321 4935 -2315
rect 5297 -2321 5355 -2315
rect 5717 -2321 5775 -2315
rect 6137 -2321 6195 -2315
rect 6557 -2321 6615 -2315
rect 6977 -2321 7035 -2315
rect 7397 -2321 7455 -2315
rect 7817 -2321 7875 -2315
rect 8237 -2321 8295 -2315
rect 467 -2591 525 -2585
rect 887 -2591 945 -2585
rect 1307 -2591 1365 -2585
rect 1727 -2591 1785 -2585
rect 2147 -2591 2205 -2585
rect 2567 -2591 2625 -2585
rect 2987 -2591 3045 -2585
rect 3407 -2591 3465 -2585
rect 3827 -2591 3885 -2585
rect 4247 -2591 4305 -2585
rect 4667 -2591 4725 -2585
rect 5087 -2591 5145 -2585
rect 5507 -2591 5565 -2585
rect 5927 -2591 5985 -2585
rect 6347 -2591 6405 -2585
rect 6767 -2591 6825 -2585
rect 7187 -2591 7245 -2585
rect 7607 -2591 7665 -2585
rect 8027 -2591 8085 -2585
rect 8447 -2591 8505 -2585
rect 467 -2625 479 -2591
rect 887 -2625 899 -2591
rect 1307 -2625 1319 -2591
rect 1727 -2625 1739 -2591
rect 2147 -2625 2159 -2591
rect 2567 -2625 2579 -2591
rect 2987 -2625 2999 -2591
rect 3407 -2625 3419 -2591
rect 3827 -2625 3839 -2591
rect 4247 -2625 4259 -2591
rect 4667 -2625 4679 -2591
rect 5087 -2625 5099 -2591
rect 5507 -2625 5519 -2591
rect 5927 -2625 5939 -2591
rect 6347 -2625 6359 -2591
rect 6767 -2625 6779 -2591
rect 7187 -2625 7199 -2591
rect 7607 -2625 7619 -2591
rect 8027 -2625 8039 -2591
rect 8447 -2625 8459 -2591
rect 467 -2631 525 -2625
rect 887 -2631 945 -2625
rect 1307 -2631 1365 -2625
rect 1727 -2631 1785 -2625
rect 2147 -2631 2205 -2625
rect 2567 -2631 2625 -2625
rect 2987 -2631 3045 -2625
rect 3407 -2631 3465 -2625
rect 3827 -2631 3885 -2625
rect 4247 -2631 4305 -2625
rect 4667 -2631 4725 -2625
rect 5087 -2631 5145 -2625
rect 5507 -2631 5565 -2625
rect 5927 -2631 5985 -2625
rect 6347 -2631 6405 -2625
rect 6767 -2631 6825 -2625
rect 7187 -2631 7245 -2625
rect 7607 -2631 7665 -2625
rect 8027 -2631 8085 -2625
rect 8447 -2631 8505 -2625
rect 257 -2721 315 -2715
rect 677 -2721 735 -2715
rect 1097 -2721 1155 -2715
rect 1517 -2721 1575 -2715
rect 1937 -2721 1995 -2715
rect 2357 -2721 2415 -2715
rect 2777 -2721 2835 -2715
rect 3197 -2721 3255 -2715
rect 3617 -2721 3675 -2715
rect 4037 -2721 4095 -2715
rect 4457 -2721 4515 -2715
rect 4877 -2721 4935 -2715
rect 5297 -2721 5355 -2715
rect 5717 -2721 5775 -2715
rect 6137 -2721 6195 -2715
rect 6557 -2721 6615 -2715
rect 6977 -2721 7035 -2715
rect 7397 -2721 7455 -2715
rect 7817 -2721 7875 -2715
rect 8237 -2721 8295 -2715
rect 257 -2755 269 -2721
rect 677 -2755 689 -2721
rect 1097 -2755 1109 -2721
rect 1517 -2755 1529 -2721
rect 1937 -2755 1949 -2721
rect 2357 -2755 2369 -2721
rect 2777 -2755 2789 -2721
rect 3197 -2755 3209 -2721
rect 3617 -2755 3629 -2721
rect 4037 -2755 4049 -2721
rect 4457 -2755 4469 -2721
rect 4877 -2755 4889 -2721
rect 5297 -2755 5309 -2721
rect 5717 -2755 5729 -2721
rect 6137 -2755 6149 -2721
rect 6557 -2755 6569 -2721
rect 6977 -2755 6989 -2721
rect 7397 -2755 7409 -2721
rect 7817 -2755 7829 -2721
rect 8237 -2755 8249 -2721
rect 257 -2761 315 -2755
rect 677 -2761 735 -2755
rect 1097 -2761 1155 -2755
rect 1517 -2761 1575 -2755
rect 1937 -2761 1995 -2755
rect 2357 -2761 2415 -2755
rect 2777 -2761 2835 -2755
rect 3197 -2761 3255 -2755
rect 3617 -2761 3675 -2755
rect 4037 -2761 4095 -2755
rect 4457 -2761 4515 -2755
rect 4877 -2761 4935 -2755
rect 5297 -2761 5355 -2755
rect 5717 -2761 5775 -2755
rect 6137 -2761 6195 -2755
rect 6557 -2761 6615 -2755
rect 6977 -2761 7035 -2755
rect 7397 -2761 7455 -2755
rect 7817 -2761 7875 -2755
rect 8237 -2761 8295 -2755
rect 467 -3031 525 -3025
rect 887 -3031 945 -3025
rect 1307 -3031 1365 -3025
rect 1727 -3031 1785 -3025
rect 2147 -3031 2205 -3025
rect 2567 -3031 2625 -3025
rect 2987 -3031 3045 -3025
rect 3407 -3031 3465 -3025
rect 3827 -3031 3885 -3025
rect 4247 -3031 4305 -3025
rect 4667 -3031 4725 -3025
rect 5087 -3031 5145 -3025
rect 5507 -3031 5565 -3025
rect 5927 -3031 5985 -3025
rect 6347 -3031 6405 -3025
rect 6767 -3031 6825 -3025
rect 7187 -3031 7245 -3025
rect 7607 -3031 7665 -3025
rect 8027 -3031 8085 -3025
rect 8447 -3031 8505 -3025
rect 467 -3065 479 -3031
rect 887 -3065 899 -3031
rect 1307 -3065 1319 -3031
rect 1727 -3065 1739 -3031
rect 2147 -3065 2159 -3031
rect 2567 -3065 2579 -3031
rect 2987 -3065 2999 -3031
rect 3407 -3065 3419 -3031
rect 3827 -3065 3839 -3031
rect 4247 -3065 4259 -3031
rect 4667 -3065 4679 -3031
rect 5087 -3065 5099 -3031
rect 5507 -3065 5519 -3031
rect 5927 -3065 5939 -3031
rect 6347 -3065 6359 -3031
rect 6767 -3065 6779 -3031
rect 7187 -3065 7199 -3031
rect 7607 -3065 7619 -3031
rect 8027 -3065 8039 -3031
rect 8447 -3065 8459 -3031
rect 467 -3071 525 -3065
rect 887 -3071 945 -3065
rect 1307 -3071 1365 -3065
rect 1727 -3071 1785 -3065
rect 2147 -3071 2205 -3065
rect 2567 -3071 2625 -3065
rect 2987 -3071 3045 -3065
rect 3407 -3071 3465 -3065
rect 3827 -3071 3885 -3065
rect 4247 -3071 4305 -3065
rect 4667 -3071 4725 -3065
rect 5087 -3071 5145 -3065
rect 5507 -3071 5565 -3065
rect 5927 -3071 5985 -3065
rect 6347 -3071 6405 -3065
rect 6767 -3071 6825 -3065
rect 7187 -3071 7245 -3065
rect 7607 -3071 7665 -3065
rect 8027 -3071 8085 -3065
rect 8447 -3071 8505 -3065
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_0
timestamp 1654572275
transform 1 0 4381 0 1 187
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_1
timestamp 1654572275
transform 1 0 4381 0 1 -253
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_2
timestamp 1654572275
transform 1 0 4381 0 1 -693
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_3
timestamp 1654572275
transform 1 0 4381 0 1 -1133
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_4
timestamp 1654572275
transform 1 0 4381 0 1 -1573
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_5
timestamp 1654572275
transform 1 0 4381 0 1 -2013
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_6
timestamp 1654572275
transform 1 0 4381 0 1 -2453
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_7
timestamp 1654572275
transform 1 0 4381 0 1 -2893
box -4382 -188 4382 188
<< end >>
