* NGSPICE file created from comparator_flat.ext - technology: sky130A

.subckt comparator_flat clk ip in outp outn VDD VSS
X0 VSS outp a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=3.6639e+12p pd=3.788e+07u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X1 VDD sky130_fd_sc_hd__nand2_4_1/A outn VDD sky130_fd_pr__pfet_01v8_hvt ad=5.351e+12p pd=5.194e+07u as=1.08e+12p ps=1.016e+07u w=1e+06u l=150000u
X2 VDD a_177_3251# sky130_fd_sc_hd__nand2_4_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X3 outn sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=6.375e+11p pd=6.55e+06u as=0p ps=0u w=500000u l=150000u
X5 VDD clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.4e+11p ps=6.56e+06u w=500000u l=150000u
X6 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=3.24e+06u as=8.05e+11p ps=8.22e+06u w=500000u l=150000u
X7 a_282_408# in a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=1.5015e+12p pd=1.504e+07u as=8.05e+11p ps=8.22e+06u w=500000u l=150000u
X8 VSS outp a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VDD sky130_fd_sc_hd__buf_2_0/A a_721_3251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X10 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X11 a_1067_3524# sky130_fd_sc_hd__nand2_4_1/A outn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X12 outp sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=0p ps=0u w=1e+06u l=150000u
X13 VSS a_177_3251# sky130_fd_sc_hd__nand2_4_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X14 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X15 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=3.1e+11p pd=3.24e+06u as=0p ps=0u w=500000u l=150000u
X16 VDD outp outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 outn outp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 outp sky130_fd_sc_hd__nand2_4_0/A a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=8.645e+11p ps=9.16e+06u w=650000u l=150000u
X19 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X20 outn outp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VDD sky130_fd_sc_hd__buf_2_1/A a_177_3251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X22 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X23 a_475_1219# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X24 VDD outn outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VDD sky130_fd_sc_hd__nand2_4_1/A outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VSS a_721_3251# sky130_fd_sc_hd__nand2_4_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X27 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X29 a_282_408# ip a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X30 a_282_408# ip a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X31 a_n16_2554# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X32 a_475_1219# in a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X33 a_282_408# in a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X34 VSS VSS a_n16_2554# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X35 a_203_3524# outn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X37 a_n16_2554# ip a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X38 outn sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VDD sky130_fd_sc_hd__nand2_4_0/A outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VSS sky130_fd_sc_hd__buf_2_1/A a_177_3251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X42 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X43 outp sky130_fd_sc_hd__nand2_4_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 sky130_fd_sc_hd__buf_2_1/A clk VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X45 sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X46 VDD a_721_3251# sky130_fd_sc_hd__nand2_4_1/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X47 VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X48 a_203_3524# sky130_fd_sc_hd__nand2_4_0/A outp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X49 VDD clk a_n16_2554# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
X50 a_475_1219# clk VDD VDD sky130_fd_pr__pfet_01v8 ad=1.425e+11p pd=1.57e+06u as=0p ps=0u w=500000u l=150000u
X51 a_n16_2554# ip a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X52 outp sky130_fd_sc_hd__nand2_4_0/A a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X53 a_1067_3524# outp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X54 outp outn VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 VDD outn outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 outn sky130_fd_sc_hd__nand2_4_1/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X58 VSS VSS a_475_1219# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X59 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X60 a_n16_2554# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X61 outp outn VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 VSS outn a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X63 a_203_3524# outn VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X64 VDD sky130_fd_sc_hd__nand2_4_0/A outp VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_1067_3524# sky130_fd_sc_hd__nand2_4_1/A outn VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X66 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X67 VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X68 outn sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X69 a_282_408# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X70 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X71 VDD outp outn VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 VSS outn a_203_3524# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X73 sky130_fd_sc_hd__nand2_4_1/A a_721_3251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 VDD VDD sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X75 a_475_1219# in a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X76 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X77 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X78 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X79 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X80 VSS clk a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X81 a_203_3524# sky130_fd_sc_hd__nand2_4_0/A outp VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X82 a_475_1219# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X83 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X84 a_1067_3524# outp VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X85 VSS sky130_fd_sc_hd__buf_2_0/A a_721_3251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X86 a_282_408# clk VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
X87 VSS VSS a_282_408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=510000u l=150000u
C0 a_721_3251# sky130_fd_sc_hd__buf_2_0/A 0.26fF
C1 a_721_3251# outp 0.02fF
C2 sky130_fd_sc_hd__nand2_4_1/A a_1067_3524# 0.14fF
C3 a_n16_2554# sky130_fd_sc_hd__buf_2_1/A 1.44fF
C4 sky130_fd_sc_hd__nand2_4_1/A a_475_1219# 0.00fF
C5 sky130_fd_sc_hd__buf_2_0/A clk 0.04fF
C6 a_475_1219# a_n16_2554# 1.23fF
C7 a_203_3524# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C8 in a_n16_2554# 0.32fF
C9 a_475_1219# sky130_fd_sc_hd__buf_2_1/A 0.65fF
C10 ip a_n16_2554# 0.97fF
C11 in sky130_fd_sc_hd__buf_2_1/A 0.15fF
C12 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_1/A 0.10fF
C13 ip sky130_fd_sc_hd__buf_2_1/A 0.22fF
C14 VDD sky130_fd_sc_hd__nand2_4_1/A 0.74fF
C15 sky130_fd_sc_hd__nand2_4_0/A a_n16_2554# 0.00fF
C16 a_203_3524# a_1067_3524# 0.03fF
C17 in a_475_1219# 1.03fF
C18 a_n16_2554# a_282_408# 0.71fF
C19 VDD a_n16_2554# 0.44fF
C20 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__buf_2_1/A 0.07fF
C21 ip a_475_1219# 0.29fF
C22 a_177_3251# a_n16_2554# 0.00fF
C23 sky130_fd_sc_hd__nand2_4_0/A a_1067_3524# 0.01fF
C24 a_282_408# sky130_fd_sc_hd__buf_2_1/A 0.09fF
C25 VDD sky130_fd_sc_hd__buf_2_1/A 3.63fF
C26 ip in 0.93fF
C27 outn sky130_fd_sc_hd__nand2_4_1/A 0.54fF
C28 VDD a_1067_3524# 0.08fF
C29 a_177_3251# sky130_fd_sc_hd__buf_2_1/A 0.26fF
C30 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__nand2_4_1/A 0.07fF
C31 outp sky130_fd_sc_hd__nand2_4_1/A 0.19fF
C32 sky130_fd_sc_hd__nand2_4_0/A a_475_1219# 0.00fF
C33 a_721_3251# sky130_fd_sc_hd__nand2_4_1/A 0.32fF
C34 a_475_1219# a_282_408# 0.73fF
C35 sky130_fd_sc_hd__buf_2_0/A a_n16_2554# 0.91fF
C36 VDD a_475_1219# 0.30fF
C37 sky130_fd_sc_hd__nand2_4_0/A a_203_3524# 0.16fF
C38 in a_282_408# 0.28fF
C39 VDD in 0.04fF
C40 outn sky130_fd_sc_hd__buf_2_1/A 0.05fF
C41 a_721_3251# a_n16_2554# 0.00fF
C42 a_177_3251# a_475_1219# 0.00fF
C43 a_203_3524# VDD 0.08fF
C44 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A 5.69fF
C45 outp sky130_fd_sc_hd__buf_2_1/A 0.05fF
C46 outn a_1067_3524# 0.52fF
C47 ip a_282_408# 0.24fF
C48 ip VDD 0.04fF
C49 a_721_3251# sky130_fd_sc_hd__buf_2_1/A 0.02fF
C50 outp a_1067_3524# 0.39fF
C51 a_203_3524# a_177_3251# 0.02fF
C52 clk a_n16_2554# 0.15fF
C53 a_721_3251# a_1067_3524# 0.02fF
C54 sky130_fd_sc_hd__nand2_4_0/A VDD 0.80fF
C55 sky130_fd_sc_hd__buf_2_0/A a_475_1219# 1.33fF
C56 a_203_3524# outn 0.41fF
C57 clk sky130_fd_sc_hd__buf_2_1/A 0.05fF
C58 sky130_fd_sc_hd__buf_2_0/A in 0.21fF
C59 VDD a_282_408# 0.02fF
C60 a_721_3251# a_475_1219# 0.00fF
C61 sky130_fd_sc_hd__nand2_4_0/A a_177_3251# 0.32fF
C62 a_203_3524# outp 0.60fF
C63 sky130_fd_sc_hd__buf_2_0/A ip 0.17fF
C64 VDD a_177_3251# 0.49fF
C65 sky130_fd_sc_hd__nand2_4_0/A outn 0.19fF
C66 clk a_475_1219# 0.13fF
C67 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__buf_2_0/A 0.02fF
C68 sky130_fd_sc_hd__nand2_4_0/A outp 0.56fF
C69 in clk 0.07fF
C70 outn VDD 2.31fF
C71 sky130_fd_sc_hd__buf_2_0/A a_282_408# 0.09fF
C72 sky130_fd_sc_hd__buf_2_0/A VDD 3.75fF
C73 outp VDD 2.29fF
C74 ip clk 0.09fF
C75 outn a_177_3251# 0.02fF
C76 a_721_3251# VDD 0.47fF
C77 sky130_fd_sc_hd__buf_2_0/A a_177_3251# 0.02fF
C78 outp a_177_3251# 0.04fF
C79 a_721_3251# a_177_3251# 0.06fF
C80 sky130_fd_sc_hd__nand2_4_1/A a_n16_2554# 0.00fF
C81 clk a_282_408# 0.48fF
C82 VDD clk 0.56fF
C83 outn sky130_fd_sc_hd__buf_2_0/A 0.04fF
C84 outn outp 1.74fF
C85 outp sky130_fd_sc_hd__buf_2_0/A 0.05fF
C86 outn a_721_3251# 0.04fF
C87 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__buf_2_1/A 0.01fF
C88 clk VSS 2.24fF
C89 in VSS 1.70fF
C90 ip VSS 1.89fF
C91 a_282_408# VSS 1.97fF
C92 a_475_1219# VSS 1.53fF
C93 a_n16_2554# VSS 1.70fF
C94 sky130_fd_sc_hd__buf_2_0/A VSS 2.01fF
C95 sky130_fd_sc_hd__buf_2_1/A VSS 1.88fF
C96 a_721_3251# VSS 0.40fF
C97 a_177_3251# VSS 0.43fF
C98 sky130_fd_sc_hd__nand2_4_1/A VSS 0.68fF
C99 sky130_fd_sc_hd__nand2_4_0/A VSS 0.69fF
C100 a_1067_3524# VSS 0.99fF
C101 outp VSS 1.48fF
C102 outn VSS 1.46fF
C103 a_203_3524# VSS 1.07fF
C104 VDD VSS 7.99fF
.ends

