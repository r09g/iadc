magic
tech sky130A
magscale 1 2
timestamp 1653697205
<< nwell >>
rect 7004 2195 8298 2845
rect 16004 2195 17298 2845
rect 7004 395 8298 1045
rect 16004 395 17298 1045
rect -7664 -7309 3823 -1120
rect 7004 -1405 8298 -755
rect 16004 -1405 17298 -755
rect 7004 -3205 8298 -2555
rect 16004 -3205 17298 -2555
rect 7004 -5005 8298 -4355
rect 16004 -5005 17298 -4355
rect 7004 -6805 8298 -6155
rect 16004 -6805 17298 -6155
<< pwell >>
rect 7004 1731 8298 2193
rect 16004 1731 17298 2193
rect 7004 -69 8298 393
rect 16004 -69 17298 393
rect 7004 -1869 8298 -1407
rect 16004 -1869 17298 -1407
rect 7004 -3669 8298 -3207
rect 16004 -3669 17298 -3207
rect 7004 -5469 8298 -5007
rect 16004 -5469 17298 -5007
rect 7004 -7269 8298 -6807
rect 16004 -7269 17298 -6807
rect -7664 -17642 13838 -7439
<< nmos >>
rect 7204 1941 7234 2045
rect 7300 1941 7330 2045
rect 7396 1941 7426 2045
rect 7492 1941 7522 2045
rect 7588 1941 7618 2045
rect 7684 1941 7714 2045
rect 7780 1941 7810 2045
rect 7876 1941 7906 2045
rect 7972 1941 8002 2045
rect 8068 1941 8098 2045
rect 16204 1941 16234 2045
rect 16300 1941 16330 2045
rect 16396 1941 16426 2045
rect 16492 1941 16522 2045
rect 16588 1941 16618 2045
rect 16684 1941 16714 2045
rect 16780 1941 16810 2045
rect 16876 1941 16906 2045
rect 16972 1941 17002 2045
rect 17068 1941 17098 2045
rect 7204 141 7234 245
rect 7300 141 7330 245
rect 7396 141 7426 245
rect 7492 141 7522 245
rect 7588 141 7618 245
rect 7684 141 7714 245
rect 7780 141 7810 245
rect 7876 141 7906 245
rect 7972 141 8002 245
rect 8068 141 8098 245
rect 16204 141 16234 245
rect 16300 141 16330 245
rect 16396 141 16426 245
rect 16492 141 16522 245
rect 16588 141 16618 245
rect 16684 141 16714 245
rect 16780 141 16810 245
rect 16876 141 16906 245
rect 16972 141 17002 245
rect 17068 141 17098 245
rect 7204 -1659 7234 -1555
rect 7300 -1659 7330 -1555
rect 7396 -1659 7426 -1555
rect 7492 -1659 7522 -1555
rect 7588 -1659 7618 -1555
rect 7684 -1659 7714 -1555
rect 7780 -1659 7810 -1555
rect 7876 -1659 7906 -1555
rect 7972 -1659 8002 -1555
rect 8068 -1659 8098 -1555
rect 16204 -1659 16234 -1555
rect 16300 -1659 16330 -1555
rect 16396 -1659 16426 -1555
rect 16492 -1659 16522 -1555
rect 16588 -1659 16618 -1555
rect 16684 -1659 16714 -1555
rect 16780 -1659 16810 -1555
rect 16876 -1659 16906 -1555
rect 16972 -1659 17002 -1555
rect 17068 -1659 17098 -1555
rect 7204 -3459 7234 -3355
rect 7300 -3459 7330 -3355
rect 7396 -3459 7426 -3355
rect 7492 -3459 7522 -3355
rect 7588 -3459 7618 -3355
rect 7684 -3459 7714 -3355
rect 7780 -3459 7810 -3355
rect 7876 -3459 7906 -3355
rect 7972 -3459 8002 -3355
rect 8068 -3459 8098 -3355
rect 16204 -3459 16234 -3355
rect 16300 -3459 16330 -3355
rect 16396 -3459 16426 -3355
rect 16492 -3459 16522 -3355
rect 16588 -3459 16618 -3355
rect 16684 -3459 16714 -3355
rect 16780 -3459 16810 -3355
rect 16876 -3459 16906 -3355
rect 16972 -3459 17002 -3355
rect 17068 -3459 17098 -3355
rect 7204 -5259 7234 -5155
rect 7300 -5259 7330 -5155
rect 7396 -5259 7426 -5155
rect 7492 -5259 7522 -5155
rect 7588 -5259 7618 -5155
rect 7684 -5259 7714 -5155
rect 7780 -5259 7810 -5155
rect 7876 -5259 7906 -5155
rect 7972 -5259 8002 -5155
rect 8068 -5259 8098 -5155
rect 16204 -5259 16234 -5155
rect 16300 -5259 16330 -5155
rect 16396 -5259 16426 -5155
rect 16492 -5259 16522 -5155
rect 16588 -5259 16618 -5155
rect 16684 -5259 16714 -5155
rect 16780 -5259 16810 -5155
rect 16876 -5259 16906 -5155
rect 16972 -5259 17002 -5155
rect 17068 -5259 17098 -5155
rect 7204 -7059 7234 -6955
rect 7300 -7059 7330 -6955
rect 7396 -7059 7426 -6955
rect 7492 -7059 7522 -6955
rect 7588 -7059 7618 -6955
rect 7684 -7059 7714 -6955
rect 7780 -7059 7810 -6955
rect 7876 -7059 7906 -6955
rect 7972 -7059 8002 -6955
rect 8068 -7059 8098 -6955
rect 16204 -7059 16234 -6955
rect 16300 -7059 16330 -6955
rect 16396 -7059 16426 -6955
rect 16492 -7059 16522 -6955
rect 16588 -7059 16618 -6955
rect 16684 -7059 16714 -6955
rect 16780 -7059 16810 -6955
rect 16876 -7059 16906 -6955
rect 16972 -7059 17002 -6955
rect 17068 -7059 17098 -6955
rect -2127 -8400 -2007 -8120
rect -1949 -8400 -1829 -8120
rect -1771 -8400 -1651 -8120
rect -1593 -8400 -1473 -8120
rect -1415 -8400 -1295 -8120
rect -1237 -8400 -1117 -8120
rect -1059 -8400 -939 -8120
rect -881 -8400 -761 -8120
rect -703 -8400 -583 -8120
rect -525 -8400 -405 -8120
rect -347 -8400 -227 -8120
rect -169 -8400 -49 -8120
rect 9 -8400 129 -8120
rect 187 -8400 307 -8120
rect 365 -8400 485 -8120
rect 543 -8400 663 -8120
rect 721 -8400 841 -8120
rect 899 -8400 1019 -8120
rect 1077 -8400 1197 -8120
rect 1255 -8400 1375 -8120
rect 1433 -8400 1553 -8120
rect 1611 -8400 1731 -8120
rect 1789 -8400 1909 -8120
rect 1967 -8400 2087 -8120
rect 2145 -8400 2265 -8120
rect 2323 -8400 2443 -8120
rect 2501 -8400 2621 -8120
rect 2679 -8400 2799 -8120
rect 2857 -8400 2977 -8120
rect 3035 -8400 3155 -8120
rect 3213 -8400 3333 -8120
rect 3391 -8400 3511 -8120
rect 3569 -8400 3689 -8120
rect 3747 -8400 3867 -8120
rect 3925 -8400 4045 -8120
rect -2127 -9400 -2007 -9120
rect -1949 -9400 -1829 -9120
rect -1771 -9400 -1651 -9120
rect -1593 -9400 -1473 -9120
rect -1415 -9400 -1295 -9120
rect -1237 -9400 -1117 -9120
rect -1059 -9400 -939 -9120
rect -881 -9400 -761 -9120
rect -703 -9400 -583 -9120
rect -525 -9400 -405 -9120
rect -347 -9400 -227 -9120
rect -169 -9400 -49 -9120
rect 9 -9400 129 -9120
rect 187 -9400 307 -9120
rect 365 -9400 485 -9120
rect 543 -9400 663 -9120
rect 721 -9400 841 -9120
rect 899 -9400 1019 -9120
rect 1077 -9400 1197 -9120
rect 1255 -9400 1375 -9120
rect 1433 -9400 1553 -9120
rect 1611 -9400 1731 -9120
rect 1789 -9400 1909 -9120
rect 1967 -9400 2087 -9120
rect 2145 -9400 2265 -9120
rect 2323 -9400 2443 -9120
rect 2501 -9400 2621 -9120
rect 2679 -9400 2799 -9120
rect 2857 -9400 2977 -9120
rect 3035 -9400 3155 -9120
rect 3213 -9400 3333 -9120
rect 3391 -9400 3511 -9120
rect 3569 -9400 3689 -9120
rect 3747 -9400 3867 -9120
rect 3925 -9400 4045 -9120
rect 6558 -9162 6678 -8882
rect 6736 -9162 6856 -8882
rect 6914 -9162 7034 -8882
rect 7092 -9162 7212 -8882
rect 7270 -9162 7390 -8882
rect 7448 -9162 7568 -8882
rect 7626 -9162 7746 -8882
rect 7804 -9162 7924 -8882
rect 7982 -9162 8102 -8882
rect 8160 -9162 8280 -8882
rect 8338 -9162 8458 -8882
rect 8516 -9162 8636 -8882
rect 8694 -9162 8814 -8882
rect 8872 -9162 8992 -8882
rect 9050 -9162 9170 -8882
rect 9228 -9162 9348 -8882
rect 10818 -9192 10938 -8912
rect 11110 -9192 11230 -8912
rect 11402 -9192 11522 -8912
rect 11694 -9192 11814 -8912
rect 11986 -9192 12106 -8912
rect 12278 -9192 12398 -8912
rect 12570 -9192 12690 -8912
rect 6558 -10062 6678 -9782
rect 6736 -10062 6856 -9782
rect 6914 -10062 7034 -9782
rect 7092 -10062 7212 -9782
rect 7270 -10062 7390 -9782
rect 7448 -10062 7568 -9782
rect 7626 -10062 7746 -9782
rect 7804 -10062 7924 -9782
rect 7982 -10062 8102 -9782
rect 8160 -10062 8280 -9782
rect 8338 -10062 8458 -9782
rect 8516 -10062 8636 -9782
rect 8694 -10062 8814 -9782
rect 8872 -10062 8992 -9782
rect 9050 -10062 9170 -9782
rect 9228 -10062 9348 -9782
rect 10818 -9962 10938 -9682
rect 11110 -9962 11230 -9682
rect 11402 -9962 11522 -9682
rect 11694 -9962 11814 -9682
rect 11986 -9962 12106 -9682
rect 12278 -9962 12398 -9682
rect 12570 -9962 12690 -9682
rect -2127 -10400 -2007 -10120
rect -1949 -10400 -1829 -10120
rect -1771 -10400 -1651 -10120
rect -1593 -10400 -1473 -10120
rect -1415 -10400 -1295 -10120
rect -1237 -10400 -1117 -10120
rect -1059 -10400 -939 -10120
rect -881 -10400 -761 -10120
rect -703 -10400 -583 -10120
rect -525 -10400 -405 -10120
rect -347 -10400 -227 -10120
rect -169 -10400 -49 -10120
rect 9 -10400 129 -10120
rect 187 -10400 307 -10120
rect 365 -10400 485 -10120
rect 543 -10400 663 -10120
rect 721 -10400 841 -10120
rect 899 -10400 1019 -10120
rect 1077 -10400 1197 -10120
rect 1255 -10400 1375 -10120
rect 1433 -10400 1553 -10120
rect 1611 -10400 1731 -10120
rect 1789 -10400 1909 -10120
rect 1967 -10400 2087 -10120
rect 2145 -10400 2265 -10120
rect 2323 -10400 2443 -10120
rect 2501 -10400 2621 -10120
rect 2679 -10400 2799 -10120
rect 2857 -10400 2977 -10120
rect 3035 -10400 3155 -10120
rect 3213 -10400 3333 -10120
rect 3391 -10400 3511 -10120
rect 3569 -10400 3689 -10120
rect 3747 -10400 3867 -10120
rect 3925 -10400 4045 -10120
rect 6558 -10962 6678 -10682
rect 6736 -10962 6856 -10682
rect 6914 -10962 7034 -10682
rect 7092 -10962 7212 -10682
rect 7270 -10962 7390 -10682
rect 7448 -10962 7568 -10682
rect 7626 -10962 7746 -10682
rect 7804 -10962 7924 -10682
rect 7982 -10962 8102 -10682
rect 8160 -10962 8280 -10682
rect 8338 -10962 8458 -10682
rect 8516 -10962 8636 -10682
rect 8694 -10962 8814 -10682
rect 8872 -10962 8992 -10682
rect 9050 -10962 9170 -10682
rect 9228 -10962 9348 -10682
rect 10818 -10732 10938 -10452
rect 11110 -10732 11230 -10452
rect 11402 -10732 11522 -10452
rect 11694 -10732 11814 -10452
rect 11986 -10732 12106 -10452
rect 12278 -10732 12398 -10452
rect 12570 -10732 12690 -10452
rect -2127 -11400 -2007 -11120
rect -1949 -11400 -1829 -11120
rect -1771 -11400 -1651 -11120
rect -1593 -11400 -1473 -11120
rect -1415 -11400 -1295 -11120
rect -1237 -11400 -1117 -11120
rect -1059 -11400 -939 -11120
rect -881 -11400 -761 -11120
rect -703 -11400 -583 -11120
rect -525 -11400 -405 -11120
rect -347 -11400 -227 -11120
rect -169 -11400 -49 -11120
rect 9 -11400 129 -11120
rect 187 -11400 307 -11120
rect 365 -11400 485 -11120
rect 543 -11400 663 -11120
rect 721 -11400 841 -11120
rect 899 -11400 1019 -11120
rect 1077 -11400 1197 -11120
rect 1255 -11400 1375 -11120
rect 1433 -11400 1553 -11120
rect 1611 -11400 1731 -11120
rect 1789 -11400 1909 -11120
rect 1967 -11400 2087 -11120
rect 2145 -11400 2265 -11120
rect 2323 -11400 2443 -11120
rect 2501 -11400 2621 -11120
rect 2679 -11400 2799 -11120
rect 2857 -11400 2977 -11120
rect 3035 -11400 3155 -11120
rect 3213 -11400 3333 -11120
rect 3391 -11400 3511 -11120
rect 3569 -11400 3689 -11120
rect 3747 -11400 3867 -11120
rect 3925 -11400 4045 -11120
rect 10818 -11502 10938 -11222
rect 11110 -11502 11230 -11222
rect 11402 -11502 11522 -11222
rect 11694 -11502 11814 -11222
rect 11986 -11502 12106 -11222
rect 12278 -11502 12398 -11222
rect 12570 -11502 12690 -11222
rect 6558 -11862 6678 -11582
rect 6736 -11862 6856 -11582
rect 6914 -11862 7034 -11582
rect 7092 -11862 7212 -11582
rect 7270 -11862 7390 -11582
rect 7448 -11862 7568 -11582
rect 7626 -11862 7746 -11582
rect 7804 -11862 7924 -11582
rect 7982 -11862 8102 -11582
rect 8160 -11862 8280 -11582
rect 8338 -11862 8458 -11582
rect 8516 -11862 8636 -11582
rect 8694 -11862 8814 -11582
rect 8872 -11862 8992 -11582
rect 9050 -11862 9170 -11582
rect 9228 -11862 9348 -11582
rect -2127 -12400 -2007 -12120
rect -1949 -12400 -1829 -12120
rect -1771 -12400 -1651 -12120
rect -1593 -12400 -1473 -12120
rect -1415 -12400 -1295 -12120
rect -1237 -12400 -1117 -12120
rect -1059 -12400 -939 -12120
rect -881 -12400 -761 -12120
rect -703 -12400 -583 -12120
rect -525 -12400 -405 -12120
rect -347 -12400 -227 -12120
rect -169 -12400 -49 -12120
rect 9 -12400 129 -12120
rect 187 -12400 307 -12120
rect 365 -12400 485 -12120
rect 543 -12400 663 -12120
rect 721 -12400 841 -12120
rect 899 -12400 1019 -12120
rect 1077 -12400 1197 -12120
rect 1255 -12400 1375 -12120
rect 1433 -12400 1553 -12120
rect 1611 -12400 1731 -12120
rect 1789 -12400 1909 -12120
rect 1967 -12400 2087 -12120
rect 2145 -12400 2265 -12120
rect 2323 -12400 2443 -12120
rect 2501 -12400 2621 -12120
rect 2679 -12400 2799 -12120
rect 2857 -12400 2977 -12120
rect 3035 -12400 3155 -12120
rect 3213 -12400 3333 -12120
rect 3391 -12400 3511 -12120
rect 3569 -12400 3689 -12120
rect 3747 -12400 3867 -12120
rect 3925 -12400 4045 -12120
rect -2127 -13400 -2007 -13120
rect -1949 -13400 -1829 -13120
rect -1771 -13400 -1651 -13120
rect -1593 -13400 -1473 -13120
rect -1415 -13400 -1295 -13120
rect -1237 -13400 -1117 -13120
rect -1059 -13400 -939 -13120
rect -881 -13400 -761 -13120
rect -703 -13400 -583 -13120
rect -525 -13400 -405 -13120
rect -347 -13400 -227 -13120
rect -169 -13400 -49 -13120
rect 9 -13400 129 -13120
rect 187 -13400 307 -13120
rect 365 -13400 485 -13120
rect 543 -13400 663 -13120
rect 721 -13400 841 -13120
rect 899 -13400 1019 -13120
rect 1077 -13400 1197 -13120
rect 1255 -13400 1375 -13120
rect 1433 -13400 1553 -13120
rect 1611 -13400 1731 -13120
rect 1789 -13400 1909 -13120
rect 1967 -13400 2087 -13120
rect 2145 -13400 2265 -13120
rect 2323 -13400 2443 -13120
rect 2501 -13400 2621 -13120
rect 2679 -13400 2799 -13120
rect 2857 -13400 2977 -13120
rect 3035 -13400 3155 -13120
rect 3213 -13400 3333 -13120
rect 3391 -13400 3511 -13120
rect 3569 -13400 3689 -13120
rect 3747 -13400 3867 -13120
rect 3925 -13400 4045 -13120
rect -5982 -14662 -5862 -14382
rect -5804 -14662 -5684 -14382
rect -5626 -14662 -5506 -14382
rect -5448 -14662 -5328 -14382
rect -5270 -14662 -5150 -14382
rect -5092 -14662 -4972 -14382
rect -4914 -14662 -4794 -14382
rect -4736 -14662 -4616 -14382
rect -4558 -14662 -4438 -14382
rect -4380 -14662 -4260 -14382
rect -4202 -14662 -4082 -14382
rect -2127 -14400 -2007 -14120
rect -1949 -14400 -1829 -14120
rect -1771 -14400 -1651 -14120
rect -1593 -14400 -1473 -14120
rect -1415 -14400 -1295 -14120
rect -1237 -14400 -1117 -14120
rect -1059 -14400 -939 -14120
rect -881 -14400 -761 -14120
rect -703 -14400 -583 -14120
rect -525 -14400 -405 -14120
rect -347 -14400 -227 -14120
rect -169 -14400 -49 -14120
rect 9 -14400 129 -14120
rect 187 -14400 307 -14120
rect 365 -14400 485 -14120
rect 543 -14400 663 -14120
rect 721 -14400 841 -14120
rect 899 -14400 1019 -14120
rect 1077 -14400 1197 -14120
rect 1255 -14400 1375 -14120
rect 1433 -14400 1553 -14120
rect 1611 -14400 1731 -14120
rect 1789 -14400 1909 -14120
rect 1967 -14400 2087 -14120
rect 2145 -14400 2265 -14120
rect 2323 -14400 2443 -14120
rect 2501 -14400 2621 -14120
rect 2679 -14400 2799 -14120
rect 2857 -14400 2977 -14120
rect 3035 -14400 3155 -14120
rect 3213 -14400 3333 -14120
rect 3391 -14400 3511 -14120
rect 3569 -14400 3689 -14120
rect 3747 -14400 3867 -14120
rect 3925 -14400 4045 -14120
rect 5623 -14400 5743 -14120
rect 5801 -14400 5921 -14120
rect 5979 -14400 6099 -14120
rect 6157 -14400 6277 -14120
rect 6335 -14400 6455 -14120
rect 6513 -14400 6633 -14120
rect 6691 -14400 6811 -14120
rect 6869 -14400 6989 -14120
rect 7047 -14400 7167 -14120
rect 7225 -14400 7345 -14120
rect 7403 -14400 7523 -14120
rect 7581 -14400 7701 -14120
rect 7759 -14400 7879 -14120
rect 7937 -14400 8057 -14120
rect 8115 -14400 8235 -14120
rect 8293 -14400 8413 -14120
rect 8471 -14400 8591 -14120
rect 8649 -14400 8769 -14120
rect 8827 -14400 8947 -14120
rect 9005 -14400 9125 -14120
rect 9183 -14400 9303 -14120
rect 9361 -14400 9481 -14120
rect 9539 -14400 9659 -14120
rect 9717 -14400 9837 -14120
rect 9895 -14400 10015 -14120
rect 10073 -14400 10193 -14120
rect 10251 -14400 10371 -14120
rect 10429 -14400 10549 -14120
rect 10607 -14400 10727 -14120
rect 10785 -14400 10905 -14120
rect 10963 -14400 11083 -14120
rect 11141 -14400 11261 -14120
rect 11319 -14400 11439 -14120
rect 11497 -14400 11617 -14120
rect 11675 -14400 11795 -14120
rect 11853 -14400 11973 -14120
rect 12031 -14400 12151 -14120
rect 12209 -14400 12329 -14120
rect 12387 -14400 12507 -14120
rect 12565 -14400 12685 -14120
rect -5982 -15362 -5862 -15082
rect -5804 -15362 -5684 -15082
rect -5626 -15362 -5506 -15082
rect -5448 -15362 -5328 -15082
rect -5270 -15362 -5150 -15082
rect -5092 -15362 -4972 -15082
rect -4914 -15362 -4794 -15082
rect -4736 -15362 -4616 -15082
rect -4558 -15362 -4438 -15082
rect -4380 -15362 -4260 -15082
rect -4202 -15362 -4082 -15082
rect -2127 -15400 -2007 -15120
rect -1949 -15400 -1829 -15120
rect -1771 -15400 -1651 -15120
rect -1593 -15400 -1473 -15120
rect -1415 -15400 -1295 -15120
rect -1237 -15400 -1117 -15120
rect -1059 -15400 -939 -15120
rect -881 -15400 -761 -15120
rect -703 -15400 -583 -15120
rect -525 -15400 -405 -15120
rect -347 -15400 -227 -15120
rect -169 -15400 -49 -15120
rect 9 -15400 129 -15120
rect 187 -15400 307 -15120
rect 365 -15400 485 -15120
rect 543 -15400 663 -15120
rect 721 -15400 841 -15120
rect 899 -15400 1019 -15120
rect 1077 -15400 1197 -15120
rect 1255 -15400 1375 -15120
rect 1433 -15400 1553 -15120
rect 1611 -15400 1731 -15120
rect 1789 -15400 1909 -15120
rect 1967 -15400 2087 -15120
rect 2145 -15400 2265 -15120
rect 2323 -15400 2443 -15120
rect 2501 -15400 2621 -15120
rect 2679 -15400 2799 -15120
rect 2857 -15400 2977 -15120
rect 3035 -15400 3155 -15120
rect 3213 -15400 3333 -15120
rect 3391 -15400 3511 -15120
rect 3569 -15400 3689 -15120
rect 3747 -15400 3867 -15120
rect 3925 -15400 4045 -15120
rect 5623 -15400 5743 -15120
rect 5801 -15400 5921 -15120
rect 5979 -15400 6099 -15120
rect 6157 -15400 6277 -15120
rect 6335 -15400 6455 -15120
rect 6513 -15400 6633 -15120
rect 6691 -15400 6811 -15120
rect 6869 -15400 6989 -15120
rect 7047 -15400 7167 -15120
rect 7225 -15400 7345 -15120
rect 7403 -15400 7523 -15120
rect 7581 -15400 7701 -15120
rect 7759 -15400 7879 -15120
rect 7937 -15400 8057 -15120
rect 8115 -15400 8235 -15120
rect 8293 -15400 8413 -15120
rect 8471 -15400 8591 -15120
rect 8649 -15400 8769 -15120
rect 8827 -15400 8947 -15120
rect 9005 -15400 9125 -15120
rect 9183 -15400 9303 -15120
rect 9361 -15400 9481 -15120
rect 9539 -15400 9659 -15120
rect 9717 -15400 9837 -15120
rect 9895 -15400 10015 -15120
rect 10073 -15400 10193 -15120
rect 10251 -15400 10371 -15120
rect 10429 -15400 10549 -15120
rect 10607 -15400 10727 -15120
rect 10785 -15400 10905 -15120
rect 10963 -15400 11083 -15120
rect 11141 -15400 11261 -15120
rect 11319 -15400 11439 -15120
rect 11497 -15400 11617 -15120
rect 11675 -15400 11795 -15120
rect 11853 -15400 11973 -15120
rect 12031 -15400 12151 -15120
rect 12209 -15400 12329 -15120
rect 12387 -15400 12507 -15120
rect 12565 -15400 12685 -15120
rect -5982 -16062 -5862 -15782
rect -5804 -16062 -5684 -15782
rect -5626 -16062 -5506 -15782
rect -5448 -16062 -5328 -15782
rect -5270 -16062 -5150 -15782
rect -5092 -16062 -4972 -15782
rect -4914 -16062 -4794 -15782
rect -4736 -16062 -4616 -15782
rect -4558 -16062 -4438 -15782
rect -4380 -16062 -4260 -15782
rect -4202 -16062 -4082 -15782
rect -2127 -16400 -2007 -16120
rect -1949 -16400 -1829 -16120
rect -1771 -16400 -1651 -16120
rect -1593 -16400 -1473 -16120
rect -1415 -16400 -1295 -16120
rect -1237 -16400 -1117 -16120
rect -1059 -16400 -939 -16120
rect -881 -16400 -761 -16120
rect -703 -16400 -583 -16120
rect -525 -16400 -405 -16120
rect -347 -16400 -227 -16120
rect -169 -16400 -49 -16120
rect 9 -16400 129 -16120
rect 187 -16400 307 -16120
rect 365 -16400 485 -16120
rect 543 -16400 663 -16120
rect 721 -16400 841 -16120
rect 899 -16400 1019 -16120
rect 1077 -16400 1197 -16120
rect 1255 -16400 1375 -16120
rect 1433 -16400 1553 -16120
rect 1611 -16400 1731 -16120
rect 1789 -16400 1909 -16120
rect 1967 -16400 2087 -16120
rect 2145 -16400 2265 -16120
rect 2323 -16400 2443 -16120
rect 2501 -16400 2621 -16120
rect 2679 -16400 2799 -16120
rect 2857 -16400 2977 -16120
rect 3035 -16400 3155 -16120
rect 3213 -16400 3333 -16120
rect 3391 -16400 3511 -16120
rect 3569 -16400 3689 -16120
rect 3747 -16400 3867 -16120
rect 3925 -16400 4045 -16120
rect 5623 -16400 5743 -16120
rect 5801 -16400 5921 -16120
rect 5979 -16400 6099 -16120
rect 6157 -16400 6277 -16120
rect 6335 -16400 6455 -16120
rect 6513 -16400 6633 -16120
rect 6691 -16400 6811 -16120
rect 6869 -16400 6989 -16120
rect 7047 -16400 7167 -16120
rect 7225 -16400 7345 -16120
rect 7403 -16400 7523 -16120
rect 7581 -16400 7701 -16120
rect 7759 -16400 7879 -16120
rect 7937 -16400 8057 -16120
rect 8115 -16400 8235 -16120
rect 8293 -16400 8413 -16120
rect 8471 -16400 8591 -16120
rect 8649 -16400 8769 -16120
rect 8827 -16400 8947 -16120
rect 9005 -16400 9125 -16120
rect 9183 -16400 9303 -16120
rect 9361 -16400 9481 -16120
rect 9539 -16400 9659 -16120
rect 9717 -16400 9837 -16120
rect 9895 -16400 10015 -16120
rect 10073 -16400 10193 -16120
rect 10251 -16400 10371 -16120
rect 10429 -16400 10549 -16120
rect 10607 -16400 10727 -16120
rect 10785 -16400 10905 -16120
rect 10963 -16400 11083 -16120
rect 11141 -16400 11261 -16120
rect 11319 -16400 11439 -16120
rect 11497 -16400 11617 -16120
rect 11675 -16400 11795 -16120
rect 11853 -16400 11973 -16120
rect 12031 -16400 12151 -16120
rect 12209 -16400 12329 -16120
rect 12387 -16400 12507 -16120
rect 12565 -16400 12685 -16120
rect -5982 -16762 -5862 -16482
rect -5804 -16762 -5684 -16482
rect -5626 -16762 -5506 -16482
rect -5448 -16762 -5328 -16482
rect -5270 -16762 -5150 -16482
rect -5092 -16762 -4972 -16482
rect -4914 -16762 -4794 -16482
rect -4736 -16762 -4616 -16482
rect -4558 -16762 -4438 -16482
rect -4380 -16762 -4260 -16482
rect -4202 -16762 -4082 -16482
<< pmos >>
rect 7204 2353 7234 2625
rect 7300 2353 7330 2625
rect 7396 2353 7426 2625
rect 7492 2353 7522 2625
rect 7588 2353 7618 2625
rect 7684 2353 7714 2625
rect 7780 2353 7810 2625
rect 7876 2353 7906 2625
rect 7972 2353 8002 2625
rect 8068 2353 8098 2625
rect 16204 2353 16234 2625
rect 16300 2353 16330 2625
rect 16396 2353 16426 2625
rect 16492 2353 16522 2625
rect 16588 2353 16618 2625
rect 16684 2353 16714 2625
rect 16780 2353 16810 2625
rect 16876 2353 16906 2625
rect 16972 2353 17002 2625
rect 17068 2353 17098 2625
rect 7204 553 7234 825
rect 7300 553 7330 825
rect 7396 553 7426 825
rect 7492 553 7522 825
rect 7588 553 7618 825
rect 7684 553 7714 825
rect 7780 553 7810 825
rect 7876 553 7906 825
rect 7972 553 8002 825
rect 8068 553 8098 825
rect 16204 553 16234 825
rect 16300 553 16330 825
rect 16396 553 16426 825
rect 16492 553 16522 825
rect 16588 553 16618 825
rect 16684 553 16714 825
rect 16780 553 16810 825
rect 16876 553 16906 825
rect 16972 553 17002 825
rect 17068 553 17098 825
rect 7204 -1247 7234 -975
rect 7300 -1247 7330 -975
rect 7396 -1247 7426 -975
rect 7492 -1247 7522 -975
rect 7588 -1247 7618 -975
rect 7684 -1247 7714 -975
rect 7780 -1247 7810 -975
rect 7876 -1247 7906 -975
rect 7972 -1247 8002 -975
rect 8068 -1247 8098 -975
rect 16204 -1247 16234 -975
rect 16300 -1247 16330 -975
rect 16396 -1247 16426 -975
rect 16492 -1247 16522 -975
rect 16588 -1247 16618 -975
rect 16684 -1247 16714 -975
rect 16780 -1247 16810 -975
rect 16876 -1247 16906 -975
rect 16972 -1247 17002 -975
rect 17068 -1247 17098 -975
rect -1408 -3152 -1288 -2872
rect -1230 -3152 -1110 -2872
rect -1052 -3152 -932 -2872
rect -874 -3152 -754 -2872
rect -696 -3152 -576 -2872
rect -518 -3152 -398 -2872
rect -340 -3152 -220 -2872
rect -162 -3152 -42 -2872
rect 16 -3152 136 -2872
rect 194 -3152 314 -2872
rect 372 -3152 492 -2872
rect 550 -3152 670 -2872
rect 728 -3152 848 -2872
rect 906 -3152 1026 -2872
rect 1084 -3152 1204 -2872
rect 1262 -3152 1382 -2872
rect 1440 -3152 1560 -2872
rect 1618 -3152 1738 -2872
rect 1796 -3152 1916 -2872
rect 1974 -3152 2094 -2872
rect 2152 -3152 2272 -2872
rect 2330 -3152 2450 -2872
rect 2508 -3152 2628 -2872
rect -1408 -4052 -1288 -3772
rect -1230 -4052 -1110 -3772
rect -1052 -4052 -932 -3772
rect -874 -4052 -754 -3772
rect -696 -4052 -576 -3772
rect -518 -4052 -398 -3772
rect -340 -4052 -220 -3772
rect -162 -4052 -42 -3772
rect 16 -4052 136 -3772
rect 194 -4052 314 -3772
rect 372 -4052 492 -3772
rect 550 -4052 670 -3772
rect 728 -4052 848 -3772
rect 906 -4052 1026 -3772
rect 1084 -4052 1204 -3772
rect 1262 -4052 1382 -3772
rect 1440 -4052 1560 -3772
rect 1618 -4052 1738 -3772
rect 1796 -4052 1916 -3772
rect 1974 -4052 2094 -3772
rect 2152 -4052 2272 -3772
rect 2330 -4052 2450 -3772
rect 2508 -4052 2628 -3772
rect -1408 -4952 -1288 -4672
rect -1230 -4952 -1110 -4672
rect -1052 -4952 -932 -4672
rect -874 -4952 -754 -4672
rect -696 -4952 -576 -4672
rect -518 -4952 -398 -4672
rect -340 -4952 -220 -4672
rect -162 -4952 -42 -4672
rect 16 -4952 136 -4672
rect 194 -4952 314 -4672
rect 372 -4952 492 -4672
rect 550 -4952 670 -4672
rect 728 -4952 848 -4672
rect 906 -4952 1026 -4672
rect 1084 -4952 1204 -4672
rect 1262 -4952 1382 -4672
rect 1440 -4952 1560 -4672
rect 1618 -4952 1738 -4672
rect 1796 -4952 1916 -4672
rect 1974 -4952 2094 -4672
rect 2152 -4952 2272 -4672
rect 2330 -4952 2450 -4672
rect 2508 -4952 2628 -4672
rect -1408 -5852 -1288 -5572
rect -1230 -5852 -1110 -5572
rect -1052 -5852 -932 -5572
rect -874 -5852 -754 -5572
rect -696 -5852 -576 -5572
rect -518 -5852 -398 -5572
rect -340 -5852 -220 -5572
rect -162 -5852 -42 -5572
rect 16 -5852 136 -5572
rect 194 -5852 314 -5572
rect 372 -5852 492 -5572
rect 550 -5852 670 -5572
rect 728 -5852 848 -5572
rect 906 -5852 1026 -5572
rect 1084 -5852 1204 -5572
rect 1262 -5852 1382 -5572
rect 1440 -5852 1560 -5572
rect 1618 -5852 1738 -5572
rect 1796 -5852 1916 -5572
rect 1974 -5852 2094 -5572
rect 2152 -5852 2272 -5572
rect 2330 -5852 2450 -5572
rect 2508 -5852 2628 -5572
rect 7204 -3047 7234 -2775
rect 7300 -3047 7330 -2775
rect 7396 -3047 7426 -2775
rect 7492 -3047 7522 -2775
rect 7588 -3047 7618 -2775
rect 7684 -3047 7714 -2775
rect 7780 -3047 7810 -2775
rect 7876 -3047 7906 -2775
rect 7972 -3047 8002 -2775
rect 8068 -3047 8098 -2775
rect 16204 -3047 16234 -2775
rect 16300 -3047 16330 -2775
rect 16396 -3047 16426 -2775
rect 16492 -3047 16522 -2775
rect 16588 -3047 16618 -2775
rect 16684 -3047 16714 -2775
rect 16780 -3047 16810 -2775
rect 16876 -3047 16906 -2775
rect 16972 -3047 17002 -2775
rect 17068 -3047 17098 -2775
rect 7204 -4847 7234 -4575
rect 7300 -4847 7330 -4575
rect 7396 -4847 7426 -4575
rect 7492 -4847 7522 -4575
rect 7588 -4847 7618 -4575
rect 7684 -4847 7714 -4575
rect 7780 -4847 7810 -4575
rect 7876 -4847 7906 -4575
rect 7972 -4847 8002 -4575
rect 8068 -4847 8098 -4575
rect 16204 -4847 16234 -4575
rect 16300 -4847 16330 -4575
rect 16396 -4847 16426 -4575
rect 16492 -4847 16522 -4575
rect 16588 -4847 16618 -4575
rect 16684 -4847 16714 -4575
rect 16780 -4847 16810 -4575
rect 16876 -4847 16906 -4575
rect 16972 -4847 17002 -4575
rect 17068 -4847 17098 -4575
rect 7204 -6647 7234 -6375
rect 7300 -6647 7330 -6375
rect 7396 -6647 7426 -6375
rect 7492 -6647 7522 -6375
rect 7588 -6647 7618 -6375
rect 7684 -6647 7714 -6375
rect 7780 -6647 7810 -6375
rect 7876 -6647 7906 -6375
rect 7972 -6647 8002 -6375
rect 8068 -6647 8098 -6375
rect 16204 -6647 16234 -6375
rect 16300 -6647 16330 -6375
rect 16396 -6647 16426 -6375
rect 16492 -6647 16522 -6375
rect 16588 -6647 16618 -6375
rect 16684 -6647 16714 -6375
rect 16780 -6647 16810 -6375
rect 16876 -6647 16906 -6375
rect 16972 -6647 17002 -6375
rect 17068 -6647 17098 -6375
<< pmoslvt >>
rect -6256 -2400 -6136 -2120
rect -6078 -2400 -5958 -2120
rect -5900 -2400 -5780 -2120
rect -5722 -2400 -5602 -2120
rect -5544 -2400 -5424 -2120
rect -5366 -2400 -5246 -2120
rect -5188 -2400 -5068 -2120
rect -5010 -2400 -4890 -2120
rect -4832 -2400 -4712 -2120
rect -4654 -2400 -4534 -2120
rect -4476 -2400 -4356 -2120
rect -4298 -2400 -4178 -2120
rect -4120 -2400 -4000 -2120
rect -3942 -2400 -3822 -2120
rect -3764 -2400 -3644 -2120
rect -3586 -2400 -3466 -2120
rect -6256 -3270 -6136 -2990
rect -6078 -3270 -5958 -2990
rect -5900 -3270 -5780 -2990
rect -5722 -3270 -5602 -2990
rect -5544 -3270 -5424 -2990
rect -5366 -3270 -5246 -2990
rect -5188 -3270 -5068 -2990
rect -5010 -3270 -4890 -2990
rect -4832 -3270 -4712 -2990
rect -4654 -3270 -4534 -2990
rect -4476 -3270 -4356 -2990
rect -4298 -3270 -4178 -2990
rect -4120 -3270 -4000 -2990
rect -3942 -3270 -3822 -2990
rect -3764 -3270 -3644 -2990
rect -3586 -3270 -3466 -2990
rect -6256 -4140 -6136 -3860
rect -6078 -4140 -5958 -3860
rect -5900 -4140 -5780 -3860
rect -5722 -4140 -5602 -3860
rect -5544 -4140 -5424 -3860
rect -5366 -4140 -5246 -3860
rect -5188 -4140 -5068 -3860
rect -5010 -4140 -4890 -3860
rect -4832 -4140 -4712 -3860
rect -4654 -4140 -4534 -3860
rect -4476 -4140 -4356 -3860
rect -4298 -4140 -4178 -3860
rect -4120 -4140 -4000 -3860
rect -3942 -4140 -3822 -3860
rect -3764 -4140 -3644 -3860
rect -3586 -4140 -3466 -3860
rect -6256 -5010 -6136 -4730
rect -6078 -5010 -5958 -4730
rect -5900 -5010 -5780 -4730
rect -5722 -5010 -5602 -4730
rect -5544 -5010 -5424 -4730
rect -5366 -5010 -5246 -4730
rect -5188 -5010 -5068 -4730
rect -5010 -5010 -4890 -4730
rect -4832 -5010 -4712 -4730
rect -4654 -5010 -4534 -4730
rect -4476 -5010 -4356 -4730
rect -4298 -5010 -4178 -4730
rect -4120 -5010 -4000 -4730
rect -3942 -5010 -3822 -4730
rect -3764 -5010 -3644 -4730
rect -3586 -5010 -3466 -4730
rect -6256 -5880 -6136 -5600
rect -6078 -5880 -5958 -5600
rect -5900 -5880 -5780 -5600
rect -5722 -5880 -5602 -5600
rect -5544 -5880 -5424 -5600
rect -5366 -5880 -5246 -5600
rect -5188 -5880 -5068 -5600
rect -5010 -5880 -4890 -5600
rect -4832 -5880 -4712 -5600
rect -4654 -5880 -4534 -5600
rect -4476 -5880 -4356 -5600
rect -4298 -5880 -4178 -5600
rect -4120 -5880 -4000 -5600
rect -3942 -5880 -3822 -5600
rect -3764 -5880 -3644 -5600
rect -3586 -5880 -3466 -5600
<< nmoslvt >>
rect -5582 -8142 -5462 -7862
rect -5404 -8142 -5284 -7862
rect -5226 -8142 -5106 -7862
rect -5048 -8142 -4928 -7862
rect -4870 -8142 -4750 -7862
rect -4692 -8142 -4572 -7862
rect -4514 -8142 -4394 -7862
rect -4336 -8142 -4216 -7862
rect -4158 -8142 -4038 -7862
rect -5582 -8692 -5462 -8412
rect -5404 -8692 -5284 -8412
rect -5226 -8692 -5106 -8412
rect -5048 -8692 -4928 -8412
rect -4870 -8692 -4750 -8412
rect -4692 -8692 -4572 -8412
rect -4514 -8692 -4394 -8412
rect -4336 -8692 -4216 -8412
rect -4158 -8692 -4038 -8412
rect -5582 -9242 -5462 -8962
rect -5404 -9242 -5284 -8962
rect -5226 -9242 -5106 -8962
rect -5048 -9242 -4928 -8962
rect -4870 -9242 -4750 -8962
rect -4692 -9242 -4572 -8962
rect -4514 -9242 -4394 -8962
rect -4336 -9242 -4216 -8962
rect -4158 -9242 -4038 -8962
rect -5582 -9792 -5462 -9512
rect -5404 -9792 -5284 -9512
rect -5226 -9792 -5106 -9512
rect -5048 -9792 -4928 -9512
rect -4870 -9792 -4750 -9512
rect -4692 -9792 -4572 -9512
rect -4514 -9792 -4394 -9512
rect -4336 -9792 -4216 -9512
rect -4158 -9792 -4038 -9512
rect -5582 -10342 -5462 -10062
rect -5404 -10342 -5284 -10062
rect -5226 -10342 -5106 -10062
rect -5048 -10342 -4928 -10062
rect -4870 -10342 -4750 -10062
rect -4692 -10342 -4572 -10062
rect -4514 -10342 -4394 -10062
rect -4336 -10342 -4216 -10062
rect -4158 -10342 -4038 -10062
rect -5582 -10892 -5462 -10612
rect -5404 -10892 -5284 -10612
rect -5226 -10892 -5106 -10612
rect -5048 -10892 -4928 -10612
rect -4870 -10892 -4750 -10612
rect -4692 -10892 -4572 -10612
rect -4514 -10892 -4394 -10612
rect -4336 -10892 -4216 -10612
rect -4158 -10892 -4038 -10612
rect -5582 -11442 -5462 -11162
rect -5404 -11442 -5284 -11162
rect -5226 -11442 -5106 -11162
rect -5048 -11442 -4928 -11162
rect -4870 -11442 -4750 -11162
rect -4692 -11442 -4572 -11162
rect -4514 -11442 -4394 -11162
rect -4336 -11442 -4216 -11162
rect -4158 -11442 -4038 -11162
rect -5582 -11992 -5462 -11712
rect -5404 -11992 -5284 -11712
rect -5226 -11992 -5106 -11712
rect -5048 -11992 -4928 -11712
rect -4870 -11992 -4750 -11712
rect -4692 -11992 -4572 -11712
rect -4514 -11992 -4394 -11712
rect -4336 -11992 -4216 -11712
rect -4158 -11992 -4038 -11712
rect -5871 -12940 -5829 -12700
rect -5621 -12940 -5579 -12700
rect -5371 -12940 -5329 -12700
rect -5121 -12940 -5079 -12700
rect -4871 -12940 -4829 -12700
rect -4621 -12940 -4579 -12700
rect -4371 -12940 -4329 -12700
rect -4121 -12940 -4079 -12700
rect -5871 -13620 -5829 -13380
rect -5621 -13620 -5579 -13380
rect -5371 -13620 -5329 -13380
rect -5121 -13620 -5079 -13380
rect -4871 -13620 -4829 -13380
rect -4621 -13620 -4579 -13380
rect -4371 -13620 -4329 -13380
rect -4121 -13620 -4079 -13380
<< ndiff >>
rect 7142 2033 7204 2045
rect 7142 1953 7154 2033
rect 7188 1953 7204 2033
rect 7142 1941 7204 1953
rect 7234 2033 7300 2045
rect 7234 1953 7250 2033
rect 7284 1953 7300 2033
rect 7234 1941 7300 1953
rect 7330 2033 7396 2045
rect 7330 1953 7346 2033
rect 7380 1953 7396 2033
rect 7330 1941 7396 1953
rect 7426 2033 7492 2045
rect 7426 1953 7442 2033
rect 7476 1953 7492 2033
rect 7426 1941 7492 1953
rect 7522 2033 7588 2045
rect 7522 1953 7538 2033
rect 7572 1953 7588 2033
rect 7522 1941 7588 1953
rect 7618 2033 7684 2045
rect 7618 1953 7634 2033
rect 7668 1953 7684 2033
rect 7618 1941 7684 1953
rect 7714 2033 7780 2045
rect 7714 1953 7730 2033
rect 7764 1953 7780 2033
rect 7714 1941 7780 1953
rect 7810 2033 7876 2045
rect 7810 1953 7826 2033
rect 7860 1953 7876 2033
rect 7810 1941 7876 1953
rect 7906 2033 7972 2045
rect 7906 1953 7922 2033
rect 7956 1953 7972 2033
rect 7906 1941 7972 1953
rect 8002 2033 8068 2045
rect 8002 1953 8018 2033
rect 8052 1953 8068 2033
rect 8002 1941 8068 1953
rect 8098 2033 8160 2045
rect 8098 1953 8114 2033
rect 8148 1953 8160 2033
rect 8098 1941 8160 1953
rect 16142 2033 16204 2045
rect 16142 1953 16154 2033
rect 16188 1953 16204 2033
rect 16142 1941 16204 1953
rect 16234 2033 16300 2045
rect 16234 1953 16250 2033
rect 16284 1953 16300 2033
rect 16234 1941 16300 1953
rect 16330 2033 16396 2045
rect 16330 1953 16346 2033
rect 16380 1953 16396 2033
rect 16330 1941 16396 1953
rect 16426 2033 16492 2045
rect 16426 1953 16442 2033
rect 16476 1953 16492 2033
rect 16426 1941 16492 1953
rect 16522 2033 16588 2045
rect 16522 1953 16538 2033
rect 16572 1953 16588 2033
rect 16522 1941 16588 1953
rect 16618 2033 16684 2045
rect 16618 1953 16634 2033
rect 16668 1953 16684 2033
rect 16618 1941 16684 1953
rect 16714 2033 16780 2045
rect 16714 1953 16730 2033
rect 16764 1953 16780 2033
rect 16714 1941 16780 1953
rect 16810 2033 16876 2045
rect 16810 1953 16826 2033
rect 16860 1953 16876 2033
rect 16810 1941 16876 1953
rect 16906 2033 16972 2045
rect 16906 1953 16922 2033
rect 16956 1953 16972 2033
rect 16906 1941 16972 1953
rect 17002 2033 17068 2045
rect 17002 1953 17018 2033
rect 17052 1953 17068 2033
rect 17002 1941 17068 1953
rect 17098 2033 17160 2045
rect 17098 1953 17114 2033
rect 17148 1953 17160 2033
rect 17098 1941 17160 1953
rect 7142 233 7204 245
rect 7142 153 7154 233
rect 7188 153 7204 233
rect 7142 141 7204 153
rect 7234 233 7300 245
rect 7234 153 7250 233
rect 7284 153 7300 233
rect 7234 141 7300 153
rect 7330 233 7396 245
rect 7330 153 7346 233
rect 7380 153 7396 233
rect 7330 141 7396 153
rect 7426 233 7492 245
rect 7426 153 7442 233
rect 7476 153 7492 233
rect 7426 141 7492 153
rect 7522 233 7588 245
rect 7522 153 7538 233
rect 7572 153 7588 233
rect 7522 141 7588 153
rect 7618 233 7684 245
rect 7618 153 7634 233
rect 7668 153 7684 233
rect 7618 141 7684 153
rect 7714 233 7780 245
rect 7714 153 7730 233
rect 7764 153 7780 233
rect 7714 141 7780 153
rect 7810 233 7876 245
rect 7810 153 7826 233
rect 7860 153 7876 233
rect 7810 141 7876 153
rect 7906 233 7972 245
rect 7906 153 7922 233
rect 7956 153 7972 233
rect 7906 141 7972 153
rect 8002 233 8068 245
rect 8002 153 8018 233
rect 8052 153 8068 233
rect 8002 141 8068 153
rect 8098 233 8160 245
rect 8098 153 8114 233
rect 8148 153 8160 233
rect 8098 141 8160 153
rect 16142 233 16204 245
rect 16142 153 16154 233
rect 16188 153 16204 233
rect 16142 141 16204 153
rect 16234 233 16300 245
rect 16234 153 16250 233
rect 16284 153 16300 233
rect 16234 141 16300 153
rect 16330 233 16396 245
rect 16330 153 16346 233
rect 16380 153 16396 233
rect 16330 141 16396 153
rect 16426 233 16492 245
rect 16426 153 16442 233
rect 16476 153 16492 233
rect 16426 141 16492 153
rect 16522 233 16588 245
rect 16522 153 16538 233
rect 16572 153 16588 233
rect 16522 141 16588 153
rect 16618 233 16684 245
rect 16618 153 16634 233
rect 16668 153 16684 233
rect 16618 141 16684 153
rect 16714 233 16780 245
rect 16714 153 16730 233
rect 16764 153 16780 233
rect 16714 141 16780 153
rect 16810 233 16876 245
rect 16810 153 16826 233
rect 16860 153 16876 233
rect 16810 141 16876 153
rect 16906 233 16972 245
rect 16906 153 16922 233
rect 16956 153 16972 233
rect 16906 141 16972 153
rect 17002 233 17068 245
rect 17002 153 17018 233
rect 17052 153 17068 233
rect 17002 141 17068 153
rect 17098 233 17160 245
rect 17098 153 17114 233
rect 17148 153 17160 233
rect 17098 141 17160 153
rect 7142 -1567 7204 -1555
rect 7142 -1647 7154 -1567
rect 7188 -1647 7204 -1567
rect 7142 -1659 7204 -1647
rect 7234 -1567 7300 -1555
rect 7234 -1647 7250 -1567
rect 7284 -1647 7300 -1567
rect 7234 -1659 7300 -1647
rect 7330 -1567 7396 -1555
rect 7330 -1647 7346 -1567
rect 7380 -1647 7396 -1567
rect 7330 -1659 7396 -1647
rect 7426 -1567 7492 -1555
rect 7426 -1647 7442 -1567
rect 7476 -1647 7492 -1567
rect 7426 -1659 7492 -1647
rect 7522 -1567 7588 -1555
rect 7522 -1647 7538 -1567
rect 7572 -1647 7588 -1567
rect 7522 -1659 7588 -1647
rect 7618 -1567 7684 -1555
rect 7618 -1647 7634 -1567
rect 7668 -1647 7684 -1567
rect 7618 -1659 7684 -1647
rect 7714 -1567 7780 -1555
rect 7714 -1647 7730 -1567
rect 7764 -1647 7780 -1567
rect 7714 -1659 7780 -1647
rect 7810 -1567 7876 -1555
rect 7810 -1647 7826 -1567
rect 7860 -1647 7876 -1567
rect 7810 -1659 7876 -1647
rect 7906 -1567 7972 -1555
rect 7906 -1647 7922 -1567
rect 7956 -1647 7972 -1567
rect 7906 -1659 7972 -1647
rect 8002 -1567 8068 -1555
rect 8002 -1647 8018 -1567
rect 8052 -1647 8068 -1567
rect 8002 -1659 8068 -1647
rect 8098 -1567 8160 -1555
rect 8098 -1647 8114 -1567
rect 8148 -1647 8160 -1567
rect 8098 -1659 8160 -1647
rect 16142 -1567 16204 -1555
rect 16142 -1647 16154 -1567
rect 16188 -1647 16204 -1567
rect 16142 -1659 16204 -1647
rect 16234 -1567 16300 -1555
rect 16234 -1647 16250 -1567
rect 16284 -1647 16300 -1567
rect 16234 -1659 16300 -1647
rect 16330 -1567 16396 -1555
rect 16330 -1647 16346 -1567
rect 16380 -1647 16396 -1567
rect 16330 -1659 16396 -1647
rect 16426 -1567 16492 -1555
rect 16426 -1647 16442 -1567
rect 16476 -1647 16492 -1567
rect 16426 -1659 16492 -1647
rect 16522 -1567 16588 -1555
rect 16522 -1647 16538 -1567
rect 16572 -1647 16588 -1567
rect 16522 -1659 16588 -1647
rect 16618 -1567 16684 -1555
rect 16618 -1647 16634 -1567
rect 16668 -1647 16684 -1567
rect 16618 -1659 16684 -1647
rect 16714 -1567 16780 -1555
rect 16714 -1647 16730 -1567
rect 16764 -1647 16780 -1567
rect 16714 -1659 16780 -1647
rect 16810 -1567 16876 -1555
rect 16810 -1647 16826 -1567
rect 16860 -1647 16876 -1567
rect 16810 -1659 16876 -1647
rect 16906 -1567 16972 -1555
rect 16906 -1647 16922 -1567
rect 16956 -1647 16972 -1567
rect 16906 -1659 16972 -1647
rect 17002 -1567 17068 -1555
rect 17002 -1647 17018 -1567
rect 17052 -1647 17068 -1567
rect 17002 -1659 17068 -1647
rect 17098 -1567 17160 -1555
rect 17098 -1647 17114 -1567
rect 17148 -1647 17160 -1567
rect 17098 -1659 17160 -1647
rect 7142 -3367 7204 -3355
rect 7142 -3447 7154 -3367
rect 7188 -3447 7204 -3367
rect 7142 -3459 7204 -3447
rect 7234 -3367 7300 -3355
rect 7234 -3447 7250 -3367
rect 7284 -3447 7300 -3367
rect 7234 -3459 7300 -3447
rect 7330 -3367 7396 -3355
rect 7330 -3447 7346 -3367
rect 7380 -3447 7396 -3367
rect 7330 -3459 7396 -3447
rect 7426 -3367 7492 -3355
rect 7426 -3447 7442 -3367
rect 7476 -3447 7492 -3367
rect 7426 -3459 7492 -3447
rect 7522 -3367 7588 -3355
rect 7522 -3447 7538 -3367
rect 7572 -3447 7588 -3367
rect 7522 -3459 7588 -3447
rect 7618 -3367 7684 -3355
rect 7618 -3447 7634 -3367
rect 7668 -3447 7684 -3367
rect 7618 -3459 7684 -3447
rect 7714 -3367 7780 -3355
rect 7714 -3447 7730 -3367
rect 7764 -3447 7780 -3367
rect 7714 -3459 7780 -3447
rect 7810 -3367 7876 -3355
rect 7810 -3447 7826 -3367
rect 7860 -3447 7876 -3367
rect 7810 -3459 7876 -3447
rect 7906 -3367 7972 -3355
rect 7906 -3447 7922 -3367
rect 7956 -3447 7972 -3367
rect 7906 -3459 7972 -3447
rect 8002 -3367 8068 -3355
rect 8002 -3447 8018 -3367
rect 8052 -3447 8068 -3367
rect 8002 -3459 8068 -3447
rect 8098 -3367 8160 -3355
rect 8098 -3447 8114 -3367
rect 8148 -3447 8160 -3367
rect 8098 -3459 8160 -3447
rect 16142 -3367 16204 -3355
rect 16142 -3447 16154 -3367
rect 16188 -3447 16204 -3367
rect 16142 -3459 16204 -3447
rect 16234 -3367 16300 -3355
rect 16234 -3447 16250 -3367
rect 16284 -3447 16300 -3367
rect 16234 -3459 16300 -3447
rect 16330 -3367 16396 -3355
rect 16330 -3447 16346 -3367
rect 16380 -3447 16396 -3367
rect 16330 -3459 16396 -3447
rect 16426 -3367 16492 -3355
rect 16426 -3447 16442 -3367
rect 16476 -3447 16492 -3367
rect 16426 -3459 16492 -3447
rect 16522 -3367 16588 -3355
rect 16522 -3447 16538 -3367
rect 16572 -3447 16588 -3367
rect 16522 -3459 16588 -3447
rect 16618 -3367 16684 -3355
rect 16618 -3447 16634 -3367
rect 16668 -3447 16684 -3367
rect 16618 -3459 16684 -3447
rect 16714 -3367 16780 -3355
rect 16714 -3447 16730 -3367
rect 16764 -3447 16780 -3367
rect 16714 -3459 16780 -3447
rect 16810 -3367 16876 -3355
rect 16810 -3447 16826 -3367
rect 16860 -3447 16876 -3367
rect 16810 -3459 16876 -3447
rect 16906 -3367 16972 -3355
rect 16906 -3447 16922 -3367
rect 16956 -3447 16972 -3367
rect 16906 -3459 16972 -3447
rect 17002 -3367 17068 -3355
rect 17002 -3447 17018 -3367
rect 17052 -3447 17068 -3367
rect 17002 -3459 17068 -3447
rect 17098 -3367 17160 -3355
rect 17098 -3447 17114 -3367
rect 17148 -3447 17160 -3367
rect 17098 -3459 17160 -3447
rect 7142 -5167 7204 -5155
rect 7142 -5247 7154 -5167
rect 7188 -5247 7204 -5167
rect 7142 -5259 7204 -5247
rect 7234 -5167 7300 -5155
rect 7234 -5247 7250 -5167
rect 7284 -5247 7300 -5167
rect 7234 -5259 7300 -5247
rect 7330 -5167 7396 -5155
rect 7330 -5247 7346 -5167
rect 7380 -5247 7396 -5167
rect 7330 -5259 7396 -5247
rect 7426 -5167 7492 -5155
rect 7426 -5247 7442 -5167
rect 7476 -5247 7492 -5167
rect 7426 -5259 7492 -5247
rect 7522 -5167 7588 -5155
rect 7522 -5247 7538 -5167
rect 7572 -5247 7588 -5167
rect 7522 -5259 7588 -5247
rect 7618 -5167 7684 -5155
rect 7618 -5247 7634 -5167
rect 7668 -5247 7684 -5167
rect 7618 -5259 7684 -5247
rect 7714 -5167 7780 -5155
rect 7714 -5247 7730 -5167
rect 7764 -5247 7780 -5167
rect 7714 -5259 7780 -5247
rect 7810 -5167 7876 -5155
rect 7810 -5247 7826 -5167
rect 7860 -5247 7876 -5167
rect 7810 -5259 7876 -5247
rect 7906 -5167 7972 -5155
rect 7906 -5247 7922 -5167
rect 7956 -5247 7972 -5167
rect 7906 -5259 7972 -5247
rect 8002 -5167 8068 -5155
rect 8002 -5247 8018 -5167
rect 8052 -5247 8068 -5167
rect 8002 -5259 8068 -5247
rect 8098 -5167 8160 -5155
rect 8098 -5247 8114 -5167
rect 8148 -5247 8160 -5167
rect 8098 -5259 8160 -5247
rect 16142 -5167 16204 -5155
rect 16142 -5247 16154 -5167
rect 16188 -5247 16204 -5167
rect 16142 -5259 16204 -5247
rect 16234 -5167 16300 -5155
rect 16234 -5247 16250 -5167
rect 16284 -5247 16300 -5167
rect 16234 -5259 16300 -5247
rect 16330 -5167 16396 -5155
rect 16330 -5247 16346 -5167
rect 16380 -5247 16396 -5167
rect 16330 -5259 16396 -5247
rect 16426 -5167 16492 -5155
rect 16426 -5247 16442 -5167
rect 16476 -5247 16492 -5167
rect 16426 -5259 16492 -5247
rect 16522 -5167 16588 -5155
rect 16522 -5247 16538 -5167
rect 16572 -5247 16588 -5167
rect 16522 -5259 16588 -5247
rect 16618 -5167 16684 -5155
rect 16618 -5247 16634 -5167
rect 16668 -5247 16684 -5167
rect 16618 -5259 16684 -5247
rect 16714 -5167 16780 -5155
rect 16714 -5247 16730 -5167
rect 16764 -5247 16780 -5167
rect 16714 -5259 16780 -5247
rect 16810 -5167 16876 -5155
rect 16810 -5247 16826 -5167
rect 16860 -5247 16876 -5167
rect 16810 -5259 16876 -5247
rect 16906 -5167 16972 -5155
rect 16906 -5247 16922 -5167
rect 16956 -5247 16972 -5167
rect 16906 -5259 16972 -5247
rect 17002 -5167 17068 -5155
rect 17002 -5247 17018 -5167
rect 17052 -5247 17068 -5167
rect 17002 -5259 17068 -5247
rect 17098 -5167 17160 -5155
rect 17098 -5247 17114 -5167
rect 17148 -5247 17160 -5167
rect 17098 -5259 17160 -5247
rect 7142 -6967 7204 -6955
rect 7142 -7047 7154 -6967
rect 7188 -7047 7204 -6967
rect 7142 -7059 7204 -7047
rect 7234 -6967 7300 -6955
rect 7234 -7047 7250 -6967
rect 7284 -7047 7300 -6967
rect 7234 -7059 7300 -7047
rect 7330 -6967 7396 -6955
rect 7330 -7047 7346 -6967
rect 7380 -7047 7396 -6967
rect 7330 -7059 7396 -7047
rect 7426 -6967 7492 -6955
rect 7426 -7047 7442 -6967
rect 7476 -7047 7492 -6967
rect 7426 -7059 7492 -7047
rect 7522 -6967 7588 -6955
rect 7522 -7047 7538 -6967
rect 7572 -7047 7588 -6967
rect 7522 -7059 7588 -7047
rect 7618 -6967 7684 -6955
rect 7618 -7047 7634 -6967
rect 7668 -7047 7684 -6967
rect 7618 -7059 7684 -7047
rect 7714 -6967 7780 -6955
rect 7714 -7047 7730 -6967
rect 7764 -7047 7780 -6967
rect 7714 -7059 7780 -7047
rect 7810 -6967 7876 -6955
rect 7810 -7047 7826 -6967
rect 7860 -7047 7876 -6967
rect 7810 -7059 7876 -7047
rect 7906 -6967 7972 -6955
rect 7906 -7047 7922 -6967
rect 7956 -7047 7972 -6967
rect 7906 -7059 7972 -7047
rect 8002 -6967 8068 -6955
rect 8002 -7047 8018 -6967
rect 8052 -7047 8068 -6967
rect 8002 -7059 8068 -7047
rect 8098 -6967 8160 -6955
rect 8098 -7047 8114 -6967
rect 8148 -7047 8160 -6967
rect 8098 -7059 8160 -7047
rect 16142 -6967 16204 -6955
rect 16142 -7047 16154 -6967
rect 16188 -7047 16204 -6967
rect 16142 -7059 16204 -7047
rect 16234 -6967 16300 -6955
rect 16234 -7047 16250 -6967
rect 16284 -7047 16300 -6967
rect 16234 -7059 16300 -7047
rect 16330 -6967 16396 -6955
rect 16330 -7047 16346 -6967
rect 16380 -7047 16396 -6967
rect 16330 -7059 16396 -7047
rect 16426 -6967 16492 -6955
rect 16426 -7047 16442 -6967
rect 16476 -7047 16492 -6967
rect 16426 -7059 16492 -7047
rect 16522 -6967 16588 -6955
rect 16522 -7047 16538 -6967
rect 16572 -7047 16588 -6967
rect 16522 -7059 16588 -7047
rect 16618 -6967 16684 -6955
rect 16618 -7047 16634 -6967
rect 16668 -7047 16684 -6967
rect 16618 -7059 16684 -7047
rect 16714 -6967 16780 -6955
rect 16714 -7047 16730 -6967
rect 16764 -7047 16780 -6967
rect 16714 -7059 16780 -7047
rect 16810 -6967 16876 -6955
rect 16810 -7047 16826 -6967
rect 16860 -7047 16876 -6967
rect 16810 -7059 16876 -7047
rect 16906 -6967 16972 -6955
rect 16906 -7047 16922 -6967
rect 16956 -7047 16972 -6967
rect 16906 -7059 16972 -7047
rect 17002 -6967 17068 -6955
rect 17002 -7047 17018 -6967
rect 17052 -7047 17068 -6967
rect 17002 -7059 17068 -7047
rect 17098 -6967 17160 -6955
rect 17098 -7047 17114 -6967
rect 17148 -7047 17160 -6967
rect 17098 -7059 17160 -7047
rect -5640 -7874 -5582 -7862
rect -5640 -8130 -5628 -7874
rect -5594 -8130 -5582 -7874
rect -5640 -8142 -5582 -8130
rect -5462 -7874 -5404 -7862
rect -5462 -8130 -5450 -7874
rect -5416 -8130 -5404 -7874
rect -5462 -8142 -5404 -8130
rect -5284 -7874 -5226 -7862
rect -5284 -8130 -5272 -7874
rect -5238 -8130 -5226 -7874
rect -5284 -8142 -5226 -8130
rect -5106 -7874 -5048 -7862
rect -5106 -8130 -5094 -7874
rect -5060 -8130 -5048 -7874
rect -5106 -8142 -5048 -8130
rect -4928 -7874 -4870 -7862
rect -4928 -8130 -4916 -7874
rect -4882 -8130 -4870 -7874
rect -4928 -8142 -4870 -8130
rect -4750 -7874 -4692 -7862
rect -4750 -8130 -4738 -7874
rect -4704 -8130 -4692 -7874
rect -4750 -8142 -4692 -8130
rect -4572 -7874 -4514 -7862
rect -4572 -8130 -4560 -7874
rect -4526 -8130 -4514 -7874
rect -4572 -8142 -4514 -8130
rect -4394 -7874 -4336 -7862
rect -4394 -8130 -4382 -7874
rect -4348 -8130 -4336 -7874
rect -4394 -8142 -4336 -8130
rect -4216 -7874 -4158 -7862
rect -4216 -8130 -4204 -7874
rect -4170 -8130 -4158 -7874
rect -4216 -8142 -4158 -8130
rect -4038 -7874 -3980 -7862
rect -4038 -8130 -4026 -7874
rect -3992 -8130 -3980 -7874
rect -4038 -8142 -3980 -8130
rect -2185 -8132 -2127 -8120
rect -2185 -8388 -2173 -8132
rect -2139 -8388 -2127 -8132
rect -2185 -8400 -2127 -8388
rect -2007 -8132 -1949 -8120
rect -2007 -8388 -1995 -8132
rect -1961 -8388 -1949 -8132
rect -2007 -8400 -1949 -8388
rect -1829 -8132 -1771 -8120
rect -1829 -8388 -1817 -8132
rect -1783 -8388 -1771 -8132
rect -1829 -8400 -1771 -8388
rect -1651 -8132 -1593 -8120
rect -1651 -8388 -1639 -8132
rect -1605 -8388 -1593 -8132
rect -1651 -8400 -1593 -8388
rect -1473 -8132 -1415 -8120
rect -1473 -8388 -1461 -8132
rect -1427 -8388 -1415 -8132
rect -1473 -8400 -1415 -8388
rect -1295 -8132 -1237 -8120
rect -1295 -8388 -1283 -8132
rect -1249 -8388 -1237 -8132
rect -1295 -8400 -1237 -8388
rect -1117 -8132 -1059 -8120
rect -1117 -8388 -1105 -8132
rect -1071 -8388 -1059 -8132
rect -1117 -8400 -1059 -8388
rect -939 -8132 -881 -8120
rect -939 -8388 -927 -8132
rect -893 -8388 -881 -8132
rect -939 -8400 -881 -8388
rect -761 -8132 -703 -8120
rect -761 -8388 -749 -8132
rect -715 -8388 -703 -8132
rect -761 -8400 -703 -8388
rect -583 -8132 -525 -8120
rect -583 -8388 -571 -8132
rect -537 -8388 -525 -8132
rect -583 -8400 -525 -8388
rect -405 -8132 -347 -8120
rect -405 -8388 -393 -8132
rect -359 -8388 -347 -8132
rect -405 -8400 -347 -8388
rect -227 -8132 -169 -8120
rect -227 -8388 -215 -8132
rect -181 -8388 -169 -8132
rect -227 -8400 -169 -8388
rect -49 -8132 9 -8120
rect -49 -8388 -37 -8132
rect -3 -8388 9 -8132
rect -49 -8400 9 -8388
rect 129 -8132 187 -8120
rect 129 -8388 141 -8132
rect 175 -8388 187 -8132
rect 129 -8400 187 -8388
rect 307 -8132 365 -8120
rect 307 -8388 319 -8132
rect 353 -8388 365 -8132
rect 307 -8400 365 -8388
rect 485 -8132 543 -8120
rect 485 -8388 497 -8132
rect 531 -8388 543 -8132
rect 485 -8400 543 -8388
rect 663 -8132 721 -8120
rect 663 -8388 675 -8132
rect 709 -8388 721 -8132
rect 663 -8400 721 -8388
rect 841 -8132 899 -8120
rect 841 -8388 853 -8132
rect 887 -8388 899 -8132
rect 841 -8400 899 -8388
rect 1019 -8132 1077 -8120
rect 1019 -8388 1031 -8132
rect 1065 -8388 1077 -8132
rect 1019 -8400 1077 -8388
rect 1197 -8132 1255 -8120
rect 1197 -8388 1209 -8132
rect 1243 -8388 1255 -8132
rect 1197 -8400 1255 -8388
rect 1375 -8132 1433 -8120
rect 1375 -8388 1387 -8132
rect 1421 -8388 1433 -8132
rect 1375 -8400 1433 -8388
rect 1553 -8132 1611 -8120
rect 1553 -8388 1565 -8132
rect 1599 -8388 1611 -8132
rect 1553 -8400 1611 -8388
rect 1731 -8132 1789 -8120
rect 1731 -8388 1743 -8132
rect 1777 -8388 1789 -8132
rect 1731 -8400 1789 -8388
rect 1909 -8132 1967 -8120
rect 1909 -8388 1921 -8132
rect 1955 -8388 1967 -8132
rect 1909 -8400 1967 -8388
rect 2087 -8132 2145 -8120
rect 2087 -8388 2099 -8132
rect 2133 -8388 2145 -8132
rect 2087 -8400 2145 -8388
rect 2265 -8132 2323 -8120
rect 2265 -8388 2277 -8132
rect 2311 -8388 2323 -8132
rect 2265 -8400 2323 -8388
rect 2443 -8132 2501 -8120
rect 2443 -8388 2455 -8132
rect 2489 -8388 2501 -8132
rect 2443 -8400 2501 -8388
rect 2621 -8132 2679 -8120
rect 2621 -8388 2633 -8132
rect 2667 -8388 2679 -8132
rect 2621 -8400 2679 -8388
rect 2799 -8132 2857 -8120
rect 2799 -8388 2811 -8132
rect 2845 -8388 2857 -8132
rect 2799 -8400 2857 -8388
rect 2977 -8132 3035 -8120
rect 2977 -8388 2989 -8132
rect 3023 -8388 3035 -8132
rect 2977 -8400 3035 -8388
rect 3155 -8132 3213 -8120
rect 3155 -8388 3167 -8132
rect 3201 -8388 3213 -8132
rect 3155 -8400 3213 -8388
rect 3333 -8132 3391 -8120
rect 3333 -8388 3345 -8132
rect 3379 -8388 3391 -8132
rect 3333 -8400 3391 -8388
rect 3511 -8132 3569 -8120
rect 3511 -8388 3523 -8132
rect 3557 -8388 3569 -8132
rect 3511 -8400 3569 -8388
rect 3689 -8132 3747 -8120
rect 3689 -8388 3701 -8132
rect 3735 -8388 3747 -8132
rect 3689 -8400 3747 -8388
rect 3867 -8132 3925 -8120
rect 3867 -8388 3879 -8132
rect 3913 -8388 3925 -8132
rect 3867 -8400 3925 -8388
rect 4045 -8132 4103 -8120
rect 4045 -8388 4057 -8132
rect 4091 -8388 4103 -8132
rect 4045 -8400 4103 -8388
rect -5640 -8424 -5582 -8412
rect -5640 -8680 -5628 -8424
rect -5594 -8680 -5582 -8424
rect -5640 -8692 -5582 -8680
rect -5462 -8424 -5404 -8412
rect -5462 -8680 -5450 -8424
rect -5416 -8680 -5404 -8424
rect -5462 -8692 -5404 -8680
rect -5284 -8424 -5226 -8412
rect -5284 -8680 -5272 -8424
rect -5238 -8680 -5226 -8424
rect -5284 -8692 -5226 -8680
rect -5106 -8424 -5048 -8412
rect -5106 -8680 -5094 -8424
rect -5060 -8680 -5048 -8424
rect -5106 -8692 -5048 -8680
rect -4928 -8424 -4870 -8412
rect -4928 -8680 -4916 -8424
rect -4882 -8680 -4870 -8424
rect -4928 -8692 -4870 -8680
rect -4750 -8424 -4692 -8412
rect -4750 -8680 -4738 -8424
rect -4704 -8680 -4692 -8424
rect -4750 -8692 -4692 -8680
rect -4572 -8424 -4514 -8412
rect -4572 -8680 -4560 -8424
rect -4526 -8680 -4514 -8424
rect -4572 -8692 -4514 -8680
rect -4394 -8424 -4336 -8412
rect -4394 -8680 -4382 -8424
rect -4348 -8680 -4336 -8424
rect -4394 -8692 -4336 -8680
rect -4216 -8424 -4158 -8412
rect -4216 -8680 -4204 -8424
rect -4170 -8680 -4158 -8424
rect -4216 -8692 -4158 -8680
rect -4038 -8424 -3980 -8412
rect -4038 -8680 -4026 -8424
rect -3992 -8680 -3980 -8424
rect -4038 -8692 -3980 -8680
rect 6500 -8894 6558 -8882
rect -5640 -8974 -5582 -8962
rect -5640 -9230 -5628 -8974
rect -5594 -9230 -5582 -8974
rect -5640 -9242 -5582 -9230
rect -5462 -8974 -5404 -8962
rect -5462 -9230 -5450 -8974
rect -5416 -9230 -5404 -8974
rect -5462 -9242 -5404 -9230
rect -5284 -8974 -5226 -8962
rect -5284 -9230 -5272 -8974
rect -5238 -9230 -5226 -8974
rect -5284 -9242 -5226 -9230
rect -5106 -8974 -5048 -8962
rect -5106 -9230 -5094 -8974
rect -5060 -9230 -5048 -8974
rect -5106 -9242 -5048 -9230
rect -4928 -8974 -4870 -8962
rect -4928 -9230 -4916 -8974
rect -4882 -9230 -4870 -8974
rect -4928 -9242 -4870 -9230
rect -4750 -8974 -4692 -8962
rect -4750 -9230 -4738 -8974
rect -4704 -9230 -4692 -8974
rect -4750 -9242 -4692 -9230
rect -4572 -8974 -4514 -8962
rect -4572 -9230 -4560 -8974
rect -4526 -9230 -4514 -8974
rect -4572 -9242 -4514 -9230
rect -4394 -8974 -4336 -8962
rect -4394 -9230 -4382 -8974
rect -4348 -9230 -4336 -8974
rect -4394 -9242 -4336 -9230
rect -4216 -8974 -4158 -8962
rect -4216 -9230 -4204 -8974
rect -4170 -9230 -4158 -8974
rect -4216 -9242 -4158 -9230
rect -4038 -8974 -3980 -8962
rect -4038 -9230 -4026 -8974
rect -3992 -9230 -3980 -8974
rect -4038 -9242 -3980 -9230
rect -2185 -9132 -2127 -9120
rect -2185 -9388 -2173 -9132
rect -2139 -9388 -2127 -9132
rect -2185 -9400 -2127 -9388
rect -2007 -9132 -1949 -9120
rect -2007 -9388 -1995 -9132
rect -1961 -9388 -1949 -9132
rect -2007 -9400 -1949 -9388
rect -1829 -9132 -1771 -9120
rect -1829 -9388 -1817 -9132
rect -1783 -9388 -1771 -9132
rect -1829 -9400 -1771 -9388
rect -1651 -9132 -1593 -9120
rect -1651 -9388 -1639 -9132
rect -1605 -9388 -1593 -9132
rect -1651 -9400 -1593 -9388
rect -1473 -9132 -1415 -9120
rect -1473 -9388 -1461 -9132
rect -1427 -9388 -1415 -9132
rect -1473 -9400 -1415 -9388
rect -1295 -9132 -1237 -9120
rect -1295 -9388 -1283 -9132
rect -1249 -9388 -1237 -9132
rect -1295 -9400 -1237 -9388
rect -1117 -9132 -1059 -9120
rect -1117 -9388 -1105 -9132
rect -1071 -9388 -1059 -9132
rect -1117 -9400 -1059 -9388
rect -939 -9132 -881 -9120
rect -939 -9388 -927 -9132
rect -893 -9388 -881 -9132
rect -939 -9400 -881 -9388
rect -761 -9132 -703 -9120
rect -761 -9388 -749 -9132
rect -715 -9388 -703 -9132
rect -761 -9400 -703 -9388
rect -583 -9132 -525 -9120
rect -583 -9388 -571 -9132
rect -537 -9388 -525 -9132
rect -583 -9400 -525 -9388
rect -405 -9132 -347 -9120
rect -405 -9388 -393 -9132
rect -359 -9388 -347 -9132
rect -405 -9400 -347 -9388
rect -227 -9132 -169 -9120
rect -227 -9388 -215 -9132
rect -181 -9388 -169 -9132
rect -227 -9400 -169 -9388
rect -49 -9132 9 -9120
rect -49 -9388 -37 -9132
rect -3 -9388 9 -9132
rect -49 -9400 9 -9388
rect 129 -9132 187 -9120
rect 129 -9388 141 -9132
rect 175 -9388 187 -9132
rect 129 -9400 187 -9388
rect 307 -9132 365 -9120
rect 307 -9388 319 -9132
rect 353 -9388 365 -9132
rect 307 -9400 365 -9388
rect 485 -9132 543 -9120
rect 485 -9388 497 -9132
rect 531 -9388 543 -9132
rect 485 -9400 543 -9388
rect 663 -9132 721 -9120
rect 663 -9388 675 -9132
rect 709 -9388 721 -9132
rect 663 -9400 721 -9388
rect 841 -9132 899 -9120
rect 841 -9388 853 -9132
rect 887 -9388 899 -9132
rect 841 -9400 899 -9388
rect 1019 -9132 1077 -9120
rect 1019 -9388 1031 -9132
rect 1065 -9388 1077 -9132
rect 1019 -9400 1077 -9388
rect 1197 -9132 1255 -9120
rect 1197 -9388 1209 -9132
rect 1243 -9388 1255 -9132
rect 1197 -9400 1255 -9388
rect 1375 -9132 1433 -9120
rect 1375 -9388 1387 -9132
rect 1421 -9388 1433 -9132
rect 1375 -9400 1433 -9388
rect 1553 -9132 1611 -9120
rect 1553 -9388 1565 -9132
rect 1599 -9388 1611 -9132
rect 1553 -9400 1611 -9388
rect 1731 -9132 1789 -9120
rect 1731 -9388 1743 -9132
rect 1777 -9388 1789 -9132
rect 1731 -9400 1789 -9388
rect 1909 -9132 1967 -9120
rect 1909 -9388 1921 -9132
rect 1955 -9388 1967 -9132
rect 1909 -9400 1967 -9388
rect 2087 -9132 2145 -9120
rect 2087 -9388 2099 -9132
rect 2133 -9388 2145 -9132
rect 2087 -9400 2145 -9388
rect 2265 -9132 2323 -9120
rect 2265 -9388 2277 -9132
rect 2311 -9388 2323 -9132
rect 2265 -9400 2323 -9388
rect 2443 -9132 2501 -9120
rect 2443 -9388 2455 -9132
rect 2489 -9388 2501 -9132
rect 2443 -9400 2501 -9388
rect 2621 -9132 2679 -9120
rect 2621 -9388 2633 -9132
rect 2667 -9388 2679 -9132
rect 2621 -9400 2679 -9388
rect 2799 -9132 2857 -9120
rect 2799 -9388 2811 -9132
rect 2845 -9388 2857 -9132
rect 2799 -9400 2857 -9388
rect 2977 -9132 3035 -9120
rect 2977 -9388 2989 -9132
rect 3023 -9388 3035 -9132
rect 2977 -9400 3035 -9388
rect 3155 -9132 3213 -9120
rect 3155 -9388 3167 -9132
rect 3201 -9388 3213 -9132
rect 3155 -9400 3213 -9388
rect 3333 -9132 3391 -9120
rect 3333 -9388 3345 -9132
rect 3379 -9388 3391 -9132
rect 3333 -9400 3391 -9388
rect 3511 -9132 3569 -9120
rect 3511 -9388 3523 -9132
rect 3557 -9388 3569 -9132
rect 3511 -9400 3569 -9388
rect 3689 -9132 3747 -9120
rect 3689 -9388 3701 -9132
rect 3735 -9388 3747 -9132
rect 3689 -9400 3747 -9388
rect 3867 -9132 3925 -9120
rect 3867 -9388 3879 -9132
rect 3913 -9388 3925 -9132
rect 3867 -9400 3925 -9388
rect 4045 -9132 4103 -9120
rect 4045 -9388 4057 -9132
rect 4091 -9388 4103 -9132
rect 6500 -9150 6512 -8894
rect 6546 -9150 6558 -8894
rect 6500 -9162 6558 -9150
rect 6678 -8894 6736 -8882
rect 6678 -9150 6690 -8894
rect 6724 -9150 6736 -8894
rect 6678 -9162 6736 -9150
rect 6856 -8894 6914 -8882
rect 6856 -9150 6868 -8894
rect 6902 -9150 6914 -8894
rect 6856 -9162 6914 -9150
rect 7034 -8894 7092 -8882
rect 7034 -9150 7046 -8894
rect 7080 -9150 7092 -8894
rect 7034 -9162 7092 -9150
rect 7212 -8894 7270 -8882
rect 7212 -9150 7224 -8894
rect 7258 -9150 7270 -8894
rect 7212 -9162 7270 -9150
rect 7390 -8894 7448 -8882
rect 7390 -9150 7402 -8894
rect 7436 -9150 7448 -8894
rect 7390 -9162 7448 -9150
rect 7568 -8894 7626 -8882
rect 7568 -9150 7580 -8894
rect 7614 -9150 7626 -8894
rect 7568 -9162 7626 -9150
rect 7746 -8894 7804 -8882
rect 7746 -9150 7758 -8894
rect 7792 -9150 7804 -8894
rect 7746 -9162 7804 -9150
rect 7924 -8894 7982 -8882
rect 7924 -9150 7936 -8894
rect 7970 -9150 7982 -8894
rect 7924 -9162 7982 -9150
rect 8102 -8894 8160 -8882
rect 8102 -9150 8114 -8894
rect 8148 -9150 8160 -8894
rect 8102 -9162 8160 -9150
rect 8280 -8894 8338 -8882
rect 8280 -9150 8292 -8894
rect 8326 -9150 8338 -8894
rect 8280 -9162 8338 -9150
rect 8458 -8894 8516 -8882
rect 8458 -9150 8470 -8894
rect 8504 -9150 8516 -8894
rect 8458 -9162 8516 -9150
rect 8636 -8894 8694 -8882
rect 8636 -9150 8648 -8894
rect 8682 -9150 8694 -8894
rect 8636 -9162 8694 -9150
rect 8814 -8894 8872 -8882
rect 8814 -9150 8826 -8894
rect 8860 -9150 8872 -8894
rect 8814 -9162 8872 -9150
rect 8992 -8894 9050 -8882
rect 8992 -9150 9004 -8894
rect 9038 -9150 9050 -8894
rect 8992 -9162 9050 -9150
rect 9170 -8894 9228 -8882
rect 9170 -9150 9182 -8894
rect 9216 -9150 9228 -8894
rect 9170 -9162 9228 -9150
rect 9348 -8894 9406 -8882
rect 9348 -9150 9360 -8894
rect 9394 -9150 9406 -8894
rect 9348 -9162 9406 -9150
rect 10760 -8924 10818 -8912
rect 4045 -9400 4103 -9388
rect 10760 -9180 10772 -8924
rect 10806 -9180 10818 -8924
rect 10760 -9192 10818 -9180
rect 10938 -8924 10996 -8912
rect 10938 -9180 10950 -8924
rect 10984 -9180 10996 -8924
rect 10938 -9192 10996 -9180
rect 11052 -8924 11110 -8912
rect 11052 -9180 11064 -8924
rect 11098 -9180 11110 -8924
rect 11052 -9192 11110 -9180
rect 11230 -8924 11288 -8912
rect 11230 -9180 11242 -8924
rect 11276 -9180 11288 -8924
rect 11230 -9192 11288 -9180
rect 11344 -8924 11402 -8912
rect 11344 -9180 11356 -8924
rect 11390 -9180 11402 -8924
rect 11344 -9192 11402 -9180
rect 11522 -8924 11580 -8912
rect 11522 -9180 11534 -8924
rect 11568 -9180 11580 -8924
rect 11522 -9192 11580 -9180
rect 11636 -8924 11694 -8912
rect 11636 -9180 11648 -8924
rect 11682 -9180 11694 -8924
rect 11636 -9192 11694 -9180
rect 11814 -8924 11872 -8912
rect 11814 -9180 11826 -8924
rect 11860 -9180 11872 -8924
rect 11814 -9192 11872 -9180
rect 11928 -8924 11986 -8912
rect 11928 -9180 11940 -8924
rect 11974 -9180 11986 -8924
rect 11928 -9192 11986 -9180
rect 12106 -8924 12164 -8912
rect 12106 -9180 12118 -8924
rect 12152 -9180 12164 -8924
rect 12106 -9192 12164 -9180
rect 12220 -8924 12278 -8912
rect 12220 -9180 12232 -8924
rect 12266 -9180 12278 -8924
rect 12220 -9192 12278 -9180
rect 12398 -8924 12456 -8912
rect 12398 -9180 12410 -8924
rect 12444 -9180 12456 -8924
rect 12398 -9192 12456 -9180
rect 12512 -8924 12570 -8912
rect 12512 -9180 12524 -8924
rect 12558 -9180 12570 -8924
rect 12512 -9192 12570 -9180
rect 12690 -8924 12748 -8912
rect 12690 -9180 12702 -8924
rect 12736 -9180 12748 -8924
rect 12690 -9192 12748 -9180
rect -5640 -9524 -5582 -9512
rect -5640 -9780 -5628 -9524
rect -5594 -9780 -5582 -9524
rect -5640 -9792 -5582 -9780
rect -5462 -9524 -5404 -9512
rect -5462 -9780 -5450 -9524
rect -5416 -9780 -5404 -9524
rect -5462 -9792 -5404 -9780
rect -5284 -9524 -5226 -9512
rect -5284 -9780 -5272 -9524
rect -5238 -9780 -5226 -9524
rect -5284 -9792 -5226 -9780
rect -5106 -9524 -5048 -9512
rect -5106 -9780 -5094 -9524
rect -5060 -9780 -5048 -9524
rect -5106 -9792 -5048 -9780
rect -4928 -9524 -4870 -9512
rect -4928 -9780 -4916 -9524
rect -4882 -9780 -4870 -9524
rect -4928 -9792 -4870 -9780
rect -4750 -9524 -4692 -9512
rect -4750 -9780 -4738 -9524
rect -4704 -9780 -4692 -9524
rect -4750 -9792 -4692 -9780
rect -4572 -9524 -4514 -9512
rect -4572 -9780 -4560 -9524
rect -4526 -9780 -4514 -9524
rect -4572 -9792 -4514 -9780
rect -4394 -9524 -4336 -9512
rect -4394 -9780 -4382 -9524
rect -4348 -9780 -4336 -9524
rect -4394 -9792 -4336 -9780
rect -4216 -9524 -4158 -9512
rect -4216 -9780 -4204 -9524
rect -4170 -9780 -4158 -9524
rect -4216 -9792 -4158 -9780
rect -4038 -9524 -3980 -9512
rect -4038 -9780 -4026 -9524
rect -3992 -9780 -3980 -9524
rect 10760 -9694 10818 -9682
rect -4038 -9792 -3980 -9780
rect 6500 -9794 6558 -9782
rect -5640 -10074 -5582 -10062
rect -5640 -10330 -5628 -10074
rect -5594 -10330 -5582 -10074
rect -5640 -10342 -5582 -10330
rect -5462 -10074 -5404 -10062
rect -5462 -10330 -5450 -10074
rect -5416 -10330 -5404 -10074
rect -5462 -10342 -5404 -10330
rect -5284 -10074 -5226 -10062
rect -5284 -10330 -5272 -10074
rect -5238 -10330 -5226 -10074
rect -5284 -10342 -5226 -10330
rect -5106 -10074 -5048 -10062
rect -5106 -10330 -5094 -10074
rect -5060 -10330 -5048 -10074
rect -5106 -10342 -5048 -10330
rect -4928 -10074 -4870 -10062
rect -4928 -10330 -4916 -10074
rect -4882 -10330 -4870 -10074
rect -4928 -10342 -4870 -10330
rect -4750 -10074 -4692 -10062
rect -4750 -10330 -4738 -10074
rect -4704 -10330 -4692 -10074
rect -4750 -10342 -4692 -10330
rect -4572 -10074 -4514 -10062
rect -4572 -10330 -4560 -10074
rect -4526 -10330 -4514 -10074
rect -4572 -10342 -4514 -10330
rect -4394 -10074 -4336 -10062
rect -4394 -10330 -4382 -10074
rect -4348 -10330 -4336 -10074
rect -4394 -10342 -4336 -10330
rect -4216 -10074 -4158 -10062
rect -4216 -10330 -4204 -10074
rect -4170 -10330 -4158 -10074
rect -4216 -10342 -4158 -10330
rect -4038 -10074 -3980 -10062
rect -4038 -10330 -4026 -10074
rect -3992 -10330 -3980 -10074
rect 6500 -10050 6512 -9794
rect 6546 -10050 6558 -9794
rect 6500 -10062 6558 -10050
rect 6678 -9794 6736 -9782
rect 6678 -10050 6690 -9794
rect 6724 -10050 6736 -9794
rect 6678 -10062 6736 -10050
rect 6856 -9794 6914 -9782
rect 6856 -10050 6868 -9794
rect 6902 -10050 6914 -9794
rect 6856 -10062 6914 -10050
rect 7034 -9794 7092 -9782
rect 7034 -10050 7046 -9794
rect 7080 -10050 7092 -9794
rect 7034 -10062 7092 -10050
rect 7212 -9794 7270 -9782
rect 7212 -10050 7224 -9794
rect 7258 -10050 7270 -9794
rect 7212 -10062 7270 -10050
rect 7390 -9794 7448 -9782
rect 7390 -10050 7402 -9794
rect 7436 -10050 7448 -9794
rect 7390 -10062 7448 -10050
rect 7568 -9794 7626 -9782
rect 7568 -10050 7580 -9794
rect 7614 -10050 7626 -9794
rect 7568 -10062 7626 -10050
rect 7746 -9794 7804 -9782
rect 7746 -10050 7758 -9794
rect 7792 -10050 7804 -9794
rect 7746 -10062 7804 -10050
rect 7924 -9794 7982 -9782
rect 7924 -10050 7936 -9794
rect 7970 -10050 7982 -9794
rect 7924 -10062 7982 -10050
rect 8102 -9794 8160 -9782
rect 8102 -10050 8114 -9794
rect 8148 -10050 8160 -9794
rect 8102 -10062 8160 -10050
rect 8280 -9794 8338 -9782
rect 8280 -10050 8292 -9794
rect 8326 -10050 8338 -9794
rect 8280 -10062 8338 -10050
rect 8458 -9794 8516 -9782
rect 8458 -10050 8470 -9794
rect 8504 -10050 8516 -9794
rect 8458 -10062 8516 -10050
rect 8636 -9794 8694 -9782
rect 8636 -10050 8648 -9794
rect 8682 -10050 8694 -9794
rect 8636 -10062 8694 -10050
rect 8814 -9794 8872 -9782
rect 8814 -10050 8826 -9794
rect 8860 -10050 8872 -9794
rect 8814 -10062 8872 -10050
rect 8992 -9794 9050 -9782
rect 8992 -10050 9004 -9794
rect 9038 -10050 9050 -9794
rect 8992 -10062 9050 -10050
rect 9170 -9794 9228 -9782
rect 9170 -10050 9182 -9794
rect 9216 -10050 9228 -9794
rect 9170 -10062 9228 -10050
rect 9348 -9794 9406 -9782
rect 9348 -10050 9360 -9794
rect 9394 -10050 9406 -9794
rect 10760 -9950 10772 -9694
rect 10806 -9950 10818 -9694
rect 10760 -9962 10818 -9950
rect 10938 -9694 10996 -9682
rect 10938 -9950 10950 -9694
rect 10984 -9950 10996 -9694
rect 10938 -9962 10996 -9950
rect 11052 -9694 11110 -9682
rect 11052 -9950 11064 -9694
rect 11098 -9950 11110 -9694
rect 11052 -9962 11110 -9950
rect 11230 -9694 11288 -9682
rect 11230 -9950 11242 -9694
rect 11276 -9950 11288 -9694
rect 11230 -9962 11288 -9950
rect 11344 -9694 11402 -9682
rect 11344 -9950 11356 -9694
rect 11390 -9950 11402 -9694
rect 11344 -9962 11402 -9950
rect 11522 -9694 11580 -9682
rect 11522 -9950 11534 -9694
rect 11568 -9950 11580 -9694
rect 11522 -9962 11580 -9950
rect 11636 -9694 11694 -9682
rect 11636 -9950 11648 -9694
rect 11682 -9950 11694 -9694
rect 11636 -9962 11694 -9950
rect 11814 -9694 11872 -9682
rect 11814 -9950 11826 -9694
rect 11860 -9950 11872 -9694
rect 11814 -9962 11872 -9950
rect 11928 -9694 11986 -9682
rect 11928 -9950 11940 -9694
rect 11974 -9950 11986 -9694
rect 11928 -9962 11986 -9950
rect 12106 -9694 12164 -9682
rect 12106 -9950 12118 -9694
rect 12152 -9950 12164 -9694
rect 12106 -9962 12164 -9950
rect 12220 -9694 12278 -9682
rect 12220 -9950 12232 -9694
rect 12266 -9950 12278 -9694
rect 12220 -9962 12278 -9950
rect 12398 -9694 12456 -9682
rect 12398 -9950 12410 -9694
rect 12444 -9950 12456 -9694
rect 12398 -9962 12456 -9950
rect 12512 -9694 12570 -9682
rect 12512 -9950 12524 -9694
rect 12558 -9950 12570 -9694
rect 12512 -9962 12570 -9950
rect 12690 -9694 12748 -9682
rect 12690 -9950 12702 -9694
rect 12736 -9950 12748 -9694
rect 12690 -9962 12748 -9950
rect 9348 -10062 9406 -10050
rect -4038 -10342 -3980 -10330
rect -2185 -10132 -2127 -10120
rect -2185 -10388 -2173 -10132
rect -2139 -10388 -2127 -10132
rect -2185 -10400 -2127 -10388
rect -2007 -10132 -1949 -10120
rect -2007 -10388 -1995 -10132
rect -1961 -10388 -1949 -10132
rect -2007 -10400 -1949 -10388
rect -1829 -10132 -1771 -10120
rect -1829 -10388 -1817 -10132
rect -1783 -10388 -1771 -10132
rect -1829 -10400 -1771 -10388
rect -1651 -10132 -1593 -10120
rect -1651 -10388 -1639 -10132
rect -1605 -10388 -1593 -10132
rect -1651 -10400 -1593 -10388
rect -1473 -10132 -1415 -10120
rect -1473 -10388 -1461 -10132
rect -1427 -10388 -1415 -10132
rect -1473 -10400 -1415 -10388
rect -1295 -10132 -1237 -10120
rect -1295 -10388 -1283 -10132
rect -1249 -10388 -1237 -10132
rect -1295 -10400 -1237 -10388
rect -1117 -10132 -1059 -10120
rect -1117 -10388 -1105 -10132
rect -1071 -10388 -1059 -10132
rect -1117 -10400 -1059 -10388
rect -939 -10132 -881 -10120
rect -939 -10388 -927 -10132
rect -893 -10388 -881 -10132
rect -939 -10400 -881 -10388
rect -761 -10132 -703 -10120
rect -761 -10388 -749 -10132
rect -715 -10388 -703 -10132
rect -761 -10400 -703 -10388
rect -583 -10132 -525 -10120
rect -583 -10388 -571 -10132
rect -537 -10388 -525 -10132
rect -583 -10400 -525 -10388
rect -405 -10132 -347 -10120
rect -405 -10388 -393 -10132
rect -359 -10388 -347 -10132
rect -405 -10400 -347 -10388
rect -227 -10132 -169 -10120
rect -227 -10388 -215 -10132
rect -181 -10388 -169 -10132
rect -227 -10400 -169 -10388
rect -49 -10132 9 -10120
rect -49 -10388 -37 -10132
rect -3 -10388 9 -10132
rect -49 -10400 9 -10388
rect 129 -10132 187 -10120
rect 129 -10388 141 -10132
rect 175 -10388 187 -10132
rect 129 -10400 187 -10388
rect 307 -10132 365 -10120
rect 307 -10388 319 -10132
rect 353 -10388 365 -10132
rect 307 -10400 365 -10388
rect 485 -10132 543 -10120
rect 485 -10388 497 -10132
rect 531 -10388 543 -10132
rect 485 -10400 543 -10388
rect 663 -10132 721 -10120
rect 663 -10388 675 -10132
rect 709 -10388 721 -10132
rect 663 -10400 721 -10388
rect 841 -10132 899 -10120
rect 841 -10388 853 -10132
rect 887 -10388 899 -10132
rect 841 -10400 899 -10388
rect 1019 -10132 1077 -10120
rect 1019 -10388 1031 -10132
rect 1065 -10388 1077 -10132
rect 1019 -10400 1077 -10388
rect 1197 -10132 1255 -10120
rect 1197 -10388 1209 -10132
rect 1243 -10388 1255 -10132
rect 1197 -10400 1255 -10388
rect 1375 -10132 1433 -10120
rect 1375 -10388 1387 -10132
rect 1421 -10388 1433 -10132
rect 1375 -10400 1433 -10388
rect 1553 -10132 1611 -10120
rect 1553 -10388 1565 -10132
rect 1599 -10388 1611 -10132
rect 1553 -10400 1611 -10388
rect 1731 -10132 1789 -10120
rect 1731 -10388 1743 -10132
rect 1777 -10388 1789 -10132
rect 1731 -10400 1789 -10388
rect 1909 -10132 1967 -10120
rect 1909 -10388 1921 -10132
rect 1955 -10388 1967 -10132
rect 1909 -10400 1967 -10388
rect 2087 -10132 2145 -10120
rect 2087 -10388 2099 -10132
rect 2133 -10388 2145 -10132
rect 2087 -10400 2145 -10388
rect 2265 -10132 2323 -10120
rect 2265 -10388 2277 -10132
rect 2311 -10388 2323 -10132
rect 2265 -10400 2323 -10388
rect 2443 -10132 2501 -10120
rect 2443 -10388 2455 -10132
rect 2489 -10388 2501 -10132
rect 2443 -10400 2501 -10388
rect 2621 -10132 2679 -10120
rect 2621 -10388 2633 -10132
rect 2667 -10388 2679 -10132
rect 2621 -10400 2679 -10388
rect 2799 -10132 2857 -10120
rect 2799 -10388 2811 -10132
rect 2845 -10388 2857 -10132
rect 2799 -10400 2857 -10388
rect 2977 -10132 3035 -10120
rect 2977 -10388 2989 -10132
rect 3023 -10388 3035 -10132
rect 2977 -10400 3035 -10388
rect 3155 -10132 3213 -10120
rect 3155 -10388 3167 -10132
rect 3201 -10388 3213 -10132
rect 3155 -10400 3213 -10388
rect 3333 -10132 3391 -10120
rect 3333 -10388 3345 -10132
rect 3379 -10388 3391 -10132
rect 3333 -10400 3391 -10388
rect 3511 -10132 3569 -10120
rect 3511 -10388 3523 -10132
rect 3557 -10388 3569 -10132
rect 3511 -10400 3569 -10388
rect 3689 -10132 3747 -10120
rect 3689 -10388 3701 -10132
rect 3735 -10388 3747 -10132
rect 3689 -10400 3747 -10388
rect 3867 -10132 3925 -10120
rect 3867 -10388 3879 -10132
rect 3913 -10388 3925 -10132
rect 3867 -10400 3925 -10388
rect 4045 -10132 4103 -10120
rect 4045 -10388 4057 -10132
rect 4091 -10388 4103 -10132
rect 4045 -10400 4103 -10388
rect 10760 -10464 10818 -10452
rect -5640 -10624 -5582 -10612
rect -5640 -10880 -5628 -10624
rect -5594 -10880 -5582 -10624
rect -5640 -10892 -5582 -10880
rect -5462 -10624 -5404 -10612
rect -5462 -10880 -5450 -10624
rect -5416 -10880 -5404 -10624
rect -5462 -10892 -5404 -10880
rect -5284 -10624 -5226 -10612
rect -5284 -10880 -5272 -10624
rect -5238 -10880 -5226 -10624
rect -5284 -10892 -5226 -10880
rect -5106 -10624 -5048 -10612
rect -5106 -10880 -5094 -10624
rect -5060 -10880 -5048 -10624
rect -5106 -10892 -5048 -10880
rect -4928 -10624 -4870 -10612
rect -4928 -10880 -4916 -10624
rect -4882 -10880 -4870 -10624
rect -4928 -10892 -4870 -10880
rect -4750 -10624 -4692 -10612
rect -4750 -10880 -4738 -10624
rect -4704 -10880 -4692 -10624
rect -4750 -10892 -4692 -10880
rect -4572 -10624 -4514 -10612
rect -4572 -10880 -4560 -10624
rect -4526 -10880 -4514 -10624
rect -4572 -10892 -4514 -10880
rect -4394 -10624 -4336 -10612
rect -4394 -10880 -4382 -10624
rect -4348 -10880 -4336 -10624
rect -4394 -10892 -4336 -10880
rect -4216 -10624 -4158 -10612
rect -4216 -10880 -4204 -10624
rect -4170 -10880 -4158 -10624
rect -4216 -10892 -4158 -10880
rect -4038 -10624 -3980 -10612
rect -4038 -10880 -4026 -10624
rect -3992 -10880 -3980 -10624
rect -4038 -10892 -3980 -10880
rect 6500 -10694 6558 -10682
rect 6500 -10950 6512 -10694
rect 6546 -10950 6558 -10694
rect 6500 -10962 6558 -10950
rect 6678 -10694 6736 -10682
rect 6678 -10950 6690 -10694
rect 6724 -10950 6736 -10694
rect 6678 -10962 6736 -10950
rect 6856 -10694 6914 -10682
rect 6856 -10950 6868 -10694
rect 6902 -10950 6914 -10694
rect 6856 -10962 6914 -10950
rect 7034 -10694 7092 -10682
rect 7034 -10950 7046 -10694
rect 7080 -10950 7092 -10694
rect 7034 -10962 7092 -10950
rect 7212 -10694 7270 -10682
rect 7212 -10950 7224 -10694
rect 7258 -10950 7270 -10694
rect 7212 -10962 7270 -10950
rect 7390 -10694 7448 -10682
rect 7390 -10950 7402 -10694
rect 7436 -10950 7448 -10694
rect 7390 -10962 7448 -10950
rect 7568 -10694 7626 -10682
rect 7568 -10950 7580 -10694
rect 7614 -10950 7626 -10694
rect 7568 -10962 7626 -10950
rect 7746 -10694 7804 -10682
rect 7746 -10950 7758 -10694
rect 7792 -10950 7804 -10694
rect 7746 -10962 7804 -10950
rect 7924 -10694 7982 -10682
rect 7924 -10950 7936 -10694
rect 7970 -10950 7982 -10694
rect 7924 -10962 7982 -10950
rect 8102 -10694 8160 -10682
rect 8102 -10950 8114 -10694
rect 8148 -10950 8160 -10694
rect 8102 -10962 8160 -10950
rect 8280 -10694 8338 -10682
rect 8280 -10950 8292 -10694
rect 8326 -10950 8338 -10694
rect 8280 -10962 8338 -10950
rect 8458 -10694 8516 -10682
rect 8458 -10950 8470 -10694
rect 8504 -10950 8516 -10694
rect 8458 -10962 8516 -10950
rect 8636 -10694 8694 -10682
rect 8636 -10950 8648 -10694
rect 8682 -10950 8694 -10694
rect 8636 -10962 8694 -10950
rect 8814 -10694 8872 -10682
rect 8814 -10950 8826 -10694
rect 8860 -10950 8872 -10694
rect 8814 -10962 8872 -10950
rect 8992 -10694 9050 -10682
rect 8992 -10950 9004 -10694
rect 9038 -10950 9050 -10694
rect 8992 -10962 9050 -10950
rect 9170 -10694 9228 -10682
rect 9170 -10950 9182 -10694
rect 9216 -10950 9228 -10694
rect 9170 -10962 9228 -10950
rect 9348 -10694 9406 -10682
rect 9348 -10950 9360 -10694
rect 9394 -10950 9406 -10694
rect 10760 -10720 10772 -10464
rect 10806 -10720 10818 -10464
rect 10760 -10732 10818 -10720
rect 10938 -10464 10996 -10452
rect 10938 -10720 10950 -10464
rect 10984 -10720 10996 -10464
rect 10938 -10732 10996 -10720
rect 11052 -10464 11110 -10452
rect 11052 -10720 11064 -10464
rect 11098 -10720 11110 -10464
rect 11052 -10732 11110 -10720
rect 11230 -10464 11288 -10452
rect 11230 -10720 11242 -10464
rect 11276 -10720 11288 -10464
rect 11230 -10732 11288 -10720
rect 11344 -10464 11402 -10452
rect 11344 -10720 11356 -10464
rect 11390 -10720 11402 -10464
rect 11344 -10732 11402 -10720
rect 11522 -10464 11580 -10452
rect 11522 -10720 11534 -10464
rect 11568 -10720 11580 -10464
rect 11522 -10732 11580 -10720
rect 11636 -10464 11694 -10452
rect 11636 -10720 11648 -10464
rect 11682 -10720 11694 -10464
rect 11636 -10732 11694 -10720
rect 11814 -10464 11872 -10452
rect 11814 -10720 11826 -10464
rect 11860 -10720 11872 -10464
rect 11814 -10732 11872 -10720
rect 11928 -10464 11986 -10452
rect 11928 -10720 11940 -10464
rect 11974 -10720 11986 -10464
rect 11928 -10732 11986 -10720
rect 12106 -10464 12164 -10452
rect 12106 -10720 12118 -10464
rect 12152 -10720 12164 -10464
rect 12106 -10732 12164 -10720
rect 12220 -10464 12278 -10452
rect 12220 -10720 12232 -10464
rect 12266 -10720 12278 -10464
rect 12220 -10732 12278 -10720
rect 12398 -10464 12456 -10452
rect 12398 -10720 12410 -10464
rect 12444 -10720 12456 -10464
rect 12398 -10732 12456 -10720
rect 12512 -10464 12570 -10452
rect 12512 -10720 12524 -10464
rect 12558 -10720 12570 -10464
rect 12512 -10732 12570 -10720
rect 12690 -10464 12748 -10452
rect 12690 -10720 12702 -10464
rect 12736 -10720 12748 -10464
rect 12690 -10732 12748 -10720
rect 9348 -10962 9406 -10950
rect -2185 -11132 -2127 -11120
rect -5640 -11174 -5582 -11162
rect -5640 -11430 -5628 -11174
rect -5594 -11430 -5582 -11174
rect -5640 -11442 -5582 -11430
rect -5462 -11174 -5404 -11162
rect -5462 -11430 -5450 -11174
rect -5416 -11430 -5404 -11174
rect -5462 -11442 -5404 -11430
rect -5284 -11174 -5226 -11162
rect -5284 -11430 -5272 -11174
rect -5238 -11430 -5226 -11174
rect -5284 -11442 -5226 -11430
rect -5106 -11174 -5048 -11162
rect -5106 -11430 -5094 -11174
rect -5060 -11430 -5048 -11174
rect -5106 -11442 -5048 -11430
rect -4928 -11174 -4870 -11162
rect -4928 -11430 -4916 -11174
rect -4882 -11430 -4870 -11174
rect -4928 -11442 -4870 -11430
rect -4750 -11174 -4692 -11162
rect -4750 -11430 -4738 -11174
rect -4704 -11430 -4692 -11174
rect -4750 -11442 -4692 -11430
rect -4572 -11174 -4514 -11162
rect -4572 -11430 -4560 -11174
rect -4526 -11430 -4514 -11174
rect -4572 -11442 -4514 -11430
rect -4394 -11174 -4336 -11162
rect -4394 -11430 -4382 -11174
rect -4348 -11430 -4336 -11174
rect -4394 -11442 -4336 -11430
rect -4216 -11174 -4158 -11162
rect -4216 -11430 -4204 -11174
rect -4170 -11430 -4158 -11174
rect -4216 -11442 -4158 -11430
rect -4038 -11174 -3980 -11162
rect -4038 -11430 -4026 -11174
rect -3992 -11430 -3980 -11174
rect -4038 -11442 -3980 -11430
rect -2185 -11388 -2173 -11132
rect -2139 -11388 -2127 -11132
rect -2185 -11400 -2127 -11388
rect -2007 -11132 -1949 -11120
rect -2007 -11388 -1995 -11132
rect -1961 -11388 -1949 -11132
rect -2007 -11400 -1949 -11388
rect -1829 -11132 -1771 -11120
rect -1829 -11388 -1817 -11132
rect -1783 -11388 -1771 -11132
rect -1829 -11400 -1771 -11388
rect -1651 -11132 -1593 -11120
rect -1651 -11388 -1639 -11132
rect -1605 -11388 -1593 -11132
rect -1651 -11400 -1593 -11388
rect -1473 -11132 -1415 -11120
rect -1473 -11388 -1461 -11132
rect -1427 -11388 -1415 -11132
rect -1473 -11400 -1415 -11388
rect -1295 -11132 -1237 -11120
rect -1295 -11388 -1283 -11132
rect -1249 -11388 -1237 -11132
rect -1295 -11400 -1237 -11388
rect -1117 -11132 -1059 -11120
rect -1117 -11388 -1105 -11132
rect -1071 -11388 -1059 -11132
rect -1117 -11400 -1059 -11388
rect -939 -11132 -881 -11120
rect -939 -11388 -927 -11132
rect -893 -11388 -881 -11132
rect -939 -11400 -881 -11388
rect -761 -11132 -703 -11120
rect -761 -11388 -749 -11132
rect -715 -11388 -703 -11132
rect -761 -11400 -703 -11388
rect -583 -11132 -525 -11120
rect -583 -11388 -571 -11132
rect -537 -11388 -525 -11132
rect -583 -11400 -525 -11388
rect -405 -11132 -347 -11120
rect -405 -11388 -393 -11132
rect -359 -11388 -347 -11132
rect -405 -11400 -347 -11388
rect -227 -11132 -169 -11120
rect -227 -11388 -215 -11132
rect -181 -11388 -169 -11132
rect -227 -11400 -169 -11388
rect -49 -11132 9 -11120
rect -49 -11388 -37 -11132
rect -3 -11388 9 -11132
rect -49 -11400 9 -11388
rect 129 -11132 187 -11120
rect 129 -11388 141 -11132
rect 175 -11388 187 -11132
rect 129 -11400 187 -11388
rect 307 -11132 365 -11120
rect 307 -11388 319 -11132
rect 353 -11388 365 -11132
rect 307 -11400 365 -11388
rect 485 -11132 543 -11120
rect 485 -11388 497 -11132
rect 531 -11388 543 -11132
rect 485 -11400 543 -11388
rect 663 -11132 721 -11120
rect 663 -11388 675 -11132
rect 709 -11388 721 -11132
rect 663 -11400 721 -11388
rect 841 -11132 899 -11120
rect 841 -11388 853 -11132
rect 887 -11388 899 -11132
rect 841 -11400 899 -11388
rect 1019 -11132 1077 -11120
rect 1019 -11388 1031 -11132
rect 1065 -11388 1077 -11132
rect 1019 -11400 1077 -11388
rect 1197 -11132 1255 -11120
rect 1197 -11388 1209 -11132
rect 1243 -11388 1255 -11132
rect 1197 -11400 1255 -11388
rect 1375 -11132 1433 -11120
rect 1375 -11388 1387 -11132
rect 1421 -11388 1433 -11132
rect 1375 -11400 1433 -11388
rect 1553 -11132 1611 -11120
rect 1553 -11388 1565 -11132
rect 1599 -11388 1611 -11132
rect 1553 -11400 1611 -11388
rect 1731 -11132 1789 -11120
rect 1731 -11388 1743 -11132
rect 1777 -11388 1789 -11132
rect 1731 -11400 1789 -11388
rect 1909 -11132 1967 -11120
rect 1909 -11388 1921 -11132
rect 1955 -11388 1967 -11132
rect 1909 -11400 1967 -11388
rect 2087 -11132 2145 -11120
rect 2087 -11388 2099 -11132
rect 2133 -11388 2145 -11132
rect 2087 -11400 2145 -11388
rect 2265 -11132 2323 -11120
rect 2265 -11388 2277 -11132
rect 2311 -11388 2323 -11132
rect 2265 -11400 2323 -11388
rect 2443 -11132 2501 -11120
rect 2443 -11388 2455 -11132
rect 2489 -11388 2501 -11132
rect 2443 -11400 2501 -11388
rect 2621 -11132 2679 -11120
rect 2621 -11388 2633 -11132
rect 2667 -11388 2679 -11132
rect 2621 -11400 2679 -11388
rect 2799 -11132 2857 -11120
rect 2799 -11388 2811 -11132
rect 2845 -11388 2857 -11132
rect 2799 -11400 2857 -11388
rect 2977 -11132 3035 -11120
rect 2977 -11388 2989 -11132
rect 3023 -11388 3035 -11132
rect 2977 -11400 3035 -11388
rect 3155 -11132 3213 -11120
rect 3155 -11388 3167 -11132
rect 3201 -11388 3213 -11132
rect 3155 -11400 3213 -11388
rect 3333 -11132 3391 -11120
rect 3333 -11388 3345 -11132
rect 3379 -11388 3391 -11132
rect 3333 -11400 3391 -11388
rect 3511 -11132 3569 -11120
rect 3511 -11388 3523 -11132
rect 3557 -11388 3569 -11132
rect 3511 -11400 3569 -11388
rect 3689 -11132 3747 -11120
rect 3689 -11388 3701 -11132
rect 3735 -11388 3747 -11132
rect 3689 -11400 3747 -11388
rect 3867 -11132 3925 -11120
rect 3867 -11388 3879 -11132
rect 3913 -11388 3925 -11132
rect 3867 -11400 3925 -11388
rect 4045 -11132 4103 -11120
rect 4045 -11388 4057 -11132
rect 4091 -11388 4103 -11132
rect 4045 -11400 4103 -11388
rect 10760 -11234 10818 -11222
rect 10760 -11490 10772 -11234
rect 10806 -11490 10818 -11234
rect 10760 -11502 10818 -11490
rect 10938 -11234 10996 -11222
rect 10938 -11490 10950 -11234
rect 10984 -11490 10996 -11234
rect 10938 -11502 10996 -11490
rect 11052 -11234 11110 -11222
rect 11052 -11490 11064 -11234
rect 11098 -11490 11110 -11234
rect 11052 -11502 11110 -11490
rect 11230 -11234 11288 -11222
rect 11230 -11490 11242 -11234
rect 11276 -11490 11288 -11234
rect 11230 -11502 11288 -11490
rect 11344 -11234 11402 -11222
rect 11344 -11490 11356 -11234
rect 11390 -11490 11402 -11234
rect 11344 -11502 11402 -11490
rect 11522 -11234 11580 -11222
rect 11522 -11490 11534 -11234
rect 11568 -11490 11580 -11234
rect 11522 -11502 11580 -11490
rect 11636 -11234 11694 -11222
rect 11636 -11490 11648 -11234
rect 11682 -11490 11694 -11234
rect 11636 -11502 11694 -11490
rect 11814 -11234 11872 -11222
rect 11814 -11490 11826 -11234
rect 11860 -11490 11872 -11234
rect 11814 -11502 11872 -11490
rect 11928 -11234 11986 -11222
rect 11928 -11490 11940 -11234
rect 11974 -11490 11986 -11234
rect 11928 -11502 11986 -11490
rect 12106 -11234 12164 -11222
rect 12106 -11490 12118 -11234
rect 12152 -11490 12164 -11234
rect 12106 -11502 12164 -11490
rect 12220 -11234 12278 -11222
rect 12220 -11490 12232 -11234
rect 12266 -11490 12278 -11234
rect 12220 -11502 12278 -11490
rect 12398 -11234 12456 -11222
rect 12398 -11490 12410 -11234
rect 12444 -11490 12456 -11234
rect 12398 -11502 12456 -11490
rect 12512 -11234 12570 -11222
rect 12512 -11490 12524 -11234
rect 12558 -11490 12570 -11234
rect 12512 -11502 12570 -11490
rect 12690 -11234 12748 -11222
rect 12690 -11490 12702 -11234
rect 12736 -11490 12748 -11234
rect 12690 -11502 12748 -11490
rect 6500 -11594 6558 -11582
rect -5640 -11724 -5582 -11712
rect -5640 -11980 -5628 -11724
rect -5594 -11980 -5582 -11724
rect -5640 -11992 -5582 -11980
rect -5462 -11724 -5404 -11712
rect -5462 -11980 -5450 -11724
rect -5416 -11980 -5404 -11724
rect -5462 -11992 -5404 -11980
rect -5284 -11724 -5226 -11712
rect -5284 -11980 -5272 -11724
rect -5238 -11980 -5226 -11724
rect -5284 -11992 -5226 -11980
rect -5106 -11724 -5048 -11712
rect -5106 -11980 -5094 -11724
rect -5060 -11980 -5048 -11724
rect -5106 -11992 -5048 -11980
rect -4928 -11724 -4870 -11712
rect -4928 -11980 -4916 -11724
rect -4882 -11980 -4870 -11724
rect -4928 -11992 -4870 -11980
rect -4750 -11724 -4692 -11712
rect -4750 -11980 -4738 -11724
rect -4704 -11980 -4692 -11724
rect -4750 -11992 -4692 -11980
rect -4572 -11724 -4514 -11712
rect -4572 -11980 -4560 -11724
rect -4526 -11980 -4514 -11724
rect -4572 -11992 -4514 -11980
rect -4394 -11724 -4336 -11712
rect -4394 -11980 -4382 -11724
rect -4348 -11980 -4336 -11724
rect -4394 -11992 -4336 -11980
rect -4216 -11724 -4158 -11712
rect -4216 -11980 -4204 -11724
rect -4170 -11980 -4158 -11724
rect -4216 -11992 -4158 -11980
rect -4038 -11724 -3980 -11712
rect -4038 -11980 -4026 -11724
rect -3992 -11980 -3980 -11724
rect 6500 -11850 6512 -11594
rect 6546 -11850 6558 -11594
rect 6500 -11862 6558 -11850
rect 6678 -11594 6736 -11582
rect 6678 -11850 6690 -11594
rect 6724 -11850 6736 -11594
rect 6678 -11862 6736 -11850
rect 6856 -11594 6914 -11582
rect 6856 -11850 6868 -11594
rect 6902 -11850 6914 -11594
rect 6856 -11862 6914 -11850
rect 7034 -11594 7092 -11582
rect 7034 -11850 7046 -11594
rect 7080 -11850 7092 -11594
rect 7034 -11862 7092 -11850
rect 7212 -11594 7270 -11582
rect 7212 -11850 7224 -11594
rect 7258 -11850 7270 -11594
rect 7212 -11862 7270 -11850
rect 7390 -11594 7448 -11582
rect 7390 -11850 7402 -11594
rect 7436 -11850 7448 -11594
rect 7390 -11862 7448 -11850
rect 7568 -11594 7626 -11582
rect 7568 -11850 7580 -11594
rect 7614 -11850 7626 -11594
rect 7568 -11862 7626 -11850
rect 7746 -11594 7804 -11582
rect 7746 -11850 7758 -11594
rect 7792 -11850 7804 -11594
rect 7746 -11862 7804 -11850
rect 7924 -11594 7982 -11582
rect 7924 -11850 7936 -11594
rect 7970 -11850 7982 -11594
rect 7924 -11862 7982 -11850
rect 8102 -11594 8160 -11582
rect 8102 -11850 8114 -11594
rect 8148 -11850 8160 -11594
rect 8102 -11862 8160 -11850
rect 8280 -11594 8338 -11582
rect 8280 -11850 8292 -11594
rect 8326 -11850 8338 -11594
rect 8280 -11862 8338 -11850
rect 8458 -11594 8516 -11582
rect 8458 -11850 8470 -11594
rect 8504 -11850 8516 -11594
rect 8458 -11862 8516 -11850
rect 8636 -11594 8694 -11582
rect 8636 -11850 8648 -11594
rect 8682 -11850 8694 -11594
rect 8636 -11862 8694 -11850
rect 8814 -11594 8872 -11582
rect 8814 -11850 8826 -11594
rect 8860 -11850 8872 -11594
rect 8814 -11862 8872 -11850
rect 8992 -11594 9050 -11582
rect 8992 -11850 9004 -11594
rect 9038 -11850 9050 -11594
rect 8992 -11862 9050 -11850
rect 9170 -11594 9228 -11582
rect 9170 -11850 9182 -11594
rect 9216 -11850 9228 -11594
rect 9170 -11862 9228 -11850
rect 9348 -11594 9406 -11582
rect 9348 -11850 9360 -11594
rect 9394 -11850 9406 -11594
rect 9348 -11862 9406 -11850
rect -4038 -11992 -3980 -11980
rect -2185 -12132 -2127 -12120
rect -2185 -12388 -2173 -12132
rect -2139 -12388 -2127 -12132
rect -2185 -12400 -2127 -12388
rect -2007 -12132 -1949 -12120
rect -2007 -12388 -1995 -12132
rect -1961 -12388 -1949 -12132
rect -2007 -12400 -1949 -12388
rect -1829 -12132 -1771 -12120
rect -1829 -12388 -1817 -12132
rect -1783 -12388 -1771 -12132
rect -1829 -12400 -1771 -12388
rect -1651 -12132 -1593 -12120
rect -1651 -12388 -1639 -12132
rect -1605 -12388 -1593 -12132
rect -1651 -12400 -1593 -12388
rect -1473 -12132 -1415 -12120
rect -1473 -12388 -1461 -12132
rect -1427 -12388 -1415 -12132
rect -1473 -12400 -1415 -12388
rect -1295 -12132 -1237 -12120
rect -1295 -12388 -1283 -12132
rect -1249 -12388 -1237 -12132
rect -1295 -12400 -1237 -12388
rect -1117 -12132 -1059 -12120
rect -1117 -12388 -1105 -12132
rect -1071 -12388 -1059 -12132
rect -1117 -12400 -1059 -12388
rect -939 -12132 -881 -12120
rect -939 -12388 -927 -12132
rect -893 -12388 -881 -12132
rect -939 -12400 -881 -12388
rect -761 -12132 -703 -12120
rect -761 -12388 -749 -12132
rect -715 -12388 -703 -12132
rect -761 -12400 -703 -12388
rect -583 -12132 -525 -12120
rect -583 -12388 -571 -12132
rect -537 -12388 -525 -12132
rect -583 -12400 -525 -12388
rect -405 -12132 -347 -12120
rect -405 -12388 -393 -12132
rect -359 -12388 -347 -12132
rect -405 -12400 -347 -12388
rect -227 -12132 -169 -12120
rect -227 -12388 -215 -12132
rect -181 -12388 -169 -12132
rect -227 -12400 -169 -12388
rect -49 -12132 9 -12120
rect -49 -12388 -37 -12132
rect -3 -12388 9 -12132
rect -49 -12400 9 -12388
rect 129 -12132 187 -12120
rect 129 -12388 141 -12132
rect 175 -12388 187 -12132
rect 129 -12400 187 -12388
rect 307 -12132 365 -12120
rect 307 -12388 319 -12132
rect 353 -12388 365 -12132
rect 307 -12400 365 -12388
rect 485 -12132 543 -12120
rect 485 -12388 497 -12132
rect 531 -12388 543 -12132
rect 485 -12400 543 -12388
rect 663 -12132 721 -12120
rect 663 -12388 675 -12132
rect 709 -12388 721 -12132
rect 663 -12400 721 -12388
rect 841 -12132 899 -12120
rect 841 -12388 853 -12132
rect 887 -12388 899 -12132
rect 841 -12400 899 -12388
rect 1019 -12132 1077 -12120
rect 1019 -12388 1031 -12132
rect 1065 -12388 1077 -12132
rect 1019 -12400 1077 -12388
rect 1197 -12132 1255 -12120
rect 1197 -12388 1209 -12132
rect 1243 -12388 1255 -12132
rect 1197 -12400 1255 -12388
rect 1375 -12132 1433 -12120
rect 1375 -12388 1387 -12132
rect 1421 -12388 1433 -12132
rect 1375 -12400 1433 -12388
rect 1553 -12132 1611 -12120
rect 1553 -12388 1565 -12132
rect 1599 -12388 1611 -12132
rect 1553 -12400 1611 -12388
rect 1731 -12132 1789 -12120
rect 1731 -12388 1743 -12132
rect 1777 -12388 1789 -12132
rect 1731 -12400 1789 -12388
rect 1909 -12132 1967 -12120
rect 1909 -12388 1921 -12132
rect 1955 -12388 1967 -12132
rect 1909 -12400 1967 -12388
rect 2087 -12132 2145 -12120
rect 2087 -12388 2099 -12132
rect 2133 -12388 2145 -12132
rect 2087 -12400 2145 -12388
rect 2265 -12132 2323 -12120
rect 2265 -12388 2277 -12132
rect 2311 -12388 2323 -12132
rect 2265 -12400 2323 -12388
rect 2443 -12132 2501 -12120
rect 2443 -12388 2455 -12132
rect 2489 -12388 2501 -12132
rect 2443 -12400 2501 -12388
rect 2621 -12132 2679 -12120
rect 2621 -12388 2633 -12132
rect 2667 -12388 2679 -12132
rect 2621 -12400 2679 -12388
rect 2799 -12132 2857 -12120
rect 2799 -12388 2811 -12132
rect 2845 -12388 2857 -12132
rect 2799 -12400 2857 -12388
rect 2977 -12132 3035 -12120
rect 2977 -12388 2989 -12132
rect 3023 -12388 3035 -12132
rect 2977 -12400 3035 -12388
rect 3155 -12132 3213 -12120
rect 3155 -12388 3167 -12132
rect 3201 -12388 3213 -12132
rect 3155 -12400 3213 -12388
rect 3333 -12132 3391 -12120
rect 3333 -12388 3345 -12132
rect 3379 -12388 3391 -12132
rect 3333 -12400 3391 -12388
rect 3511 -12132 3569 -12120
rect 3511 -12388 3523 -12132
rect 3557 -12388 3569 -12132
rect 3511 -12400 3569 -12388
rect 3689 -12132 3747 -12120
rect 3689 -12388 3701 -12132
rect 3735 -12388 3747 -12132
rect 3689 -12400 3747 -12388
rect 3867 -12132 3925 -12120
rect 3867 -12388 3879 -12132
rect 3913 -12388 3925 -12132
rect 3867 -12400 3925 -12388
rect 4045 -12132 4103 -12120
rect 4045 -12388 4057 -12132
rect 4091 -12388 4103 -12132
rect 4045 -12400 4103 -12388
rect -5929 -12712 -5871 -12700
rect -5929 -12928 -5917 -12712
rect -5883 -12928 -5871 -12712
rect -5929 -12940 -5871 -12928
rect -5829 -12712 -5771 -12700
rect -5829 -12928 -5817 -12712
rect -5783 -12928 -5771 -12712
rect -5829 -12940 -5771 -12928
rect -5679 -12712 -5621 -12700
rect -5679 -12928 -5667 -12712
rect -5633 -12928 -5621 -12712
rect -5679 -12940 -5621 -12928
rect -5579 -12712 -5521 -12700
rect -5579 -12928 -5567 -12712
rect -5533 -12928 -5521 -12712
rect -5579 -12940 -5521 -12928
rect -5429 -12712 -5371 -12700
rect -5429 -12928 -5417 -12712
rect -5383 -12928 -5371 -12712
rect -5429 -12940 -5371 -12928
rect -5329 -12712 -5271 -12700
rect -5329 -12928 -5317 -12712
rect -5283 -12928 -5271 -12712
rect -5329 -12940 -5271 -12928
rect -5179 -12712 -5121 -12700
rect -5179 -12928 -5167 -12712
rect -5133 -12928 -5121 -12712
rect -5179 -12940 -5121 -12928
rect -5079 -12712 -5021 -12700
rect -5079 -12928 -5067 -12712
rect -5033 -12928 -5021 -12712
rect -5079 -12940 -5021 -12928
rect -4929 -12712 -4871 -12700
rect -4929 -12928 -4917 -12712
rect -4883 -12928 -4871 -12712
rect -4929 -12940 -4871 -12928
rect -4829 -12712 -4771 -12700
rect -4829 -12928 -4817 -12712
rect -4783 -12928 -4771 -12712
rect -4829 -12940 -4771 -12928
rect -4679 -12712 -4621 -12700
rect -4679 -12928 -4667 -12712
rect -4633 -12928 -4621 -12712
rect -4679 -12940 -4621 -12928
rect -4579 -12712 -4521 -12700
rect -4579 -12928 -4567 -12712
rect -4533 -12928 -4521 -12712
rect -4579 -12940 -4521 -12928
rect -4429 -12712 -4371 -12700
rect -4429 -12928 -4417 -12712
rect -4383 -12928 -4371 -12712
rect -4429 -12940 -4371 -12928
rect -4329 -12712 -4271 -12700
rect -4329 -12928 -4317 -12712
rect -4283 -12928 -4271 -12712
rect -4329 -12940 -4271 -12928
rect -4179 -12712 -4121 -12700
rect -4179 -12928 -4167 -12712
rect -4133 -12928 -4121 -12712
rect -4179 -12940 -4121 -12928
rect -4079 -12712 -4021 -12700
rect -4079 -12928 -4067 -12712
rect -4033 -12928 -4021 -12712
rect -4079 -12940 -4021 -12928
rect -2185 -13132 -2127 -13120
rect -5929 -13392 -5871 -13380
rect -5929 -13608 -5917 -13392
rect -5883 -13608 -5871 -13392
rect -5929 -13620 -5871 -13608
rect -5829 -13392 -5771 -13380
rect -5829 -13608 -5817 -13392
rect -5783 -13608 -5771 -13392
rect -5829 -13620 -5771 -13608
rect -5679 -13392 -5621 -13380
rect -5679 -13608 -5667 -13392
rect -5633 -13608 -5621 -13392
rect -5679 -13620 -5621 -13608
rect -5579 -13392 -5521 -13380
rect -5579 -13608 -5567 -13392
rect -5533 -13608 -5521 -13392
rect -5579 -13620 -5521 -13608
rect -5429 -13392 -5371 -13380
rect -5429 -13608 -5417 -13392
rect -5383 -13608 -5371 -13392
rect -5429 -13620 -5371 -13608
rect -5329 -13392 -5271 -13380
rect -5329 -13608 -5317 -13392
rect -5283 -13608 -5271 -13392
rect -5329 -13620 -5271 -13608
rect -5179 -13392 -5121 -13380
rect -5179 -13608 -5167 -13392
rect -5133 -13608 -5121 -13392
rect -5179 -13620 -5121 -13608
rect -5079 -13392 -5021 -13380
rect -5079 -13608 -5067 -13392
rect -5033 -13608 -5021 -13392
rect -5079 -13620 -5021 -13608
rect -4929 -13392 -4871 -13380
rect -4929 -13608 -4917 -13392
rect -4883 -13608 -4871 -13392
rect -4929 -13620 -4871 -13608
rect -4829 -13392 -4771 -13380
rect -4829 -13608 -4817 -13392
rect -4783 -13608 -4771 -13392
rect -4829 -13620 -4771 -13608
rect -4679 -13392 -4621 -13380
rect -4679 -13608 -4667 -13392
rect -4633 -13608 -4621 -13392
rect -4679 -13620 -4621 -13608
rect -4579 -13392 -4521 -13380
rect -4579 -13608 -4567 -13392
rect -4533 -13608 -4521 -13392
rect -4579 -13620 -4521 -13608
rect -4429 -13392 -4371 -13380
rect -4429 -13608 -4417 -13392
rect -4383 -13608 -4371 -13392
rect -4429 -13620 -4371 -13608
rect -4329 -13392 -4271 -13380
rect -4329 -13608 -4317 -13392
rect -4283 -13608 -4271 -13392
rect -4329 -13620 -4271 -13608
rect -4179 -13392 -4121 -13380
rect -4179 -13608 -4167 -13392
rect -4133 -13608 -4121 -13392
rect -4179 -13620 -4121 -13608
rect -4079 -13392 -4021 -13380
rect -4079 -13608 -4067 -13392
rect -4033 -13608 -4021 -13392
rect -2185 -13388 -2173 -13132
rect -2139 -13388 -2127 -13132
rect -2185 -13400 -2127 -13388
rect -2007 -13132 -1949 -13120
rect -2007 -13388 -1995 -13132
rect -1961 -13388 -1949 -13132
rect -2007 -13400 -1949 -13388
rect -1829 -13132 -1771 -13120
rect -1829 -13388 -1817 -13132
rect -1783 -13388 -1771 -13132
rect -1829 -13400 -1771 -13388
rect -1651 -13132 -1593 -13120
rect -1651 -13388 -1639 -13132
rect -1605 -13388 -1593 -13132
rect -1651 -13400 -1593 -13388
rect -1473 -13132 -1415 -13120
rect -1473 -13388 -1461 -13132
rect -1427 -13388 -1415 -13132
rect -1473 -13400 -1415 -13388
rect -1295 -13132 -1237 -13120
rect -1295 -13388 -1283 -13132
rect -1249 -13388 -1237 -13132
rect -1295 -13400 -1237 -13388
rect -1117 -13132 -1059 -13120
rect -1117 -13388 -1105 -13132
rect -1071 -13388 -1059 -13132
rect -1117 -13400 -1059 -13388
rect -939 -13132 -881 -13120
rect -939 -13388 -927 -13132
rect -893 -13388 -881 -13132
rect -939 -13400 -881 -13388
rect -761 -13132 -703 -13120
rect -761 -13388 -749 -13132
rect -715 -13388 -703 -13132
rect -761 -13400 -703 -13388
rect -583 -13132 -525 -13120
rect -583 -13388 -571 -13132
rect -537 -13388 -525 -13132
rect -583 -13400 -525 -13388
rect -405 -13132 -347 -13120
rect -405 -13388 -393 -13132
rect -359 -13388 -347 -13132
rect -405 -13400 -347 -13388
rect -227 -13132 -169 -13120
rect -227 -13388 -215 -13132
rect -181 -13388 -169 -13132
rect -227 -13400 -169 -13388
rect -49 -13132 9 -13120
rect -49 -13388 -37 -13132
rect -3 -13388 9 -13132
rect -49 -13400 9 -13388
rect 129 -13132 187 -13120
rect 129 -13388 141 -13132
rect 175 -13388 187 -13132
rect 129 -13400 187 -13388
rect 307 -13132 365 -13120
rect 307 -13388 319 -13132
rect 353 -13388 365 -13132
rect 307 -13400 365 -13388
rect 485 -13132 543 -13120
rect 485 -13388 497 -13132
rect 531 -13388 543 -13132
rect 485 -13400 543 -13388
rect 663 -13132 721 -13120
rect 663 -13388 675 -13132
rect 709 -13388 721 -13132
rect 663 -13400 721 -13388
rect 841 -13132 899 -13120
rect 841 -13388 853 -13132
rect 887 -13388 899 -13132
rect 841 -13400 899 -13388
rect 1019 -13132 1077 -13120
rect 1019 -13388 1031 -13132
rect 1065 -13388 1077 -13132
rect 1019 -13400 1077 -13388
rect 1197 -13132 1255 -13120
rect 1197 -13388 1209 -13132
rect 1243 -13388 1255 -13132
rect 1197 -13400 1255 -13388
rect 1375 -13132 1433 -13120
rect 1375 -13388 1387 -13132
rect 1421 -13388 1433 -13132
rect 1375 -13400 1433 -13388
rect 1553 -13132 1611 -13120
rect 1553 -13388 1565 -13132
rect 1599 -13388 1611 -13132
rect 1553 -13400 1611 -13388
rect 1731 -13132 1789 -13120
rect 1731 -13388 1743 -13132
rect 1777 -13388 1789 -13132
rect 1731 -13400 1789 -13388
rect 1909 -13132 1967 -13120
rect 1909 -13388 1921 -13132
rect 1955 -13388 1967 -13132
rect 1909 -13400 1967 -13388
rect 2087 -13132 2145 -13120
rect 2087 -13388 2099 -13132
rect 2133 -13388 2145 -13132
rect 2087 -13400 2145 -13388
rect 2265 -13132 2323 -13120
rect 2265 -13388 2277 -13132
rect 2311 -13388 2323 -13132
rect 2265 -13400 2323 -13388
rect 2443 -13132 2501 -13120
rect 2443 -13388 2455 -13132
rect 2489 -13388 2501 -13132
rect 2443 -13400 2501 -13388
rect 2621 -13132 2679 -13120
rect 2621 -13388 2633 -13132
rect 2667 -13388 2679 -13132
rect 2621 -13400 2679 -13388
rect 2799 -13132 2857 -13120
rect 2799 -13388 2811 -13132
rect 2845 -13388 2857 -13132
rect 2799 -13400 2857 -13388
rect 2977 -13132 3035 -13120
rect 2977 -13388 2989 -13132
rect 3023 -13388 3035 -13132
rect 2977 -13400 3035 -13388
rect 3155 -13132 3213 -13120
rect 3155 -13388 3167 -13132
rect 3201 -13388 3213 -13132
rect 3155 -13400 3213 -13388
rect 3333 -13132 3391 -13120
rect 3333 -13388 3345 -13132
rect 3379 -13388 3391 -13132
rect 3333 -13400 3391 -13388
rect 3511 -13132 3569 -13120
rect 3511 -13388 3523 -13132
rect 3557 -13388 3569 -13132
rect 3511 -13400 3569 -13388
rect 3689 -13132 3747 -13120
rect 3689 -13388 3701 -13132
rect 3735 -13388 3747 -13132
rect 3689 -13400 3747 -13388
rect 3867 -13132 3925 -13120
rect 3867 -13388 3879 -13132
rect 3913 -13388 3925 -13132
rect 3867 -13400 3925 -13388
rect 4045 -13132 4103 -13120
rect 4045 -13388 4057 -13132
rect 4091 -13388 4103 -13132
rect 4045 -13400 4103 -13388
rect -4079 -13620 -4021 -13608
rect -2185 -14132 -2127 -14120
rect -6040 -14394 -5982 -14382
rect -6040 -14650 -6028 -14394
rect -5994 -14650 -5982 -14394
rect -6040 -14662 -5982 -14650
rect -5862 -14394 -5804 -14382
rect -5862 -14650 -5850 -14394
rect -5816 -14650 -5804 -14394
rect -5862 -14662 -5804 -14650
rect -5684 -14394 -5626 -14382
rect -5684 -14650 -5672 -14394
rect -5638 -14650 -5626 -14394
rect -5684 -14662 -5626 -14650
rect -5506 -14394 -5448 -14382
rect -5506 -14650 -5494 -14394
rect -5460 -14650 -5448 -14394
rect -5506 -14662 -5448 -14650
rect -5328 -14394 -5270 -14382
rect -5328 -14650 -5316 -14394
rect -5282 -14650 -5270 -14394
rect -5328 -14662 -5270 -14650
rect -5150 -14394 -5092 -14382
rect -5150 -14650 -5138 -14394
rect -5104 -14650 -5092 -14394
rect -5150 -14662 -5092 -14650
rect -4972 -14394 -4914 -14382
rect -4972 -14650 -4960 -14394
rect -4926 -14650 -4914 -14394
rect -4972 -14662 -4914 -14650
rect -4794 -14394 -4736 -14382
rect -4794 -14650 -4782 -14394
rect -4748 -14650 -4736 -14394
rect -4794 -14662 -4736 -14650
rect -4616 -14394 -4558 -14382
rect -4616 -14650 -4604 -14394
rect -4570 -14650 -4558 -14394
rect -4616 -14662 -4558 -14650
rect -4438 -14394 -4380 -14382
rect -4438 -14650 -4426 -14394
rect -4392 -14650 -4380 -14394
rect -4438 -14662 -4380 -14650
rect -4260 -14394 -4202 -14382
rect -4260 -14650 -4248 -14394
rect -4214 -14650 -4202 -14394
rect -4260 -14662 -4202 -14650
rect -4082 -14394 -4024 -14382
rect -4082 -14650 -4070 -14394
rect -4036 -14650 -4024 -14394
rect -2185 -14388 -2173 -14132
rect -2139 -14388 -2127 -14132
rect -2185 -14400 -2127 -14388
rect -2007 -14132 -1949 -14120
rect -2007 -14388 -1995 -14132
rect -1961 -14388 -1949 -14132
rect -2007 -14400 -1949 -14388
rect -1829 -14132 -1771 -14120
rect -1829 -14388 -1817 -14132
rect -1783 -14388 -1771 -14132
rect -1829 -14400 -1771 -14388
rect -1651 -14132 -1593 -14120
rect -1651 -14388 -1639 -14132
rect -1605 -14388 -1593 -14132
rect -1651 -14400 -1593 -14388
rect -1473 -14132 -1415 -14120
rect -1473 -14388 -1461 -14132
rect -1427 -14388 -1415 -14132
rect -1473 -14400 -1415 -14388
rect -1295 -14132 -1237 -14120
rect -1295 -14388 -1283 -14132
rect -1249 -14388 -1237 -14132
rect -1295 -14400 -1237 -14388
rect -1117 -14132 -1059 -14120
rect -1117 -14388 -1105 -14132
rect -1071 -14388 -1059 -14132
rect -1117 -14400 -1059 -14388
rect -939 -14132 -881 -14120
rect -939 -14388 -927 -14132
rect -893 -14388 -881 -14132
rect -939 -14400 -881 -14388
rect -761 -14132 -703 -14120
rect -761 -14388 -749 -14132
rect -715 -14388 -703 -14132
rect -761 -14400 -703 -14388
rect -583 -14132 -525 -14120
rect -583 -14388 -571 -14132
rect -537 -14388 -525 -14132
rect -583 -14400 -525 -14388
rect -405 -14132 -347 -14120
rect -405 -14388 -393 -14132
rect -359 -14388 -347 -14132
rect -405 -14400 -347 -14388
rect -227 -14132 -169 -14120
rect -227 -14388 -215 -14132
rect -181 -14388 -169 -14132
rect -227 -14400 -169 -14388
rect -49 -14132 9 -14120
rect -49 -14388 -37 -14132
rect -3 -14388 9 -14132
rect -49 -14400 9 -14388
rect 129 -14132 187 -14120
rect 129 -14388 141 -14132
rect 175 -14388 187 -14132
rect 129 -14400 187 -14388
rect 307 -14132 365 -14120
rect 307 -14388 319 -14132
rect 353 -14388 365 -14132
rect 307 -14400 365 -14388
rect 485 -14132 543 -14120
rect 485 -14388 497 -14132
rect 531 -14388 543 -14132
rect 485 -14400 543 -14388
rect 663 -14132 721 -14120
rect 663 -14388 675 -14132
rect 709 -14388 721 -14132
rect 663 -14400 721 -14388
rect 841 -14132 899 -14120
rect 841 -14388 853 -14132
rect 887 -14388 899 -14132
rect 841 -14400 899 -14388
rect 1019 -14132 1077 -14120
rect 1019 -14388 1031 -14132
rect 1065 -14388 1077 -14132
rect 1019 -14400 1077 -14388
rect 1197 -14132 1255 -14120
rect 1197 -14388 1209 -14132
rect 1243 -14388 1255 -14132
rect 1197 -14400 1255 -14388
rect 1375 -14132 1433 -14120
rect 1375 -14388 1387 -14132
rect 1421 -14388 1433 -14132
rect 1375 -14400 1433 -14388
rect 1553 -14132 1611 -14120
rect 1553 -14388 1565 -14132
rect 1599 -14388 1611 -14132
rect 1553 -14400 1611 -14388
rect 1731 -14132 1789 -14120
rect 1731 -14388 1743 -14132
rect 1777 -14388 1789 -14132
rect 1731 -14400 1789 -14388
rect 1909 -14132 1967 -14120
rect 1909 -14388 1921 -14132
rect 1955 -14388 1967 -14132
rect 1909 -14400 1967 -14388
rect 2087 -14132 2145 -14120
rect 2087 -14388 2099 -14132
rect 2133 -14388 2145 -14132
rect 2087 -14400 2145 -14388
rect 2265 -14132 2323 -14120
rect 2265 -14388 2277 -14132
rect 2311 -14388 2323 -14132
rect 2265 -14400 2323 -14388
rect 2443 -14132 2501 -14120
rect 2443 -14388 2455 -14132
rect 2489 -14388 2501 -14132
rect 2443 -14400 2501 -14388
rect 2621 -14132 2679 -14120
rect 2621 -14388 2633 -14132
rect 2667 -14388 2679 -14132
rect 2621 -14400 2679 -14388
rect 2799 -14132 2857 -14120
rect 2799 -14388 2811 -14132
rect 2845 -14388 2857 -14132
rect 2799 -14400 2857 -14388
rect 2977 -14132 3035 -14120
rect 2977 -14388 2989 -14132
rect 3023 -14388 3035 -14132
rect 2977 -14400 3035 -14388
rect 3155 -14132 3213 -14120
rect 3155 -14388 3167 -14132
rect 3201 -14388 3213 -14132
rect 3155 -14400 3213 -14388
rect 3333 -14132 3391 -14120
rect 3333 -14388 3345 -14132
rect 3379 -14388 3391 -14132
rect 3333 -14400 3391 -14388
rect 3511 -14132 3569 -14120
rect 3511 -14388 3523 -14132
rect 3557 -14388 3569 -14132
rect 3511 -14400 3569 -14388
rect 3689 -14132 3747 -14120
rect 3689 -14388 3701 -14132
rect 3735 -14388 3747 -14132
rect 3689 -14400 3747 -14388
rect 3867 -14132 3925 -14120
rect 3867 -14388 3879 -14132
rect 3913 -14388 3925 -14132
rect 3867 -14400 3925 -14388
rect 4045 -14132 4103 -14120
rect 4045 -14388 4057 -14132
rect 4091 -14388 4103 -14132
rect 4045 -14400 4103 -14388
rect 5565 -14132 5623 -14120
rect 5565 -14388 5577 -14132
rect 5611 -14388 5623 -14132
rect 5565 -14400 5623 -14388
rect 5743 -14132 5801 -14120
rect 5743 -14388 5755 -14132
rect 5789 -14388 5801 -14132
rect 5743 -14400 5801 -14388
rect 5921 -14132 5979 -14120
rect 5921 -14388 5933 -14132
rect 5967 -14388 5979 -14132
rect 5921 -14400 5979 -14388
rect 6099 -14132 6157 -14120
rect 6099 -14388 6111 -14132
rect 6145 -14388 6157 -14132
rect 6099 -14400 6157 -14388
rect 6277 -14132 6335 -14120
rect 6277 -14388 6289 -14132
rect 6323 -14388 6335 -14132
rect 6277 -14400 6335 -14388
rect 6455 -14132 6513 -14120
rect 6455 -14388 6467 -14132
rect 6501 -14388 6513 -14132
rect 6455 -14400 6513 -14388
rect 6633 -14132 6691 -14120
rect 6633 -14388 6645 -14132
rect 6679 -14388 6691 -14132
rect 6633 -14400 6691 -14388
rect 6811 -14132 6869 -14120
rect 6811 -14388 6823 -14132
rect 6857 -14388 6869 -14132
rect 6811 -14400 6869 -14388
rect 6989 -14132 7047 -14120
rect 6989 -14388 7001 -14132
rect 7035 -14388 7047 -14132
rect 6989 -14400 7047 -14388
rect 7167 -14132 7225 -14120
rect 7167 -14388 7179 -14132
rect 7213 -14388 7225 -14132
rect 7167 -14400 7225 -14388
rect 7345 -14132 7403 -14120
rect 7345 -14388 7357 -14132
rect 7391 -14388 7403 -14132
rect 7345 -14400 7403 -14388
rect 7523 -14132 7581 -14120
rect 7523 -14388 7535 -14132
rect 7569 -14388 7581 -14132
rect 7523 -14400 7581 -14388
rect 7701 -14132 7759 -14120
rect 7701 -14388 7713 -14132
rect 7747 -14388 7759 -14132
rect 7701 -14400 7759 -14388
rect 7879 -14132 7937 -14120
rect 7879 -14388 7891 -14132
rect 7925 -14388 7937 -14132
rect 7879 -14400 7937 -14388
rect 8057 -14132 8115 -14120
rect 8057 -14388 8069 -14132
rect 8103 -14388 8115 -14132
rect 8057 -14400 8115 -14388
rect 8235 -14132 8293 -14120
rect 8235 -14388 8247 -14132
rect 8281 -14388 8293 -14132
rect 8235 -14400 8293 -14388
rect 8413 -14132 8471 -14120
rect 8413 -14388 8425 -14132
rect 8459 -14388 8471 -14132
rect 8413 -14400 8471 -14388
rect 8591 -14132 8649 -14120
rect 8591 -14388 8603 -14132
rect 8637 -14388 8649 -14132
rect 8591 -14400 8649 -14388
rect 8769 -14132 8827 -14120
rect 8769 -14388 8781 -14132
rect 8815 -14388 8827 -14132
rect 8769 -14400 8827 -14388
rect 8947 -14132 9005 -14120
rect 8947 -14388 8959 -14132
rect 8993 -14388 9005 -14132
rect 8947 -14400 9005 -14388
rect 9125 -14132 9183 -14120
rect 9125 -14388 9137 -14132
rect 9171 -14388 9183 -14132
rect 9125 -14400 9183 -14388
rect 9303 -14132 9361 -14120
rect 9303 -14388 9315 -14132
rect 9349 -14388 9361 -14132
rect 9303 -14400 9361 -14388
rect 9481 -14132 9539 -14120
rect 9481 -14388 9493 -14132
rect 9527 -14388 9539 -14132
rect 9481 -14400 9539 -14388
rect 9659 -14132 9717 -14120
rect 9659 -14388 9671 -14132
rect 9705 -14388 9717 -14132
rect 9659 -14400 9717 -14388
rect 9837 -14132 9895 -14120
rect 9837 -14388 9849 -14132
rect 9883 -14388 9895 -14132
rect 9837 -14400 9895 -14388
rect 10015 -14132 10073 -14120
rect 10015 -14388 10027 -14132
rect 10061 -14388 10073 -14132
rect 10015 -14400 10073 -14388
rect 10193 -14132 10251 -14120
rect 10193 -14388 10205 -14132
rect 10239 -14388 10251 -14132
rect 10193 -14400 10251 -14388
rect 10371 -14132 10429 -14120
rect 10371 -14388 10383 -14132
rect 10417 -14388 10429 -14132
rect 10371 -14400 10429 -14388
rect 10549 -14132 10607 -14120
rect 10549 -14388 10561 -14132
rect 10595 -14388 10607 -14132
rect 10549 -14400 10607 -14388
rect 10727 -14132 10785 -14120
rect 10727 -14388 10739 -14132
rect 10773 -14388 10785 -14132
rect 10727 -14400 10785 -14388
rect 10905 -14132 10963 -14120
rect 10905 -14388 10917 -14132
rect 10951 -14388 10963 -14132
rect 10905 -14400 10963 -14388
rect 11083 -14132 11141 -14120
rect 11083 -14388 11095 -14132
rect 11129 -14388 11141 -14132
rect 11083 -14400 11141 -14388
rect 11261 -14132 11319 -14120
rect 11261 -14388 11273 -14132
rect 11307 -14388 11319 -14132
rect 11261 -14400 11319 -14388
rect 11439 -14132 11497 -14120
rect 11439 -14388 11451 -14132
rect 11485 -14388 11497 -14132
rect 11439 -14400 11497 -14388
rect 11617 -14132 11675 -14120
rect 11617 -14388 11629 -14132
rect 11663 -14388 11675 -14132
rect 11617 -14400 11675 -14388
rect 11795 -14132 11853 -14120
rect 11795 -14388 11807 -14132
rect 11841 -14388 11853 -14132
rect 11795 -14400 11853 -14388
rect 11973 -14132 12031 -14120
rect 11973 -14388 11985 -14132
rect 12019 -14388 12031 -14132
rect 11973 -14400 12031 -14388
rect 12151 -14132 12209 -14120
rect 12151 -14388 12163 -14132
rect 12197 -14388 12209 -14132
rect 12151 -14400 12209 -14388
rect 12329 -14132 12387 -14120
rect 12329 -14388 12341 -14132
rect 12375 -14388 12387 -14132
rect 12329 -14400 12387 -14388
rect 12507 -14132 12565 -14120
rect 12507 -14388 12519 -14132
rect 12553 -14388 12565 -14132
rect 12507 -14400 12565 -14388
rect 12685 -14132 12743 -14120
rect 12685 -14388 12697 -14132
rect 12731 -14388 12743 -14132
rect 12685 -14400 12743 -14388
rect -4082 -14662 -4024 -14650
rect -6040 -15094 -5982 -15082
rect -6040 -15350 -6028 -15094
rect -5994 -15350 -5982 -15094
rect -6040 -15362 -5982 -15350
rect -5862 -15094 -5804 -15082
rect -5862 -15350 -5850 -15094
rect -5816 -15350 -5804 -15094
rect -5862 -15362 -5804 -15350
rect -5684 -15094 -5626 -15082
rect -5684 -15350 -5672 -15094
rect -5638 -15350 -5626 -15094
rect -5684 -15362 -5626 -15350
rect -5506 -15094 -5448 -15082
rect -5506 -15350 -5494 -15094
rect -5460 -15350 -5448 -15094
rect -5506 -15362 -5448 -15350
rect -5328 -15094 -5270 -15082
rect -5328 -15350 -5316 -15094
rect -5282 -15350 -5270 -15094
rect -5328 -15362 -5270 -15350
rect -5150 -15094 -5092 -15082
rect -5150 -15350 -5138 -15094
rect -5104 -15350 -5092 -15094
rect -5150 -15362 -5092 -15350
rect -4972 -15094 -4914 -15082
rect -4972 -15350 -4960 -15094
rect -4926 -15350 -4914 -15094
rect -4972 -15362 -4914 -15350
rect -4794 -15094 -4736 -15082
rect -4794 -15350 -4782 -15094
rect -4748 -15350 -4736 -15094
rect -4794 -15362 -4736 -15350
rect -4616 -15094 -4558 -15082
rect -4616 -15350 -4604 -15094
rect -4570 -15350 -4558 -15094
rect -4616 -15362 -4558 -15350
rect -4438 -15094 -4380 -15082
rect -4438 -15350 -4426 -15094
rect -4392 -15350 -4380 -15094
rect -4438 -15362 -4380 -15350
rect -4260 -15094 -4202 -15082
rect -4260 -15350 -4248 -15094
rect -4214 -15350 -4202 -15094
rect -4260 -15362 -4202 -15350
rect -4082 -15094 -4024 -15082
rect -4082 -15350 -4070 -15094
rect -4036 -15350 -4024 -15094
rect -2185 -15132 -2127 -15120
rect -4082 -15362 -4024 -15350
rect -2185 -15388 -2173 -15132
rect -2139 -15388 -2127 -15132
rect -2185 -15400 -2127 -15388
rect -2007 -15132 -1949 -15120
rect -2007 -15388 -1995 -15132
rect -1961 -15388 -1949 -15132
rect -2007 -15400 -1949 -15388
rect -1829 -15132 -1771 -15120
rect -1829 -15388 -1817 -15132
rect -1783 -15388 -1771 -15132
rect -1829 -15400 -1771 -15388
rect -1651 -15132 -1593 -15120
rect -1651 -15388 -1639 -15132
rect -1605 -15388 -1593 -15132
rect -1651 -15400 -1593 -15388
rect -1473 -15132 -1415 -15120
rect -1473 -15388 -1461 -15132
rect -1427 -15388 -1415 -15132
rect -1473 -15400 -1415 -15388
rect -1295 -15132 -1237 -15120
rect -1295 -15388 -1283 -15132
rect -1249 -15388 -1237 -15132
rect -1295 -15400 -1237 -15388
rect -1117 -15132 -1059 -15120
rect -1117 -15388 -1105 -15132
rect -1071 -15388 -1059 -15132
rect -1117 -15400 -1059 -15388
rect -939 -15132 -881 -15120
rect -939 -15388 -927 -15132
rect -893 -15388 -881 -15132
rect -939 -15400 -881 -15388
rect -761 -15132 -703 -15120
rect -761 -15388 -749 -15132
rect -715 -15388 -703 -15132
rect -761 -15400 -703 -15388
rect -583 -15132 -525 -15120
rect -583 -15388 -571 -15132
rect -537 -15388 -525 -15132
rect -583 -15400 -525 -15388
rect -405 -15132 -347 -15120
rect -405 -15388 -393 -15132
rect -359 -15388 -347 -15132
rect -405 -15400 -347 -15388
rect -227 -15132 -169 -15120
rect -227 -15388 -215 -15132
rect -181 -15388 -169 -15132
rect -227 -15400 -169 -15388
rect -49 -15132 9 -15120
rect -49 -15388 -37 -15132
rect -3 -15388 9 -15132
rect -49 -15400 9 -15388
rect 129 -15132 187 -15120
rect 129 -15388 141 -15132
rect 175 -15388 187 -15132
rect 129 -15400 187 -15388
rect 307 -15132 365 -15120
rect 307 -15388 319 -15132
rect 353 -15388 365 -15132
rect 307 -15400 365 -15388
rect 485 -15132 543 -15120
rect 485 -15388 497 -15132
rect 531 -15388 543 -15132
rect 485 -15400 543 -15388
rect 663 -15132 721 -15120
rect 663 -15388 675 -15132
rect 709 -15388 721 -15132
rect 663 -15400 721 -15388
rect 841 -15132 899 -15120
rect 841 -15388 853 -15132
rect 887 -15388 899 -15132
rect 841 -15400 899 -15388
rect 1019 -15132 1077 -15120
rect 1019 -15388 1031 -15132
rect 1065 -15388 1077 -15132
rect 1019 -15400 1077 -15388
rect 1197 -15132 1255 -15120
rect 1197 -15388 1209 -15132
rect 1243 -15388 1255 -15132
rect 1197 -15400 1255 -15388
rect 1375 -15132 1433 -15120
rect 1375 -15388 1387 -15132
rect 1421 -15388 1433 -15132
rect 1375 -15400 1433 -15388
rect 1553 -15132 1611 -15120
rect 1553 -15388 1565 -15132
rect 1599 -15388 1611 -15132
rect 1553 -15400 1611 -15388
rect 1731 -15132 1789 -15120
rect 1731 -15388 1743 -15132
rect 1777 -15388 1789 -15132
rect 1731 -15400 1789 -15388
rect 1909 -15132 1967 -15120
rect 1909 -15388 1921 -15132
rect 1955 -15388 1967 -15132
rect 1909 -15400 1967 -15388
rect 2087 -15132 2145 -15120
rect 2087 -15388 2099 -15132
rect 2133 -15388 2145 -15132
rect 2087 -15400 2145 -15388
rect 2265 -15132 2323 -15120
rect 2265 -15388 2277 -15132
rect 2311 -15388 2323 -15132
rect 2265 -15400 2323 -15388
rect 2443 -15132 2501 -15120
rect 2443 -15388 2455 -15132
rect 2489 -15388 2501 -15132
rect 2443 -15400 2501 -15388
rect 2621 -15132 2679 -15120
rect 2621 -15388 2633 -15132
rect 2667 -15388 2679 -15132
rect 2621 -15400 2679 -15388
rect 2799 -15132 2857 -15120
rect 2799 -15388 2811 -15132
rect 2845 -15388 2857 -15132
rect 2799 -15400 2857 -15388
rect 2977 -15132 3035 -15120
rect 2977 -15388 2989 -15132
rect 3023 -15388 3035 -15132
rect 2977 -15400 3035 -15388
rect 3155 -15132 3213 -15120
rect 3155 -15388 3167 -15132
rect 3201 -15388 3213 -15132
rect 3155 -15400 3213 -15388
rect 3333 -15132 3391 -15120
rect 3333 -15388 3345 -15132
rect 3379 -15388 3391 -15132
rect 3333 -15400 3391 -15388
rect 3511 -15132 3569 -15120
rect 3511 -15388 3523 -15132
rect 3557 -15388 3569 -15132
rect 3511 -15400 3569 -15388
rect 3689 -15132 3747 -15120
rect 3689 -15388 3701 -15132
rect 3735 -15388 3747 -15132
rect 3689 -15400 3747 -15388
rect 3867 -15132 3925 -15120
rect 3867 -15388 3879 -15132
rect 3913 -15388 3925 -15132
rect 3867 -15400 3925 -15388
rect 4045 -15132 4103 -15120
rect 4045 -15388 4057 -15132
rect 4091 -15388 4103 -15132
rect 4045 -15400 4103 -15388
rect 5565 -15132 5623 -15120
rect 5565 -15388 5577 -15132
rect 5611 -15388 5623 -15132
rect 5565 -15400 5623 -15388
rect 5743 -15132 5801 -15120
rect 5743 -15388 5755 -15132
rect 5789 -15388 5801 -15132
rect 5743 -15400 5801 -15388
rect 5921 -15132 5979 -15120
rect 5921 -15388 5933 -15132
rect 5967 -15388 5979 -15132
rect 5921 -15400 5979 -15388
rect 6099 -15132 6157 -15120
rect 6099 -15388 6111 -15132
rect 6145 -15388 6157 -15132
rect 6099 -15400 6157 -15388
rect 6277 -15132 6335 -15120
rect 6277 -15388 6289 -15132
rect 6323 -15388 6335 -15132
rect 6277 -15400 6335 -15388
rect 6455 -15132 6513 -15120
rect 6455 -15388 6467 -15132
rect 6501 -15388 6513 -15132
rect 6455 -15400 6513 -15388
rect 6633 -15132 6691 -15120
rect 6633 -15388 6645 -15132
rect 6679 -15388 6691 -15132
rect 6633 -15400 6691 -15388
rect 6811 -15132 6869 -15120
rect 6811 -15388 6823 -15132
rect 6857 -15388 6869 -15132
rect 6811 -15400 6869 -15388
rect 6989 -15132 7047 -15120
rect 6989 -15388 7001 -15132
rect 7035 -15388 7047 -15132
rect 6989 -15400 7047 -15388
rect 7167 -15132 7225 -15120
rect 7167 -15388 7179 -15132
rect 7213 -15388 7225 -15132
rect 7167 -15400 7225 -15388
rect 7345 -15132 7403 -15120
rect 7345 -15388 7357 -15132
rect 7391 -15388 7403 -15132
rect 7345 -15400 7403 -15388
rect 7523 -15132 7581 -15120
rect 7523 -15388 7535 -15132
rect 7569 -15388 7581 -15132
rect 7523 -15400 7581 -15388
rect 7701 -15132 7759 -15120
rect 7701 -15388 7713 -15132
rect 7747 -15388 7759 -15132
rect 7701 -15400 7759 -15388
rect 7879 -15132 7937 -15120
rect 7879 -15388 7891 -15132
rect 7925 -15388 7937 -15132
rect 7879 -15400 7937 -15388
rect 8057 -15132 8115 -15120
rect 8057 -15388 8069 -15132
rect 8103 -15388 8115 -15132
rect 8057 -15400 8115 -15388
rect 8235 -15132 8293 -15120
rect 8235 -15388 8247 -15132
rect 8281 -15388 8293 -15132
rect 8235 -15400 8293 -15388
rect 8413 -15132 8471 -15120
rect 8413 -15388 8425 -15132
rect 8459 -15388 8471 -15132
rect 8413 -15400 8471 -15388
rect 8591 -15132 8649 -15120
rect 8591 -15388 8603 -15132
rect 8637 -15388 8649 -15132
rect 8591 -15400 8649 -15388
rect 8769 -15132 8827 -15120
rect 8769 -15388 8781 -15132
rect 8815 -15388 8827 -15132
rect 8769 -15400 8827 -15388
rect 8947 -15132 9005 -15120
rect 8947 -15388 8959 -15132
rect 8993 -15388 9005 -15132
rect 8947 -15400 9005 -15388
rect 9125 -15132 9183 -15120
rect 9125 -15388 9137 -15132
rect 9171 -15388 9183 -15132
rect 9125 -15400 9183 -15388
rect 9303 -15132 9361 -15120
rect 9303 -15388 9315 -15132
rect 9349 -15388 9361 -15132
rect 9303 -15400 9361 -15388
rect 9481 -15132 9539 -15120
rect 9481 -15388 9493 -15132
rect 9527 -15388 9539 -15132
rect 9481 -15400 9539 -15388
rect 9659 -15132 9717 -15120
rect 9659 -15388 9671 -15132
rect 9705 -15388 9717 -15132
rect 9659 -15400 9717 -15388
rect 9837 -15132 9895 -15120
rect 9837 -15388 9849 -15132
rect 9883 -15388 9895 -15132
rect 9837 -15400 9895 -15388
rect 10015 -15132 10073 -15120
rect 10015 -15388 10027 -15132
rect 10061 -15388 10073 -15132
rect 10015 -15400 10073 -15388
rect 10193 -15132 10251 -15120
rect 10193 -15388 10205 -15132
rect 10239 -15388 10251 -15132
rect 10193 -15400 10251 -15388
rect 10371 -15132 10429 -15120
rect 10371 -15388 10383 -15132
rect 10417 -15388 10429 -15132
rect 10371 -15400 10429 -15388
rect 10549 -15132 10607 -15120
rect 10549 -15388 10561 -15132
rect 10595 -15388 10607 -15132
rect 10549 -15400 10607 -15388
rect 10727 -15132 10785 -15120
rect 10727 -15388 10739 -15132
rect 10773 -15388 10785 -15132
rect 10727 -15400 10785 -15388
rect 10905 -15132 10963 -15120
rect 10905 -15388 10917 -15132
rect 10951 -15388 10963 -15132
rect 10905 -15400 10963 -15388
rect 11083 -15132 11141 -15120
rect 11083 -15388 11095 -15132
rect 11129 -15388 11141 -15132
rect 11083 -15400 11141 -15388
rect 11261 -15132 11319 -15120
rect 11261 -15388 11273 -15132
rect 11307 -15388 11319 -15132
rect 11261 -15400 11319 -15388
rect 11439 -15132 11497 -15120
rect 11439 -15388 11451 -15132
rect 11485 -15388 11497 -15132
rect 11439 -15400 11497 -15388
rect 11617 -15132 11675 -15120
rect 11617 -15388 11629 -15132
rect 11663 -15388 11675 -15132
rect 11617 -15400 11675 -15388
rect 11795 -15132 11853 -15120
rect 11795 -15388 11807 -15132
rect 11841 -15388 11853 -15132
rect 11795 -15400 11853 -15388
rect 11973 -15132 12031 -15120
rect 11973 -15388 11985 -15132
rect 12019 -15388 12031 -15132
rect 11973 -15400 12031 -15388
rect 12151 -15132 12209 -15120
rect 12151 -15388 12163 -15132
rect 12197 -15388 12209 -15132
rect 12151 -15400 12209 -15388
rect 12329 -15132 12387 -15120
rect 12329 -15388 12341 -15132
rect 12375 -15388 12387 -15132
rect 12329 -15400 12387 -15388
rect 12507 -15132 12565 -15120
rect 12507 -15388 12519 -15132
rect 12553 -15388 12565 -15132
rect 12507 -15400 12565 -15388
rect 12685 -15132 12743 -15120
rect 12685 -15388 12697 -15132
rect 12731 -15388 12743 -15132
rect 12685 -15400 12743 -15388
rect -6040 -15794 -5982 -15782
rect -6040 -16050 -6028 -15794
rect -5994 -16050 -5982 -15794
rect -6040 -16062 -5982 -16050
rect -5862 -15794 -5804 -15782
rect -5862 -16050 -5850 -15794
rect -5816 -16050 -5804 -15794
rect -5862 -16062 -5804 -16050
rect -5684 -15794 -5626 -15782
rect -5684 -16050 -5672 -15794
rect -5638 -16050 -5626 -15794
rect -5684 -16062 -5626 -16050
rect -5506 -15794 -5448 -15782
rect -5506 -16050 -5494 -15794
rect -5460 -16050 -5448 -15794
rect -5506 -16062 -5448 -16050
rect -5328 -15794 -5270 -15782
rect -5328 -16050 -5316 -15794
rect -5282 -16050 -5270 -15794
rect -5328 -16062 -5270 -16050
rect -5150 -15794 -5092 -15782
rect -5150 -16050 -5138 -15794
rect -5104 -16050 -5092 -15794
rect -5150 -16062 -5092 -16050
rect -4972 -15794 -4914 -15782
rect -4972 -16050 -4960 -15794
rect -4926 -16050 -4914 -15794
rect -4972 -16062 -4914 -16050
rect -4794 -15794 -4736 -15782
rect -4794 -16050 -4782 -15794
rect -4748 -16050 -4736 -15794
rect -4794 -16062 -4736 -16050
rect -4616 -15794 -4558 -15782
rect -4616 -16050 -4604 -15794
rect -4570 -16050 -4558 -15794
rect -4616 -16062 -4558 -16050
rect -4438 -15794 -4380 -15782
rect -4438 -16050 -4426 -15794
rect -4392 -16050 -4380 -15794
rect -4438 -16062 -4380 -16050
rect -4260 -15794 -4202 -15782
rect -4260 -16050 -4248 -15794
rect -4214 -16050 -4202 -15794
rect -4260 -16062 -4202 -16050
rect -4082 -15794 -4024 -15782
rect -4082 -16050 -4070 -15794
rect -4036 -16050 -4024 -15794
rect -4082 -16062 -4024 -16050
rect -2185 -16132 -2127 -16120
rect -2185 -16388 -2173 -16132
rect -2139 -16388 -2127 -16132
rect -2185 -16400 -2127 -16388
rect -2007 -16132 -1949 -16120
rect -2007 -16388 -1995 -16132
rect -1961 -16388 -1949 -16132
rect -2007 -16400 -1949 -16388
rect -1829 -16132 -1771 -16120
rect -1829 -16388 -1817 -16132
rect -1783 -16388 -1771 -16132
rect -1829 -16400 -1771 -16388
rect -1651 -16132 -1593 -16120
rect -1651 -16388 -1639 -16132
rect -1605 -16388 -1593 -16132
rect -1651 -16400 -1593 -16388
rect -1473 -16132 -1415 -16120
rect -1473 -16388 -1461 -16132
rect -1427 -16388 -1415 -16132
rect -1473 -16400 -1415 -16388
rect -1295 -16132 -1237 -16120
rect -1295 -16388 -1283 -16132
rect -1249 -16388 -1237 -16132
rect -1295 -16400 -1237 -16388
rect -1117 -16132 -1059 -16120
rect -1117 -16388 -1105 -16132
rect -1071 -16388 -1059 -16132
rect -1117 -16400 -1059 -16388
rect -939 -16132 -881 -16120
rect -939 -16388 -927 -16132
rect -893 -16388 -881 -16132
rect -939 -16400 -881 -16388
rect -761 -16132 -703 -16120
rect -761 -16388 -749 -16132
rect -715 -16388 -703 -16132
rect -761 -16400 -703 -16388
rect -583 -16132 -525 -16120
rect -583 -16388 -571 -16132
rect -537 -16388 -525 -16132
rect -583 -16400 -525 -16388
rect -405 -16132 -347 -16120
rect -405 -16388 -393 -16132
rect -359 -16388 -347 -16132
rect -405 -16400 -347 -16388
rect -227 -16132 -169 -16120
rect -227 -16388 -215 -16132
rect -181 -16388 -169 -16132
rect -227 -16400 -169 -16388
rect -49 -16132 9 -16120
rect -49 -16388 -37 -16132
rect -3 -16388 9 -16132
rect -49 -16400 9 -16388
rect 129 -16132 187 -16120
rect 129 -16388 141 -16132
rect 175 -16388 187 -16132
rect 129 -16400 187 -16388
rect 307 -16132 365 -16120
rect 307 -16388 319 -16132
rect 353 -16388 365 -16132
rect 307 -16400 365 -16388
rect 485 -16132 543 -16120
rect 485 -16388 497 -16132
rect 531 -16388 543 -16132
rect 485 -16400 543 -16388
rect 663 -16132 721 -16120
rect 663 -16388 675 -16132
rect 709 -16388 721 -16132
rect 663 -16400 721 -16388
rect 841 -16132 899 -16120
rect 841 -16388 853 -16132
rect 887 -16388 899 -16132
rect 841 -16400 899 -16388
rect 1019 -16132 1077 -16120
rect 1019 -16388 1031 -16132
rect 1065 -16388 1077 -16132
rect 1019 -16400 1077 -16388
rect 1197 -16132 1255 -16120
rect 1197 -16388 1209 -16132
rect 1243 -16388 1255 -16132
rect 1197 -16400 1255 -16388
rect 1375 -16132 1433 -16120
rect 1375 -16388 1387 -16132
rect 1421 -16388 1433 -16132
rect 1375 -16400 1433 -16388
rect 1553 -16132 1611 -16120
rect 1553 -16388 1565 -16132
rect 1599 -16388 1611 -16132
rect 1553 -16400 1611 -16388
rect 1731 -16132 1789 -16120
rect 1731 -16388 1743 -16132
rect 1777 -16388 1789 -16132
rect 1731 -16400 1789 -16388
rect 1909 -16132 1967 -16120
rect 1909 -16388 1921 -16132
rect 1955 -16388 1967 -16132
rect 1909 -16400 1967 -16388
rect 2087 -16132 2145 -16120
rect 2087 -16388 2099 -16132
rect 2133 -16388 2145 -16132
rect 2087 -16400 2145 -16388
rect 2265 -16132 2323 -16120
rect 2265 -16388 2277 -16132
rect 2311 -16388 2323 -16132
rect 2265 -16400 2323 -16388
rect 2443 -16132 2501 -16120
rect 2443 -16388 2455 -16132
rect 2489 -16388 2501 -16132
rect 2443 -16400 2501 -16388
rect 2621 -16132 2679 -16120
rect 2621 -16388 2633 -16132
rect 2667 -16388 2679 -16132
rect 2621 -16400 2679 -16388
rect 2799 -16132 2857 -16120
rect 2799 -16388 2811 -16132
rect 2845 -16388 2857 -16132
rect 2799 -16400 2857 -16388
rect 2977 -16132 3035 -16120
rect 2977 -16388 2989 -16132
rect 3023 -16388 3035 -16132
rect 2977 -16400 3035 -16388
rect 3155 -16132 3213 -16120
rect 3155 -16388 3167 -16132
rect 3201 -16388 3213 -16132
rect 3155 -16400 3213 -16388
rect 3333 -16132 3391 -16120
rect 3333 -16388 3345 -16132
rect 3379 -16388 3391 -16132
rect 3333 -16400 3391 -16388
rect 3511 -16132 3569 -16120
rect 3511 -16388 3523 -16132
rect 3557 -16388 3569 -16132
rect 3511 -16400 3569 -16388
rect 3689 -16132 3747 -16120
rect 3689 -16388 3701 -16132
rect 3735 -16388 3747 -16132
rect 3689 -16400 3747 -16388
rect 3867 -16132 3925 -16120
rect 3867 -16388 3879 -16132
rect 3913 -16388 3925 -16132
rect 3867 -16400 3925 -16388
rect 4045 -16132 4103 -16120
rect 4045 -16388 4057 -16132
rect 4091 -16388 4103 -16132
rect 4045 -16400 4103 -16388
rect 5565 -16132 5623 -16120
rect 5565 -16388 5577 -16132
rect 5611 -16388 5623 -16132
rect 5565 -16400 5623 -16388
rect 5743 -16132 5801 -16120
rect 5743 -16388 5755 -16132
rect 5789 -16388 5801 -16132
rect 5743 -16400 5801 -16388
rect 5921 -16132 5979 -16120
rect 5921 -16388 5933 -16132
rect 5967 -16388 5979 -16132
rect 5921 -16400 5979 -16388
rect 6099 -16132 6157 -16120
rect 6099 -16388 6111 -16132
rect 6145 -16388 6157 -16132
rect 6099 -16400 6157 -16388
rect 6277 -16132 6335 -16120
rect 6277 -16388 6289 -16132
rect 6323 -16388 6335 -16132
rect 6277 -16400 6335 -16388
rect 6455 -16132 6513 -16120
rect 6455 -16388 6467 -16132
rect 6501 -16388 6513 -16132
rect 6455 -16400 6513 -16388
rect 6633 -16132 6691 -16120
rect 6633 -16388 6645 -16132
rect 6679 -16388 6691 -16132
rect 6633 -16400 6691 -16388
rect 6811 -16132 6869 -16120
rect 6811 -16388 6823 -16132
rect 6857 -16388 6869 -16132
rect 6811 -16400 6869 -16388
rect 6989 -16132 7047 -16120
rect 6989 -16388 7001 -16132
rect 7035 -16388 7047 -16132
rect 6989 -16400 7047 -16388
rect 7167 -16132 7225 -16120
rect 7167 -16388 7179 -16132
rect 7213 -16388 7225 -16132
rect 7167 -16400 7225 -16388
rect 7345 -16132 7403 -16120
rect 7345 -16388 7357 -16132
rect 7391 -16388 7403 -16132
rect 7345 -16400 7403 -16388
rect 7523 -16132 7581 -16120
rect 7523 -16388 7535 -16132
rect 7569 -16388 7581 -16132
rect 7523 -16400 7581 -16388
rect 7701 -16132 7759 -16120
rect 7701 -16388 7713 -16132
rect 7747 -16388 7759 -16132
rect 7701 -16400 7759 -16388
rect 7879 -16132 7937 -16120
rect 7879 -16388 7891 -16132
rect 7925 -16388 7937 -16132
rect 7879 -16400 7937 -16388
rect 8057 -16132 8115 -16120
rect 8057 -16388 8069 -16132
rect 8103 -16388 8115 -16132
rect 8057 -16400 8115 -16388
rect 8235 -16132 8293 -16120
rect 8235 -16388 8247 -16132
rect 8281 -16388 8293 -16132
rect 8235 -16400 8293 -16388
rect 8413 -16132 8471 -16120
rect 8413 -16388 8425 -16132
rect 8459 -16388 8471 -16132
rect 8413 -16400 8471 -16388
rect 8591 -16132 8649 -16120
rect 8591 -16388 8603 -16132
rect 8637 -16388 8649 -16132
rect 8591 -16400 8649 -16388
rect 8769 -16132 8827 -16120
rect 8769 -16388 8781 -16132
rect 8815 -16388 8827 -16132
rect 8769 -16400 8827 -16388
rect 8947 -16132 9005 -16120
rect 8947 -16388 8959 -16132
rect 8993 -16388 9005 -16132
rect 8947 -16400 9005 -16388
rect 9125 -16132 9183 -16120
rect 9125 -16388 9137 -16132
rect 9171 -16388 9183 -16132
rect 9125 -16400 9183 -16388
rect 9303 -16132 9361 -16120
rect 9303 -16388 9315 -16132
rect 9349 -16388 9361 -16132
rect 9303 -16400 9361 -16388
rect 9481 -16132 9539 -16120
rect 9481 -16388 9493 -16132
rect 9527 -16388 9539 -16132
rect 9481 -16400 9539 -16388
rect 9659 -16132 9717 -16120
rect 9659 -16388 9671 -16132
rect 9705 -16388 9717 -16132
rect 9659 -16400 9717 -16388
rect 9837 -16132 9895 -16120
rect 9837 -16388 9849 -16132
rect 9883 -16388 9895 -16132
rect 9837 -16400 9895 -16388
rect 10015 -16132 10073 -16120
rect 10015 -16388 10027 -16132
rect 10061 -16388 10073 -16132
rect 10015 -16400 10073 -16388
rect 10193 -16132 10251 -16120
rect 10193 -16388 10205 -16132
rect 10239 -16388 10251 -16132
rect 10193 -16400 10251 -16388
rect 10371 -16132 10429 -16120
rect 10371 -16388 10383 -16132
rect 10417 -16388 10429 -16132
rect 10371 -16400 10429 -16388
rect 10549 -16132 10607 -16120
rect 10549 -16388 10561 -16132
rect 10595 -16388 10607 -16132
rect 10549 -16400 10607 -16388
rect 10727 -16132 10785 -16120
rect 10727 -16388 10739 -16132
rect 10773 -16388 10785 -16132
rect 10727 -16400 10785 -16388
rect 10905 -16132 10963 -16120
rect 10905 -16388 10917 -16132
rect 10951 -16388 10963 -16132
rect 10905 -16400 10963 -16388
rect 11083 -16132 11141 -16120
rect 11083 -16388 11095 -16132
rect 11129 -16388 11141 -16132
rect 11083 -16400 11141 -16388
rect 11261 -16132 11319 -16120
rect 11261 -16388 11273 -16132
rect 11307 -16388 11319 -16132
rect 11261 -16400 11319 -16388
rect 11439 -16132 11497 -16120
rect 11439 -16388 11451 -16132
rect 11485 -16388 11497 -16132
rect 11439 -16400 11497 -16388
rect 11617 -16132 11675 -16120
rect 11617 -16388 11629 -16132
rect 11663 -16388 11675 -16132
rect 11617 -16400 11675 -16388
rect 11795 -16132 11853 -16120
rect 11795 -16388 11807 -16132
rect 11841 -16388 11853 -16132
rect 11795 -16400 11853 -16388
rect 11973 -16132 12031 -16120
rect 11973 -16388 11985 -16132
rect 12019 -16388 12031 -16132
rect 11973 -16400 12031 -16388
rect 12151 -16132 12209 -16120
rect 12151 -16388 12163 -16132
rect 12197 -16388 12209 -16132
rect 12151 -16400 12209 -16388
rect 12329 -16132 12387 -16120
rect 12329 -16388 12341 -16132
rect 12375 -16388 12387 -16132
rect 12329 -16400 12387 -16388
rect 12507 -16132 12565 -16120
rect 12507 -16388 12519 -16132
rect 12553 -16388 12565 -16132
rect 12507 -16400 12565 -16388
rect 12685 -16132 12743 -16120
rect 12685 -16388 12697 -16132
rect 12731 -16388 12743 -16132
rect 12685 -16400 12743 -16388
rect -6040 -16494 -5982 -16482
rect -6040 -16750 -6028 -16494
rect -5994 -16750 -5982 -16494
rect -6040 -16762 -5982 -16750
rect -5862 -16494 -5804 -16482
rect -5862 -16750 -5850 -16494
rect -5816 -16750 -5804 -16494
rect -5862 -16762 -5804 -16750
rect -5684 -16494 -5626 -16482
rect -5684 -16750 -5672 -16494
rect -5638 -16750 -5626 -16494
rect -5684 -16762 -5626 -16750
rect -5506 -16494 -5448 -16482
rect -5506 -16750 -5494 -16494
rect -5460 -16750 -5448 -16494
rect -5506 -16762 -5448 -16750
rect -5328 -16494 -5270 -16482
rect -5328 -16750 -5316 -16494
rect -5282 -16750 -5270 -16494
rect -5328 -16762 -5270 -16750
rect -5150 -16494 -5092 -16482
rect -5150 -16750 -5138 -16494
rect -5104 -16750 -5092 -16494
rect -5150 -16762 -5092 -16750
rect -4972 -16494 -4914 -16482
rect -4972 -16750 -4960 -16494
rect -4926 -16750 -4914 -16494
rect -4972 -16762 -4914 -16750
rect -4794 -16494 -4736 -16482
rect -4794 -16750 -4782 -16494
rect -4748 -16750 -4736 -16494
rect -4794 -16762 -4736 -16750
rect -4616 -16494 -4558 -16482
rect -4616 -16750 -4604 -16494
rect -4570 -16750 -4558 -16494
rect -4616 -16762 -4558 -16750
rect -4438 -16494 -4380 -16482
rect -4438 -16750 -4426 -16494
rect -4392 -16750 -4380 -16494
rect -4438 -16762 -4380 -16750
rect -4260 -16494 -4202 -16482
rect -4260 -16750 -4248 -16494
rect -4214 -16750 -4202 -16494
rect -4260 -16762 -4202 -16750
rect -4082 -16494 -4024 -16482
rect -4082 -16750 -4070 -16494
rect -4036 -16750 -4024 -16494
rect -4082 -16762 -4024 -16750
<< pdiff >>
rect 7142 2613 7204 2625
rect 7142 2365 7154 2613
rect 7188 2365 7204 2613
rect 7142 2353 7204 2365
rect 7234 2613 7300 2625
rect 7234 2365 7250 2613
rect 7284 2365 7300 2613
rect 7234 2353 7300 2365
rect 7330 2613 7396 2625
rect 7330 2365 7346 2613
rect 7380 2365 7396 2613
rect 7330 2353 7396 2365
rect 7426 2613 7492 2625
rect 7426 2365 7442 2613
rect 7476 2365 7492 2613
rect 7426 2353 7492 2365
rect 7522 2613 7588 2625
rect 7522 2365 7538 2613
rect 7572 2365 7588 2613
rect 7522 2353 7588 2365
rect 7618 2613 7684 2625
rect 7618 2365 7634 2613
rect 7668 2365 7684 2613
rect 7618 2353 7684 2365
rect 7714 2613 7780 2625
rect 7714 2365 7730 2613
rect 7764 2365 7780 2613
rect 7714 2353 7780 2365
rect 7810 2613 7876 2625
rect 7810 2365 7826 2613
rect 7860 2365 7876 2613
rect 7810 2353 7876 2365
rect 7906 2613 7972 2625
rect 7906 2365 7922 2613
rect 7956 2365 7972 2613
rect 7906 2353 7972 2365
rect 8002 2613 8068 2625
rect 8002 2365 8018 2613
rect 8052 2365 8068 2613
rect 8002 2353 8068 2365
rect 8098 2613 8160 2625
rect 8098 2365 8114 2613
rect 8148 2365 8160 2613
rect 8098 2353 8160 2365
rect 16142 2613 16204 2625
rect 16142 2365 16154 2613
rect 16188 2365 16204 2613
rect 16142 2353 16204 2365
rect 16234 2613 16300 2625
rect 16234 2365 16250 2613
rect 16284 2365 16300 2613
rect 16234 2353 16300 2365
rect 16330 2613 16396 2625
rect 16330 2365 16346 2613
rect 16380 2365 16396 2613
rect 16330 2353 16396 2365
rect 16426 2613 16492 2625
rect 16426 2365 16442 2613
rect 16476 2365 16492 2613
rect 16426 2353 16492 2365
rect 16522 2613 16588 2625
rect 16522 2365 16538 2613
rect 16572 2365 16588 2613
rect 16522 2353 16588 2365
rect 16618 2613 16684 2625
rect 16618 2365 16634 2613
rect 16668 2365 16684 2613
rect 16618 2353 16684 2365
rect 16714 2613 16780 2625
rect 16714 2365 16730 2613
rect 16764 2365 16780 2613
rect 16714 2353 16780 2365
rect 16810 2613 16876 2625
rect 16810 2365 16826 2613
rect 16860 2365 16876 2613
rect 16810 2353 16876 2365
rect 16906 2613 16972 2625
rect 16906 2365 16922 2613
rect 16956 2365 16972 2613
rect 16906 2353 16972 2365
rect 17002 2613 17068 2625
rect 17002 2365 17018 2613
rect 17052 2365 17068 2613
rect 17002 2353 17068 2365
rect 17098 2613 17160 2625
rect 17098 2365 17114 2613
rect 17148 2365 17160 2613
rect 17098 2353 17160 2365
rect 7142 813 7204 825
rect 7142 565 7154 813
rect 7188 565 7204 813
rect 7142 553 7204 565
rect 7234 813 7300 825
rect 7234 565 7250 813
rect 7284 565 7300 813
rect 7234 553 7300 565
rect 7330 813 7396 825
rect 7330 565 7346 813
rect 7380 565 7396 813
rect 7330 553 7396 565
rect 7426 813 7492 825
rect 7426 565 7442 813
rect 7476 565 7492 813
rect 7426 553 7492 565
rect 7522 813 7588 825
rect 7522 565 7538 813
rect 7572 565 7588 813
rect 7522 553 7588 565
rect 7618 813 7684 825
rect 7618 565 7634 813
rect 7668 565 7684 813
rect 7618 553 7684 565
rect 7714 813 7780 825
rect 7714 565 7730 813
rect 7764 565 7780 813
rect 7714 553 7780 565
rect 7810 813 7876 825
rect 7810 565 7826 813
rect 7860 565 7876 813
rect 7810 553 7876 565
rect 7906 813 7972 825
rect 7906 565 7922 813
rect 7956 565 7972 813
rect 7906 553 7972 565
rect 8002 813 8068 825
rect 8002 565 8018 813
rect 8052 565 8068 813
rect 8002 553 8068 565
rect 8098 813 8160 825
rect 8098 565 8114 813
rect 8148 565 8160 813
rect 8098 553 8160 565
rect 16142 813 16204 825
rect 16142 565 16154 813
rect 16188 565 16204 813
rect 16142 553 16204 565
rect 16234 813 16300 825
rect 16234 565 16250 813
rect 16284 565 16300 813
rect 16234 553 16300 565
rect 16330 813 16396 825
rect 16330 565 16346 813
rect 16380 565 16396 813
rect 16330 553 16396 565
rect 16426 813 16492 825
rect 16426 565 16442 813
rect 16476 565 16492 813
rect 16426 553 16492 565
rect 16522 813 16588 825
rect 16522 565 16538 813
rect 16572 565 16588 813
rect 16522 553 16588 565
rect 16618 813 16684 825
rect 16618 565 16634 813
rect 16668 565 16684 813
rect 16618 553 16684 565
rect 16714 813 16780 825
rect 16714 565 16730 813
rect 16764 565 16780 813
rect 16714 553 16780 565
rect 16810 813 16876 825
rect 16810 565 16826 813
rect 16860 565 16876 813
rect 16810 553 16876 565
rect 16906 813 16972 825
rect 16906 565 16922 813
rect 16956 565 16972 813
rect 16906 553 16972 565
rect 17002 813 17068 825
rect 17002 565 17018 813
rect 17052 565 17068 813
rect 17002 553 17068 565
rect 17098 813 17160 825
rect 17098 565 17114 813
rect 17148 565 17160 813
rect 17098 553 17160 565
rect 7142 -987 7204 -975
rect 7142 -1235 7154 -987
rect 7188 -1235 7204 -987
rect 7142 -1247 7204 -1235
rect 7234 -987 7300 -975
rect 7234 -1235 7250 -987
rect 7284 -1235 7300 -987
rect 7234 -1247 7300 -1235
rect 7330 -987 7396 -975
rect 7330 -1235 7346 -987
rect 7380 -1235 7396 -987
rect 7330 -1247 7396 -1235
rect 7426 -987 7492 -975
rect 7426 -1235 7442 -987
rect 7476 -1235 7492 -987
rect 7426 -1247 7492 -1235
rect 7522 -987 7588 -975
rect 7522 -1235 7538 -987
rect 7572 -1235 7588 -987
rect 7522 -1247 7588 -1235
rect 7618 -987 7684 -975
rect 7618 -1235 7634 -987
rect 7668 -1235 7684 -987
rect 7618 -1247 7684 -1235
rect 7714 -987 7780 -975
rect 7714 -1235 7730 -987
rect 7764 -1235 7780 -987
rect 7714 -1247 7780 -1235
rect 7810 -987 7876 -975
rect 7810 -1235 7826 -987
rect 7860 -1235 7876 -987
rect 7810 -1247 7876 -1235
rect 7906 -987 7972 -975
rect 7906 -1235 7922 -987
rect 7956 -1235 7972 -987
rect 7906 -1247 7972 -1235
rect 8002 -987 8068 -975
rect 8002 -1235 8018 -987
rect 8052 -1235 8068 -987
rect 8002 -1247 8068 -1235
rect 8098 -987 8160 -975
rect 8098 -1235 8114 -987
rect 8148 -1235 8160 -987
rect 8098 -1247 8160 -1235
rect 16142 -987 16204 -975
rect 16142 -1235 16154 -987
rect 16188 -1235 16204 -987
rect 16142 -1247 16204 -1235
rect 16234 -987 16300 -975
rect 16234 -1235 16250 -987
rect 16284 -1235 16300 -987
rect 16234 -1247 16300 -1235
rect 16330 -987 16396 -975
rect 16330 -1235 16346 -987
rect 16380 -1235 16396 -987
rect 16330 -1247 16396 -1235
rect 16426 -987 16492 -975
rect 16426 -1235 16442 -987
rect 16476 -1235 16492 -987
rect 16426 -1247 16492 -1235
rect 16522 -987 16588 -975
rect 16522 -1235 16538 -987
rect 16572 -1235 16588 -987
rect 16522 -1247 16588 -1235
rect 16618 -987 16684 -975
rect 16618 -1235 16634 -987
rect 16668 -1235 16684 -987
rect 16618 -1247 16684 -1235
rect 16714 -987 16780 -975
rect 16714 -1235 16730 -987
rect 16764 -1235 16780 -987
rect 16714 -1247 16780 -1235
rect 16810 -987 16876 -975
rect 16810 -1235 16826 -987
rect 16860 -1235 16876 -987
rect 16810 -1247 16876 -1235
rect 16906 -987 16972 -975
rect 16906 -1235 16922 -987
rect 16956 -1235 16972 -987
rect 16906 -1247 16972 -1235
rect 17002 -987 17068 -975
rect 17002 -1235 17018 -987
rect 17052 -1235 17068 -987
rect 17002 -1247 17068 -1235
rect 17098 -987 17160 -975
rect 17098 -1235 17114 -987
rect 17148 -1235 17160 -987
rect 17098 -1247 17160 -1235
rect -6314 -2132 -6256 -2120
rect -6314 -2388 -6302 -2132
rect -6268 -2388 -6256 -2132
rect -6314 -2400 -6256 -2388
rect -6136 -2132 -6078 -2120
rect -6136 -2388 -6124 -2132
rect -6090 -2388 -6078 -2132
rect -6136 -2400 -6078 -2388
rect -5958 -2132 -5900 -2120
rect -5958 -2388 -5946 -2132
rect -5912 -2388 -5900 -2132
rect -5958 -2400 -5900 -2388
rect -5780 -2132 -5722 -2120
rect -5780 -2388 -5768 -2132
rect -5734 -2388 -5722 -2132
rect -5780 -2400 -5722 -2388
rect -5602 -2132 -5544 -2120
rect -5602 -2388 -5590 -2132
rect -5556 -2388 -5544 -2132
rect -5602 -2400 -5544 -2388
rect -5424 -2132 -5366 -2120
rect -5424 -2388 -5412 -2132
rect -5378 -2388 -5366 -2132
rect -5424 -2400 -5366 -2388
rect -5246 -2132 -5188 -2120
rect -5246 -2388 -5234 -2132
rect -5200 -2388 -5188 -2132
rect -5246 -2400 -5188 -2388
rect -5068 -2132 -5010 -2120
rect -5068 -2388 -5056 -2132
rect -5022 -2388 -5010 -2132
rect -5068 -2400 -5010 -2388
rect -4890 -2132 -4832 -2120
rect -4890 -2388 -4878 -2132
rect -4844 -2388 -4832 -2132
rect -4890 -2400 -4832 -2388
rect -4712 -2132 -4654 -2120
rect -4712 -2388 -4700 -2132
rect -4666 -2388 -4654 -2132
rect -4712 -2400 -4654 -2388
rect -4534 -2132 -4476 -2120
rect -4534 -2388 -4522 -2132
rect -4488 -2388 -4476 -2132
rect -4534 -2400 -4476 -2388
rect -4356 -2132 -4298 -2120
rect -4356 -2388 -4344 -2132
rect -4310 -2388 -4298 -2132
rect -4356 -2400 -4298 -2388
rect -4178 -2132 -4120 -2120
rect -4178 -2388 -4166 -2132
rect -4132 -2388 -4120 -2132
rect -4178 -2400 -4120 -2388
rect -4000 -2132 -3942 -2120
rect -4000 -2388 -3988 -2132
rect -3954 -2388 -3942 -2132
rect -4000 -2400 -3942 -2388
rect -3822 -2132 -3764 -2120
rect -3822 -2388 -3810 -2132
rect -3776 -2388 -3764 -2132
rect -3822 -2400 -3764 -2388
rect -3644 -2132 -3586 -2120
rect -3644 -2388 -3632 -2132
rect -3598 -2388 -3586 -2132
rect -3644 -2400 -3586 -2388
rect -3466 -2132 -3408 -2120
rect -3466 -2388 -3454 -2132
rect -3420 -2388 -3408 -2132
rect -3466 -2400 -3408 -2388
rect -1466 -2884 -1408 -2872
rect -6314 -3002 -6256 -2990
rect -6314 -3258 -6302 -3002
rect -6268 -3258 -6256 -3002
rect -6314 -3270 -6256 -3258
rect -6136 -3002 -6078 -2990
rect -6136 -3258 -6124 -3002
rect -6090 -3258 -6078 -3002
rect -6136 -3270 -6078 -3258
rect -5958 -3002 -5900 -2990
rect -5958 -3258 -5946 -3002
rect -5912 -3258 -5900 -3002
rect -5958 -3270 -5900 -3258
rect -5780 -3002 -5722 -2990
rect -5780 -3258 -5768 -3002
rect -5734 -3258 -5722 -3002
rect -5780 -3270 -5722 -3258
rect -5602 -3002 -5544 -2990
rect -5602 -3258 -5590 -3002
rect -5556 -3258 -5544 -3002
rect -5602 -3270 -5544 -3258
rect -5424 -3002 -5366 -2990
rect -5424 -3258 -5412 -3002
rect -5378 -3258 -5366 -3002
rect -5424 -3270 -5366 -3258
rect -5246 -3002 -5188 -2990
rect -5246 -3258 -5234 -3002
rect -5200 -3258 -5188 -3002
rect -5246 -3270 -5188 -3258
rect -5068 -3002 -5010 -2990
rect -5068 -3258 -5056 -3002
rect -5022 -3258 -5010 -3002
rect -5068 -3270 -5010 -3258
rect -4890 -3002 -4832 -2990
rect -4890 -3258 -4878 -3002
rect -4844 -3258 -4832 -3002
rect -4890 -3270 -4832 -3258
rect -4712 -3002 -4654 -2990
rect -4712 -3258 -4700 -3002
rect -4666 -3258 -4654 -3002
rect -4712 -3270 -4654 -3258
rect -4534 -3002 -4476 -2990
rect -4534 -3258 -4522 -3002
rect -4488 -3258 -4476 -3002
rect -4534 -3270 -4476 -3258
rect -4356 -3002 -4298 -2990
rect -4356 -3258 -4344 -3002
rect -4310 -3258 -4298 -3002
rect -4356 -3270 -4298 -3258
rect -4178 -3002 -4120 -2990
rect -4178 -3258 -4166 -3002
rect -4132 -3258 -4120 -3002
rect -4178 -3270 -4120 -3258
rect -4000 -3002 -3942 -2990
rect -4000 -3258 -3988 -3002
rect -3954 -3258 -3942 -3002
rect -4000 -3270 -3942 -3258
rect -3822 -3002 -3764 -2990
rect -3822 -3258 -3810 -3002
rect -3776 -3258 -3764 -3002
rect -3822 -3270 -3764 -3258
rect -3644 -3002 -3586 -2990
rect -3644 -3258 -3632 -3002
rect -3598 -3258 -3586 -3002
rect -3644 -3270 -3586 -3258
rect -3466 -3002 -3408 -2990
rect -3466 -3258 -3454 -3002
rect -3420 -3258 -3408 -3002
rect -1466 -3140 -1454 -2884
rect -1420 -3140 -1408 -2884
rect -1466 -3152 -1408 -3140
rect -1288 -2884 -1230 -2872
rect -1288 -3140 -1276 -2884
rect -1242 -3140 -1230 -2884
rect -1288 -3152 -1230 -3140
rect -1110 -2884 -1052 -2872
rect -1110 -3140 -1098 -2884
rect -1064 -3140 -1052 -2884
rect -1110 -3152 -1052 -3140
rect -932 -2884 -874 -2872
rect -932 -3140 -920 -2884
rect -886 -3140 -874 -2884
rect -932 -3152 -874 -3140
rect -754 -2884 -696 -2872
rect -754 -3140 -742 -2884
rect -708 -3140 -696 -2884
rect -754 -3152 -696 -3140
rect -576 -2884 -518 -2872
rect -576 -3140 -564 -2884
rect -530 -3140 -518 -2884
rect -576 -3152 -518 -3140
rect -398 -2884 -340 -2872
rect -398 -3140 -386 -2884
rect -352 -3140 -340 -2884
rect -398 -3152 -340 -3140
rect -220 -2884 -162 -2872
rect -220 -3140 -208 -2884
rect -174 -3140 -162 -2884
rect -220 -3152 -162 -3140
rect -42 -2884 16 -2872
rect -42 -3140 -30 -2884
rect 4 -3140 16 -2884
rect -42 -3152 16 -3140
rect 136 -2884 194 -2872
rect 136 -3140 148 -2884
rect 182 -3140 194 -2884
rect 136 -3152 194 -3140
rect 314 -2884 372 -2872
rect 314 -3140 326 -2884
rect 360 -3140 372 -2884
rect 314 -3152 372 -3140
rect 492 -2884 550 -2872
rect 492 -3140 504 -2884
rect 538 -3140 550 -2884
rect 492 -3152 550 -3140
rect 670 -2884 728 -2872
rect 670 -3140 682 -2884
rect 716 -3140 728 -2884
rect 670 -3152 728 -3140
rect 848 -2884 906 -2872
rect 848 -3140 860 -2884
rect 894 -3140 906 -2884
rect 848 -3152 906 -3140
rect 1026 -2884 1084 -2872
rect 1026 -3140 1038 -2884
rect 1072 -3140 1084 -2884
rect 1026 -3152 1084 -3140
rect 1204 -2884 1262 -2872
rect 1204 -3140 1216 -2884
rect 1250 -3140 1262 -2884
rect 1204 -3152 1262 -3140
rect 1382 -2884 1440 -2872
rect 1382 -3140 1394 -2884
rect 1428 -3140 1440 -2884
rect 1382 -3152 1440 -3140
rect 1560 -2884 1618 -2872
rect 1560 -3140 1572 -2884
rect 1606 -3140 1618 -2884
rect 1560 -3152 1618 -3140
rect 1738 -2884 1796 -2872
rect 1738 -3140 1750 -2884
rect 1784 -3140 1796 -2884
rect 1738 -3152 1796 -3140
rect 1916 -2884 1974 -2872
rect 1916 -3140 1928 -2884
rect 1962 -3140 1974 -2884
rect 1916 -3152 1974 -3140
rect 2094 -2884 2152 -2872
rect 2094 -3140 2106 -2884
rect 2140 -3140 2152 -2884
rect 2094 -3152 2152 -3140
rect 2272 -2884 2330 -2872
rect 2272 -3140 2284 -2884
rect 2318 -3140 2330 -2884
rect 2272 -3152 2330 -3140
rect 2450 -2884 2508 -2872
rect 2450 -3140 2462 -2884
rect 2496 -3140 2508 -2884
rect 2450 -3152 2508 -3140
rect 2628 -2884 2686 -2872
rect 2628 -3140 2640 -2884
rect 2674 -3140 2686 -2884
rect 2628 -3152 2686 -3140
rect -3466 -3270 -3408 -3258
rect -1466 -3784 -1408 -3772
rect -6314 -3872 -6256 -3860
rect -6314 -4128 -6302 -3872
rect -6268 -4128 -6256 -3872
rect -6314 -4140 -6256 -4128
rect -6136 -3872 -6078 -3860
rect -6136 -4128 -6124 -3872
rect -6090 -4128 -6078 -3872
rect -6136 -4140 -6078 -4128
rect -5958 -3872 -5900 -3860
rect -5958 -4128 -5946 -3872
rect -5912 -4128 -5900 -3872
rect -5958 -4140 -5900 -4128
rect -5780 -3872 -5722 -3860
rect -5780 -4128 -5768 -3872
rect -5734 -4128 -5722 -3872
rect -5780 -4140 -5722 -4128
rect -5602 -3872 -5544 -3860
rect -5602 -4128 -5590 -3872
rect -5556 -4128 -5544 -3872
rect -5602 -4140 -5544 -4128
rect -5424 -3872 -5366 -3860
rect -5424 -4128 -5412 -3872
rect -5378 -4128 -5366 -3872
rect -5424 -4140 -5366 -4128
rect -5246 -3872 -5188 -3860
rect -5246 -4128 -5234 -3872
rect -5200 -4128 -5188 -3872
rect -5246 -4140 -5188 -4128
rect -5068 -3872 -5010 -3860
rect -5068 -4128 -5056 -3872
rect -5022 -4128 -5010 -3872
rect -5068 -4140 -5010 -4128
rect -4890 -3872 -4832 -3860
rect -4890 -4128 -4878 -3872
rect -4844 -4128 -4832 -3872
rect -4890 -4140 -4832 -4128
rect -4712 -3872 -4654 -3860
rect -4712 -4128 -4700 -3872
rect -4666 -4128 -4654 -3872
rect -4712 -4140 -4654 -4128
rect -4534 -3872 -4476 -3860
rect -4534 -4128 -4522 -3872
rect -4488 -4128 -4476 -3872
rect -4534 -4140 -4476 -4128
rect -4356 -3872 -4298 -3860
rect -4356 -4128 -4344 -3872
rect -4310 -4128 -4298 -3872
rect -4356 -4140 -4298 -4128
rect -4178 -3872 -4120 -3860
rect -4178 -4128 -4166 -3872
rect -4132 -4128 -4120 -3872
rect -4178 -4140 -4120 -4128
rect -4000 -3872 -3942 -3860
rect -4000 -4128 -3988 -3872
rect -3954 -4128 -3942 -3872
rect -4000 -4140 -3942 -4128
rect -3822 -3872 -3764 -3860
rect -3822 -4128 -3810 -3872
rect -3776 -4128 -3764 -3872
rect -3822 -4140 -3764 -4128
rect -3644 -3872 -3586 -3860
rect -3644 -4128 -3632 -3872
rect -3598 -4128 -3586 -3872
rect -3644 -4140 -3586 -4128
rect -3466 -3872 -3408 -3860
rect -3466 -4128 -3454 -3872
rect -3420 -4128 -3408 -3872
rect -1466 -4040 -1454 -3784
rect -1420 -4040 -1408 -3784
rect -1466 -4052 -1408 -4040
rect -1288 -3784 -1230 -3772
rect -1288 -4040 -1276 -3784
rect -1242 -4040 -1230 -3784
rect -1288 -4052 -1230 -4040
rect -1110 -3784 -1052 -3772
rect -1110 -4040 -1098 -3784
rect -1064 -4040 -1052 -3784
rect -1110 -4052 -1052 -4040
rect -932 -3784 -874 -3772
rect -932 -4040 -920 -3784
rect -886 -4040 -874 -3784
rect -932 -4052 -874 -4040
rect -754 -3784 -696 -3772
rect -754 -4040 -742 -3784
rect -708 -4040 -696 -3784
rect -754 -4052 -696 -4040
rect -576 -3784 -518 -3772
rect -576 -4040 -564 -3784
rect -530 -4040 -518 -3784
rect -576 -4052 -518 -4040
rect -398 -3784 -340 -3772
rect -398 -4040 -386 -3784
rect -352 -4040 -340 -3784
rect -398 -4052 -340 -4040
rect -220 -3784 -162 -3772
rect -220 -4040 -208 -3784
rect -174 -4040 -162 -3784
rect -220 -4052 -162 -4040
rect -42 -3784 16 -3772
rect -42 -4040 -30 -3784
rect 4 -4040 16 -3784
rect -42 -4052 16 -4040
rect 136 -3784 194 -3772
rect 136 -4040 148 -3784
rect 182 -4040 194 -3784
rect 136 -4052 194 -4040
rect 314 -3784 372 -3772
rect 314 -4040 326 -3784
rect 360 -4040 372 -3784
rect 314 -4052 372 -4040
rect 492 -3784 550 -3772
rect 492 -4040 504 -3784
rect 538 -4040 550 -3784
rect 492 -4052 550 -4040
rect 670 -3784 728 -3772
rect 670 -4040 682 -3784
rect 716 -4040 728 -3784
rect 670 -4052 728 -4040
rect 848 -3784 906 -3772
rect 848 -4040 860 -3784
rect 894 -4040 906 -3784
rect 848 -4052 906 -4040
rect 1026 -3784 1084 -3772
rect 1026 -4040 1038 -3784
rect 1072 -4040 1084 -3784
rect 1026 -4052 1084 -4040
rect 1204 -3784 1262 -3772
rect 1204 -4040 1216 -3784
rect 1250 -4040 1262 -3784
rect 1204 -4052 1262 -4040
rect 1382 -3784 1440 -3772
rect 1382 -4040 1394 -3784
rect 1428 -4040 1440 -3784
rect 1382 -4052 1440 -4040
rect 1560 -3784 1618 -3772
rect 1560 -4040 1572 -3784
rect 1606 -4040 1618 -3784
rect 1560 -4052 1618 -4040
rect 1738 -3784 1796 -3772
rect 1738 -4040 1750 -3784
rect 1784 -4040 1796 -3784
rect 1738 -4052 1796 -4040
rect 1916 -3784 1974 -3772
rect 1916 -4040 1928 -3784
rect 1962 -4040 1974 -3784
rect 1916 -4052 1974 -4040
rect 2094 -3784 2152 -3772
rect 2094 -4040 2106 -3784
rect 2140 -4040 2152 -3784
rect 2094 -4052 2152 -4040
rect 2272 -3784 2330 -3772
rect 2272 -4040 2284 -3784
rect 2318 -4040 2330 -3784
rect 2272 -4052 2330 -4040
rect 2450 -3784 2508 -3772
rect 2450 -4040 2462 -3784
rect 2496 -4040 2508 -3784
rect 2450 -4052 2508 -4040
rect 2628 -3784 2686 -3772
rect 2628 -4040 2640 -3784
rect 2674 -4040 2686 -3784
rect 2628 -4052 2686 -4040
rect -3466 -4140 -3408 -4128
rect -1466 -4684 -1408 -4672
rect -6314 -4742 -6256 -4730
rect -6314 -4998 -6302 -4742
rect -6268 -4998 -6256 -4742
rect -6314 -5010 -6256 -4998
rect -6136 -4742 -6078 -4730
rect -6136 -4998 -6124 -4742
rect -6090 -4998 -6078 -4742
rect -6136 -5010 -6078 -4998
rect -5958 -4742 -5900 -4730
rect -5958 -4998 -5946 -4742
rect -5912 -4998 -5900 -4742
rect -5958 -5010 -5900 -4998
rect -5780 -4742 -5722 -4730
rect -5780 -4998 -5768 -4742
rect -5734 -4998 -5722 -4742
rect -5780 -5010 -5722 -4998
rect -5602 -4742 -5544 -4730
rect -5602 -4998 -5590 -4742
rect -5556 -4998 -5544 -4742
rect -5602 -5010 -5544 -4998
rect -5424 -4742 -5366 -4730
rect -5424 -4998 -5412 -4742
rect -5378 -4998 -5366 -4742
rect -5424 -5010 -5366 -4998
rect -5246 -4742 -5188 -4730
rect -5246 -4998 -5234 -4742
rect -5200 -4998 -5188 -4742
rect -5246 -5010 -5188 -4998
rect -5068 -4742 -5010 -4730
rect -5068 -4998 -5056 -4742
rect -5022 -4998 -5010 -4742
rect -5068 -5010 -5010 -4998
rect -4890 -4742 -4832 -4730
rect -4890 -4998 -4878 -4742
rect -4844 -4998 -4832 -4742
rect -4890 -5010 -4832 -4998
rect -4712 -4742 -4654 -4730
rect -4712 -4998 -4700 -4742
rect -4666 -4998 -4654 -4742
rect -4712 -5010 -4654 -4998
rect -4534 -4742 -4476 -4730
rect -4534 -4998 -4522 -4742
rect -4488 -4998 -4476 -4742
rect -4534 -5010 -4476 -4998
rect -4356 -4742 -4298 -4730
rect -4356 -4998 -4344 -4742
rect -4310 -4998 -4298 -4742
rect -4356 -5010 -4298 -4998
rect -4178 -4742 -4120 -4730
rect -4178 -4998 -4166 -4742
rect -4132 -4998 -4120 -4742
rect -4178 -5010 -4120 -4998
rect -4000 -4742 -3942 -4730
rect -4000 -4998 -3988 -4742
rect -3954 -4998 -3942 -4742
rect -4000 -5010 -3942 -4998
rect -3822 -4742 -3764 -4730
rect -3822 -4998 -3810 -4742
rect -3776 -4998 -3764 -4742
rect -3822 -5010 -3764 -4998
rect -3644 -4742 -3586 -4730
rect -3644 -4998 -3632 -4742
rect -3598 -4998 -3586 -4742
rect -3644 -5010 -3586 -4998
rect -3466 -4742 -3408 -4730
rect -3466 -4998 -3454 -4742
rect -3420 -4998 -3408 -4742
rect -1466 -4940 -1454 -4684
rect -1420 -4940 -1408 -4684
rect -1466 -4952 -1408 -4940
rect -1288 -4684 -1230 -4672
rect -1288 -4940 -1276 -4684
rect -1242 -4940 -1230 -4684
rect -1288 -4952 -1230 -4940
rect -1110 -4684 -1052 -4672
rect -1110 -4940 -1098 -4684
rect -1064 -4940 -1052 -4684
rect -1110 -4952 -1052 -4940
rect -932 -4684 -874 -4672
rect -932 -4940 -920 -4684
rect -886 -4940 -874 -4684
rect -932 -4952 -874 -4940
rect -754 -4684 -696 -4672
rect -754 -4940 -742 -4684
rect -708 -4940 -696 -4684
rect -754 -4952 -696 -4940
rect -576 -4684 -518 -4672
rect -576 -4940 -564 -4684
rect -530 -4940 -518 -4684
rect -576 -4952 -518 -4940
rect -398 -4684 -340 -4672
rect -398 -4940 -386 -4684
rect -352 -4940 -340 -4684
rect -398 -4952 -340 -4940
rect -220 -4684 -162 -4672
rect -220 -4940 -208 -4684
rect -174 -4940 -162 -4684
rect -220 -4952 -162 -4940
rect -42 -4684 16 -4672
rect -42 -4940 -30 -4684
rect 4 -4940 16 -4684
rect -42 -4952 16 -4940
rect 136 -4684 194 -4672
rect 136 -4940 148 -4684
rect 182 -4940 194 -4684
rect 136 -4952 194 -4940
rect 314 -4684 372 -4672
rect 314 -4940 326 -4684
rect 360 -4940 372 -4684
rect 314 -4952 372 -4940
rect 492 -4684 550 -4672
rect 492 -4940 504 -4684
rect 538 -4940 550 -4684
rect 492 -4952 550 -4940
rect 670 -4684 728 -4672
rect 670 -4940 682 -4684
rect 716 -4940 728 -4684
rect 670 -4952 728 -4940
rect 848 -4684 906 -4672
rect 848 -4940 860 -4684
rect 894 -4940 906 -4684
rect 848 -4952 906 -4940
rect 1026 -4684 1084 -4672
rect 1026 -4940 1038 -4684
rect 1072 -4940 1084 -4684
rect 1026 -4952 1084 -4940
rect 1204 -4684 1262 -4672
rect 1204 -4940 1216 -4684
rect 1250 -4940 1262 -4684
rect 1204 -4952 1262 -4940
rect 1382 -4684 1440 -4672
rect 1382 -4940 1394 -4684
rect 1428 -4940 1440 -4684
rect 1382 -4952 1440 -4940
rect 1560 -4684 1618 -4672
rect 1560 -4940 1572 -4684
rect 1606 -4940 1618 -4684
rect 1560 -4952 1618 -4940
rect 1738 -4684 1796 -4672
rect 1738 -4940 1750 -4684
rect 1784 -4940 1796 -4684
rect 1738 -4952 1796 -4940
rect 1916 -4684 1974 -4672
rect 1916 -4940 1928 -4684
rect 1962 -4940 1974 -4684
rect 1916 -4952 1974 -4940
rect 2094 -4684 2152 -4672
rect 2094 -4940 2106 -4684
rect 2140 -4940 2152 -4684
rect 2094 -4952 2152 -4940
rect 2272 -4684 2330 -4672
rect 2272 -4940 2284 -4684
rect 2318 -4940 2330 -4684
rect 2272 -4952 2330 -4940
rect 2450 -4684 2508 -4672
rect 2450 -4940 2462 -4684
rect 2496 -4940 2508 -4684
rect 2450 -4952 2508 -4940
rect 2628 -4684 2686 -4672
rect 2628 -4940 2640 -4684
rect 2674 -4940 2686 -4684
rect 2628 -4952 2686 -4940
rect -3466 -5010 -3408 -4998
rect -1466 -5584 -1408 -5572
rect -6314 -5612 -6256 -5600
rect -6314 -5868 -6302 -5612
rect -6268 -5868 -6256 -5612
rect -6314 -5880 -6256 -5868
rect -6136 -5612 -6078 -5600
rect -6136 -5868 -6124 -5612
rect -6090 -5868 -6078 -5612
rect -6136 -5880 -6078 -5868
rect -5958 -5612 -5900 -5600
rect -5958 -5868 -5946 -5612
rect -5912 -5868 -5900 -5612
rect -5958 -5880 -5900 -5868
rect -5780 -5612 -5722 -5600
rect -5780 -5868 -5768 -5612
rect -5734 -5868 -5722 -5612
rect -5780 -5880 -5722 -5868
rect -5602 -5612 -5544 -5600
rect -5602 -5868 -5590 -5612
rect -5556 -5868 -5544 -5612
rect -5602 -5880 -5544 -5868
rect -5424 -5612 -5366 -5600
rect -5424 -5868 -5412 -5612
rect -5378 -5868 -5366 -5612
rect -5424 -5880 -5366 -5868
rect -5246 -5612 -5188 -5600
rect -5246 -5868 -5234 -5612
rect -5200 -5868 -5188 -5612
rect -5246 -5880 -5188 -5868
rect -5068 -5612 -5010 -5600
rect -5068 -5868 -5056 -5612
rect -5022 -5868 -5010 -5612
rect -5068 -5880 -5010 -5868
rect -4890 -5612 -4832 -5600
rect -4890 -5868 -4878 -5612
rect -4844 -5868 -4832 -5612
rect -4890 -5880 -4832 -5868
rect -4712 -5612 -4654 -5600
rect -4712 -5868 -4700 -5612
rect -4666 -5868 -4654 -5612
rect -4712 -5880 -4654 -5868
rect -4534 -5612 -4476 -5600
rect -4534 -5868 -4522 -5612
rect -4488 -5868 -4476 -5612
rect -4534 -5880 -4476 -5868
rect -4356 -5612 -4298 -5600
rect -4356 -5868 -4344 -5612
rect -4310 -5868 -4298 -5612
rect -4356 -5880 -4298 -5868
rect -4178 -5612 -4120 -5600
rect -4178 -5868 -4166 -5612
rect -4132 -5868 -4120 -5612
rect -4178 -5880 -4120 -5868
rect -4000 -5612 -3942 -5600
rect -4000 -5868 -3988 -5612
rect -3954 -5868 -3942 -5612
rect -4000 -5880 -3942 -5868
rect -3822 -5612 -3764 -5600
rect -3822 -5868 -3810 -5612
rect -3776 -5868 -3764 -5612
rect -3822 -5880 -3764 -5868
rect -3644 -5612 -3586 -5600
rect -3644 -5868 -3632 -5612
rect -3598 -5868 -3586 -5612
rect -3644 -5880 -3586 -5868
rect -3466 -5612 -3408 -5600
rect -3466 -5868 -3454 -5612
rect -3420 -5868 -3408 -5612
rect -1466 -5840 -1454 -5584
rect -1420 -5840 -1408 -5584
rect -1466 -5852 -1408 -5840
rect -1288 -5584 -1230 -5572
rect -1288 -5840 -1276 -5584
rect -1242 -5840 -1230 -5584
rect -1288 -5852 -1230 -5840
rect -1110 -5584 -1052 -5572
rect -1110 -5840 -1098 -5584
rect -1064 -5840 -1052 -5584
rect -1110 -5852 -1052 -5840
rect -932 -5584 -874 -5572
rect -932 -5840 -920 -5584
rect -886 -5840 -874 -5584
rect -932 -5852 -874 -5840
rect -754 -5584 -696 -5572
rect -754 -5840 -742 -5584
rect -708 -5840 -696 -5584
rect -754 -5852 -696 -5840
rect -576 -5584 -518 -5572
rect -576 -5840 -564 -5584
rect -530 -5840 -518 -5584
rect -576 -5852 -518 -5840
rect -398 -5584 -340 -5572
rect -398 -5840 -386 -5584
rect -352 -5840 -340 -5584
rect -398 -5852 -340 -5840
rect -220 -5584 -162 -5572
rect -220 -5840 -208 -5584
rect -174 -5840 -162 -5584
rect -220 -5852 -162 -5840
rect -42 -5584 16 -5572
rect -42 -5840 -30 -5584
rect 4 -5840 16 -5584
rect -42 -5852 16 -5840
rect 136 -5584 194 -5572
rect 136 -5840 148 -5584
rect 182 -5840 194 -5584
rect 136 -5852 194 -5840
rect 314 -5584 372 -5572
rect 314 -5840 326 -5584
rect 360 -5840 372 -5584
rect 314 -5852 372 -5840
rect 492 -5584 550 -5572
rect 492 -5840 504 -5584
rect 538 -5840 550 -5584
rect 492 -5852 550 -5840
rect 670 -5584 728 -5572
rect 670 -5840 682 -5584
rect 716 -5840 728 -5584
rect 670 -5852 728 -5840
rect 848 -5584 906 -5572
rect 848 -5840 860 -5584
rect 894 -5840 906 -5584
rect 848 -5852 906 -5840
rect 1026 -5584 1084 -5572
rect 1026 -5840 1038 -5584
rect 1072 -5840 1084 -5584
rect 1026 -5852 1084 -5840
rect 1204 -5584 1262 -5572
rect 1204 -5840 1216 -5584
rect 1250 -5840 1262 -5584
rect 1204 -5852 1262 -5840
rect 1382 -5584 1440 -5572
rect 1382 -5840 1394 -5584
rect 1428 -5840 1440 -5584
rect 1382 -5852 1440 -5840
rect 1560 -5584 1618 -5572
rect 1560 -5840 1572 -5584
rect 1606 -5840 1618 -5584
rect 1560 -5852 1618 -5840
rect 1738 -5584 1796 -5572
rect 1738 -5840 1750 -5584
rect 1784 -5840 1796 -5584
rect 1738 -5852 1796 -5840
rect 1916 -5584 1974 -5572
rect 1916 -5840 1928 -5584
rect 1962 -5840 1974 -5584
rect 1916 -5852 1974 -5840
rect 2094 -5584 2152 -5572
rect 2094 -5840 2106 -5584
rect 2140 -5840 2152 -5584
rect 2094 -5852 2152 -5840
rect 2272 -5584 2330 -5572
rect 2272 -5840 2284 -5584
rect 2318 -5840 2330 -5584
rect 2272 -5852 2330 -5840
rect 2450 -5584 2508 -5572
rect 2450 -5840 2462 -5584
rect 2496 -5840 2508 -5584
rect 2450 -5852 2508 -5840
rect 2628 -5584 2686 -5572
rect 2628 -5840 2640 -5584
rect 2674 -5840 2686 -5584
rect 2628 -5852 2686 -5840
rect -3466 -5880 -3408 -5868
rect 7142 -2787 7204 -2775
rect 7142 -3035 7154 -2787
rect 7188 -3035 7204 -2787
rect 7142 -3047 7204 -3035
rect 7234 -2787 7300 -2775
rect 7234 -3035 7250 -2787
rect 7284 -3035 7300 -2787
rect 7234 -3047 7300 -3035
rect 7330 -2787 7396 -2775
rect 7330 -3035 7346 -2787
rect 7380 -3035 7396 -2787
rect 7330 -3047 7396 -3035
rect 7426 -2787 7492 -2775
rect 7426 -3035 7442 -2787
rect 7476 -3035 7492 -2787
rect 7426 -3047 7492 -3035
rect 7522 -2787 7588 -2775
rect 7522 -3035 7538 -2787
rect 7572 -3035 7588 -2787
rect 7522 -3047 7588 -3035
rect 7618 -2787 7684 -2775
rect 7618 -3035 7634 -2787
rect 7668 -3035 7684 -2787
rect 7618 -3047 7684 -3035
rect 7714 -2787 7780 -2775
rect 7714 -3035 7730 -2787
rect 7764 -3035 7780 -2787
rect 7714 -3047 7780 -3035
rect 7810 -2787 7876 -2775
rect 7810 -3035 7826 -2787
rect 7860 -3035 7876 -2787
rect 7810 -3047 7876 -3035
rect 7906 -2787 7972 -2775
rect 7906 -3035 7922 -2787
rect 7956 -3035 7972 -2787
rect 7906 -3047 7972 -3035
rect 8002 -2787 8068 -2775
rect 8002 -3035 8018 -2787
rect 8052 -3035 8068 -2787
rect 8002 -3047 8068 -3035
rect 8098 -2787 8160 -2775
rect 8098 -3035 8114 -2787
rect 8148 -3035 8160 -2787
rect 8098 -3047 8160 -3035
rect 16142 -2787 16204 -2775
rect 16142 -3035 16154 -2787
rect 16188 -3035 16204 -2787
rect 16142 -3047 16204 -3035
rect 16234 -2787 16300 -2775
rect 16234 -3035 16250 -2787
rect 16284 -3035 16300 -2787
rect 16234 -3047 16300 -3035
rect 16330 -2787 16396 -2775
rect 16330 -3035 16346 -2787
rect 16380 -3035 16396 -2787
rect 16330 -3047 16396 -3035
rect 16426 -2787 16492 -2775
rect 16426 -3035 16442 -2787
rect 16476 -3035 16492 -2787
rect 16426 -3047 16492 -3035
rect 16522 -2787 16588 -2775
rect 16522 -3035 16538 -2787
rect 16572 -3035 16588 -2787
rect 16522 -3047 16588 -3035
rect 16618 -2787 16684 -2775
rect 16618 -3035 16634 -2787
rect 16668 -3035 16684 -2787
rect 16618 -3047 16684 -3035
rect 16714 -2787 16780 -2775
rect 16714 -3035 16730 -2787
rect 16764 -3035 16780 -2787
rect 16714 -3047 16780 -3035
rect 16810 -2787 16876 -2775
rect 16810 -3035 16826 -2787
rect 16860 -3035 16876 -2787
rect 16810 -3047 16876 -3035
rect 16906 -2787 16972 -2775
rect 16906 -3035 16922 -2787
rect 16956 -3035 16972 -2787
rect 16906 -3047 16972 -3035
rect 17002 -2787 17068 -2775
rect 17002 -3035 17018 -2787
rect 17052 -3035 17068 -2787
rect 17002 -3047 17068 -3035
rect 17098 -2787 17160 -2775
rect 17098 -3035 17114 -2787
rect 17148 -3035 17160 -2787
rect 17098 -3047 17160 -3035
rect 7142 -4587 7204 -4575
rect 7142 -4835 7154 -4587
rect 7188 -4835 7204 -4587
rect 7142 -4847 7204 -4835
rect 7234 -4587 7300 -4575
rect 7234 -4835 7250 -4587
rect 7284 -4835 7300 -4587
rect 7234 -4847 7300 -4835
rect 7330 -4587 7396 -4575
rect 7330 -4835 7346 -4587
rect 7380 -4835 7396 -4587
rect 7330 -4847 7396 -4835
rect 7426 -4587 7492 -4575
rect 7426 -4835 7442 -4587
rect 7476 -4835 7492 -4587
rect 7426 -4847 7492 -4835
rect 7522 -4587 7588 -4575
rect 7522 -4835 7538 -4587
rect 7572 -4835 7588 -4587
rect 7522 -4847 7588 -4835
rect 7618 -4587 7684 -4575
rect 7618 -4835 7634 -4587
rect 7668 -4835 7684 -4587
rect 7618 -4847 7684 -4835
rect 7714 -4587 7780 -4575
rect 7714 -4835 7730 -4587
rect 7764 -4835 7780 -4587
rect 7714 -4847 7780 -4835
rect 7810 -4587 7876 -4575
rect 7810 -4835 7826 -4587
rect 7860 -4835 7876 -4587
rect 7810 -4847 7876 -4835
rect 7906 -4587 7972 -4575
rect 7906 -4835 7922 -4587
rect 7956 -4835 7972 -4587
rect 7906 -4847 7972 -4835
rect 8002 -4587 8068 -4575
rect 8002 -4835 8018 -4587
rect 8052 -4835 8068 -4587
rect 8002 -4847 8068 -4835
rect 8098 -4587 8160 -4575
rect 8098 -4835 8114 -4587
rect 8148 -4835 8160 -4587
rect 8098 -4847 8160 -4835
rect 16142 -4587 16204 -4575
rect 16142 -4835 16154 -4587
rect 16188 -4835 16204 -4587
rect 16142 -4847 16204 -4835
rect 16234 -4587 16300 -4575
rect 16234 -4835 16250 -4587
rect 16284 -4835 16300 -4587
rect 16234 -4847 16300 -4835
rect 16330 -4587 16396 -4575
rect 16330 -4835 16346 -4587
rect 16380 -4835 16396 -4587
rect 16330 -4847 16396 -4835
rect 16426 -4587 16492 -4575
rect 16426 -4835 16442 -4587
rect 16476 -4835 16492 -4587
rect 16426 -4847 16492 -4835
rect 16522 -4587 16588 -4575
rect 16522 -4835 16538 -4587
rect 16572 -4835 16588 -4587
rect 16522 -4847 16588 -4835
rect 16618 -4587 16684 -4575
rect 16618 -4835 16634 -4587
rect 16668 -4835 16684 -4587
rect 16618 -4847 16684 -4835
rect 16714 -4587 16780 -4575
rect 16714 -4835 16730 -4587
rect 16764 -4835 16780 -4587
rect 16714 -4847 16780 -4835
rect 16810 -4587 16876 -4575
rect 16810 -4835 16826 -4587
rect 16860 -4835 16876 -4587
rect 16810 -4847 16876 -4835
rect 16906 -4587 16972 -4575
rect 16906 -4835 16922 -4587
rect 16956 -4835 16972 -4587
rect 16906 -4847 16972 -4835
rect 17002 -4587 17068 -4575
rect 17002 -4835 17018 -4587
rect 17052 -4835 17068 -4587
rect 17002 -4847 17068 -4835
rect 17098 -4587 17160 -4575
rect 17098 -4835 17114 -4587
rect 17148 -4835 17160 -4587
rect 17098 -4847 17160 -4835
rect 7142 -6387 7204 -6375
rect 7142 -6635 7154 -6387
rect 7188 -6635 7204 -6387
rect 7142 -6647 7204 -6635
rect 7234 -6387 7300 -6375
rect 7234 -6635 7250 -6387
rect 7284 -6635 7300 -6387
rect 7234 -6647 7300 -6635
rect 7330 -6387 7396 -6375
rect 7330 -6635 7346 -6387
rect 7380 -6635 7396 -6387
rect 7330 -6647 7396 -6635
rect 7426 -6387 7492 -6375
rect 7426 -6635 7442 -6387
rect 7476 -6635 7492 -6387
rect 7426 -6647 7492 -6635
rect 7522 -6387 7588 -6375
rect 7522 -6635 7538 -6387
rect 7572 -6635 7588 -6387
rect 7522 -6647 7588 -6635
rect 7618 -6387 7684 -6375
rect 7618 -6635 7634 -6387
rect 7668 -6635 7684 -6387
rect 7618 -6647 7684 -6635
rect 7714 -6387 7780 -6375
rect 7714 -6635 7730 -6387
rect 7764 -6635 7780 -6387
rect 7714 -6647 7780 -6635
rect 7810 -6387 7876 -6375
rect 7810 -6635 7826 -6387
rect 7860 -6635 7876 -6387
rect 7810 -6647 7876 -6635
rect 7906 -6387 7972 -6375
rect 7906 -6635 7922 -6387
rect 7956 -6635 7972 -6387
rect 7906 -6647 7972 -6635
rect 8002 -6387 8068 -6375
rect 8002 -6635 8018 -6387
rect 8052 -6635 8068 -6387
rect 8002 -6647 8068 -6635
rect 8098 -6387 8160 -6375
rect 8098 -6635 8114 -6387
rect 8148 -6635 8160 -6387
rect 8098 -6647 8160 -6635
rect 16142 -6387 16204 -6375
rect 16142 -6635 16154 -6387
rect 16188 -6635 16204 -6387
rect 16142 -6647 16204 -6635
rect 16234 -6387 16300 -6375
rect 16234 -6635 16250 -6387
rect 16284 -6635 16300 -6387
rect 16234 -6647 16300 -6635
rect 16330 -6387 16396 -6375
rect 16330 -6635 16346 -6387
rect 16380 -6635 16396 -6387
rect 16330 -6647 16396 -6635
rect 16426 -6387 16492 -6375
rect 16426 -6635 16442 -6387
rect 16476 -6635 16492 -6387
rect 16426 -6647 16492 -6635
rect 16522 -6387 16588 -6375
rect 16522 -6635 16538 -6387
rect 16572 -6635 16588 -6387
rect 16522 -6647 16588 -6635
rect 16618 -6387 16684 -6375
rect 16618 -6635 16634 -6387
rect 16668 -6635 16684 -6387
rect 16618 -6647 16684 -6635
rect 16714 -6387 16780 -6375
rect 16714 -6635 16730 -6387
rect 16764 -6635 16780 -6387
rect 16714 -6647 16780 -6635
rect 16810 -6387 16876 -6375
rect 16810 -6635 16826 -6387
rect 16860 -6635 16876 -6387
rect 16810 -6647 16876 -6635
rect 16906 -6387 16972 -6375
rect 16906 -6635 16922 -6387
rect 16956 -6635 16972 -6387
rect 16906 -6647 16972 -6635
rect 17002 -6387 17068 -6375
rect 17002 -6635 17018 -6387
rect 17052 -6635 17068 -6387
rect 17002 -6647 17068 -6635
rect 17098 -6387 17160 -6375
rect 17098 -6635 17114 -6387
rect 17148 -6635 17160 -6387
rect 17098 -6647 17160 -6635
<< ndiffc >>
rect 7154 1953 7188 2033
rect 7250 1953 7284 2033
rect 7346 1953 7380 2033
rect 7442 1953 7476 2033
rect 7538 1953 7572 2033
rect 7634 1953 7668 2033
rect 7730 1953 7764 2033
rect 7826 1953 7860 2033
rect 7922 1953 7956 2033
rect 8018 1953 8052 2033
rect 8114 1953 8148 2033
rect 16154 1953 16188 2033
rect 16250 1953 16284 2033
rect 16346 1953 16380 2033
rect 16442 1953 16476 2033
rect 16538 1953 16572 2033
rect 16634 1953 16668 2033
rect 16730 1953 16764 2033
rect 16826 1953 16860 2033
rect 16922 1953 16956 2033
rect 17018 1953 17052 2033
rect 17114 1953 17148 2033
rect 7154 153 7188 233
rect 7250 153 7284 233
rect 7346 153 7380 233
rect 7442 153 7476 233
rect 7538 153 7572 233
rect 7634 153 7668 233
rect 7730 153 7764 233
rect 7826 153 7860 233
rect 7922 153 7956 233
rect 8018 153 8052 233
rect 8114 153 8148 233
rect 16154 153 16188 233
rect 16250 153 16284 233
rect 16346 153 16380 233
rect 16442 153 16476 233
rect 16538 153 16572 233
rect 16634 153 16668 233
rect 16730 153 16764 233
rect 16826 153 16860 233
rect 16922 153 16956 233
rect 17018 153 17052 233
rect 17114 153 17148 233
rect 7154 -1647 7188 -1567
rect 7250 -1647 7284 -1567
rect 7346 -1647 7380 -1567
rect 7442 -1647 7476 -1567
rect 7538 -1647 7572 -1567
rect 7634 -1647 7668 -1567
rect 7730 -1647 7764 -1567
rect 7826 -1647 7860 -1567
rect 7922 -1647 7956 -1567
rect 8018 -1647 8052 -1567
rect 8114 -1647 8148 -1567
rect 16154 -1647 16188 -1567
rect 16250 -1647 16284 -1567
rect 16346 -1647 16380 -1567
rect 16442 -1647 16476 -1567
rect 16538 -1647 16572 -1567
rect 16634 -1647 16668 -1567
rect 16730 -1647 16764 -1567
rect 16826 -1647 16860 -1567
rect 16922 -1647 16956 -1567
rect 17018 -1647 17052 -1567
rect 17114 -1647 17148 -1567
rect 7154 -3447 7188 -3367
rect 7250 -3447 7284 -3367
rect 7346 -3447 7380 -3367
rect 7442 -3447 7476 -3367
rect 7538 -3447 7572 -3367
rect 7634 -3447 7668 -3367
rect 7730 -3447 7764 -3367
rect 7826 -3447 7860 -3367
rect 7922 -3447 7956 -3367
rect 8018 -3447 8052 -3367
rect 8114 -3447 8148 -3367
rect 16154 -3447 16188 -3367
rect 16250 -3447 16284 -3367
rect 16346 -3447 16380 -3367
rect 16442 -3447 16476 -3367
rect 16538 -3447 16572 -3367
rect 16634 -3447 16668 -3367
rect 16730 -3447 16764 -3367
rect 16826 -3447 16860 -3367
rect 16922 -3447 16956 -3367
rect 17018 -3447 17052 -3367
rect 17114 -3447 17148 -3367
rect 7154 -5247 7188 -5167
rect 7250 -5247 7284 -5167
rect 7346 -5247 7380 -5167
rect 7442 -5247 7476 -5167
rect 7538 -5247 7572 -5167
rect 7634 -5247 7668 -5167
rect 7730 -5247 7764 -5167
rect 7826 -5247 7860 -5167
rect 7922 -5247 7956 -5167
rect 8018 -5247 8052 -5167
rect 8114 -5247 8148 -5167
rect 16154 -5247 16188 -5167
rect 16250 -5247 16284 -5167
rect 16346 -5247 16380 -5167
rect 16442 -5247 16476 -5167
rect 16538 -5247 16572 -5167
rect 16634 -5247 16668 -5167
rect 16730 -5247 16764 -5167
rect 16826 -5247 16860 -5167
rect 16922 -5247 16956 -5167
rect 17018 -5247 17052 -5167
rect 17114 -5247 17148 -5167
rect 7154 -7047 7188 -6967
rect 7250 -7047 7284 -6967
rect 7346 -7047 7380 -6967
rect 7442 -7047 7476 -6967
rect 7538 -7047 7572 -6967
rect 7634 -7047 7668 -6967
rect 7730 -7047 7764 -6967
rect 7826 -7047 7860 -6967
rect 7922 -7047 7956 -6967
rect 8018 -7047 8052 -6967
rect 8114 -7047 8148 -6967
rect 16154 -7047 16188 -6967
rect 16250 -7047 16284 -6967
rect 16346 -7047 16380 -6967
rect 16442 -7047 16476 -6967
rect 16538 -7047 16572 -6967
rect 16634 -7047 16668 -6967
rect 16730 -7047 16764 -6967
rect 16826 -7047 16860 -6967
rect 16922 -7047 16956 -6967
rect 17018 -7047 17052 -6967
rect 17114 -7047 17148 -6967
rect -5628 -8130 -5594 -7874
rect -5450 -8130 -5416 -7874
rect -5272 -8130 -5238 -7874
rect -5094 -8130 -5060 -7874
rect -4916 -8130 -4882 -7874
rect -4738 -8130 -4704 -7874
rect -4560 -8130 -4526 -7874
rect -4382 -8130 -4348 -7874
rect -4204 -8130 -4170 -7874
rect -4026 -8130 -3992 -7874
rect -2173 -8388 -2139 -8132
rect -1995 -8388 -1961 -8132
rect -1817 -8388 -1783 -8132
rect -1639 -8388 -1605 -8132
rect -1461 -8388 -1427 -8132
rect -1283 -8388 -1249 -8132
rect -1105 -8388 -1071 -8132
rect -927 -8388 -893 -8132
rect -749 -8388 -715 -8132
rect -571 -8388 -537 -8132
rect -393 -8388 -359 -8132
rect -215 -8388 -181 -8132
rect -37 -8388 -3 -8132
rect 141 -8388 175 -8132
rect 319 -8388 353 -8132
rect 497 -8388 531 -8132
rect 675 -8388 709 -8132
rect 853 -8388 887 -8132
rect 1031 -8388 1065 -8132
rect 1209 -8388 1243 -8132
rect 1387 -8388 1421 -8132
rect 1565 -8388 1599 -8132
rect 1743 -8388 1777 -8132
rect 1921 -8388 1955 -8132
rect 2099 -8388 2133 -8132
rect 2277 -8388 2311 -8132
rect 2455 -8388 2489 -8132
rect 2633 -8388 2667 -8132
rect 2811 -8388 2845 -8132
rect 2989 -8388 3023 -8132
rect 3167 -8388 3201 -8132
rect 3345 -8388 3379 -8132
rect 3523 -8388 3557 -8132
rect 3701 -8388 3735 -8132
rect 3879 -8388 3913 -8132
rect 4057 -8388 4091 -8132
rect -5628 -8680 -5594 -8424
rect -5450 -8680 -5416 -8424
rect -5272 -8680 -5238 -8424
rect -5094 -8680 -5060 -8424
rect -4916 -8680 -4882 -8424
rect -4738 -8680 -4704 -8424
rect -4560 -8680 -4526 -8424
rect -4382 -8680 -4348 -8424
rect -4204 -8680 -4170 -8424
rect -4026 -8680 -3992 -8424
rect -5628 -9230 -5594 -8974
rect -5450 -9230 -5416 -8974
rect -5272 -9230 -5238 -8974
rect -5094 -9230 -5060 -8974
rect -4916 -9230 -4882 -8974
rect -4738 -9230 -4704 -8974
rect -4560 -9230 -4526 -8974
rect -4382 -9230 -4348 -8974
rect -4204 -9230 -4170 -8974
rect -4026 -9230 -3992 -8974
rect -2173 -9388 -2139 -9132
rect -1995 -9388 -1961 -9132
rect -1817 -9388 -1783 -9132
rect -1639 -9388 -1605 -9132
rect -1461 -9388 -1427 -9132
rect -1283 -9388 -1249 -9132
rect -1105 -9388 -1071 -9132
rect -927 -9388 -893 -9132
rect -749 -9388 -715 -9132
rect -571 -9388 -537 -9132
rect -393 -9388 -359 -9132
rect -215 -9388 -181 -9132
rect -37 -9388 -3 -9132
rect 141 -9388 175 -9132
rect 319 -9388 353 -9132
rect 497 -9388 531 -9132
rect 675 -9388 709 -9132
rect 853 -9388 887 -9132
rect 1031 -9388 1065 -9132
rect 1209 -9388 1243 -9132
rect 1387 -9388 1421 -9132
rect 1565 -9388 1599 -9132
rect 1743 -9388 1777 -9132
rect 1921 -9388 1955 -9132
rect 2099 -9388 2133 -9132
rect 2277 -9388 2311 -9132
rect 2455 -9388 2489 -9132
rect 2633 -9388 2667 -9132
rect 2811 -9388 2845 -9132
rect 2989 -9388 3023 -9132
rect 3167 -9388 3201 -9132
rect 3345 -9388 3379 -9132
rect 3523 -9388 3557 -9132
rect 3701 -9388 3735 -9132
rect 3879 -9388 3913 -9132
rect 4057 -9388 4091 -9132
rect 6512 -9150 6546 -8894
rect 6690 -9150 6724 -8894
rect 6868 -9150 6902 -8894
rect 7046 -9150 7080 -8894
rect 7224 -9150 7258 -8894
rect 7402 -9150 7436 -8894
rect 7580 -9150 7614 -8894
rect 7758 -9150 7792 -8894
rect 7936 -9150 7970 -8894
rect 8114 -9150 8148 -8894
rect 8292 -9150 8326 -8894
rect 8470 -9150 8504 -8894
rect 8648 -9150 8682 -8894
rect 8826 -9150 8860 -8894
rect 9004 -9150 9038 -8894
rect 9182 -9150 9216 -8894
rect 9360 -9150 9394 -8894
rect 10772 -9180 10806 -8924
rect 10950 -9180 10984 -8924
rect 11064 -9180 11098 -8924
rect 11242 -9180 11276 -8924
rect 11356 -9180 11390 -8924
rect 11534 -9180 11568 -8924
rect 11648 -9180 11682 -8924
rect 11826 -9180 11860 -8924
rect 11940 -9180 11974 -8924
rect 12118 -9180 12152 -8924
rect 12232 -9180 12266 -8924
rect 12410 -9180 12444 -8924
rect 12524 -9180 12558 -8924
rect 12702 -9180 12736 -8924
rect -5628 -9780 -5594 -9524
rect -5450 -9780 -5416 -9524
rect -5272 -9780 -5238 -9524
rect -5094 -9780 -5060 -9524
rect -4916 -9780 -4882 -9524
rect -4738 -9780 -4704 -9524
rect -4560 -9780 -4526 -9524
rect -4382 -9780 -4348 -9524
rect -4204 -9780 -4170 -9524
rect -4026 -9780 -3992 -9524
rect -5628 -10330 -5594 -10074
rect -5450 -10330 -5416 -10074
rect -5272 -10330 -5238 -10074
rect -5094 -10330 -5060 -10074
rect -4916 -10330 -4882 -10074
rect -4738 -10330 -4704 -10074
rect -4560 -10330 -4526 -10074
rect -4382 -10330 -4348 -10074
rect -4204 -10330 -4170 -10074
rect -4026 -10330 -3992 -10074
rect 6512 -10050 6546 -9794
rect 6690 -10050 6724 -9794
rect 6868 -10050 6902 -9794
rect 7046 -10050 7080 -9794
rect 7224 -10050 7258 -9794
rect 7402 -10050 7436 -9794
rect 7580 -10050 7614 -9794
rect 7758 -10050 7792 -9794
rect 7936 -10050 7970 -9794
rect 8114 -10050 8148 -9794
rect 8292 -10050 8326 -9794
rect 8470 -10050 8504 -9794
rect 8648 -10050 8682 -9794
rect 8826 -10050 8860 -9794
rect 9004 -10050 9038 -9794
rect 9182 -10050 9216 -9794
rect 9360 -10050 9394 -9794
rect 10772 -9950 10806 -9694
rect 10950 -9950 10984 -9694
rect 11064 -9950 11098 -9694
rect 11242 -9950 11276 -9694
rect 11356 -9950 11390 -9694
rect 11534 -9950 11568 -9694
rect 11648 -9950 11682 -9694
rect 11826 -9950 11860 -9694
rect 11940 -9950 11974 -9694
rect 12118 -9950 12152 -9694
rect 12232 -9950 12266 -9694
rect 12410 -9950 12444 -9694
rect 12524 -9950 12558 -9694
rect 12702 -9950 12736 -9694
rect -2173 -10388 -2139 -10132
rect -1995 -10388 -1961 -10132
rect -1817 -10388 -1783 -10132
rect -1639 -10388 -1605 -10132
rect -1461 -10388 -1427 -10132
rect -1283 -10388 -1249 -10132
rect -1105 -10388 -1071 -10132
rect -927 -10388 -893 -10132
rect -749 -10388 -715 -10132
rect -571 -10388 -537 -10132
rect -393 -10388 -359 -10132
rect -215 -10388 -181 -10132
rect -37 -10388 -3 -10132
rect 141 -10388 175 -10132
rect 319 -10388 353 -10132
rect 497 -10388 531 -10132
rect 675 -10388 709 -10132
rect 853 -10388 887 -10132
rect 1031 -10388 1065 -10132
rect 1209 -10388 1243 -10132
rect 1387 -10388 1421 -10132
rect 1565 -10388 1599 -10132
rect 1743 -10388 1777 -10132
rect 1921 -10388 1955 -10132
rect 2099 -10388 2133 -10132
rect 2277 -10388 2311 -10132
rect 2455 -10388 2489 -10132
rect 2633 -10388 2667 -10132
rect 2811 -10388 2845 -10132
rect 2989 -10388 3023 -10132
rect 3167 -10388 3201 -10132
rect 3345 -10388 3379 -10132
rect 3523 -10388 3557 -10132
rect 3701 -10388 3735 -10132
rect 3879 -10388 3913 -10132
rect 4057 -10388 4091 -10132
rect -5628 -10880 -5594 -10624
rect -5450 -10880 -5416 -10624
rect -5272 -10880 -5238 -10624
rect -5094 -10880 -5060 -10624
rect -4916 -10880 -4882 -10624
rect -4738 -10880 -4704 -10624
rect -4560 -10880 -4526 -10624
rect -4382 -10880 -4348 -10624
rect -4204 -10880 -4170 -10624
rect -4026 -10880 -3992 -10624
rect 6512 -10950 6546 -10694
rect 6690 -10950 6724 -10694
rect 6868 -10950 6902 -10694
rect 7046 -10950 7080 -10694
rect 7224 -10950 7258 -10694
rect 7402 -10950 7436 -10694
rect 7580 -10950 7614 -10694
rect 7758 -10950 7792 -10694
rect 7936 -10950 7970 -10694
rect 8114 -10950 8148 -10694
rect 8292 -10950 8326 -10694
rect 8470 -10950 8504 -10694
rect 8648 -10950 8682 -10694
rect 8826 -10950 8860 -10694
rect 9004 -10950 9038 -10694
rect 9182 -10950 9216 -10694
rect 9360 -10950 9394 -10694
rect 10772 -10720 10806 -10464
rect 10950 -10720 10984 -10464
rect 11064 -10720 11098 -10464
rect 11242 -10720 11276 -10464
rect 11356 -10720 11390 -10464
rect 11534 -10720 11568 -10464
rect 11648 -10720 11682 -10464
rect 11826 -10720 11860 -10464
rect 11940 -10720 11974 -10464
rect 12118 -10720 12152 -10464
rect 12232 -10720 12266 -10464
rect 12410 -10720 12444 -10464
rect 12524 -10720 12558 -10464
rect 12702 -10720 12736 -10464
rect -5628 -11430 -5594 -11174
rect -5450 -11430 -5416 -11174
rect -5272 -11430 -5238 -11174
rect -5094 -11430 -5060 -11174
rect -4916 -11430 -4882 -11174
rect -4738 -11430 -4704 -11174
rect -4560 -11430 -4526 -11174
rect -4382 -11430 -4348 -11174
rect -4204 -11430 -4170 -11174
rect -4026 -11430 -3992 -11174
rect -2173 -11388 -2139 -11132
rect -1995 -11388 -1961 -11132
rect -1817 -11388 -1783 -11132
rect -1639 -11388 -1605 -11132
rect -1461 -11388 -1427 -11132
rect -1283 -11388 -1249 -11132
rect -1105 -11388 -1071 -11132
rect -927 -11388 -893 -11132
rect -749 -11388 -715 -11132
rect -571 -11388 -537 -11132
rect -393 -11388 -359 -11132
rect -215 -11388 -181 -11132
rect -37 -11388 -3 -11132
rect 141 -11388 175 -11132
rect 319 -11388 353 -11132
rect 497 -11388 531 -11132
rect 675 -11388 709 -11132
rect 853 -11388 887 -11132
rect 1031 -11388 1065 -11132
rect 1209 -11388 1243 -11132
rect 1387 -11388 1421 -11132
rect 1565 -11388 1599 -11132
rect 1743 -11388 1777 -11132
rect 1921 -11388 1955 -11132
rect 2099 -11388 2133 -11132
rect 2277 -11388 2311 -11132
rect 2455 -11388 2489 -11132
rect 2633 -11388 2667 -11132
rect 2811 -11388 2845 -11132
rect 2989 -11388 3023 -11132
rect 3167 -11388 3201 -11132
rect 3345 -11388 3379 -11132
rect 3523 -11388 3557 -11132
rect 3701 -11388 3735 -11132
rect 3879 -11388 3913 -11132
rect 4057 -11388 4091 -11132
rect 10772 -11490 10806 -11234
rect 10950 -11490 10984 -11234
rect 11064 -11490 11098 -11234
rect 11242 -11490 11276 -11234
rect 11356 -11490 11390 -11234
rect 11534 -11490 11568 -11234
rect 11648 -11490 11682 -11234
rect 11826 -11490 11860 -11234
rect 11940 -11490 11974 -11234
rect 12118 -11490 12152 -11234
rect 12232 -11490 12266 -11234
rect 12410 -11490 12444 -11234
rect 12524 -11490 12558 -11234
rect 12702 -11490 12736 -11234
rect -5628 -11980 -5594 -11724
rect -5450 -11980 -5416 -11724
rect -5272 -11980 -5238 -11724
rect -5094 -11980 -5060 -11724
rect -4916 -11980 -4882 -11724
rect -4738 -11980 -4704 -11724
rect -4560 -11980 -4526 -11724
rect -4382 -11980 -4348 -11724
rect -4204 -11980 -4170 -11724
rect -4026 -11980 -3992 -11724
rect 6512 -11850 6546 -11594
rect 6690 -11850 6724 -11594
rect 6868 -11850 6902 -11594
rect 7046 -11850 7080 -11594
rect 7224 -11850 7258 -11594
rect 7402 -11850 7436 -11594
rect 7580 -11850 7614 -11594
rect 7758 -11850 7792 -11594
rect 7936 -11850 7970 -11594
rect 8114 -11850 8148 -11594
rect 8292 -11850 8326 -11594
rect 8470 -11850 8504 -11594
rect 8648 -11850 8682 -11594
rect 8826 -11850 8860 -11594
rect 9004 -11850 9038 -11594
rect 9182 -11850 9216 -11594
rect 9360 -11850 9394 -11594
rect -2173 -12388 -2139 -12132
rect -1995 -12388 -1961 -12132
rect -1817 -12388 -1783 -12132
rect -1639 -12388 -1605 -12132
rect -1461 -12388 -1427 -12132
rect -1283 -12388 -1249 -12132
rect -1105 -12388 -1071 -12132
rect -927 -12388 -893 -12132
rect -749 -12388 -715 -12132
rect -571 -12388 -537 -12132
rect -393 -12388 -359 -12132
rect -215 -12388 -181 -12132
rect -37 -12388 -3 -12132
rect 141 -12388 175 -12132
rect 319 -12388 353 -12132
rect 497 -12388 531 -12132
rect 675 -12388 709 -12132
rect 853 -12388 887 -12132
rect 1031 -12388 1065 -12132
rect 1209 -12388 1243 -12132
rect 1387 -12388 1421 -12132
rect 1565 -12388 1599 -12132
rect 1743 -12388 1777 -12132
rect 1921 -12388 1955 -12132
rect 2099 -12388 2133 -12132
rect 2277 -12388 2311 -12132
rect 2455 -12388 2489 -12132
rect 2633 -12388 2667 -12132
rect 2811 -12388 2845 -12132
rect 2989 -12388 3023 -12132
rect 3167 -12388 3201 -12132
rect 3345 -12388 3379 -12132
rect 3523 -12388 3557 -12132
rect 3701 -12388 3735 -12132
rect 3879 -12388 3913 -12132
rect 4057 -12388 4091 -12132
rect -5917 -12928 -5883 -12712
rect -5817 -12928 -5783 -12712
rect -5667 -12928 -5633 -12712
rect -5567 -12928 -5533 -12712
rect -5417 -12928 -5383 -12712
rect -5317 -12928 -5283 -12712
rect -5167 -12928 -5133 -12712
rect -5067 -12928 -5033 -12712
rect -4917 -12928 -4883 -12712
rect -4817 -12928 -4783 -12712
rect -4667 -12928 -4633 -12712
rect -4567 -12928 -4533 -12712
rect -4417 -12928 -4383 -12712
rect -4317 -12928 -4283 -12712
rect -4167 -12928 -4133 -12712
rect -4067 -12928 -4033 -12712
rect -5917 -13608 -5883 -13392
rect -5817 -13608 -5783 -13392
rect -5667 -13608 -5633 -13392
rect -5567 -13608 -5533 -13392
rect -5417 -13608 -5383 -13392
rect -5317 -13608 -5283 -13392
rect -5167 -13608 -5133 -13392
rect -5067 -13608 -5033 -13392
rect -4917 -13608 -4883 -13392
rect -4817 -13608 -4783 -13392
rect -4667 -13608 -4633 -13392
rect -4567 -13608 -4533 -13392
rect -4417 -13608 -4383 -13392
rect -4317 -13608 -4283 -13392
rect -4167 -13608 -4133 -13392
rect -4067 -13608 -4033 -13392
rect -2173 -13388 -2139 -13132
rect -1995 -13388 -1961 -13132
rect -1817 -13388 -1783 -13132
rect -1639 -13388 -1605 -13132
rect -1461 -13388 -1427 -13132
rect -1283 -13388 -1249 -13132
rect -1105 -13388 -1071 -13132
rect -927 -13388 -893 -13132
rect -749 -13388 -715 -13132
rect -571 -13388 -537 -13132
rect -393 -13388 -359 -13132
rect -215 -13388 -181 -13132
rect -37 -13388 -3 -13132
rect 141 -13388 175 -13132
rect 319 -13388 353 -13132
rect 497 -13388 531 -13132
rect 675 -13388 709 -13132
rect 853 -13388 887 -13132
rect 1031 -13388 1065 -13132
rect 1209 -13388 1243 -13132
rect 1387 -13388 1421 -13132
rect 1565 -13388 1599 -13132
rect 1743 -13388 1777 -13132
rect 1921 -13388 1955 -13132
rect 2099 -13388 2133 -13132
rect 2277 -13388 2311 -13132
rect 2455 -13388 2489 -13132
rect 2633 -13388 2667 -13132
rect 2811 -13388 2845 -13132
rect 2989 -13388 3023 -13132
rect 3167 -13388 3201 -13132
rect 3345 -13388 3379 -13132
rect 3523 -13388 3557 -13132
rect 3701 -13388 3735 -13132
rect 3879 -13388 3913 -13132
rect 4057 -13388 4091 -13132
rect -6028 -14650 -5994 -14394
rect -5850 -14650 -5816 -14394
rect -5672 -14650 -5638 -14394
rect -5494 -14650 -5460 -14394
rect -5316 -14650 -5282 -14394
rect -5138 -14650 -5104 -14394
rect -4960 -14650 -4926 -14394
rect -4782 -14650 -4748 -14394
rect -4604 -14650 -4570 -14394
rect -4426 -14650 -4392 -14394
rect -4248 -14650 -4214 -14394
rect -4070 -14650 -4036 -14394
rect -2173 -14388 -2139 -14132
rect -1995 -14388 -1961 -14132
rect -1817 -14388 -1783 -14132
rect -1639 -14388 -1605 -14132
rect -1461 -14388 -1427 -14132
rect -1283 -14388 -1249 -14132
rect -1105 -14388 -1071 -14132
rect -927 -14388 -893 -14132
rect -749 -14388 -715 -14132
rect -571 -14388 -537 -14132
rect -393 -14388 -359 -14132
rect -215 -14388 -181 -14132
rect -37 -14388 -3 -14132
rect 141 -14388 175 -14132
rect 319 -14388 353 -14132
rect 497 -14388 531 -14132
rect 675 -14388 709 -14132
rect 853 -14388 887 -14132
rect 1031 -14388 1065 -14132
rect 1209 -14388 1243 -14132
rect 1387 -14388 1421 -14132
rect 1565 -14388 1599 -14132
rect 1743 -14388 1777 -14132
rect 1921 -14388 1955 -14132
rect 2099 -14388 2133 -14132
rect 2277 -14388 2311 -14132
rect 2455 -14388 2489 -14132
rect 2633 -14388 2667 -14132
rect 2811 -14388 2845 -14132
rect 2989 -14388 3023 -14132
rect 3167 -14388 3201 -14132
rect 3345 -14388 3379 -14132
rect 3523 -14388 3557 -14132
rect 3701 -14388 3735 -14132
rect 3879 -14388 3913 -14132
rect 4057 -14388 4091 -14132
rect 5577 -14388 5611 -14132
rect 5755 -14388 5789 -14132
rect 5933 -14388 5967 -14132
rect 6111 -14388 6145 -14132
rect 6289 -14388 6323 -14132
rect 6467 -14388 6501 -14132
rect 6645 -14388 6679 -14132
rect 6823 -14388 6857 -14132
rect 7001 -14388 7035 -14132
rect 7179 -14388 7213 -14132
rect 7357 -14388 7391 -14132
rect 7535 -14388 7569 -14132
rect 7713 -14388 7747 -14132
rect 7891 -14388 7925 -14132
rect 8069 -14388 8103 -14132
rect 8247 -14388 8281 -14132
rect 8425 -14388 8459 -14132
rect 8603 -14388 8637 -14132
rect 8781 -14388 8815 -14132
rect 8959 -14388 8993 -14132
rect 9137 -14388 9171 -14132
rect 9315 -14388 9349 -14132
rect 9493 -14388 9527 -14132
rect 9671 -14388 9705 -14132
rect 9849 -14388 9883 -14132
rect 10027 -14388 10061 -14132
rect 10205 -14388 10239 -14132
rect 10383 -14388 10417 -14132
rect 10561 -14388 10595 -14132
rect 10739 -14388 10773 -14132
rect 10917 -14388 10951 -14132
rect 11095 -14388 11129 -14132
rect 11273 -14388 11307 -14132
rect 11451 -14388 11485 -14132
rect 11629 -14388 11663 -14132
rect 11807 -14388 11841 -14132
rect 11985 -14388 12019 -14132
rect 12163 -14388 12197 -14132
rect 12341 -14388 12375 -14132
rect 12519 -14388 12553 -14132
rect 12697 -14388 12731 -14132
rect -6028 -15350 -5994 -15094
rect -5850 -15350 -5816 -15094
rect -5672 -15350 -5638 -15094
rect -5494 -15350 -5460 -15094
rect -5316 -15350 -5282 -15094
rect -5138 -15350 -5104 -15094
rect -4960 -15350 -4926 -15094
rect -4782 -15350 -4748 -15094
rect -4604 -15350 -4570 -15094
rect -4426 -15350 -4392 -15094
rect -4248 -15350 -4214 -15094
rect -4070 -15350 -4036 -15094
rect -2173 -15388 -2139 -15132
rect -1995 -15388 -1961 -15132
rect -1817 -15388 -1783 -15132
rect -1639 -15388 -1605 -15132
rect -1461 -15388 -1427 -15132
rect -1283 -15388 -1249 -15132
rect -1105 -15388 -1071 -15132
rect -927 -15388 -893 -15132
rect -749 -15388 -715 -15132
rect -571 -15388 -537 -15132
rect -393 -15388 -359 -15132
rect -215 -15388 -181 -15132
rect -37 -15388 -3 -15132
rect 141 -15388 175 -15132
rect 319 -15388 353 -15132
rect 497 -15388 531 -15132
rect 675 -15388 709 -15132
rect 853 -15388 887 -15132
rect 1031 -15388 1065 -15132
rect 1209 -15388 1243 -15132
rect 1387 -15388 1421 -15132
rect 1565 -15388 1599 -15132
rect 1743 -15388 1777 -15132
rect 1921 -15388 1955 -15132
rect 2099 -15388 2133 -15132
rect 2277 -15388 2311 -15132
rect 2455 -15388 2489 -15132
rect 2633 -15388 2667 -15132
rect 2811 -15388 2845 -15132
rect 2989 -15388 3023 -15132
rect 3167 -15388 3201 -15132
rect 3345 -15388 3379 -15132
rect 3523 -15388 3557 -15132
rect 3701 -15388 3735 -15132
rect 3879 -15388 3913 -15132
rect 4057 -15388 4091 -15132
rect 5577 -15388 5611 -15132
rect 5755 -15388 5789 -15132
rect 5933 -15388 5967 -15132
rect 6111 -15388 6145 -15132
rect 6289 -15388 6323 -15132
rect 6467 -15388 6501 -15132
rect 6645 -15388 6679 -15132
rect 6823 -15388 6857 -15132
rect 7001 -15388 7035 -15132
rect 7179 -15388 7213 -15132
rect 7357 -15388 7391 -15132
rect 7535 -15388 7569 -15132
rect 7713 -15388 7747 -15132
rect 7891 -15388 7925 -15132
rect 8069 -15388 8103 -15132
rect 8247 -15388 8281 -15132
rect 8425 -15388 8459 -15132
rect 8603 -15388 8637 -15132
rect 8781 -15388 8815 -15132
rect 8959 -15388 8993 -15132
rect 9137 -15388 9171 -15132
rect 9315 -15388 9349 -15132
rect 9493 -15388 9527 -15132
rect 9671 -15388 9705 -15132
rect 9849 -15388 9883 -15132
rect 10027 -15388 10061 -15132
rect 10205 -15388 10239 -15132
rect 10383 -15388 10417 -15132
rect 10561 -15388 10595 -15132
rect 10739 -15388 10773 -15132
rect 10917 -15388 10951 -15132
rect 11095 -15388 11129 -15132
rect 11273 -15388 11307 -15132
rect 11451 -15388 11485 -15132
rect 11629 -15388 11663 -15132
rect 11807 -15388 11841 -15132
rect 11985 -15388 12019 -15132
rect 12163 -15388 12197 -15132
rect 12341 -15388 12375 -15132
rect 12519 -15388 12553 -15132
rect 12697 -15388 12731 -15132
rect -6028 -16050 -5994 -15794
rect -5850 -16050 -5816 -15794
rect -5672 -16050 -5638 -15794
rect -5494 -16050 -5460 -15794
rect -5316 -16050 -5282 -15794
rect -5138 -16050 -5104 -15794
rect -4960 -16050 -4926 -15794
rect -4782 -16050 -4748 -15794
rect -4604 -16050 -4570 -15794
rect -4426 -16050 -4392 -15794
rect -4248 -16050 -4214 -15794
rect -4070 -16050 -4036 -15794
rect -2173 -16388 -2139 -16132
rect -1995 -16388 -1961 -16132
rect -1817 -16388 -1783 -16132
rect -1639 -16388 -1605 -16132
rect -1461 -16388 -1427 -16132
rect -1283 -16388 -1249 -16132
rect -1105 -16388 -1071 -16132
rect -927 -16388 -893 -16132
rect -749 -16388 -715 -16132
rect -571 -16388 -537 -16132
rect -393 -16388 -359 -16132
rect -215 -16388 -181 -16132
rect -37 -16388 -3 -16132
rect 141 -16388 175 -16132
rect 319 -16388 353 -16132
rect 497 -16388 531 -16132
rect 675 -16388 709 -16132
rect 853 -16388 887 -16132
rect 1031 -16388 1065 -16132
rect 1209 -16388 1243 -16132
rect 1387 -16388 1421 -16132
rect 1565 -16388 1599 -16132
rect 1743 -16388 1777 -16132
rect 1921 -16388 1955 -16132
rect 2099 -16388 2133 -16132
rect 2277 -16388 2311 -16132
rect 2455 -16388 2489 -16132
rect 2633 -16388 2667 -16132
rect 2811 -16388 2845 -16132
rect 2989 -16388 3023 -16132
rect 3167 -16388 3201 -16132
rect 3345 -16388 3379 -16132
rect 3523 -16388 3557 -16132
rect 3701 -16388 3735 -16132
rect 3879 -16388 3913 -16132
rect 4057 -16388 4091 -16132
rect 5577 -16388 5611 -16132
rect 5755 -16388 5789 -16132
rect 5933 -16388 5967 -16132
rect 6111 -16388 6145 -16132
rect 6289 -16388 6323 -16132
rect 6467 -16388 6501 -16132
rect 6645 -16388 6679 -16132
rect 6823 -16388 6857 -16132
rect 7001 -16388 7035 -16132
rect 7179 -16388 7213 -16132
rect 7357 -16388 7391 -16132
rect 7535 -16388 7569 -16132
rect 7713 -16388 7747 -16132
rect 7891 -16388 7925 -16132
rect 8069 -16388 8103 -16132
rect 8247 -16388 8281 -16132
rect 8425 -16388 8459 -16132
rect 8603 -16388 8637 -16132
rect 8781 -16388 8815 -16132
rect 8959 -16388 8993 -16132
rect 9137 -16388 9171 -16132
rect 9315 -16388 9349 -16132
rect 9493 -16388 9527 -16132
rect 9671 -16388 9705 -16132
rect 9849 -16388 9883 -16132
rect 10027 -16388 10061 -16132
rect 10205 -16388 10239 -16132
rect 10383 -16388 10417 -16132
rect 10561 -16388 10595 -16132
rect 10739 -16388 10773 -16132
rect 10917 -16388 10951 -16132
rect 11095 -16388 11129 -16132
rect 11273 -16388 11307 -16132
rect 11451 -16388 11485 -16132
rect 11629 -16388 11663 -16132
rect 11807 -16388 11841 -16132
rect 11985 -16388 12019 -16132
rect 12163 -16388 12197 -16132
rect 12341 -16388 12375 -16132
rect 12519 -16388 12553 -16132
rect 12697 -16388 12731 -16132
rect -6028 -16750 -5994 -16494
rect -5850 -16750 -5816 -16494
rect -5672 -16750 -5638 -16494
rect -5494 -16750 -5460 -16494
rect -5316 -16750 -5282 -16494
rect -5138 -16750 -5104 -16494
rect -4960 -16750 -4926 -16494
rect -4782 -16750 -4748 -16494
rect -4604 -16750 -4570 -16494
rect -4426 -16750 -4392 -16494
rect -4248 -16750 -4214 -16494
rect -4070 -16750 -4036 -16494
<< pdiffc >>
rect 7154 2365 7188 2613
rect 7250 2365 7284 2613
rect 7346 2365 7380 2613
rect 7442 2365 7476 2613
rect 7538 2365 7572 2613
rect 7634 2365 7668 2613
rect 7730 2365 7764 2613
rect 7826 2365 7860 2613
rect 7922 2365 7956 2613
rect 8018 2365 8052 2613
rect 8114 2365 8148 2613
rect 16154 2365 16188 2613
rect 16250 2365 16284 2613
rect 16346 2365 16380 2613
rect 16442 2365 16476 2613
rect 16538 2365 16572 2613
rect 16634 2365 16668 2613
rect 16730 2365 16764 2613
rect 16826 2365 16860 2613
rect 16922 2365 16956 2613
rect 17018 2365 17052 2613
rect 17114 2365 17148 2613
rect 7154 565 7188 813
rect 7250 565 7284 813
rect 7346 565 7380 813
rect 7442 565 7476 813
rect 7538 565 7572 813
rect 7634 565 7668 813
rect 7730 565 7764 813
rect 7826 565 7860 813
rect 7922 565 7956 813
rect 8018 565 8052 813
rect 8114 565 8148 813
rect 16154 565 16188 813
rect 16250 565 16284 813
rect 16346 565 16380 813
rect 16442 565 16476 813
rect 16538 565 16572 813
rect 16634 565 16668 813
rect 16730 565 16764 813
rect 16826 565 16860 813
rect 16922 565 16956 813
rect 17018 565 17052 813
rect 17114 565 17148 813
rect 7154 -1235 7188 -987
rect 7250 -1235 7284 -987
rect 7346 -1235 7380 -987
rect 7442 -1235 7476 -987
rect 7538 -1235 7572 -987
rect 7634 -1235 7668 -987
rect 7730 -1235 7764 -987
rect 7826 -1235 7860 -987
rect 7922 -1235 7956 -987
rect 8018 -1235 8052 -987
rect 8114 -1235 8148 -987
rect 16154 -1235 16188 -987
rect 16250 -1235 16284 -987
rect 16346 -1235 16380 -987
rect 16442 -1235 16476 -987
rect 16538 -1235 16572 -987
rect 16634 -1235 16668 -987
rect 16730 -1235 16764 -987
rect 16826 -1235 16860 -987
rect 16922 -1235 16956 -987
rect 17018 -1235 17052 -987
rect 17114 -1235 17148 -987
rect -6302 -2388 -6268 -2132
rect -6124 -2388 -6090 -2132
rect -5946 -2388 -5912 -2132
rect -5768 -2388 -5734 -2132
rect -5590 -2388 -5556 -2132
rect -5412 -2388 -5378 -2132
rect -5234 -2388 -5200 -2132
rect -5056 -2388 -5022 -2132
rect -4878 -2388 -4844 -2132
rect -4700 -2388 -4666 -2132
rect -4522 -2388 -4488 -2132
rect -4344 -2388 -4310 -2132
rect -4166 -2388 -4132 -2132
rect -3988 -2388 -3954 -2132
rect -3810 -2388 -3776 -2132
rect -3632 -2388 -3598 -2132
rect -3454 -2388 -3420 -2132
rect -6302 -3258 -6268 -3002
rect -6124 -3258 -6090 -3002
rect -5946 -3258 -5912 -3002
rect -5768 -3258 -5734 -3002
rect -5590 -3258 -5556 -3002
rect -5412 -3258 -5378 -3002
rect -5234 -3258 -5200 -3002
rect -5056 -3258 -5022 -3002
rect -4878 -3258 -4844 -3002
rect -4700 -3258 -4666 -3002
rect -4522 -3258 -4488 -3002
rect -4344 -3258 -4310 -3002
rect -4166 -3258 -4132 -3002
rect -3988 -3258 -3954 -3002
rect -3810 -3258 -3776 -3002
rect -3632 -3258 -3598 -3002
rect -3454 -3258 -3420 -3002
rect -1454 -3140 -1420 -2884
rect -1276 -3140 -1242 -2884
rect -1098 -3140 -1064 -2884
rect -920 -3140 -886 -2884
rect -742 -3140 -708 -2884
rect -564 -3140 -530 -2884
rect -386 -3140 -352 -2884
rect -208 -3140 -174 -2884
rect -30 -3140 4 -2884
rect 148 -3140 182 -2884
rect 326 -3140 360 -2884
rect 504 -3140 538 -2884
rect 682 -3140 716 -2884
rect 860 -3140 894 -2884
rect 1038 -3140 1072 -2884
rect 1216 -3140 1250 -2884
rect 1394 -3140 1428 -2884
rect 1572 -3140 1606 -2884
rect 1750 -3140 1784 -2884
rect 1928 -3140 1962 -2884
rect 2106 -3140 2140 -2884
rect 2284 -3140 2318 -2884
rect 2462 -3140 2496 -2884
rect 2640 -3140 2674 -2884
rect -6302 -4128 -6268 -3872
rect -6124 -4128 -6090 -3872
rect -5946 -4128 -5912 -3872
rect -5768 -4128 -5734 -3872
rect -5590 -4128 -5556 -3872
rect -5412 -4128 -5378 -3872
rect -5234 -4128 -5200 -3872
rect -5056 -4128 -5022 -3872
rect -4878 -4128 -4844 -3872
rect -4700 -4128 -4666 -3872
rect -4522 -4128 -4488 -3872
rect -4344 -4128 -4310 -3872
rect -4166 -4128 -4132 -3872
rect -3988 -4128 -3954 -3872
rect -3810 -4128 -3776 -3872
rect -3632 -4128 -3598 -3872
rect -3454 -4128 -3420 -3872
rect -1454 -4040 -1420 -3784
rect -1276 -4040 -1242 -3784
rect -1098 -4040 -1064 -3784
rect -920 -4040 -886 -3784
rect -742 -4040 -708 -3784
rect -564 -4040 -530 -3784
rect -386 -4040 -352 -3784
rect -208 -4040 -174 -3784
rect -30 -4040 4 -3784
rect 148 -4040 182 -3784
rect 326 -4040 360 -3784
rect 504 -4040 538 -3784
rect 682 -4040 716 -3784
rect 860 -4040 894 -3784
rect 1038 -4040 1072 -3784
rect 1216 -4040 1250 -3784
rect 1394 -4040 1428 -3784
rect 1572 -4040 1606 -3784
rect 1750 -4040 1784 -3784
rect 1928 -4040 1962 -3784
rect 2106 -4040 2140 -3784
rect 2284 -4040 2318 -3784
rect 2462 -4040 2496 -3784
rect 2640 -4040 2674 -3784
rect -6302 -4998 -6268 -4742
rect -6124 -4998 -6090 -4742
rect -5946 -4998 -5912 -4742
rect -5768 -4998 -5734 -4742
rect -5590 -4998 -5556 -4742
rect -5412 -4998 -5378 -4742
rect -5234 -4998 -5200 -4742
rect -5056 -4998 -5022 -4742
rect -4878 -4998 -4844 -4742
rect -4700 -4998 -4666 -4742
rect -4522 -4998 -4488 -4742
rect -4344 -4998 -4310 -4742
rect -4166 -4998 -4132 -4742
rect -3988 -4998 -3954 -4742
rect -3810 -4998 -3776 -4742
rect -3632 -4998 -3598 -4742
rect -3454 -4998 -3420 -4742
rect -1454 -4940 -1420 -4684
rect -1276 -4940 -1242 -4684
rect -1098 -4940 -1064 -4684
rect -920 -4940 -886 -4684
rect -742 -4940 -708 -4684
rect -564 -4940 -530 -4684
rect -386 -4940 -352 -4684
rect -208 -4940 -174 -4684
rect -30 -4940 4 -4684
rect 148 -4940 182 -4684
rect 326 -4940 360 -4684
rect 504 -4940 538 -4684
rect 682 -4940 716 -4684
rect 860 -4940 894 -4684
rect 1038 -4940 1072 -4684
rect 1216 -4940 1250 -4684
rect 1394 -4940 1428 -4684
rect 1572 -4940 1606 -4684
rect 1750 -4940 1784 -4684
rect 1928 -4940 1962 -4684
rect 2106 -4940 2140 -4684
rect 2284 -4940 2318 -4684
rect 2462 -4940 2496 -4684
rect 2640 -4940 2674 -4684
rect -6302 -5868 -6268 -5612
rect -6124 -5868 -6090 -5612
rect -5946 -5868 -5912 -5612
rect -5768 -5868 -5734 -5612
rect -5590 -5868 -5556 -5612
rect -5412 -5868 -5378 -5612
rect -5234 -5868 -5200 -5612
rect -5056 -5868 -5022 -5612
rect -4878 -5868 -4844 -5612
rect -4700 -5868 -4666 -5612
rect -4522 -5868 -4488 -5612
rect -4344 -5868 -4310 -5612
rect -4166 -5868 -4132 -5612
rect -3988 -5868 -3954 -5612
rect -3810 -5868 -3776 -5612
rect -3632 -5868 -3598 -5612
rect -3454 -5868 -3420 -5612
rect -1454 -5840 -1420 -5584
rect -1276 -5840 -1242 -5584
rect -1098 -5840 -1064 -5584
rect -920 -5840 -886 -5584
rect -742 -5840 -708 -5584
rect -564 -5840 -530 -5584
rect -386 -5840 -352 -5584
rect -208 -5840 -174 -5584
rect -30 -5840 4 -5584
rect 148 -5840 182 -5584
rect 326 -5840 360 -5584
rect 504 -5840 538 -5584
rect 682 -5840 716 -5584
rect 860 -5840 894 -5584
rect 1038 -5840 1072 -5584
rect 1216 -5840 1250 -5584
rect 1394 -5840 1428 -5584
rect 1572 -5840 1606 -5584
rect 1750 -5840 1784 -5584
rect 1928 -5840 1962 -5584
rect 2106 -5840 2140 -5584
rect 2284 -5840 2318 -5584
rect 2462 -5840 2496 -5584
rect 2640 -5840 2674 -5584
rect 7154 -3035 7188 -2787
rect 7250 -3035 7284 -2787
rect 7346 -3035 7380 -2787
rect 7442 -3035 7476 -2787
rect 7538 -3035 7572 -2787
rect 7634 -3035 7668 -2787
rect 7730 -3035 7764 -2787
rect 7826 -3035 7860 -2787
rect 7922 -3035 7956 -2787
rect 8018 -3035 8052 -2787
rect 8114 -3035 8148 -2787
rect 16154 -3035 16188 -2787
rect 16250 -3035 16284 -2787
rect 16346 -3035 16380 -2787
rect 16442 -3035 16476 -2787
rect 16538 -3035 16572 -2787
rect 16634 -3035 16668 -2787
rect 16730 -3035 16764 -2787
rect 16826 -3035 16860 -2787
rect 16922 -3035 16956 -2787
rect 17018 -3035 17052 -2787
rect 17114 -3035 17148 -2787
rect 7154 -4835 7188 -4587
rect 7250 -4835 7284 -4587
rect 7346 -4835 7380 -4587
rect 7442 -4835 7476 -4587
rect 7538 -4835 7572 -4587
rect 7634 -4835 7668 -4587
rect 7730 -4835 7764 -4587
rect 7826 -4835 7860 -4587
rect 7922 -4835 7956 -4587
rect 8018 -4835 8052 -4587
rect 8114 -4835 8148 -4587
rect 16154 -4835 16188 -4587
rect 16250 -4835 16284 -4587
rect 16346 -4835 16380 -4587
rect 16442 -4835 16476 -4587
rect 16538 -4835 16572 -4587
rect 16634 -4835 16668 -4587
rect 16730 -4835 16764 -4587
rect 16826 -4835 16860 -4587
rect 16922 -4835 16956 -4587
rect 17018 -4835 17052 -4587
rect 17114 -4835 17148 -4587
rect 7154 -6635 7188 -6387
rect 7250 -6635 7284 -6387
rect 7346 -6635 7380 -6387
rect 7442 -6635 7476 -6387
rect 7538 -6635 7572 -6387
rect 7634 -6635 7668 -6387
rect 7730 -6635 7764 -6387
rect 7826 -6635 7860 -6387
rect 7922 -6635 7956 -6387
rect 8018 -6635 8052 -6387
rect 8114 -6635 8148 -6387
rect 16154 -6635 16188 -6387
rect 16250 -6635 16284 -6387
rect 16346 -6635 16380 -6387
rect 16442 -6635 16476 -6387
rect 16538 -6635 16572 -6387
rect 16634 -6635 16668 -6387
rect 16730 -6635 16764 -6387
rect 16826 -6635 16860 -6387
rect 16922 -6635 16956 -6387
rect 17018 -6635 17052 -6387
rect 17114 -6635 17148 -6387
<< psubdiff >>
rect 7040 2123 7136 2157
rect 8166 2123 8262 2157
rect 7040 2061 7074 2123
rect 8228 2061 8262 2123
rect 7040 1801 7074 1863
rect 8228 1801 8262 1863
rect 7040 1767 7136 1801
rect 8166 1767 8262 1801
rect 16040 2123 16136 2157
rect 17166 2123 17262 2157
rect 16040 2061 16074 2123
rect 17228 2061 17262 2123
rect 16040 1801 16074 1863
rect 17228 1801 17262 1863
rect 16040 1767 16136 1801
rect 17166 1767 17262 1801
rect 7040 323 7136 357
rect 8166 323 8262 357
rect 7040 261 7074 323
rect 8228 261 8262 323
rect 7040 1 7074 63
rect 8228 1 8262 63
rect 7040 -33 7136 1
rect 8166 -33 8262 1
rect 16040 323 16136 357
rect 17166 323 17262 357
rect 16040 261 16074 323
rect 17228 261 17262 323
rect 16040 1 16074 63
rect 17228 1 17262 63
rect 16040 -33 16136 1
rect 17166 -33 17262 1
rect 7040 -1477 7136 -1443
rect 8166 -1477 8262 -1443
rect 7040 -1539 7074 -1477
rect 8228 -1539 8262 -1477
rect 7040 -1799 7074 -1737
rect 8228 -1799 8262 -1737
rect 7040 -1833 7136 -1799
rect 8166 -1833 8262 -1799
rect 16040 -1477 16136 -1443
rect 17166 -1477 17262 -1443
rect 16040 -1539 16074 -1477
rect 17228 -1539 17262 -1477
rect 16040 -1799 16074 -1737
rect 17228 -1799 17262 -1737
rect 16040 -1833 16136 -1799
rect 17166 -1833 17262 -1799
rect 7040 -3277 7136 -3243
rect 8166 -3277 8262 -3243
rect 7040 -3339 7074 -3277
rect 8228 -3339 8262 -3277
rect 7040 -3599 7074 -3537
rect 8228 -3599 8262 -3537
rect 7040 -3633 7136 -3599
rect 8166 -3633 8262 -3599
rect 16040 -3277 16136 -3243
rect 17166 -3277 17262 -3243
rect 16040 -3339 16074 -3277
rect 17228 -3339 17262 -3277
rect 16040 -3599 16074 -3537
rect 17228 -3599 17262 -3537
rect 16040 -3633 16136 -3599
rect 17166 -3633 17262 -3599
rect 7040 -5077 7136 -5043
rect 8166 -5077 8262 -5043
rect 7040 -5139 7074 -5077
rect 8228 -5139 8262 -5077
rect 7040 -5399 7074 -5337
rect 8228 -5399 8262 -5337
rect 7040 -5433 7136 -5399
rect 8166 -5433 8262 -5399
rect 16040 -5077 16136 -5043
rect 17166 -5077 17262 -5043
rect 16040 -5139 16074 -5077
rect 17228 -5139 17262 -5077
rect 16040 -5399 16074 -5337
rect 17228 -5399 17262 -5337
rect 16040 -5433 16136 -5399
rect 17166 -5433 17262 -5399
rect 7040 -6877 7136 -6843
rect 8166 -6877 8262 -6843
rect 7040 -6939 7074 -6877
rect 8228 -6939 8262 -6877
rect 7040 -7199 7074 -7137
rect 8228 -7199 8262 -7137
rect 7040 -7233 7136 -7199
rect 8166 -7233 8262 -7199
rect 16040 -6877 16136 -6843
rect 17166 -6877 17262 -6843
rect 16040 -6939 16074 -6877
rect 17228 -6939 17262 -6877
rect 16040 -7199 16074 -7137
rect 17228 -7199 17262 -7137
rect 16040 -7233 16136 -7199
rect 17166 -7233 17262 -7199
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect 13619 -7731 13719 -7621
rect -3009 -9276 -2783 -9252
rect -3009 -9454 -2985 -9276
rect -2807 -9454 -2783 -9276
rect 9958 -9191 10184 -9167
rect 9958 -9369 9982 -9191
rect 10160 -9369 10184 -9191
rect 9958 -9393 10184 -9369
rect -3009 -9478 -2783 -9454
rect -3009 -11276 -2783 -11252
rect -3009 -11454 -2985 -11276
rect -2807 -11454 -2783 -11276
rect 5662 -11151 5888 -11127
rect 5662 -11329 5686 -11151
rect 5864 -11329 5888 -11151
rect 5662 -11353 5888 -11329
rect 9958 -11191 10184 -11167
rect 9958 -11369 9982 -11191
rect 10160 -11369 10184 -11191
rect 9958 -11393 10184 -11369
rect -3009 -11478 -2783 -11454
rect 8413 -12554 8639 -12530
rect 8413 -12732 8437 -12554
rect 8615 -12732 8639 -12554
rect 8413 -12756 8639 -12732
rect 11413 -12554 11639 -12530
rect 11413 -12732 11437 -12554
rect 11615 -12732 11639 -12554
rect 11413 -12756 11639 -12732
rect -3009 -13276 -2783 -13252
rect -3009 -13454 -2985 -13276
rect -2807 -13454 -2783 -13276
rect -3009 -13478 -2783 -13454
rect 4519 -14869 4745 -14845
rect 4519 -15047 4543 -14869
rect 4721 -15047 4745 -14869
rect 4519 -15071 4745 -15047
rect -3009 -15276 -2783 -15252
rect -3009 -15454 -2985 -15276
rect -2807 -15454 -2783 -15276
rect -3009 -15478 -2783 -15454
rect -7605 -17459 -7505 -17268
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< nsubdiff >>
rect 7040 2775 7136 2809
rect 8166 2775 8262 2809
rect 7040 2713 7074 2775
rect 8228 2713 8262 2775
rect 7040 2265 7074 2327
rect 8228 2265 8262 2327
rect 7040 2231 7136 2265
rect 8166 2231 8262 2265
rect 16040 2775 16136 2809
rect 17166 2775 17262 2809
rect 16040 2713 16074 2775
rect 17228 2713 17262 2775
rect 16040 2265 16074 2327
rect 17228 2265 17262 2327
rect 16040 2231 16136 2265
rect 17166 2231 17262 2265
rect 7040 975 7136 1009
rect 8166 975 8262 1009
rect 7040 913 7074 975
rect 8228 913 8262 975
rect 7040 465 7074 527
rect 8228 465 8262 527
rect 7040 431 7136 465
rect 8166 431 8262 465
rect 16040 975 16136 1009
rect 17166 975 17262 1009
rect 16040 913 16074 975
rect 17228 913 17262 975
rect 16040 465 16074 527
rect 17228 465 17262 527
rect 16040 431 16136 465
rect 17166 431 17262 465
rect 7040 -825 7136 -791
rect 8166 -825 8262 -791
rect 7040 -887 7074 -825
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect 3610 -1520 3703 -1353
rect 8228 -887 8262 -825
rect 7040 -1335 7074 -1273
rect 8228 -1335 8262 -1273
rect 7040 -1369 7136 -1335
rect 8166 -1369 8262 -1335
rect 16040 -825 16136 -791
rect 17166 -825 17262 -791
rect 16040 -887 16074 -825
rect 17228 -887 17262 -825
rect 16040 -1335 16074 -1273
rect 17228 -1335 17262 -1273
rect 16040 -1369 16136 -1335
rect 17166 -1369 17262 -1335
rect -2210 -3043 -1984 -3019
rect -2210 -3221 -2186 -3043
rect -2008 -3221 -1984 -3043
rect -2210 -3245 -1984 -3221
rect -3058 -5662 -2832 -5638
rect -3058 -5840 -3034 -5662
rect -2856 -5840 -2832 -5662
rect -3058 -5864 -2832 -5840
rect -7605 -7140 -7512 -6976
rect 7040 -2625 7136 -2591
rect 8166 -2625 8262 -2591
rect 7040 -2687 7074 -2625
rect 8228 -2687 8262 -2625
rect 7040 -3135 7074 -3073
rect 8228 -3135 8262 -3073
rect 7040 -3169 7136 -3135
rect 8166 -3169 8262 -3135
rect 16040 -2625 16136 -2591
rect 17166 -2625 17262 -2591
rect 16040 -2687 16074 -2625
rect 17228 -2687 17262 -2625
rect 16040 -3135 16074 -3073
rect 17228 -3135 17262 -3073
rect 16040 -3169 16136 -3135
rect 17166 -3169 17262 -3135
rect 7040 -4425 7136 -4391
rect 8166 -4425 8262 -4391
rect 7040 -4487 7074 -4425
rect 8228 -4487 8262 -4425
rect 7040 -4935 7074 -4873
rect 8228 -4935 8262 -4873
rect 7040 -4969 7136 -4935
rect 8166 -4969 8262 -4935
rect 16040 -4425 16136 -4391
rect 17166 -4425 17262 -4391
rect 16040 -4487 16074 -4425
rect 17228 -4487 17262 -4425
rect 16040 -4935 16074 -4873
rect 17228 -4935 17262 -4873
rect 16040 -4969 16136 -4935
rect 17166 -4969 17262 -4935
rect 7040 -6225 7136 -6191
rect 8166 -6225 8262 -6191
rect 7040 -6287 7074 -6225
rect 8228 -6287 8262 -6225
rect 7040 -6735 7074 -6673
rect 8228 -6735 8262 -6673
rect 7040 -6769 7136 -6735
rect 8166 -6769 8262 -6735
rect 16040 -6225 16136 -6191
rect 17166 -6225 17262 -6191
rect 16040 -6287 16074 -6225
rect 17228 -6287 17262 -6225
rect 16040 -6735 16074 -6673
rect 17228 -6735 17262 -6673
rect 16040 -6769 16136 -6735
rect 17166 -6769 17262 -6735
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
<< psubdiffcont >>
rect 7136 2123 8166 2157
rect 7040 1863 7074 2061
rect 8228 1863 8262 2061
rect 7136 1767 8166 1801
rect 16136 2123 17166 2157
rect 16040 1863 16074 2061
rect 17228 1863 17262 2061
rect 16136 1767 17166 1801
rect 7136 323 8166 357
rect 7040 63 7074 261
rect 8228 63 8262 261
rect 7136 -33 8166 1
rect 16136 323 17166 357
rect 16040 63 16074 261
rect 17228 63 17262 261
rect 16136 -33 17166 1
rect 7136 -1477 8166 -1443
rect 7040 -1737 7074 -1539
rect 8228 -1737 8262 -1539
rect 7136 -1833 8166 -1799
rect 16136 -1477 17166 -1443
rect 16040 -1737 16074 -1539
rect 17228 -1737 17262 -1539
rect 16136 -1833 17166 -1799
rect 7136 -3277 8166 -3243
rect 7040 -3537 7074 -3339
rect 8228 -3537 8262 -3339
rect 7136 -3633 8166 -3599
rect 16136 -3277 17166 -3243
rect 16040 -3537 16074 -3339
rect 17228 -3537 17262 -3339
rect 16136 -3633 17166 -3599
rect 7136 -5077 8166 -5043
rect 7040 -5337 7074 -5139
rect 8228 -5337 8262 -5139
rect 7136 -5433 8166 -5399
rect 16136 -5077 17166 -5043
rect 16040 -5337 16074 -5139
rect 17228 -5337 17262 -5139
rect 16136 -5433 17166 -5399
rect 7136 -6877 8166 -6843
rect 7040 -7137 7074 -6939
rect 8228 -7137 8262 -6939
rect 7136 -7233 8166 -7199
rect 16136 -6877 17166 -6843
rect 16040 -7137 16074 -6939
rect 17228 -7137 17262 -6939
rect 16136 -7233 17166 -7199
rect -7264 -7621 13443 -7521
rect -7605 -17268 -7505 -7850
rect -2985 -9454 -2807 -9276
rect 9982 -9369 10160 -9191
rect -2985 -11454 -2807 -11276
rect 5686 -11329 5864 -11151
rect 9982 -11369 10160 -11191
rect 8437 -12732 8615 -12554
rect 11437 -12732 11615 -12554
rect -2985 -13454 -2807 -13276
rect 4543 -15047 4721 -14869
rect -2985 -15454 -2807 -15276
rect 13619 -17149 13719 -7731
rect -7323 -17559 13384 -17459
<< nsubdiffcont >>
rect 7136 2775 8166 2809
rect 7040 2327 7074 2713
rect 8228 2327 8262 2713
rect 7136 2231 8166 2265
rect 16136 2775 17166 2809
rect 16040 2327 16074 2713
rect 17228 2327 17262 2713
rect 16136 2231 17166 2265
rect 7136 975 8166 1009
rect 7040 527 7074 913
rect 8228 527 8262 913
rect 7136 431 8166 465
rect 16136 975 17166 1009
rect 16040 527 16074 913
rect 17228 527 17262 913
rect 16136 431 17166 465
rect 7136 -825 8166 -791
rect -7379 -1353 3329 -1260
rect -7605 -6976 -7512 -1507
rect 7040 -1273 7074 -887
rect 8228 -1273 8262 -887
rect 7136 -1369 8166 -1335
rect 16136 -825 17166 -791
rect 16040 -1273 16074 -887
rect 17228 -1273 17262 -887
rect 16136 -1369 17166 -1335
rect -2186 -3221 -2008 -3043
rect -3034 -5840 -2856 -5662
rect 3610 -6989 3703 -1520
rect 7136 -2625 8166 -2591
rect 7040 -3073 7074 -2687
rect 8228 -3073 8262 -2687
rect 7136 -3169 8166 -3135
rect 16136 -2625 17166 -2591
rect 16040 -3073 16074 -2687
rect 17228 -3073 17262 -2687
rect 16136 -3169 17166 -3135
rect 7136 -4425 8166 -4391
rect 7040 -4873 7074 -4487
rect 8228 -4873 8262 -4487
rect 7136 -4969 8166 -4935
rect 16136 -4425 17166 -4391
rect 16040 -4873 16074 -4487
rect 17228 -4873 17262 -4487
rect 16136 -4969 17166 -4935
rect 7136 -6225 8166 -6191
rect 7040 -6673 7074 -6287
rect 8228 -6673 8262 -6287
rect 7136 -6769 8166 -6735
rect 16136 -6225 17166 -6191
rect 16040 -6673 16074 -6287
rect 17228 -6673 17262 -6287
rect 16136 -6769 17166 -6735
rect -7282 -7233 3426 -7140
<< poly >>
rect 7138 2707 8164 2723
rect 7138 2673 7154 2707
rect 7188 2673 7346 2707
rect 7380 2673 7538 2707
rect 7572 2673 7730 2707
rect 7764 2673 7922 2707
rect 7956 2673 8114 2707
rect 8148 2673 8164 2707
rect 7138 2657 8164 2673
rect 7204 2625 7234 2657
rect 7300 2625 7330 2657
rect 7396 2625 7426 2657
rect 7492 2625 7522 2657
rect 7588 2625 7618 2657
rect 7684 2625 7714 2657
rect 7780 2625 7810 2657
rect 7876 2625 7906 2657
rect 7972 2625 8002 2657
rect 8068 2625 8098 2657
rect 7204 2327 7234 2353
rect 7300 2327 7330 2353
rect 7396 2327 7426 2353
rect 7492 2327 7522 2353
rect 7588 2327 7618 2353
rect 7684 2327 7714 2353
rect 7780 2327 7810 2353
rect 7876 2327 7906 2353
rect 7972 2327 8002 2353
rect 8068 2327 8098 2353
rect 16138 2707 17164 2723
rect 16138 2673 16154 2707
rect 16188 2673 16346 2707
rect 16380 2673 16538 2707
rect 16572 2673 16730 2707
rect 16764 2673 16922 2707
rect 16956 2673 17114 2707
rect 17148 2673 17164 2707
rect 16138 2657 17164 2673
rect 16204 2625 16234 2657
rect 16300 2625 16330 2657
rect 16396 2625 16426 2657
rect 16492 2625 16522 2657
rect 16588 2625 16618 2657
rect 16684 2625 16714 2657
rect 16780 2625 16810 2657
rect 16876 2625 16906 2657
rect 16972 2625 17002 2657
rect 17068 2625 17098 2657
rect 16204 2327 16234 2353
rect 16300 2327 16330 2353
rect 16396 2327 16426 2353
rect 16492 2327 16522 2353
rect 16588 2327 16618 2353
rect 16684 2327 16714 2353
rect 16780 2327 16810 2353
rect 16876 2327 16906 2353
rect 16972 2327 17002 2353
rect 17068 2327 17098 2353
rect 7204 2045 7234 2071
rect 7300 2045 7330 2071
rect 7396 2045 7426 2071
rect 7492 2045 7522 2071
rect 7588 2045 7618 2071
rect 7684 2045 7714 2071
rect 7780 2045 7810 2071
rect 7876 2045 7906 2071
rect 7972 2045 8002 2071
rect 8068 2045 8098 2071
rect 7204 1919 7234 1941
rect 7300 1919 7330 1941
rect 7396 1919 7426 1941
rect 7492 1919 7522 1941
rect 7588 1919 7618 1941
rect 7684 1919 7714 1941
rect 7780 1919 7810 1941
rect 7876 1919 7906 1941
rect 7972 1919 8002 1941
rect 8068 1919 8098 1941
rect 7138 1899 8164 1919
rect 7138 1865 7154 1899
rect 7188 1865 7346 1899
rect 7380 1865 7538 1899
rect 7572 1865 7730 1899
rect 7764 1865 7922 1899
rect 7956 1865 8114 1899
rect 8148 1865 8164 1899
rect 7138 1853 8164 1865
rect 16204 2045 16234 2071
rect 16300 2045 16330 2071
rect 16396 2045 16426 2071
rect 16492 2045 16522 2071
rect 16588 2045 16618 2071
rect 16684 2045 16714 2071
rect 16780 2045 16810 2071
rect 16876 2045 16906 2071
rect 16972 2045 17002 2071
rect 17068 2045 17098 2071
rect 16204 1919 16234 1941
rect 16300 1919 16330 1941
rect 16396 1919 16426 1941
rect 16492 1919 16522 1941
rect 16588 1919 16618 1941
rect 16684 1919 16714 1941
rect 16780 1919 16810 1941
rect 16876 1919 16906 1941
rect 16972 1919 17002 1941
rect 17068 1919 17098 1941
rect 16138 1899 17164 1919
rect 16138 1865 16154 1899
rect 16188 1865 16346 1899
rect 16380 1865 16538 1899
rect 16572 1865 16730 1899
rect 16764 1865 16922 1899
rect 16956 1865 17114 1899
rect 17148 1865 17164 1899
rect 16138 1853 17164 1865
rect 7138 907 8164 923
rect 7138 873 7154 907
rect 7188 873 7346 907
rect 7380 873 7538 907
rect 7572 873 7730 907
rect 7764 873 7922 907
rect 7956 873 8114 907
rect 8148 873 8164 907
rect 7138 857 8164 873
rect 7204 825 7234 857
rect 7300 825 7330 857
rect 7396 825 7426 857
rect 7492 825 7522 857
rect 7588 825 7618 857
rect 7684 825 7714 857
rect 7780 825 7810 857
rect 7876 825 7906 857
rect 7972 825 8002 857
rect 8068 825 8098 857
rect 7204 527 7234 553
rect 7300 527 7330 553
rect 7396 527 7426 553
rect 7492 527 7522 553
rect 7588 527 7618 553
rect 7684 527 7714 553
rect 7780 527 7810 553
rect 7876 527 7906 553
rect 7972 527 8002 553
rect 8068 527 8098 553
rect 16138 907 17164 923
rect 16138 873 16154 907
rect 16188 873 16346 907
rect 16380 873 16538 907
rect 16572 873 16730 907
rect 16764 873 16922 907
rect 16956 873 17114 907
rect 17148 873 17164 907
rect 16138 857 17164 873
rect 16204 825 16234 857
rect 16300 825 16330 857
rect 16396 825 16426 857
rect 16492 825 16522 857
rect 16588 825 16618 857
rect 16684 825 16714 857
rect 16780 825 16810 857
rect 16876 825 16906 857
rect 16972 825 17002 857
rect 17068 825 17098 857
rect 16204 527 16234 553
rect 16300 527 16330 553
rect 16396 527 16426 553
rect 16492 527 16522 553
rect 16588 527 16618 553
rect 16684 527 16714 553
rect 16780 527 16810 553
rect 16876 527 16906 553
rect 16972 527 17002 553
rect 17068 527 17098 553
rect 7204 245 7234 271
rect 7300 245 7330 271
rect 7396 245 7426 271
rect 7492 245 7522 271
rect 7588 245 7618 271
rect 7684 245 7714 271
rect 7780 245 7810 271
rect 7876 245 7906 271
rect 7972 245 8002 271
rect 8068 245 8098 271
rect 7204 119 7234 141
rect 7300 119 7330 141
rect 7396 119 7426 141
rect 7492 119 7522 141
rect 7588 119 7618 141
rect 7684 119 7714 141
rect 7780 119 7810 141
rect 7876 119 7906 141
rect 7972 119 8002 141
rect 8068 119 8098 141
rect 7138 99 8164 119
rect 7138 65 7154 99
rect 7188 65 7346 99
rect 7380 65 7538 99
rect 7572 65 7730 99
rect 7764 65 7922 99
rect 7956 65 8114 99
rect 8148 65 8164 99
rect 7138 53 8164 65
rect 16204 245 16234 271
rect 16300 245 16330 271
rect 16396 245 16426 271
rect 16492 245 16522 271
rect 16588 245 16618 271
rect 16684 245 16714 271
rect 16780 245 16810 271
rect 16876 245 16906 271
rect 16972 245 17002 271
rect 17068 245 17098 271
rect 16204 119 16234 141
rect 16300 119 16330 141
rect 16396 119 16426 141
rect 16492 119 16522 141
rect 16588 119 16618 141
rect 16684 119 16714 141
rect 16780 119 16810 141
rect 16876 119 16906 141
rect 16972 119 17002 141
rect 17068 119 17098 141
rect 16138 99 17164 119
rect 16138 65 16154 99
rect 16188 65 16346 99
rect 16380 65 16538 99
rect 16572 65 16730 99
rect 16764 65 16922 99
rect 16956 65 17114 99
rect 17148 65 17164 99
rect 16138 53 17164 65
rect 7138 -893 8164 -877
rect 7138 -927 7154 -893
rect 7188 -927 7346 -893
rect 7380 -927 7538 -893
rect 7572 -927 7730 -893
rect 7764 -927 7922 -893
rect 7956 -927 8114 -893
rect 8148 -927 8164 -893
rect 7138 -943 8164 -927
rect 7204 -975 7234 -943
rect 7300 -975 7330 -943
rect 7396 -975 7426 -943
rect 7492 -975 7522 -943
rect 7588 -975 7618 -943
rect 7684 -975 7714 -943
rect 7780 -975 7810 -943
rect 7876 -975 7906 -943
rect 7972 -975 8002 -943
rect 8068 -975 8098 -943
rect 7204 -1273 7234 -1247
rect 7300 -1273 7330 -1247
rect 7396 -1273 7426 -1247
rect 7492 -1273 7522 -1247
rect 7588 -1273 7618 -1247
rect 7684 -1273 7714 -1247
rect 7780 -1273 7810 -1247
rect 7876 -1273 7906 -1247
rect 7972 -1273 8002 -1247
rect 8068 -1273 8098 -1247
rect 16138 -893 17164 -877
rect 16138 -927 16154 -893
rect 16188 -927 16346 -893
rect 16380 -927 16538 -893
rect 16572 -927 16730 -893
rect 16764 -927 16922 -893
rect 16956 -927 17114 -893
rect 17148 -927 17164 -893
rect 16138 -943 17164 -927
rect 16204 -975 16234 -943
rect 16300 -975 16330 -943
rect 16396 -975 16426 -943
rect 16492 -975 16522 -943
rect 16588 -975 16618 -943
rect 16684 -975 16714 -943
rect 16780 -975 16810 -943
rect 16876 -975 16906 -943
rect 16972 -975 17002 -943
rect 17068 -975 17098 -943
rect 16204 -1273 16234 -1247
rect 16300 -1273 16330 -1247
rect 16396 -1273 16426 -1247
rect 16492 -1273 16522 -1247
rect 16588 -1273 16618 -1247
rect 16684 -1273 16714 -1247
rect 16780 -1273 16810 -1247
rect 16876 -1273 16906 -1247
rect 16972 -1273 17002 -1247
rect 17068 -1273 17098 -1247
rect -6234 -2039 -6158 -2023
rect -6234 -2055 -6218 -2039
rect -6256 -2073 -6218 -2055
rect -6174 -2055 -6158 -2039
rect -6056 -2039 -5980 -2023
rect -6056 -2055 -6040 -2039
rect -6174 -2073 -6136 -2055
rect -6256 -2120 -6136 -2073
rect -6078 -2073 -6040 -2055
rect -5996 -2055 -5980 -2039
rect -5878 -2039 -5802 -2023
rect -5878 -2055 -5862 -2039
rect -5996 -2073 -5958 -2055
rect -6078 -2120 -5958 -2073
rect -5900 -2073 -5862 -2055
rect -5818 -2055 -5802 -2039
rect -5700 -2039 -5624 -2023
rect -5700 -2055 -5684 -2039
rect -5818 -2073 -5780 -2055
rect -5900 -2120 -5780 -2073
rect -5722 -2073 -5684 -2055
rect -5640 -2055 -5624 -2039
rect -5522 -2039 -5446 -2023
rect -5522 -2055 -5506 -2039
rect -5640 -2073 -5602 -2055
rect -5722 -2120 -5602 -2073
rect -5544 -2073 -5506 -2055
rect -5462 -2055 -5446 -2039
rect -5344 -2039 -5268 -2023
rect -5344 -2055 -5328 -2039
rect -5462 -2073 -5424 -2055
rect -5544 -2120 -5424 -2073
rect -5366 -2073 -5328 -2055
rect -5284 -2055 -5268 -2039
rect -5166 -2039 -5090 -2023
rect -5166 -2055 -5150 -2039
rect -5284 -2073 -5246 -2055
rect -5366 -2120 -5246 -2073
rect -5188 -2073 -5150 -2055
rect -5106 -2055 -5090 -2039
rect -4988 -2039 -4912 -2023
rect -4988 -2055 -4972 -2039
rect -5106 -2073 -5068 -2055
rect -5188 -2120 -5068 -2073
rect -5010 -2073 -4972 -2055
rect -4928 -2055 -4912 -2039
rect -4810 -2039 -4734 -2023
rect -4810 -2055 -4794 -2039
rect -4928 -2073 -4890 -2055
rect -5010 -2120 -4890 -2073
rect -4832 -2073 -4794 -2055
rect -4750 -2055 -4734 -2039
rect -4632 -2039 -4556 -2023
rect -4632 -2055 -4616 -2039
rect -4750 -2073 -4712 -2055
rect -4832 -2120 -4712 -2073
rect -4654 -2073 -4616 -2055
rect -4572 -2055 -4556 -2039
rect -4454 -2039 -4378 -2023
rect -4454 -2055 -4438 -2039
rect -4572 -2073 -4534 -2055
rect -4654 -2120 -4534 -2073
rect -4476 -2073 -4438 -2055
rect -4394 -2055 -4378 -2039
rect -4276 -2039 -4200 -2023
rect -4276 -2055 -4260 -2039
rect -4394 -2073 -4356 -2055
rect -4476 -2120 -4356 -2073
rect -4298 -2073 -4260 -2055
rect -4216 -2055 -4200 -2039
rect -4098 -2039 -4022 -2023
rect -4098 -2055 -4082 -2039
rect -4216 -2073 -4178 -2055
rect -4298 -2120 -4178 -2073
rect -4120 -2073 -4082 -2055
rect -4038 -2055 -4022 -2039
rect -3920 -2039 -3844 -2023
rect -3920 -2055 -3904 -2039
rect -4038 -2073 -4000 -2055
rect -4120 -2120 -4000 -2073
rect -3942 -2073 -3904 -2055
rect -3860 -2055 -3844 -2039
rect -3742 -2039 -3666 -2023
rect -3742 -2055 -3726 -2039
rect -3860 -2073 -3822 -2055
rect -3942 -2120 -3822 -2073
rect -3764 -2073 -3726 -2055
rect -3682 -2055 -3666 -2039
rect -3564 -2039 -3488 -2023
rect -3564 -2055 -3548 -2039
rect -3682 -2073 -3644 -2055
rect -3764 -2120 -3644 -2073
rect -3586 -2073 -3548 -2055
rect -3504 -2055 -3488 -2039
rect -3504 -2073 -3466 -2055
rect -3586 -2120 -3466 -2073
rect -6256 -2447 -6136 -2400
rect -6256 -2465 -6218 -2447
rect -6234 -2481 -6218 -2465
rect -6174 -2465 -6136 -2447
rect -6078 -2447 -5958 -2400
rect -6078 -2465 -6040 -2447
rect -6174 -2481 -6158 -2465
rect -6234 -2497 -6158 -2481
rect -6056 -2481 -6040 -2465
rect -5996 -2465 -5958 -2447
rect -5900 -2447 -5780 -2400
rect -5900 -2465 -5862 -2447
rect -5996 -2481 -5980 -2465
rect -6056 -2497 -5980 -2481
rect -5878 -2481 -5862 -2465
rect -5818 -2465 -5780 -2447
rect -5722 -2447 -5602 -2400
rect -5722 -2465 -5684 -2447
rect -5818 -2481 -5802 -2465
rect -5878 -2497 -5802 -2481
rect -5700 -2481 -5684 -2465
rect -5640 -2465 -5602 -2447
rect -5544 -2447 -5424 -2400
rect -5544 -2465 -5506 -2447
rect -5640 -2481 -5624 -2465
rect -5700 -2497 -5624 -2481
rect -5522 -2481 -5506 -2465
rect -5462 -2465 -5424 -2447
rect -5366 -2447 -5246 -2400
rect -5366 -2465 -5328 -2447
rect -5462 -2481 -5446 -2465
rect -5522 -2497 -5446 -2481
rect -5344 -2481 -5328 -2465
rect -5284 -2465 -5246 -2447
rect -5188 -2447 -5068 -2400
rect -5188 -2465 -5150 -2447
rect -5284 -2481 -5268 -2465
rect -5344 -2497 -5268 -2481
rect -5166 -2481 -5150 -2465
rect -5106 -2465 -5068 -2447
rect -5010 -2447 -4890 -2400
rect -5010 -2465 -4972 -2447
rect -5106 -2481 -5090 -2465
rect -5166 -2497 -5090 -2481
rect -4988 -2481 -4972 -2465
rect -4928 -2465 -4890 -2447
rect -4832 -2447 -4712 -2400
rect -4832 -2465 -4794 -2447
rect -4928 -2481 -4912 -2465
rect -4988 -2497 -4912 -2481
rect -4810 -2481 -4794 -2465
rect -4750 -2465 -4712 -2447
rect -4654 -2447 -4534 -2400
rect -4654 -2465 -4616 -2447
rect -4750 -2481 -4734 -2465
rect -4810 -2497 -4734 -2481
rect -4632 -2481 -4616 -2465
rect -4572 -2465 -4534 -2447
rect -4476 -2447 -4356 -2400
rect -4476 -2465 -4438 -2447
rect -4572 -2481 -4556 -2465
rect -4632 -2497 -4556 -2481
rect -4454 -2481 -4438 -2465
rect -4394 -2465 -4356 -2447
rect -4298 -2447 -4178 -2400
rect -4298 -2465 -4260 -2447
rect -4394 -2481 -4378 -2465
rect -4454 -2497 -4378 -2481
rect -4276 -2481 -4260 -2465
rect -4216 -2465 -4178 -2447
rect -4120 -2447 -4000 -2400
rect -4120 -2465 -4082 -2447
rect -4216 -2481 -4200 -2465
rect -4276 -2497 -4200 -2481
rect -4098 -2481 -4082 -2465
rect -4038 -2465 -4000 -2447
rect -3942 -2447 -3822 -2400
rect -3942 -2465 -3904 -2447
rect -4038 -2481 -4022 -2465
rect -4098 -2497 -4022 -2481
rect -3920 -2481 -3904 -2465
rect -3860 -2465 -3822 -2447
rect -3764 -2447 -3644 -2400
rect -3764 -2465 -3726 -2447
rect -3860 -2481 -3844 -2465
rect -3920 -2497 -3844 -2481
rect -3742 -2481 -3726 -2465
rect -3682 -2465 -3644 -2447
rect -3586 -2447 -3466 -2400
rect -3586 -2465 -3548 -2447
rect -3682 -2481 -3666 -2465
rect -3742 -2497 -3666 -2481
rect -3564 -2481 -3548 -2465
rect -3504 -2465 -3466 -2447
rect -3504 -2481 -3488 -2465
rect -3564 -2497 -3488 -2481
rect -1386 -2791 -1310 -2775
rect -1386 -2807 -1370 -2791
rect -1408 -2825 -1370 -2807
rect -1326 -2807 -1310 -2791
rect -1208 -2791 -1132 -2775
rect -1208 -2807 -1192 -2791
rect -1326 -2825 -1288 -2807
rect -1408 -2872 -1288 -2825
rect -1230 -2825 -1192 -2807
rect -1148 -2807 -1132 -2791
rect -1030 -2791 -954 -2775
rect -1030 -2807 -1014 -2791
rect -1148 -2825 -1110 -2807
rect -1230 -2872 -1110 -2825
rect -1052 -2825 -1014 -2807
rect -970 -2807 -954 -2791
rect -852 -2791 -776 -2775
rect -852 -2807 -836 -2791
rect -970 -2825 -932 -2807
rect -1052 -2872 -932 -2825
rect -874 -2825 -836 -2807
rect -792 -2807 -776 -2791
rect -674 -2791 -598 -2775
rect -674 -2807 -658 -2791
rect -792 -2825 -754 -2807
rect -874 -2872 -754 -2825
rect -696 -2825 -658 -2807
rect -614 -2807 -598 -2791
rect -496 -2791 -420 -2775
rect -496 -2807 -480 -2791
rect -614 -2825 -576 -2807
rect -696 -2872 -576 -2825
rect -518 -2825 -480 -2807
rect -436 -2807 -420 -2791
rect -318 -2791 -242 -2775
rect -318 -2807 -302 -2791
rect -436 -2825 -398 -2807
rect -518 -2872 -398 -2825
rect -340 -2825 -302 -2807
rect -258 -2807 -242 -2791
rect -140 -2791 -64 -2775
rect -140 -2807 -124 -2791
rect -258 -2825 -220 -2807
rect -340 -2872 -220 -2825
rect -162 -2825 -124 -2807
rect -80 -2807 -64 -2791
rect 38 -2791 114 -2775
rect 38 -2807 54 -2791
rect -80 -2825 -42 -2807
rect -162 -2872 -42 -2825
rect 16 -2825 54 -2807
rect 98 -2807 114 -2791
rect 216 -2791 292 -2775
rect 216 -2807 232 -2791
rect 98 -2825 136 -2807
rect 16 -2872 136 -2825
rect 194 -2825 232 -2807
rect 276 -2807 292 -2791
rect 394 -2791 470 -2775
rect 394 -2807 410 -2791
rect 276 -2825 314 -2807
rect 194 -2872 314 -2825
rect 372 -2825 410 -2807
rect 454 -2807 470 -2791
rect 572 -2791 648 -2775
rect 572 -2807 588 -2791
rect 454 -2825 492 -2807
rect 372 -2872 492 -2825
rect 550 -2825 588 -2807
rect 632 -2807 648 -2791
rect 750 -2791 826 -2775
rect 750 -2807 766 -2791
rect 632 -2825 670 -2807
rect 550 -2872 670 -2825
rect 728 -2825 766 -2807
rect 810 -2807 826 -2791
rect 928 -2791 1004 -2775
rect 928 -2807 944 -2791
rect 810 -2825 848 -2807
rect 728 -2872 848 -2825
rect 906 -2825 944 -2807
rect 988 -2807 1004 -2791
rect 1106 -2791 1182 -2775
rect 1106 -2807 1122 -2791
rect 988 -2825 1026 -2807
rect 906 -2872 1026 -2825
rect 1084 -2825 1122 -2807
rect 1166 -2807 1182 -2791
rect 1284 -2791 1360 -2775
rect 1284 -2807 1300 -2791
rect 1166 -2825 1204 -2807
rect 1084 -2872 1204 -2825
rect 1262 -2825 1300 -2807
rect 1344 -2807 1360 -2791
rect 1462 -2791 1538 -2775
rect 1462 -2807 1478 -2791
rect 1344 -2825 1382 -2807
rect 1262 -2872 1382 -2825
rect 1440 -2825 1478 -2807
rect 1522 -2807 1538 -2791
rect 1640 -2791 1716 -2775
rect 1640 -2807 1656 -2791
rect 1522 -2825 1560 -2807
rect 1440 -2872 1560 -2825
rect 1618 -2825 1656 -2807
rect 1700 -2807 1716 -2791
rect 1818 -2791 1894 -2775
rect 1818 -2807 1834 -2791
rect 1700 -2825 1738 -2807
rect 1618 -2872 1738 -2825
rect 1796 -2825 1834 -2807
rect 1878 -2807 1894 -2791
rect 1996 -2791 2072 -2775
rect 1996 -2807 2012 -2791
rect 1878 -2825 1916 -2807
rect 1796 -2872 1916 -2825
rect 1974 -2825 2012 -2807
rect 2056 -2807 2072 -2791
rect 2174 -2791 2250 -2775
rect 2174 -2807 2190 -2791
rect 2056 -2825 2094 -2807
rect 1974 -2872 2094 -2825
rect 2152 -2825 2190 -2807
rect 2234 -2807 2250 -2791
rect 2352 -2791 2428 -2775
rect 2352 -2807 2368 -2791
rect 2234 -2825 2272 -2807
rect 2152 -2872 2272 -2825
rect 2330 -2825 2368 -2807
rect 2412 -2807 2428 -2791
rect 2530 -2791 2606 -2775
rect 2530 -2807 2546 -2791
rect 2412 -2825 2450 -2807
rect 2330 -2872 2450 -2825
rect 2508 -2825 2546 -2807
rect 2590 -2807 2606 -2791
rect 2590 -2825 2628 -2807
rect 2508 -2872 2628 -2825
rect -6234 -2909 -6158 -2893
rect -6234 -2925 -6218 -2909
rect -6256 -2943 -6218 -2925
rect -6174 -2925 -6158 -2909
rect -6056 -2909 -5980 -2893
rect -6056 -2925 -6040 -2909
rect -6174 -2943 -6136 -2925
rect -6256 -2990 -6136 -2943
rect -6078 -2943 -6040 -2925
rect -5996 -2925 -5980 -2909
rect -5878 -2909 -5802 -2893
rect -5878 -2925 -5862 -2909
rect -5996 -2943 -5958 -2925
rect -6078 -2990 -5958 -2943
rect -5900 -2943 -5862 -2925
rect -5818 -2925 -5802 -2909
rect -5700 -2909 -5624 -2893
rect -5700 -2925 -5684 -2909
rect -5818 -2943 -5780 -2925
rect -5900 -2990 -5780 -2943
rect -5722 -2943 -5684 -2925
rect -5640 -2925 -5624 -2909
rect -5522 -2909 -5446 -2893
rect -5522 -2925 -5506 -2909
rect -5640 -2943 -5602 -2925
rect -5722 -2990 -5602 -2943
rect -5544 -2943 -5506 -2925
rect -5462 -2925 -5446 -2909
rect -5344 -2909 -5268 -2893
rect -5344 -2925 -5328 -2909
rect -5462 -2943 -5424 -2925
rect -5544 -2990 -5424 -2943
rect -5366 -2943 -5328 -2925
rect -5284 -2925 -5268 -2909
rect -5166 -2909 -5090 -2893
rect -5166 -2925 -5150 -2909
rect -5284 -2943 -5246 -2925
rect -5366 -2990 -5246 -2943
rect -5188 -2943 -5150 -2925
rect -5106 -2925 -5090 -2909
rect -4988 -2909 -4912 -2893
rect -4988 -2925 -4972 -2909
rect -5106 -2943 -5068 -2925
rect -5188 -2990 -5068 -2943
rect -5010 -2943 -4972 -2925
rect -4928 -2925 -4912 -2909
rect -4810 -2909 -4734 -2893
rect -4810 -2925 -4794 -2909
rect -4928 -2943 -4890 -2925
rect -5010 -2990 -4890 -2943
rect -4832 -2943 -4794 -2925
rect -4750 -2925 -4734 -2909
rect -4632 -2909 -4556 -2893
rect -4632 -2925 -4616 -2909
rect -4750 -2943 -4712 -2925
rect -4832 -2990 -4712 -2943
rect -4654 -2943 -4616 -2925
rect -4572 -2925 -4556 -2909
rect -4454 -2909 -4378 -2893
rect -4454 -2925 -4438 -2909
rect -4572 -2943 -4534 -2925
rect -4654 -2990 -4534 -2943
rect -4476 -2943 -4438 -2925
rect -4394 -2925 -4378 -2909
rect -4276 -2909 -4200 -2893
rect -4276 -2925 -4260 -2909
rect -4394 -2943 -4356 -2925
rect -4476 -2990 -4356 -2943
rect -4298 -2943 -4260 -2925
rect -4216 -2925 -4200 -2909
rect -4098 -2909 -4022 -2893
rect -4098 -2925 -4082 -2909
rect -4216 -2943 -4178 -2925
rect -4298 -2990 -4178 -2943
rect -4120 -2943 -4082 -2925
rect -4038 -2925 -4022 -2909
rect -3920 -2909 -3844 -2893
rect -3920 -2925 -3904 -2909
rect -4038 -2943 -4000 -2925
rect -4120 -2990 -4000 -2943
rect -3942 -2943 -3904 -2925
rect -3860 -2925 -3844 -2909
rect -3742 -2909 -3666 -2893
rect -3742 -2925 -3726 -2909
rect -3860 -2943 -3822 -2925
rect -3942 -2990 -3822 -2943
rect -3764 -2943 -3726 -2925
rect -3682 -2925 -3666 -2909
rect -3564 -2909 -3488 -2893
rect -3564 -2925 -3548 -2909
rect -3682 -2943 -3644 -2925
rect -3764 -2990 -3644 -2943
rect -3586 -2943 -3548 -2925
rect -3504 -2925 -3488 -2909
rect -3504 -2943 -3466 -2925
rect -3586 -2990 -3466 -2943
rect -1408 -3199 -1288 -3152
rect -1408 -3217 -1370 -3199
rect -1386 -3233 -1370 -3217
rect -1326 -3217 -1288 -3199
rect -1230 -3199 -1110 -3152
rect -1230 -3217 -1192 -3199
rect -1326 -3233 -1310 -3217
rect -1386 -3249 -1310 -3233
rect -1208 -3233 -1192 -3217
rect -1148 -3217 -1110 -3199
rect -1052 -3199 -932 -3152
rect -1052 -3217 -1014 -3199
rect -1148 -3233 -1132 -3217
rect -1208 -3249 -1132 -3233
rect -1030 -3233 -1014 -3217
rect -970 -3217 -932 -3199
rect -874 -3199 -754 -3152
rect -874 -3217 -836 -3199
rect -970 -3233 -954 -3217
rect -1030 -3249 -954 -3233
rect -852 -3233 -836 -3217
rect -792 -3217 -754 -3199
rect -696 -3199 -576 -3152
rect -696 -3217 -658 -3199
rect -792 -3233 -776 -3217
rect -852 -3249 -776 -3233
rect -674 -3233 -658 -3217
rect -614 -3217 -576 -3199
rect -518 -3199 -398 -3152
rect -518 -3217 -480 -3199
rect -614 -3233 -598 -3217
rect -674 -3249 -598 -3233
rect -496 -3233 -480 -3217
rect -436 -3217 -398 -3199
rect -340 -3199 -220 -3152
rect -340 -3217 -302 -3199
rect -436 -3233 -420 -3217
rect -496 -3249 -420 -3233
rect -318 -3233 -302 -3217
rect -258 -3217 -220 -3199
rect -162 -3199 -42 -3152
rect -162 -3217 -124 -3199
rect -258 -3233 -242 -3217
rect -318 -3249 -242 -3233
rect -140 -3233 -124 -3217
rect -80 -3217 -42 -3199
rect 16 -3199 136 -3152
rect 16 -3217 54 -3199
rect -80 -3233 -64 -3217
rect -140 -3249 -64 -3233
rect 38 -3233 54 -3217
rect 98 -3217 136 -3199
rect 194 -3199 314 -3152
rect 194 -3217 232 -3199
rect 98 -3233 114 -3217
rect 38 -3249 114 -3233
rect 216 -3233 232 -3217
rect 276 -3217 314 -3199
rect 372 -3199 492 -3152
rect 372 -3217 410 -3199
rect 276 -3233 292 -3217
rect 216 -3249 292 -3233
rect 394 -3233 410 -3217
rect 454 -3217 492 -3199
rect 550 -3199 670 -3152
rect 550 -3217 588 -3199
rect 454 -3233 470 -3217
rect 394 -3249 470 -3233
rect 572 -3233 588 -3217
rect 632 -3217 670 -3199
rect 728 -3199 848 -3152
rect 728 -3217 766 -3199
rect 632 -3233 648 -3217
rect 572 -3249 648 -3233
rect 750 -3233 766 -3217
rect 810 -3217 848 -3199
rect 906 -3199 1026 -3152
rect 906 -3217 944 -3199
rect 810 -3233 826 -3217
rect 750 -3249 826 -3233
rect 928 -3233 944 -3217
rect 988 -3217 1026 -3199
rect 1084 -3199 1204 -3152
rect 1084 -3217 1122 -3199
rect 988 -3233 1004 -3217
rect 928 -3249 1004 -3233
rect 1106 -3233 1122 -3217
rect 1166 -3217 1204 -3199
rect 1262 -3199 1382 -3152
rect 1262 -3217 1300 -3199
rect 1166 -3233 1182 -3217
rect 1106 -3249 1182 -3233
rect 1284 -3233 1300 -3217
rect 1344 -3217 1382 -3199
rect 1440 -3199 1560 -3152
rect 1440 -3217 1478 -3199
rect 1344 -3233 1360 -3217
rect 1284 -3249 1360 -3233
rect 1462 -3233 1478 -3217
rect 1522 -3217 1560 -3199
rect 1618 -3199 1738 -3152
rect 1618 -3217 1656 -3199
rect 1522 -3233 1538 -3217
rect 1462 -3249 1538 -3233
rect 1640 -3233 1656 -3217
rect 1700 -3217 1738 -3199
rect 1796 -3199 1916 -3152
rect 1796 -3217 1834 -3199
rect 1700 -3233 1716 -3217
rect 1640 -3249 1716 -3233
rect 1818 -3233 1834 -3217
rect 1878 -3217 1916 -3199
rect 1974 -3199 2094 -3152
rect 1974 -3217 2012 -3199
rect 1878 -3233 1894 -3217
rect 1818 -3249 1894 -3233
rect 1996 -3233 2012 -3217
rect 2056 -3217 2094 -3199
rect 2152 -3199 2272 -3152
rect 2152 -3217 2190 -3199
rect 2056 -3233 2072 -3217
rect 1996 -3249 2072 -3233
rect 2174 -3233 2190 -3217
rect 2234 -3217 2272 -3199
rect 2330 -3199 2450 -3152
rect 2330 -3217 2368 -3199
rect 2234 -3233 2250 -3217
rect 2174 -3249 2250 -3233
rect 2352 -3233 2368 -3217
rect 2412 -3217 2450 -3199
rect 2508 -3199 2628 -3152
rect 2508 -3217 2546 -3199
rect 2412 -3233 2428 -3217
rect 2352 -3249 2428 -3233
rect 2530 -3233 2546 -3217
rect 2590 -3217 2628 -3199
rect 2590 -3233 2606 -3217
rect 2530 -3249 2606 -3233
rect -6256 -3317 -6136 -3270
rect -6256 -3335 -6218 -3317
rect -6234 -3351 -6218 -3335
rect -6174 -3335 -6136 -3317
rect -6078 -3317 -5958 -3270
rect -6078 -3335 -6040 -3317
rect -6174 -3351 -6158 -3335
rect -6234 -3367 -6158 -3351
rect -6056 -3351 -6040 -3335
rect -5996 -3335 -5958 -3317
rect -5900 -3317 -5780 -3270
rect -5900 -3335 -5862 -3317
rect -5996 -3351 -5980 -3335
rect -6056 -3367 -5980 -3351
rect -5878 -3351 -5862 -3335
rect -5818 -3335 -5780 -3317
rect -5722 -3317 -5602 -3270
rect -5722 -3335 -5684 -3317
rect -5818 -3351 -5802 -3335
rect -5878 -3367 -5802 -3351
rect -5700 -3351 -5684 -3335
rect -5640 -3335 -5602 -3317
rect -5544 -3317 -5424 -3270
rect -5544 -3335 -5506 -3317
rect -5640 -3351 -5624 -3335
rect -5700 -3367 -5624 -3351
rect -5522 -3351 -5506 -3335
rect -5462 -3335 -5424 -3317
rect -5366 -3317 -5246 -3270
rect -5366 -3335 -5328 -3317
rect -5462 -3351 -5446 -3335
rect -5522 -3367 -5446 -3351
rect -5344 -3351 -5328 -3335
rect -5284 -3335 -5246 -3317
rect -5188 -3317 -5068 -3270
rect -5188 -3335 -5150 -3317
rect -5284 -3351 -5268 -3335
rect -5344 -3367 -5268 -3351
rect -5166 -3351 -5150 -3335
rect -5106 -3335 -5068 -3317
rect -5010 -3317 -4890 -3270
rect -5010 -3335 -4972 -3317
rect -5106 -3351 -5090 -3335
rect -5166 -3367 -5090 -3351
rect -4988 -3351 -4972 -3335
rect -4928 -3335 -4890 -3317
rect -4832 -3317 -4712 -3270
rect -4832 -3335 -4794 -3317
rect -4928 -3351 -4912 -3335
rect -4988 -3367 -4912 -3351
rect -4810 -3351 -4794 -3335
rect -4750 -3335 -4712 -3317
rect -4654 -3317 -4534 -3270
rect -4654 -3335 -4616 -3317
rect -4750 -3351 -4734 -3335
rect -4810 -3367 -4734 -3351
rect -4632 -3351 -4616 -3335
rect -4572 -3335 -4534 -3317
rect -4476 -3317 -4356 -3270
rect -4476 -3335 -4438 -3317
rect -4572 -3351 -4556 -3335
rect -4632 -3367 -4556 -3351
rect -4454 -3351 -4438 -3335
rect -4394 -3335 -4356 -3317
rect -4298 -3317 -4178 -3270
rect -4298 -3335 -4260 -3317
rect -4394 -3351 -4378 -3335
rect -4454 -3367 -4378 -3351
rect -4276 -3351 -4260 -3335
rect -4216 -3335 -4178 -3317
rect -4120 -3317 -4000 -3270
rect -4120 -3335 -4082 -3317
rect -4216 -3351 -4200 -3335
rect -4276 -3367 -4200 -3351
rect -4098 -3351 -4082 -3335
rect -4038 -3335 -4000 -3317
rect -3942 -3317 -3822 -3270
rect -3942 -3335 -3904 -3317
rect -4038 -3351 -4022 -3335
rect -4098 -3367 -4022 -3351
rect -3920 -3351 -3904 -3335
rect -3860 -3335 -3822 -3317
rect -3764 -3317 -3644 -3270
rect -3764 -3335 -3726 -3317
rect -3860 -3351 -3844 -3335
rect -3920 -3367 -3844 -3351
rect -3742 -3351 -3726 -3335
rect -3682 -3335 -3644 -3317
rect -3586 -3317 -3466 -3270
rect -3586 -3335 -3548 -3317
rect -3682 -3351 -3666 -3335
rect -3742 -3367 -3666 -3351
rect -3564 -3351 -3548 -3335
rect -3504 -3335 -3466 -3317
rect -3504 -3351 -3488 -3335
rect -3564 -3367 -3488 -3351
rect -1386 -3691 -1310 -3675
rect -1386 -3707 -1370 -3691
rect -1408 -3725 -1370 -3707
rect -1326 -3707 -1310 -3691
rect -1208 -3691 -1132 -3675
rect -1208 -3707 -1192 -3691
rect -1326 -3725 -1288 -3707
rect -6234 -3779 -6158 -3763
rect -6234 -3795 -6218 -3779
rect -6256 -3813 -6218 -3795
rect -6174 -3795 -6158 -3779
rect -6056 -3779 -5980 -3763
rect -6056 -3795 -6040 -3779
rect -6174 -3813 -6136 -3795
rect -6256 -3860 -6136 -3813
rect -6078 -3813 -6040 -3795
rect -5996 -3795 -5980 -3779
rect -5878 -3779 -5802 -3763
rect -5878 -3795 -5862 -3779
rect -5996 -3813 -5958 -3795
rect -6078 -3860 -5958 -3813
rect -5900 -3813 -5862 -3795
rect -5818 -3795 -5802 -3779
rect -5700 -3779 -5624 -3763
rect -5700 -3795 -5684 -3779
rect -5818 -3813 -5780 -3795
rect -5900 -3860 -5780 -3813
rect -5722 -3813 -5684 -3795
rect -5640 -3795 -5624 -3779
rect -5522 -3779 -5446 -3763
rect -5522 -3795 -5506 -3779
rect -5640 -3813 -5602 -3795
rect -5722 -3860 -5602 -3813
rect -5544 -3813 -5506 -3795
rect -5462 -3795 -5446 -3779
rect -5344 -3779 -5268 -3763
rect -5344 -3795 -5328 -3779
rect -5462 -3813 -5424 -3795
rect -5544 -3860 -5424 -3813
rect -5366 -3813 -5328 -3795
rect -5284 -3795 -5268 -3779
rect -5166 -3779 -5090 -3763
rect -5166 -3795 -5150 -3779
rect -5284 -3813 -5246 -3795
rect -5366 -3860 -5246 -3813
rect -5188 -3813 -5150 -3795
rect -5106 -3795 -5090 -3779
rect -4988 -3779 -4912 -3763
rect -4988 -3795 -4972 -3779
rect -5106 -3813 -5068 -3795
rect -5188 -3860 -5068 -3813
rect -5010 -3813 -4972 -3795
rect -4928 -3795 -4912 -3779
rect -4810 -3779 -4734 -3763
rect -4810 -3795 -4794 -3779
rect -4928 -3813 -4890 -3795
rect -5010 -3860 -4890 -3813
rect -4832 -3813 -4794 -3795
rect -4750 -3795 -4734 -3779
rect -4632 -3779 -4556 -3763
rect -4632 -3795 -4616 -3779
rect -4750 -3813 -4712 -3795
rect -4832 -3860 -4712 -3813
rect -4654 -3813 -4616 -3795
rect -4572 -3795 -4556 -3779
rect -4454 -3779 -4378 -3763
rect -4454 -3795 -4438 -3779
rect -4572 -3813 -4534 -3795
rect -4654 -3860 -4534 -3813
rect -4476 -3813 -4438 -3795
rect -4394 -3795 -4378 -3779
rect -4276 -3779 -4200 -3763
rect -4276 -3795 -4260 -3779
rect -4394 -3813 -4356 -3795
rect -4476 -3860 -4356 -3813
rect -4298 -3813 -4260 -3795
rect -4216 -3795 -4200 -3779
rect -4098 -3779 -4022 -3763
rect -4098 -3795 -4082 -3779
rect -4216 -3813 -4178 -3795
rect -4298 -3860 -4178 -3813
rect -4120 -3813 -4082 -3795
rect -4038 -3795 -4022 -3779
rect -3920 -3779 -3844 -3763
rect -3920 -3795 -3904 -3779
rect -4038 -3813 -4000 -3795
rect -4120 -3860 -4000 -3813
rect -3942 -3813 -3904 -3795
rect -3860 -3795 -3844 -3779
rect -3742 -3779 -3666 -3763
rect -3742 -3795 -3726 -3779
rect -3860 -3813 -3822 -3795
rect -3942 -3860 -3822 -3813
rect -3764 -3813 -3726 -3795
rect -3682 -3795 -3666 -3779
rect -3564 -3779 -3488 -3763
rect -1408 -3772 -1288 -3725
rect -1230 -3725 -1192 -3707
rect -1148 -3707 -1132 -3691
rect -1030 -3691 -954 -3675
rect -1030 -3707 -1014 -3691
rect -1148 -3725 -1110 -3707
rect -1230 -3772 -1110 -3725
rect -1052 -3725 -1014 -3707
rect -970 -3707 -954 -3691
rect -852 -3691 -776 -3675
rect -852 -3707 -836 -3691
rect -970 -3725 -932 -3707
rect -1052 -3772 -932 -3725
rect -874 -3725 -836 -3707
rect -792 -3707 -776 -3691
rect -674 -3691 -598 -3675
rect -674 -3707 -658 -3691
rect -792 -3725 -754 -3707
rect -874 -3772 -754 -3725
rect -696 -3725 -658 -3707
rect -614 -3707 -598 -3691
rect -496 -3691 -420 -3675
rect -496 -3707 -480 -3691
rect -614 -3725 -576 -3707
rect -696 -3772 -576 -3725
rect -518 -3725 -480 -3707
rect -436 -3707 -420 -3691
rect -318 -3691 -242 -3675
rect -318 -3707 -302 -3691
rect -436 -3725 -398 -3707
rect -518 -3772 -398 -3725
rect -340 -3725 -302 -3707
rect -258 -3707 -242 -3691
rect -140 -3691 -64 -3675
rect -140 -3707 -124 -3691
rect -258 -3725 -220 -3707
rect -340 -3772 -220 -3725
rect -162 -3725 -124 -3707
rect -80 -3707 -64 -3691
rect 38 -3691 114 -3675
rect 38 -3707 54 -3691
rect -80 -3725 -42 -3707
rect -162 -3772 -42 -3725
rect 16 -3725 54 -3707
rect 98 -3707 114 -3691
rect 216 -3691 292 -3675
rect 216 -3707 232 -3691
rect 98 -3725 136 -3707
rect 16 -3772 136 -3725
rect 194 -3725 232 -3707
rect 276 -3707 292 -3691
rect 394 -3691 470 -3675
rect 394 -3707 410 -3691
rect 276 -3725 314 -3707
rect 194 -3772 314 -3725
rect 372 -3725 410 -3707
rect 454 -3707 470 -3691
rect 572 -3691 648 -3675
rect 572 -3707 588 -3691
rect 454 -3725 492 -3707
rect 372 -3772 492 -3725
rect 550 -3725 588 -3707
rect 632 -3707 648 -3691
rect 750 -3691 826 -3675
rect 750 -3707 766 -3691
rect 632 -3725 670 -3707
rect 550 -3772 670 -3725
rect 728 -3725 766 -3707
rect 810 -3707 826 -3691
rect 928 -3691 1004 -3675
rect 928 -3707 944 -3691
rect 810 -3725 848 -3707
rect 728 -3772 848 -3725
rect 906 -3725 944 -3707
rect 988 -3707 1004 -3691
rect 1106 -3691 1182 -3675
rect 1106 -3707 1122 -3691
rect 988 -3725 1026 -3707
rect 906 -3772 1026 -3725
rect 1084 -3725 1122 -3707
rect 1166 -3707 1182 -3691
rect 1284 -3691 1360 -3675
rect 1284 -3707 1300 -3691
rect 1166 -3725 1204 -3707
rect 1084 -3772 1204 -3725
rect 1262 -3725 1300 -3707
rect 1344 -3707 1360 -3691
rect 1462 -3691 1538 -3675
rect 1462 -3707 1478 -3691
rect 1344 -3725 1382 -3707
rect 1262 -3772 1382 -3725
rect 1440 -3725 1478 -3707
rect 1522 -3707 1538 -3691
rect 1640 -3691 1716 -3675
rect 1640 -3707 1656 -3691
rect 1522 -3725 1560 -3707
rect 1440 -3772 1560 -3725
rect 1618 -3725 1656 -3707
rect 1700 -3707 1716 -3691
rect 1818 -3691 1894 -3675
rect 1818 -3707 1834 -3691
rect 1700 -3725 1738 -3707
rect 1618 -3772 1738 -3725
rect 1796 -3725 1834 -3707
rect 1878 -3707 1894 -3691
rect 1996 -3691 2072 -3675
rect 1996 -3707 2012 -3691
rect 1878 -3725 1916 -3707
rect 1796 -3772 1916 -3725
rect 1974 -3725 2012 -3707
rect 2056 -3707 2072 -3691
rect 2174 -3691 2250 -3675
rect 2174 -3707 2190 -3691
rect 2056 -3725 2094 -3707
rect 1974 -3772 2094 -3725
rect 2152 -3725 2190 -3707
rect 2234 -3707 2250 -3691
rect 2352 -3691 2428 -3675
rect 2352 -3707 2368 -3691
rect 2234 -3725 2272 -3707
rect 2152 -3772 2272 -3725
rect 2330 -3725 2368 -3707
rect 2412 -3707 2428 -3691
rect 2530 -3691 2606 -3675
rect 2530 -3707 2546 -3691
rect 2412 -3725 2450 -3707
rect 2330 -3772 2450 -3725
rect 2508 -3725 2546 -3707
rect 2590 -3707 2606 -3691
rect 2590 -3725 2628 -3707
rect 2508 -3772 2628 -3725
rect -3564 -3795 -3548 -3779
rect -3682 -3813 -3644 -3795
rect -3764 -3860 -3644 -3813
rect -3586 -3813 -3548 -3795
rect -3504 -3795 -3488 -3779
rect -3504 -3813 -3466 -3795
rect -3586 -3860 -3466 -3813
rect -1408 -4099 -1288 -4052
rect -1408 -4117 -1370 -4099
rect -1386 -4133 -1370 -4117
rect -1326 -4117 -1288 -4099
rect -1230 -4099 -1110 -4052
rect -1230 -4117 -1192 -4099
rect -1326 -4133 -1310 -4117
rect -6256 -4187 -6136 -4140
rect -6256 -4205 -6218 -4187
rect -6234 -4221 -6218 -4205
rect -6174 -4205 -6136 -4187
rect -6078 -4187 -5958 -4140
rect -6078 -4205 -6040 -4187
rect -6174 -4221 -6158 -4205
rect -6234 -4237 -6158 -4221
rect -6056 -4221 -6040 -4205
rect -5996 -4205 -5958 -4187
rect -5900 -4187 -5780 -4140
rect -5900 -4205 -5862 -4187
rect -5996 -4221 -5980 -4205
rect -6056 -4237 -5980 -4221
rect -5878 -4221 -5862 -4205
rect -5818 -4205 -5780 -4187
rect -5722 -4187 -5602 -4140
rect -5722 -4205 -5684 -4187
rect -5818 -4221 -5802 -4205
rect -5878 -4237 -5802 -4221
rect -5700 -4221 -5684 -4205
rect -5640 -4205 -5602 -4187
rect -5544 -4187 -5424 -4140
rect -5544 -4205 -5506 -4187
rect -5640 -4221 -5624 -4205
rect -5700 -4237 -5624 -4221
rect -5522 -4221 -5506 -4205
rect -5462 -4205 -5424 -4187
rect -5366 -4187 -5246 -4140
rect -5366 -4205 -5328 -4187
rect -5462 -4221 -5446 -4205
rect -5522 -4237 -5446 -4221
rect -5344 -4221 -5328 -4205
rect -5284 -4205 -5246 -4187
rect -5188 -4187 -5068 -4140
rect -5188 -4205 -5150 -4187
rect -5284 -4221 -5268 -4205
rect -5344 -4237 -5268 -4221
rect -5166 -4221 -5150 -4205
rect -5106 -4205 -5068 -4187
rect -5010 -4187 -4890 -4140
rect -5010 -4205 -4972 -4187
rect -5106 -4221 -5090 -4205
rect -5166 -4237 -5090 -4221
rect -4988 -4221 -4972 -4205
rect -4928 -4205 -4890 -4187
rect -4832 -4187 -4712 -4140
rect -4832 -4205 -4794 -4187
rect -4928 -4221 -4912 -4205
rect -4988 -4237 -4912 -4221
rect -4810 -4221 -4794 -4205
rect -4750 -4205 -4712 -4187
rect -4654 -4187 -4534 -4140
rect -4654 -4205 -4616 -4187
rect -4750 -4221 -4734 -4205
rect -4810 -4237 -4734 -4221
rect -4632 -4221 -4616 -4205
rect -4572 -4205 -4534 -4187
rect -4476 -4187 -4356 -4140
rect -4476 -4205 -4438 -4187
rect -4572 -4221 -4556 -4205
rect -4632 -4237 -4556 -4221
rect -4454 -4221 -4438 -4205
rect -4394 -4205 -4356 -4187
rect -4298 -4187 -4178 -4140
rect -4298 -4205 -4260 -4187
rect -4394 -4221 -4378 -4205
rect -4454 -4237 -4378 -4221
rect -4276 -4221 -4260 -4205
rect -4216 -4205 -4178 -4187
rect -4120 -4187 -4000 -4140
rect -4120 -4205 -4082 -4187
rect -4216 -4221 -4200 -4205
rect -4276 -4237 -4200 -4221
rect -4098 -4221 -4082 -4205
rect -4038 -4205 -4000 -4187
rect -3942 -4187 -3822 -4140
rect -3942 -4205 -3904 -4187
rect -4038 -4221 -4022 -4205
rect -4098 -4237 -4022 -4221
rect -3920 -4221 -3904 -4205
rect -3860 -4205 -3822 -4187
rect -3764 -4187 -3644 -4140
rect -3764 -4205 -3726 -4187
rect -3860 -4221 -3844 -4205
rect -3920 -4237 -3844 -4221
rect -3742 -4221 -3726 -4205
rect -3682 -4205 -3644 -4187
rect -3586 -4187 -3466 -4140
rect -1386 -4149 -1310 -4133
rect -1208 -4133 -1192 -4117
rect -1148 -4117 -1110 -4099
rect -1052 -4099 -932 -4052
rect -1052 -4117 -1014 -4099
rect -1148 -4133 -1132 -4117
rect -1208 -4149 -1132 -4133
rect -1030 -4133 -1014 -4117
rect -970 -4117 -932 -4099
rect -874 -4099 -754 -4052
rect -874 -4117 -836 -4099
rect -970 -4133 -954 -4117
rect -1030 -4149 -954 -4133
rect -852 -4133 -836 -4117
rect -792 -4117 -754 -4099
rect -696 -4099 -576 -4052
rect -696 -4117 -658 -4099
rect -792 -4133 -776 -4117
rect -852 -4149 -776 -4133
rect -674 -4133 -658 -4117
rect -614 -4117 -576 -4099
rect -518 -4099 -398 -4052
rect -518 -4117 -480 -4099
rect -614 -4133 -598 -4117
rect -674 -4149 -598 -4133
rect -496 -4133 -480 -4117
rect -436 -4117 -398 -4099
rect -340 -4099 -220 -4052
rect -340 -4117 -302 -4099
rect -436 -4133 -420 -4117
rect -496 -4149 -420 -4133
rect -318 -4133 -302 -4117
rect -258 -4117 -220 -4099
rect -162 -4099 -42 -4052
rect -162 -4117 -124 -4099
rect -258 -4133 -242 -4117
rect -318 -4149 -242 -4133
rect -140 -4133 -124 -4117
rect -80 -4117 -42 -4099
rect 16 -4099 136 -4052
rect 16 -4117 54 -4099
rect -80 -4133 -64 -4117
rect -140 -4149 -64 -4133
rect 38 -4133 54 -4117
rect 98 -4117 136 -4099
rect 194 -4099 314 -4052
rect 194 -4117 232 -4099
rect 98 -4133 114 -4117
rect 38 -4149 114 -4133
rect 216 -4133 232 -4117
rect 276 -4117 314 -4099
rect 372 -4099 492 -4052
rect 372 -4117 410 -4099
rect 276 -4133 292 -4117
rect 216 -4149 292 -4133
rect 394 -4133 410 -4117
rect 454 -4117 492 -4099
rect 550 -4099 670 -4052
rect 550 -4117 588 -4099
rect 454 -4133 470 -4117
rect 394 -4149 470 -4133
rect 572 -4133 588 -4117
rect 632 -4117 670 -4099
rect 728 -4099 848 -4052
rect 728 -4117 766 -4099
rect 632 -4133 648 -4117
rect 572 -4149 648 -4133
rect 750 -4133 766 -4117
rect 810 -4117 848 -4099
rect 906 -4099 1026 -4052
rect 906 -4117 944 -4099
rect 810 -4133 826 -4117
rect 750 -4149 826 -4133
rect 928 -4133 944 -4117
rect 988 -4117 1026 -4099
rect 1084 -4099 1204 -4052
rect 1084 -4117 1122 -4099
rect 988 -4133 1004 -4117
rect 928 -4149 1004 -4133
rect 1106 -4133 1122 -4117
rect 1166 -4117 1204 -4099
rect 1262 -4099 1382 -4052
rect 1262 -4117 1300 -4099
rect 1166 -4133 1182 -4117
rect 1106 -4149 1182 -4133
rect 1284 -4133 1300 -4117
rect 1344 -4117 1382 -4099
rect 1440 -4099 1560 -4052
rect 1440 -4117 1478 -4099
rect 1344 -4133 1360 -4117
rect 1284 -4149 1360 -4133
rect 1462 -4133 1478 -4117
rect 1522 -4117 1560 -4099
rect 1618 -4099 1738 -4052
rect 1618 -4117 1656 -4099
rect 1522 -4133 1538 -4117
rect 1462 -4149 1538 -4133
rect 1640 -4133 1656 -4117
rect 1700 -4117 1738 -4099
rect 1796 -4099 1916 -4052
rect 1796 -4117 1834 -4099
rect 1700 -4133 1716 -4117
rect 1640 -4149 1716 -4133
rect 1818 -4133 1834 -4117
rect 1878 -4117 1916 -4099
rect 1974 -4099 2094 -4052
rect 1974 -4117 2012 -4099
rect 1878 -4133 1894 -4117
rect 1818 -4149 1894 -4133
rect 1996 -4133 2012 -4117
rect 2056 -4117 2094 -4099
rect 2152 -4099 2272 -4052
rect 2152 -4117 2190 -4099
rect 2056 -4133 2072 -4117
rect 1996 -4149 2072 -4133
rect 2174 -4133 2190 -4117
rect 2234 -4117 2272 -4099
rect 2330 -4099 2450 -4052
rect 2330 -4117 2368 -4099
rect 2234 -4133 2250 -4117
rect 2174 -4149 2250 -4133
rect 2352 -4133 2368 -4117
rect 2412 -4117 2450 -4099
rect 2508 -4099 2628 -4052
rect 2508 -4117 2546 -4099
rect 2412 -4133 2428 -4117
rect 2352 -4149 2428 -4133
rect 2530 -4133 2546 -4117
rect 2590 -4117 2628 -4099
rect 2590 -4133 2606 -4117
rect 2530 -4149 2606 -4133
rect -3586 -4205 -3548 -4187
rect -3682 -4221 -3666 -4205
rect -3742 -4237 -3666 -4221
rect -3564 -4221 -3548 -4205
rect -3504 -4205 -3466 -4187
rect -3504 -4221 -3488 -4205
rect -3564 -4237 -3488 -4221
rect -1386 -4591 -1310 -4575
rect -1386 -4607 -1370 -4591
rect -1408 -4625 -1370 -4607
rect -1326 -4607 -1310 -4591
rect -1208 -4591 -1132 -4575
rect -1208 -4607 -1192 -4591
rect -1326 -4625 -1288 -4607
rect -6234 -4649 -6158 -4633
rect -6234 -4665 -6218 -4649
rect -6256 -4683 -6218 -4665
rect -6174 -4665 -6158 -4649
rect -6056 -4649 -5980 -4633
rect -6056 -4665 -6040 -4649
rect -6174 -4683 -6136 -4665
rect -6256 -4730 -6136 -4683
rect -6078 -4683 -6040 -4665
rect -5996 -4665 -5980 -4649
rect -5878 -4649 -5802 -4633
rect -5878 -4665 -5862 -4649
rect -5996 -4683 -5958 -4665
rect -6078 -4730 -5958 -4683
rect -5900 -4683 -5862 -4665
rect -5818 -4665 -5802 -4649
rect -5700 -4649 -5624 -4633
rect -5700 -4665 -5684 -4649
rect -5818 -4683 -5780 -4665
rect -5900 -4730 -5780 -4683
rect -5722 -4683 -5684 -4665
rect -5640 -4665 -5624 -4649
rect -5522 -4649 -5446 -4633
rect -5522 -4665 -5506 -4649
rect -5640 -4683 -5602 -4665
rect -5722 -4730 -5602 -4683
rect -5544 -4683 -5506 -4665
rect -5462 -4665 -5446 -4649
rect -5344 -4649 -5268 -4633
rect -5344 -4665 -5328 -4649
rect -5462 -4683 -5424 -4665
rect -5544 -4730 -5424 -4683
rect -5366 -4683 -5328 -4665
rect -5284 -4665 -5268 -4649
rect -5166 -4649 -5090 -4633
rect -5166 -4665 -5150 -4649
rect -5284 -4683 -5246 -4665
rect -5366 -4730 -5246 -4683
rect -5188 -4683 -5150 -4665
rect -5106 -4665 -5090 -4649
rect -4988 -4649 -4912 -4633
rect -4988 -4665 -4972 -4649
rect -5106 -4683 -5068 -4665
rect -5188 -4730 -5068 -4683
rect -5010 -4683 -4972 -4665
rect -4928 -4665 -4912 -4649
rect -4810 -4649 -4734 -4633
rect -4810 -4665 -4794 -4649
rect -4928 -4683 -4890 -4665
rect -5010 -4730 -4890 -4683
rect -4832 -4683 -4794 -4665
rect -4750 -4665 -4734 -4649
rect -4632 -4649 -4556 -4633
rect -4632 -4665 -4616 -4649
rect -4750 -4683 -4712 -4665
rect -4832 -4730 -4712 -4683
rect -4654 -4683 -4616 -4665
rect -4572 -4665 -4556 -4649
rect -4454 -4649 -4378 -4633
rect -4454 -4665 -4438 -4649
rect -4572 -4683 -4534 -4665
rect -4654 -4730 -4534 -4683
rect -4476 -4683 -4438 -4665
rect -4394 -4665 -4378 -4649
rect -4276 -4649 -4200 -4633
rect -4276 -4665 -4260 -4649
rect -4394 -4683 -4356 -4665
rect -4476 -4730 -4356 -4683
rect -4298 -4683 -4260 -4665
rect -4216 -4665 -4200 -4649
rect -4098 -4649 -4022 -4633
rect -4098 -4665 -4082 -4649
rect -4216 -4683 -4178 -4665
rect -4298 -4730 -4178 -4683
rect -4120 -4683 -4082 -4665
rect -4038 -4665 -4022 -4649
rect -3920 -4649 -3844 -4633
rect -3920 -4665 -3904 -4649
rect -4038 -4683 -4000 -4665
rect -4120 -4730 -4000 -4683
rect -3942 -4683 -3904 -4665
rect -3860 -4665 -3844 -4649
rect -3742 -4649 -3666 -4633
rect -3742 -4665 -3726 -4649
rect -3860 -4683 -3822 -4665
rect -3942 -4730 -3822 -4683
rect -3764 -4683 -3726 -4665
rect -3682 -4665 -3666 -4649
rect -3564 -4649 -3488 -4633
rect -3564 -4665 -3548 -4649
rect -3682 -4683 -3644 -4665
rect -3764 -4730 -3644 -4683
rect -3586 -4683 -3548 -4665
rect -3504 -4665 -3488 -4649
rect -3504 -4683 -3466 -4665
rect -1408 -4672 -1288 -4625
rect -1230 -4625 -1192 -4607
rect -1148 -4607 -1132 -4591
rect -1030 -4591 -954 -4575
rect -1030 -4607 -1014 -4591
rect -1148 -4625 -1110 -4607
rect -1230 -4672 -1110 -4625
rect -1052 -4625 -1014 -4607
rect -970 -4607 -954 -4591
rect -852 -4591 -776 -4575
rect -852 -4607 -836 -4591
rect -970 -4625 -932 -4607
rect -1052 -4672 -932 -4625
rect -874 -4625 -836 -4607
rect -792 -4607 -776 -4591
rect -674 -4591 -598 -4575
rect -674 -4607 -658 -4591
rect -792 -4625 -754 -4607
rect -874 -4672 -754 -4625
rect -696 -4625 -658 -4607
rect -614 -4607 -598 -4591
rect -496 -4591 -420 -4575
rect -496 -4607 -480 -4591
rect -614 -4625 -576 -4607
rect -696 -4672 -576 -4625
rect -518 -4625 -480 -4607
rect -436 -4607 -420 -4591
rect -318 -4591 -242 -4575
rect -318 -4607 -302 -4591
rect -436 -4625 -398 -4607
rect -518 -4672 -398 -4625
rect -340 -4625 -302 -4607
rect -258 -4607 -242 -4591
rect -140 -4591 -64 -4575
rect -140 -4607 -124 -4591
rect -258 -4625 -220 -4607
rect -340 -4672 -220 -4625
rect -162 -4625 -124 -4607
rect -80 -4607 -64 -4591
rect 38 -4591 114 -4575
rect 38 -4607 54 -4591
rect -80 -4625 -42 -4607
rect -162 -4672 -42 -4625
rect 16 -4625 54 -4607
rect 98 -4607 114 -4591
rect 216 -4591 292 -4575
rect 216 -4607 232 -4591
rect 98 -4625 136 -4607
rect 16 -4672 136 -4625
rect 194 -4625 232 -4607
rect 276 -4607 292 -4591
rect 394 -4591 470 -4575
rect 394 -4607 410 -4591
rect 276 -4625 314 -4607
rect 194 -4672 314 -4625
rect 372 -4625 410 -4607
rect 454 -4607 470 -4591
rect 572 -4591 648 -4575
rect 572 -4607 588 -4591
rect 454 -4625 492 -4607
rect 372 -4672 492 -4625
rect 550 -4625 588 -4607
rect 632 -4607 648 -4591
rect 750 -4591 826 -4575
rect 750 -4607 766 -4591
rect 632 -4625 670 -4607
rect 550 -4672 670 -4625
rect 728 -4625 766 -4607
rect 810 -4607 826 -4591
rect 928 -4591 1004 -4575
rect 928 -4607 944 -4591
rect 810 -4625 848 -4607
rect 728 -4672 848 -4625
rect 906 -4625 944 -4607
rect 988 -4607 1004 -4591
rect 1106 -4591 1182 -4575
rect 1106 -4607 1122 -4591
rect 988 -4625 1026 -4607
rect 906 -4672 1026 -4625
rect 1084 -4625 1122 -4607
rect 1166 -4607 1182 -4591
rect 1284 -4591 1360 -4575
rect 1284 -4607 1300 -4591
rect 1166 -4625 1204 -4607
rect 1084 -4672 1204 -4625
rect 1262 -4625 1300 -4607
rect 1344 -4607 1360 -4591
rect 1462 -4591 1538 -4575
rect 1462 -4607 1478 -4591
rect 1344 -4625 1382 -4607
rect 1262 -4672 1382 -4625
rect 1440 -4625 1478 -4607
rect 1522 -4607 1538 -4591
rect 1640 -4591 1716 -4575
rect 1640 -4607 1656 -4591
rect 1522 -4625 1560 -4607
rect 1440 -4672 1560 -4625
rect 1618 -4625 1656 -4607
rect 1700 -4607 1716 -4591
rect 1818 -4591 1894 -4575
rect 1818 -4607 1834 -4591
rect 1700 -4625 1738 -4607
rect 1618 -4672 1738 -4625
rect 1796 -4625 1834 -4607
rect 1878 -4607 1894 -4591
rect 1996 -4591 2072 -4575
rect 1996 -4607 2012 -4591
rect 1878 -4625 1916 -4607
rect 1796 -4672 1916 -4625
rect 1974 -4625 2012 -4607
rect 2056 -4607 2072 -4591
rect 2174 -4591 2250 -4575
rect 2174 -4607 2190 -4591
rect 2056 -4625 2094 -4607
rect 1974 -4672 2094 -4625
rect 2152 -4625 2190 -4607
rect 2234 -4607 2250 -4591
rect 2352 -4591 2428 -4575
rect 2352 -4607 2368 -4591
rect 2234 -4625 2272 -4607
rect 2152 -4672 2272 -4625
rect 2330 -4625 2368 -4607
rect 2412 -4607 2428 -4591
rect 2530 -4591 2606 -4575
rect 2530 -4607 2546 -4591
rect 2412 -4625 2450 -4607
rect 2330 -4672 2450 -4625
rect 2508 -4625 2546 -4607
rect 2590 -4607 2606 -4591
rect 2590 -4625 2628 -4607
rect 2508 -4672 2628 -4625
rect -3586 -4730 -3466 -4683
rect -1408 -4999 -1288 -4952
rect -6256 -5057 -6136 -5010
rect -6256 -5075 -6218 -5057
rect -6234 -5091 -6218 -5075
rect -6174 -5075 -6136 -5057
rect -6078 -5057 -5958 -5010
rect -6078 -5075 -6040 -5057
rect -6174 -5091 -6158 -5075
rect -6234 -5107 -6158 -5091
rect -6056 -5091 -6040 -5075
rect -5996 -5075 -5958 -5057
rect -5900 -5057 -5780 -5010
rect -5900 -5075 -5862 -5057
rect -5996 -5091 -5980 -5075
rect -6056 -5107 -5980 -5091
rect -5878 -5091 -5862 -5075
rect -5818 -5075 -5780 -5057
rect -5722 -5057 -5602 -5010
rect -5722 -5075 -5684 -5057
rect -5818 -5091 -5802 -5075
rect -5878 -5107 -5802 -5091
rect -5700 -5091 -5684 -5075
rect -5640 -5075 -5602 -5057
rect -5544 -5057 -5424 -5010
rect -5544 -5075 -5506 -5057
rect -5640 -5091 -5624 -5075
rect -5700 -5107 -5624 -5091
rect -5522 -5091 -5506 -5075
rect -5462 -5075 -5424 -5057
rect -5366 -5057 -5246 -5010
rect -5366 -5075 -5328 -5057
rect -5462 -5091 -5446 -5075
rect -5522 -5107 -5446 -5091
rect -5344 -5091 -5328 -5075
rect -5284 -5075 -5246 -5057
rect -5188 -5057 -5068 -5010
rect -5188 -5075 -5150 -5057
rect -5284 -5091 -5268 -5075
rect -5344 -5107 -5268 -5091
rect -5166 -5091 -5150 -5075
rect -5106 -5075 -5068 -5057
rect -5010 -5057 -4890 -5010
rect -5010 -5075 -4972 -5057
rect -5106 -5091 -5090 -5075
rect -5166 -5107 -5090 -5091
rect -4988 -5091 -4972 -5075
rect -4928 -5075 -4890 -5057
rect -4832 -5057 -4712 -5010
rect -4832 -5075 -4794 -5057
rect -4928 -5091 -4912 -5075
rect -4988 -5107 -4912 -5091
rect -4810 -5091 -4794 -5075
rect -4750 -5075 -4712 -5057
rect -4654 -5057 -4534 -5010
rect -4654 -5075 -4616 -5057
rect -4750 -5091 -4734 -5075
rect -4810 -5107 -4734 -5091
rect -4632 -5091 -4616 -5075
rect -4572 -5075 -4534 -5057
rect -4476 -5057 -4356 -5010
rect -4476 -5075 -4438 -5057
rect -4572 -5091 -4556 -5075
rect -4632 -5107 -4556 -5091
rect -4454 -5091 -4438 -5075
rect -4394 -5075 -4356 -5057
rect -4298 -5057 -4178 -5010
rect -4298 -5075 -4260 -5057
rect -4394 -5091 -4378 -5075
rect -4454 -5107 -4378 -5091
rect -4276 -5091 -4260 -5075
rect -4216 -5075 -4178 -5057
rect -4120 -5057 -4000 -5010
rect -4120 -5075 -4082 -5057
rect -4216 -5091 -4200 -5075
rect -4276 -5107 -4200 -5091
rect -4098 -5091 -4082 -5075
rect -4038 -5075 -4000 -5057
rect -3942 -5057 -3822 -5010
rect -3942 -5075 -3904 -5057
rect -4038 -5091 -4022 -5075
rect -4098 -5107 -4022 -5091
rect -3920 -5091 -3904 -5075
rect -3860 -5075 -3822 -5057
rect -3764 -5057 -3644 -5010
rect -3764 -5075 -3726 -5057
rect -3860 -5091 -3844 -5075
rect -3920 -5107 -3844 -5091
rect -3742 -5091 -3726 -5075
rect -3682 -5075 -3644 -5057
rect -3586 -5057 -3466 -5010
rect -1408 -5017 -1370 -4999
rect -1386 -5033 -1370 -5017
rect -1326 -5017 -1288 -4999
rect -1230 -4999 -1110 -4952
rect -1230 -5017 -1192 -4999
rect -1326 -5033 -1310 -5017
rect -1386 -5049 -1310 -5033
rect -1208 -5033 -1192 -5017
rect -1148 -5017 -1110 -4999
rect -1052 -4999 -932 -4952
rect -1052 -5017 -1014 -4999
rect -1148 -5033 -1132 -5017
rect -1208 -5049 -1132 -5033
rect -1030 -5033 -1014 -5017
rect -970 -5017 -932 -4999
rect -874 -4999 -754 -4952
rect -874 -5017 -836 -4999
rect -970 -5033 -954 -5017
rect -1030 -5049 -954 -5033
rect -852 -5033 -836 -5017
rect -792 -5017 -754 -4999
rect -696 -4999 -576 -4952
rect -696 -5017 -658 -4999
rect -792 -5033 -776 -5017
rect -852 -5049 -776 -5033
rect -674 -5033 -658 -5017
rect -614 -5017 -576 -4999
rect -518 -4999 -398 -4952
rect -518 -5017 -480 -4999
rect -614 -5033 -598 -5017
rect -674 -5049 -598 -5033
rect -496 -5033 -480 -5017
rect -436 -5017 -398 -4999
rect -340 -4999 -220 -4952
rect -340 -5017 -302 -4999
rect -436 -5033 -420 -5017
rect -496 -5049 -420 -5033
rect -318 -5033 -302 -5017
rect -258 -5017 -220 -4999
rect -162 -4999 -42 -4952
rect -162 -5017 -124 -4999
rect -258 -5033 -242 -5017
rect -318 -5049 -242 -5033
rect -140 -5033 -124 -5017
rect -80 -5017 -42 -4999
rect 16 -4999 136 -4952
rect 16 -5017 54 -4999
rect -80 -5033 -64 -5017
rect -140 -5049 -64 -5033
rect 38 -5033 54 -5017
rect 98 -5017 136 -4999
rect 194 -4999 314 -4952
rect 194 -5017 232 -4999
rect 98 -5033 114 -5017
rect 38 -5049 114 -5033
rect 216 -5033 232 -5017
rect 276 -5017 314 -4999
rect 372 -4999 492 -4952
rect 372 -5017 410 -4999
rect 276 -5033 292 -5017
rect 216 -5049 292 -5033
rect 394 -5033 410 -5017
rect 454 -5017 492 -4999
rect 550 -4999 670 -4952
rect 550 -5017 588 -4999
rect 454 -5033 470 -5017
rect 394 -5049 470 -5033
rect 572 -5033 588 -5017
rect 632 -5017 670 -4999
rect 728 -4999 848 -4952
rect 728 -5017 766 -4999
rect 632 -5033 648 -5017
rect 572 -5049 648 -5033
rect 750 -5033 766 -5017
rect 810 -5017 848 -4999
rect 906 -4999 1026 -4952
rect 906 -5017 944 -4999
rect 810 -5033 826 -5017
rect 750 -5049 826 -5033
rect 928 -5033 944 -5017
rect 988 -5017 1026 -4999
rect 1084 -4999 1204 -4952
rect 1084 -5017 1122 -4999
rect 988 -5033 1004 -5017
rect 928 -5049 1004 -5033
rect 1106 -5033 1122 -5017
rect 1166 -5017 1204 -4999
rect 1262 -4999 1382 -4952
rect 1262 -5017 1300 -4999
rect 1166 -5033 1182 -5017
rect 1106 -5049 1182 -5033
rect 1284 -5033 1300 -5017
rect 1344 -5017 1382 -4999
rect 1440 -4999 1560 -4952
rect 1440 -5017 1478 -4999
rect 1344 -5033 1360 -5017
rect 1284 -5049 1360 -5033
rect 1462 -5033 1478 -5017
rect 1522 -5017 1560 -4999
rect 1618 -4999 1738 -4952
rect 1618 -5017 1656 -4999
rect 1522 -5033 1538 -5017
rect 1462 -5049 1538 -5033
rect 1640 -5033 1656 -5017
rect 1700 -5017 1738 -4999
rect 1796 -4999 1916 -4952
rect 1796 -5017 1834 -4999
rect 1700 -5033 1716 -5017
rect 1640 -5049 1716 -5033
rect 1818 -5033 1834 -5017
rect 1878 -5017 1916 -4999
rect 1974 -4999 2094 -4952
rect 1974 -5017 2012 -4999
rect 1878 -5033 1894 -5017
rect 1818 -5049 1894 -5033
rect 1996 -5033 2012 -5017
rect 2056 -5017 2094 -4999
rect 2152 -4999 2272 -4952
rect 2152 -5017 2190 -4999
rect 2056 -5033 2072 -5017
rect 1996 -5049 2072 -5033
rect 2174 -5033 2190 -5017
rect 2234 -5017 2272 -4999
rect 2330 -4999 2450 -4952
rect 2330 -5017 2368 -4999
rect 2234 -5033 2250 -5017
rect 2174 -5049 2250 -5033
rect 2352 -5033 2368 -5017
rect 2412 -5017 2450 -4999
rect 2508 -4999 2628 -4952
rect 2508 -5017 2546 -4999
rect 2412 -5033 2428 -5017
rect 2352 -5049 2428 -5033
rect 2530 -5033 2546 -5017
rect 2590 -5017 2628 -4999
rect 2590 -5033 2606 -5017
rect 2530 -5049 2606 -5033
rect -3586 -5075 -3548 -5057
rect -3682 -5091 -3666 -5075
rect -3742 -5107 -3666 -5091
rect -3564 -5091 -3548 -5075
rect -3504 -5075 -3466 -5057
rect -3504 -5091 -3488 -5075
rect -3564 -5107 -3488 -5091
rect -1386 -5491 -1310 -5475
rect -6234 -5519 -6158 -5503
rect -6234 -5535 -6218 -5519
rect -6256 -5553 -6218 -5535
rect -6174 -5535 -6158 -5519
rect -6056 -5519 -5980 -5503
rect -6056 -5535 -6040 -5519
rect -6174 -5553 -6136 -5535
rect -6256 -5600 -6136 -5553
rect -6078 -5553 -6040 -5535
rect -5996 -5535 -5980 -5519
rect -5878 -5519 -5802 -5503
rect -5878 -5535 -5862 -5519
rect -5996 -5553 -5958 -5535
rect -6078 -5600 -5958 -5553
rect -5900 -5553 -5862 -5535
rect -5818 -5535 -5802 -5519
rect -5700 -5519 -5624 -5503
rect -5700 -5535 -5684 -5519
rect -5818 -5553 -5780 -5535
rect -5900 -5600 -5780 -5553
rect -5722 -5553 -5684 -5535
rect -5640 -5535 -5624 -5519
rect -5522 -5519 -5446 -5503
rect -5522 -5535 -5506 -5519
rect -5640 -5553 -5602 -5535
rect -5722 -5600 -5602 -5553
rect -5544 -5553 -5506 -5535
rect -5462 -5535 -5446 -5519
rect -5344 -5519 -5268 -5503
rect -5344 -5535 -5328 -5519
rect -5462 -5553 -5424 -5535
rect -5544 -5600 -5424 -5553
rect -5366 -5553 -5328 -5535
rect -5284 -5535 -5268 -5519
rect -5166 -5519 -5090 -5503
rect -5166 -5535 -5150 -5519
rect -5284 -5553 -5246 -5535
rect -5366 -5600 -5246 -5553
rect -5188 -5553 -5150 -5535
rect -5106 -5535 -5090 -5519
rect -4988 -5519 -4912 -5503
rect -4988 -5535 -4972 -5519
rect -5106 -5553 -5068 -5535
rect -5188 -5600 -5068 -5553
rect -5010 -5553 -4972 -5535
rect -4928 -5535 -4912 -5519
rect -4810 -5519 -4734 -5503
rect -4810 -5535 -4794 -5519
rect -4928 -5553 -4890 -5535
rect -5010 -5600 -4890 -5553
rect -4832 -5553 -4794 -5535
rect -4750 -5535 -4734 -5519
rect -4632 -5519 -4556 -5503
rect -4632 -5535 -4616 -5519
rect -4750 -5553 -4712 -5535
rect -4832 -5600 -4712 -5553
rect -4654 -5553 -4616 -5535
rect -4572 -5535 -4556 -5519
rect -4454 -5519 -4378 -5503
rect -4454 -5535 -4438 -5519
rect -4572 -5553 -4534 -5535
rect -4654 -5600 -4534 -5553
rect -4476 -5553 -4438 -5535
rect -4394 -5535 -4378 -5519
rect -4276 -5519 -4200 -5503
rect -4276 -5535 -4260 -5519
rect -4394 -5553 -4356 -5535
rect -4476 -5600 -4356 -5553
rect -4298 -5553 -4260 -5535
rect -4216 -5535 -4200 -5519
rect -4098 -5519 -4022 -5503
rect -4098 -5535 -4082 -5519
rect -4216 -5553 -4178 -5535
rect -4298 -5600 -4178 -5553
rect -4120 -5553 -4082 -5535
rect -4038 -5535 -4022 -5519
rect -3920 -5519 -3844 -5503
rect -3920 -5535 -3904 -5519
rect -4038 -5553 -4000 -5535
rect -4120 -5600 -4000 -5553
rect -3942 -5553 -3904 -5535
rect -3860 -5535 -3844 -5519
rect -3742 -5519 -3666 -5503
rect -3742 -5535 -3726 -5519
rect -3860 -5553 -3822 -5535
rect -3942 -5600 -3822 -5553
rect -3764 -5553 -3726 -5535
rect -3682 -5535 -3666 -5519
rect -3564 -5519 -3488 -5503
rect -1386 -5507 -1370 -5491
rect -3564 -5535 -3548 -5519
rect -3682 -5553 -3644 -5535
rect -3764 -5600 -3644 -5553
rect -3586 -5553 -3548 -5535
rect -3504 -5535 -3488 -5519
rect -1408 -5525 -1370 -5507
rect -1326 -5507 -1310 -5491
rect -1208 -5491 -1132 -5475
rect -1208 -5507 -1192 -5491
rect -1326 -5525 -1288 -5507
rect -3504 -5553 -3466 -5535
rect -3586 -5600 -3466 -5553
rect -1408 -5572 -1288 -5525
rect -1230 -5525 -1192 -5507
rect -1148 -5507 -1132 -5491
rect -1030 -5491 -954 -5475
rect -1030 -5507 -1014 -5491
rect -1148 -5525 -1110 -5507
rect -1230 -5572 -1110 -5525
rect -1052 -5525 -1014 -5507
rect -970 -5507 -954 -5491
rect -852 -5491 -776 -5475
rect -852 -5507 -836 -5491
rect -970 -5525 -932 -5507
rect -1052 -5572 -932 -5525
rect -874 -5525 -836 -5507
rect -792 -5507 -776 -5491
rect -674 -5491 -598 -5475
rect -674 -5507 -658 -5491
rect -792 -5525 -754 -5507
rect -874 -5572 -754 -5525
rect -696 -5525 -658 -5507
rect -614 -5507 -598 -5491
rect -496 -5491 -420 -5475
rect -496 -5507 -480 -5491
rect -614 -5525 -576 -5507
rect -696 -5572 -576 -5525
rect -518 -5525 -480 -5507
rect -436 -5507 -420 -5491
rect -318 -5491 -242 -5475
rect -318 -5507 -302 -5491
rect -436 -5525 -398 -5507
rect -518 -5572 -398 -5525
rect -340 -5525 -302 -5507
rect -258 -5507 -242 -5491
rect -140 -5491 -64 -5475
rect -140 -5507 -124 -5491
rect -258 -5525 -220 -5507
rect -340 -5572 -220 -5525
rect -162 -5525 -124 -5507
rect -80 -5507 -64 -5491
rect 38 -5491 114 -5475
rect 38 -5507 54 -5491
rect -80 -5525 -42 -5507
rect -162 -5572 -42 -5525
rect 16 -5525 54 -5507
rect 98 -5507 114 -5491
rect 216 -5491 292 -5475
rect 216 -5507 232 -5491
rect 98 -5525 136 -5507
rect 16 -5572 136 -5525
rect 194 -5525 232 -5507
rect 276 -5507 292 -5491
rect 394 -5491 470 -5475
rect 394 -5507 410 -5491
rect 276 -5525 314 -5507
rect 194 -5572 314 -5525
rect 372 -5525 410 -5507
rect 454 -5507 470 -5491
rect 572 -5491 648 -5475
rect 572 -5507 588 -5491
rect 454 -5525 492 -5507
rect 372 -5572 492 -5525
rect 550 -5525 588 -5507
rect 632 -5507 648 -5491
rect 750 -5491 826 -5475
rect 750 -5507 766 -5491
rect 632 -5525 670 -5507
rect 550 -5572 670 -5525
rect 728 -5525 766 -5507
rect 810 -5507 826 -5491
rect 928 -5491 1004 -5475
rect 928 -5507 944 -5491
rect 810 -5525 848 -5507
rect 728 -5572 848 -5525
rect 906 -5525 944 -5507
rect 988 -5507 1004 -5491
rect 1106 -5491 1182 -5475
rect 1106 -5507 1122 -5491
rect 988 -5525 1026 -5507
rect 906 -5572 1026 -5525
rect 1084 -5525 1122 -5507
rect 1166 -5507 1182 -5491
rect 1284 -5491 1360 -5475
rect 1284 -5507 1300 -5491
rect 1166 -5525 1204 -5507
rect 1084 -5572 1204 -5525
rect 1262 -5525 1300 -5507
rect 1344 -5507 1360 -5491
rect 1462 -5491 1538 -5475
rect 1462 -5507 1478 -5491
rect 1344 -5525 1382 -5507
rect 1262 -5572 1382 -5525
rect 1440 -5525 1478 -5507
rect 1522 -5507 1538 -5491
rect 1640 -5491 1716 -5475
rect 1640 -5507 1656 -5491
rect 1522 -5525 1560 -5507
rect 1440 -5572 1560 -5525
rect 1618 -5525 1656 -5507
rect 1700 -5507 1716 -5491
rect 1818 -5491 1894 -5475
rect 1818 -5507 1834 -5491
rect 1700 -5525 1738 -5507
rect 1618 -5572 1738 -5525
rect 1796 -5525 1834 -5507
rect 1878 -5507 1894 -5491
rect 1996 -5491 2072 -5475
rect 1996 -5507 2012 -5491
rect 1878 -5525 1916 -5507
rect 1796 -5572 1916 -5525
rect 1974 -5525 2012 -5507
rect 2056 -5507 2072 -5491
rect 2174 -5491 2250 -5475
rect 2174 -5507 2190 -5491
rect 2056 -5525 2094 -5507
rect 1974 -5572 2094 -5525
rect 2152 -5525 2190 -5507
rect 2234 -5507 2250 -5491
rect 2352 -5491 2428 -5475
rect 2352 -5507 2368 -5491
rect 2234 -5525 2272 -5507
rect 2152 -5572 2272 -5525
rect 2330 -5525 2368 -5507
rect 2412 -5507 2428 -5491
rect 2530 -5491 2606 -5475
rect 2530 -5507 2546 -5491
rect 2412 -5525 2450 -5507
rect 2330 -5572 2450 -5525
rect 2508 -5525 2546 -5507
rect 2590 -5507 2606 -5491
rect 2590 -5525 2628 -5507
rect 2508 -5572 2628 -5525
rect -6256 -5927 -6136 -5880
rect -6256 -5945 -6218 -5927
rect -6234 -5961 -6218 -5945
rect -6174 -5945 -6136 -5927
rect -6078 -5927 -5958 -5880
rect -6078 -5945 -6040 -5927
rect -6174 -5961 -6158 -5945
rect -6234 -5977 -6158 -5961
rect -6056 -5961 -6040 -5945
rect -5996 -5945 -5958 -5927
rect -5900 -5927 -5780 -5880
rect -5900 -5945 -5862 -5927
rect -5996 -5961 -5980 -5945
rect -6056 -5977 -5980 -5961
rect -5878 -5961 -5862 -5945
rect -5818 -5945 -5780 -5927
rect -5722 -5927 -5602 -5880
rect -5722 -5945 -5684 -5927
rect -5818 -5961 -5802 -5945
rect -5878 -5977 -5802 -5961
rect -5700 -5961 -5684 -5945
rect -5640 -5945 -5602 -5927
rect -5544 -5927 -5424 -5880
rect -5544 -5945 -5506 -5927
rect -5640 -5961 -5624 -5945
rect -5700 -5977 -5624 -5961
rect -5522 -5961 -5506 -5945
rect -5462 -5945 -5424 -5927
rect -5366 -5927 -5246 -5880
rect -5366 -5945 -5328 -5927
rect -5462 -5961 -5446 -5945
rect -5522 -5977 -5446 -5961
rect -5344 -5961 -5328 -5945
rect -5284 -5945 -5246 -5927
rect -5188 -5927 -5068 -5880
rect -5188 -5945 -5150 -5927
rect -5284 -5961 -5268 -5945
rect -5344 -5977 -5268 -5961
rect -5166 -5961 -5150 -5945
rect -5106 -5945 -5068 -5927
rect -5010 -5927 -4890 -5880
rect -5010 -5945 -4972 -5927
rect -5106 -5961 -5090 -5945
rect -5166 -5977 -5090 -5961
rect -4988 -5961 -4972 -5945
rect -4928 -5945 -4890 -5927
rect -4832 -5927 -4712 -5880
rect -4832 -5945 -4794 -5927
rect -4928 -5961 -4912 -5945
rect -4988 -5977 -4912 -5961
rect -4810 -5961 -4794 -5945
rect -4750 -5945 -4712 -5927
rect -4654 -5927 -4534 -5880
rect -4654 -5945 -4616 -5927
rect -4750 -5961 -4734 -5945
rect -4810 -5977 -4734 -5961
rect -4632 -5961 -4616 -5945
rect -4572 -5945 -4534 -5927
rect -4476 -5927 -4356 -5880
rect -4476 -5945 -4438 -5927
rect -4572 -5961 -4556 -5945
rect -4632 -5977 -4556 -5961
rect -4454 -5961 -4438 -5945
rect -4394 -5945 -4356 -5927
rect -4298 -5927 -4178 -5880
rect -4298 -5945 -4260 -5927
rect -4394 -5961 -4378 -5945
rect -4454 -5977 -4378 -5961
rect -4276 -5961 -4260 -5945
rect -4216 -5945 -4178 -5927
rect -4120 -5927 -4000 -5880
rect -4120 -5945 -4082 -5927
rect -4216 -5961 -4200 -5945
rect -4276 -5977 -4200 -5961
rect -4098 -5961 -4082 -5945
rect -4038 -5945 -4000 -5927
rect -3942 -5927 -3822 -5880
rect -3942 -5945 -3904 -5927
rect -4038 -5961 -4022 -5945
rect -4098 -5977 -4022 -5961
rect -3920 -5961 -3904 -5945
rect -3860 -5945 -3822 -5927
rect -3764 -5927 -3644 -5880
rect -3764 -5945 -3726 -5927
rect -3860 -5961 -3844 -5945
rect -3920 -5977 -3844 -5961
rect -3742 -5961 -3726 -5945
rect -3682 -5945 -3644 -5927
rect -3586 -5927 -3466 -5880
rect -1408 -5899 -1288 -5852
rect -1408 -5917 -1370 -5899
rect -3586 -5945 -3548 -5927
rect -3682 -5961 -3666 -5945
rect -3742 -5977 -3666 -5961
rect -3564 -5961 -3548 -5945
rect -3504 -5945 -3466 -5927
rect -1386 -5933 -1370 -5917
rect -1326 -5917 -1288 -5899
rect -1230 -5899 -1110 -5852
rect -1230 -5917 -1192 -5899
rect -1326 -5933 -1310 -5917
rect -3504 -5961 -3488 -5945
rect -1386 -5949 -1310 -5933
rect -1208 -5933 -1192 -5917
rect -1148 -5917 -1110 -5899
rect -1052 -5899 -932 -5852
rect -1052 -5917 -1014 -5899
rect -1148 -5933 -1132 -5917
rect -1208 -5949 -1132 -5933
rect -1030 -5933 -1014 -5917
rect -970 -5917 -932 -5899
rect -874 -5899 -754 -5852
rect -874 -5917 -836 -5899
rect -970 -5933 -954 -5917
rect -1030 -5949 -954 -5933
rect -852 -5933 -836 -5917
rect -792 -5917 -754 -5899
rect -696 -5899 -576 -5852
rect -696 -5917 -658 -5899
rect -792 -5933 -776 -5917
rect -852 -5949 -776 -5933
rect -674 -5933 -658 -5917
rect -614 -5917 -576 -5899
rect -518 -5899 -398 -5852
rect -518 -5917 -480 -5899
rect -614 -5933 -598 -5917
rect -674 -5949 -598 -5933
rect -496 -5933 -480 -5917
rect -436 -5917 -398 -5899
rect -340 -5899 -220 -5852
rect -340 -5917 -302 -5899
rect -436 -5933 -420 -5917
rect -496 -5949 -420 -5933
rect -318 -5933 -302 -5917
rect -258 -5917 -220 -5899
rect -162 -5899 -42 -5852
rect -162 -5917 -124 -5899
rect -258 -5933 -242 -5917
rect -318 -5949 -242 -5933
rect -140 -5933 -124 -5917
rect -80 -5917 -42 -5899
rect 16 -5899 136 -5852
rect 16 -5917 54 -5899
rect -80 -5933 -64 -5917
rect -140 -5949 -64 -5933
rect 38 -5933 54 -5917
rect 98 -5917 136 -5899
rect 194 -5899 314 -5852
rect 194 -5917 232 -5899
rect 98 -5933 114 -5917
rect 38 -5949 114 -5933
rect 216 -5933 232 -5917
rect 276 -5917 314 -5899
rect 372 -5899 492 -5852
rect 372 -5917 410 -5899
rect 276 -5933 292 -5917
rect 216 -5949 292 -5933
rect 394 -5933 410 -5917
rect 454 -5917 492 -5899
rect 550 -5899 670 -5852
rect 550 -5917 588 -5899
rect 454 -5933 470 -5917
rect 394 -5949 470 -5933
rect 572 -5933 588 -5917
rect 632 -5917 670 -5899
rect 728 -5899 848 -5852
rect 728 -5917 766 -5899
rect 632 -5933 648 -5917
rect 572 -5949 648 -5933
rect 750 -5933 766 -5917
rect 810 -5917 848 -5899
rect 906 -5899 1026 -5852
rect 906 -5917 944 -5899
rect 810 -5933 826 -5917
rect 750 -5949 826 -5933
rect 928 -5933 944 -5917
rect 988 -5917 1026 -5899
rect 1084 -5899 1204 -5852
rect 1084 -5917 1122 -5899
rect 988 -5933 1004 -5917
rect 928 -5949 1004 -5933
rect 1106 -5933 1122 -5917
rect 1166 -5917 1204 -5899
rect 1262 -5899 1382 -5852
rect 1262 -5917 1300 -5899
rect 1166 -5933 1182 -5917
rect 1106 -5949 1182 -5933
rect 1284 -5933 1300 -5917
rect 1344 -5917 1382 -5899
rect 1440 -5899 1560 -5852
rect 1440 -5917 1478 -5899
rect 1344 -5933 1360 -5917
rect 1284 -5949 1360 -5933
rect 1462 -5933 1478 -5917
rect 1522 -5917 1560 -5899
rect 1618 -5899 1738 -5852
rect 1618 -5917 1656 -5899
rect 1522 -5933 1538 -5917
rect 1462 -5949 1538 -5933
rect 1640 -5933 1656 -5917
rect 1700 -5917 1738 -5899
rect 1796 -5899 1916 -5852
rect 1796 -5917 1834 -5899
rect 1700 -5933 1716 -5917
rect 1640 -5949 1716 -5933
rect 1818 -5933 1834 -5917
rect 1878 -5917 1916 -5899
rect 1974 -5899 2094 -5852
rect 1974 -5917 2012 -5899
rect 1878 -5933 1894 -5917
rect 1818 -5949 1894 -5933
rect 1996 -5933 2012 -5917
rect 2056 -5917 2094 -5899
rect 2152 -5899 2272 -5852
rect 2152 -5917 2190 -5899
rect 2056 -5933 2072 -5917
rect 1996 -5949 2072 -5933
rect 2174 -5933 2190 -5917
rect 2234 -5917 2272 -5899
rect 2330 -5899 2450 -5852
rect 2330 -5917 2368 -5899
rect 2234 -5933 2250 -5917
rect 2174 -5949 2250 -5933
rect 2352 -5933 2368 -5917
rect 2412 -5917 2450 -5899
rect 2508 -5899 2628 -5852
rect 2508 -5917 2546 -5899
rect 2412 -5933 2428 -5917
rect 2352 -5949 2428 -5933
rect 2530 -5933 2546 -5917
rect 2590 -5917 2628 -5899
rect 2590 -5933 2606 -5917
rect 2530 -5949 2606 -5933
rect -3564 -5977 -3488 -5961
rect 7204 -1555 7234 -1529
rect 7300 -1555 7330 -1529
rect 7396 -1555 7426 -1529
rect 7492 -1555 7522 -1529
rect 7588 -1555 7618 -1529
rect 7684 -1555 7714 -1529
rect 7780 -1555 7810 -1529
rect 7876 -1555 7906 -1529
rect 7972 -1555 8002 -1529
rect 8068 -1555 8098 -1529
rect 7204 -1681 7234 -1659
rect 7300 -1681 7330 -1659
rect 7396 -1681 7426 -1659
rect 7492 -1681 7522 -1659
rect 7588 -1681 7618 -1659
rect 7684 -1681 7714 -1659
rect 7780 -1681 7810 -1659
rect 7876 -1681 7906 -1659
rect 7972 -1681 8002 -1659
rect 8068 -1681 8098 -1659
rect 7138 -1701 8164 -1681
rect 7138 -1735 7154 -1701
rect 7188 -1735 7346 -1701
rect 7380 -1735 7538 -1701
rect 7572 -1735 7730 -1701
rect 7764 -1735 7922 -1701
rect 7956 -1735 8114 -1701
rect 8148 -1735 8164 -1701
rect 7138 -1747 8164 -1735
rect 16204 -1555 16234 -1529
rect 16300 -1555 16330 -1529
rect 16396 -1555 16426 -1529
rect 16492 -1555 16522 -1529
rect 16588 -1555 16618 -1529
rect 16684 -1555 16714 -1529
rect 16780 -1555 16810 -1529
rect 16876 -1555 16906 -1529
rect 16972 -1555 17002 -1529
rect 17068 -1555 17098 -1529
rect 16204 -1681 16234 -1659
rect 16300 -1681 16330 -1659
rect 16396 -1681 16426 -1659
rect 16492 -1681 16522 -1659
rect 16588 -1681 16618 -1659
rect 16684 -1681 16714 -1659
rect 16780 -1681 16810 -1659
rect 16876 -1681 16906 -1659
rect 16972 -1681 17002 -1659
rect 17068 -1681 17098 -1659
rect 16138 -1701 17164 -1681
rect 16138 -1735 16154 -1701
rect 16188 -1735 16346 -1701
rect 16380 -1735 16538 -1701
rect 16572 -1735 16730 -1701
rect 16764 -1735 16922 -1701
rect 16956 -1735 17114 -1701
rect 17148 -1735 17164 -1701
rect 16138 -1747 17164 -1735
rect 7138 -2693 8164 -2677
rect 7138 -2727 7154 -2693
rect 7188 -2727 7346 -2693
rect 7380 -2727 7538 -2693
rect 7572 -2727 7730 -2693
rect 7764 -2727 7922 -2693
rect 7956 -2727 8114 -2693
rect 8148 -2727 8164 -2693
rect 7138 -2743 8164 -2727
rect 7204 -2775 7234 -2743
rect 7300 -2775 7330 -2743
rect 7396 -2775 7426 -2743
rect 7492 -2775 7522 -2743
rect 7588 -2775 7618 -2743
rect 7684 -2775 7714 -2743
rect 7780 -2775 7810 -2743
rect 7876 -2775 7906 -2743
rect 7972 -2775 8002 -2743
rect 8068 -2775 8098 -2743
rect 7204 -3073 7234 -3047
rect 7300 -3073 7330 -3047
rect 7396 -3073 7426 -3047
rect 7492 -3073 7522 -3047
rect 7588 -3073 7618 -3047
rect 7684 -3073 7714 -3047
rect 7780 -3073 7810 -3047
rect 7876 -3073 7906 -3047
rect 7972 -3073 8002 -3047
rect 8068 -3073 8098 -3047
rect 16138 -2693 17164 -2677
rect 16138 -2727 16154 -2693
rect 16188 -2727 16346 -2693
rect 16380 -2727 16538 -2693
rect 16572 -2727 16730 -2693
rect 16764 -2727 16922 -2693
rect 16956 -2727 17114 -2693
rect 17148 -2727 17164 -2693
rect 16138 -2743 17164 -2727
rect 16204 -2775 16234 -2743
rect 16300 -2775 16330 -2743
rect 16396 -2775 16426 -2743
rect 16492 -2775 16522 -2743
rect 16588 -2775 16618 -2743
rect 16684 -2775 16714 -2743
rect 16780 -2775 16810 -2743
rect 16876 -2775 16906 -2743
rect 16972 -2775 17002 -2743
rect 17068 -2775 17098 -2743
rect 16204 -3073 16234 -3047
rect 16300 -3073 16330 -3047
rect 16396 -3073 16426 -3047
rect 16492 -3073 16522 -3047
rect 16588 -3073 16618 -3047
rect 16684 -3073 16714 -3047
rect 16780 -3073 16810 -3047
rect 16876 -3073 16906 -3047
rect 16972 -3073 17002 -3047
rect 17068 -3073 17098 -3047
rect 7204 -3355 7234 -3329
rect 7300 -3355 7330 -3329
rect 7396 -3355 7426 -3329
rect 7492 -3355 7522 -3329
rect 7588 -3355 7618 -3329
rect 7684 -3355 7714 -3329
rect 7780 -3355 7810 -3329
rect 7876 -3355 7906 -3329
rect 7972 -3355 8002 -3329
rect 8068 -3355 8098 -3329
rect 7204 -3481 7234 -3459
rect 7300 -3481 7330 -3459
rect 7396 -3481 7426 -3459
rect 7492 -3481 7522 -3459
rect 7588 -3481 7618 -3459
rect 7684 -3481 7714 -3459
rect 7780 -3481 7810 -3459
rect 7876 -3481 7906 -3459
rect 7972 -3481 8002 -3459
rect 8068 -3481 8098 -3459
rect 7138 -3501 8164 -3481
rect 7138 -3535 7154 -3501
rect 7188 -3535 7346 -3501
rect 7380 -3535 7538 -3501
rect 7572 -3535 7730 -3501
rect 7764 -3535 7922 -3501
rect 7956 -3535 8114 -3501
rect 8148 -3535 8164 -3501
rect 7138 -3547 8164 -3535
rect 16204 -3355 16234 -3329
rect 16300 -3355 16330 -3329
rect 16396 -3355 16426 -3329
rect 16492 -3355 16522 -3329
rect 16588 -3355 16618 -3329
rect 16684 -3355 16714 -3329
rect 16780 -3355 16810 -3329
rect 16876 -3355 16906 -3329
rect 16972 -3355 17002 -3329
rect 17068 -3355 17098 -3329
rect 16204 -3481 16234 -3459
rect 16300 -3481 16330 -3459
rect 16396 -3481 16426 -3459
rect 16492 -3481 16522 -3459
rect 16588 -3481 16618 -3459
rect 16684 -3481 16714 -3459
rect 16780 -3481 16810 -3459
rect 16876 -3481 16906 -3459
rect 16972 -3481 17002 -3459
rect 17068 -3481 17098 -3459
rect 16138 -3501 17164 -3481
rect 16138 -3535 16154 -3501
rect 16188 -3535 16346 -3501
rect 16380 -3535 16538 -3501
rect 16572 -3535 16730 -3501
rect 16764 -3535 16922 -3501
rect 16956 -3535 17114 -3501
rect 17148 -3535 17164 -3501
rect 16138 -3547 17164 -3535
rect 7138 -4493 8164 -4477
rect 7138 -4527 7154 -4493
rect 7188 -4527 7346 -4493
rect 7380 -4527 7538 -4493
rect 7572 -4527 7730 -4493
rect 7764 -4527 7922 -4493
rect 7956 -4527 8114 -4493
rect 8148 -4527 8164 -4493
rect 7138 -4543 8164 -4527
rect 7204 -4575 7234 -4543
rect 7300 -4575 7330 -4543
rect 7396 -4575 7426 -4543
rect 7492 -4575 7522 -4543
rect 7588 -4575 7618 -4543
rect 7684 -4575 7714 -4543
rect 7780 -4575 7810 -4543
rect 7876 -4575 7906 -4543
rect 7972 -4575 8002 -4543
rect 8068 -4575 8098 -4543
rect 7204 -4873 7234 -4847
rect 7300 -4873 7330 -4847
rect 7396 -4873 7426 -4847
rect 7492 -4873 7522 -4847
rect 7588 -4873 7618 -4847
rect 7684 -4873 7714 -4847
rect 7780 -4873 7810 -4847
rect 7876 -4873 7906 -4847
rect 7972 -4873 8002 -4847
rect 8068 -4873 8098 -4847
rect 16138 -4493 17164 -4477
rect 16138 -4527 16154 -4493
rect 16188 -4527 16346 -4493
rect 16380 -4527 16538 -4493
rect 16572 -4527 16730 -4493
rect 16764 -4527 16922 -4493
rect 16956 -4527 17114 -4493
rect 17148 -4527 17164 -4493
rect 16138 -4543 17164 -4527
rect 16204 -4575 16234 -4543
rect 16300 -4575 16330 -4543
rect 16396 -4575 16426 -4543
rect 16492 -4575 16522 -4543
rect 16588 -4575 16618 -4543
rect 16684 -4575 16714 -4543
rect 16780 -4575 16810 -4543
rect 16876 -4575 16906 -4543
rect 16972 -4575 17002 -4543
rect 17068 -4575 17098 -4543
rect 16204 -4873 16234 -4847
rect 16300 -4873 16330 -4847
rect 16396 -4873 16426 -4847
rect 16492 -4873 16522 -4847
rect 16588 -4873 16618 -4847
rect 16684 -4873 16714 -4847
rect 16780 -4873 16810 -4847
rect 16876 -4873 16906 -4847
rect 16972 -4873 17002 -4847
rect 17068 -4873 17098 -4847
rect 7204 -5155 7234 -5129
rect 7300 -5155 7330 -5129
rect 7396 -5155 7426 -5129
rect 7492 -5155 7522 -5129
rect 7588 -5155 7618 -5129
rect 7684 -5155 7714 -5129
rect 7780 -5155 7810 -5129
rect 7876 -5155 7906 -5129
rect 7972 -5155 8002 -5129
rect 8068 -5155 8098 -5129
rect 7204 -5281 7234 -5259
rect 7300 -5281 7330 -5259
rect 7396 -5281 7426 -5259
rect 7492 -5281 7522 -5259
rect 7588 -5281 7618 -5259
rect 7684 -5281 7714 -5259
rect 7780 -5281 7810 -5259
rect 7876 -5281 7906 -5259
rect 7972 -5281 8002 -5259
rect 8068 -5281 8098 -5259
rect 7138 -5301 8164 -5281
rect 7138 -5335 7154 -5301
rect 7188 -5335 7346 -5301
rect 7380 -5335 7538 -5301
rect 7572 -5335 7730 -5301
rect 7764 -5335 7922 -5301
rect 7956 -5335 8114 -5301
rect 8148 -5335 8164 -5301
rect 7138 -5347 8164 -5335
rect 16204 -5155 16234 -5129
rect 16300 -5155 16330 -5129
rect 16396 -5155 16426 -5129
rect 16492 -5155 16522 -5129
rect 16588 -5155 16618 -5129
rect 16684 -5155 16714 -5129
rect 16780 -5155 16810 -5129
rect 16876 -5155 16906 -5129
rect 16972 -5155 17002 -5129
rect 17068 -5155 17098 -5129
rect 16204 -5281 16234 -5259
rect 16300 -5281 16330 -5259
rect 16396 -5281 16426 -5259
rect 16492 -5281 16522 -5259
rect 16588 -5281 16618 -5259
rect 16684 -5281 16714 -5259
rect 16780 -5281 16810 -5259
rect 16876 -5281 16906 -5259
rect 16972 -5281 17002 -5259
rect 17068 -5281 17098 -5259
rect 16138 -5301 17164 -5281
rect 16138 -5335 16154 -5301
rect 16188 -5335 16346 -5301
rect 16380 -5335 16538 -5301
rect 16572 -5335 16730 -5301
rect 16764 -5335 16922 -5301
rect 16956 -5335 17114 -5301
rect 17148 -5335 17164 -5301
rect 16138 -5347 17164 -5335
rect 7138 -6293 8164 -6277
rect 7138 -6327 7154 -6293
rect 7188 -6327 7346 -6293
rect 7380 -6327 7538 -6293
rect 7572 -6327 7730 -6293
rect 7764 -6327 7922 -6293
rect 7956 -6327 8114 -6293
rect 8148 -6327 8164 -6293
rect 7138 -6343 8164 -6327
rect 7204 -6375 7234 -6343
rect 7300 -6375 7330 -6343
rect 7396 -6375 7426 -6343
rect 7492 -6375 7522 -6343
rect 7588 -6375 7618 -6343
rect 7684 -6375 7714 -6343
rect 7780 -6375 7810 -6343
rect 7876 -6375 7906 -6343
rect 7972 -6375 8002 -6343
rect 8068 -6375 8098 -6343
rect 7204 -6673 7234 -6647
rect 7300 -6673 7330 -6647
rect 7396 -6673 7426 -6647
rect 7492 -6673 7522 -6647
rect 7588 -6673 7618 -6647
rect 7684 -6673 7714 -6647
rect 7780 -6673 7810 -6647
rect 7876 -6673 7906 -6647
rect 7972 -6673 8002 -6647
rect 8068 -6673 8098 -6647
rect 16138 -6293 17164 -6277
rect 16138 -6327 16154 -6293
rect 16188 -6327 16346 -6293
rect 16380 -6327 16538 -6293
rect 16572 -6327 16730 -6293
rect 16764 -6327 16922 -6293
rect 16956 -6327 17114 -6293
rect 17148 -6327 17164 -6293
rect 16138 -6343 17164 -6327
rect 16204 -6375 16234 -6343
rect 16300 -6375 16330 -6343
rect 16396 -6375 16426 -6343
rect 16492 -6375 16522 -6343
rect 16588 -6375 16618 -6343
rect 16684 -6375 16714 -6343
rect 16780 -6375 16810 -6343
rect 16876 -6375 16906 -6343
rect 16972 -6375 17002 -6343
rect 17068 -6375 17098 -6343
rect 16204 -6673 16234 -6647
rect 16300 -6673 16330 -6647
rect 16396 -6673 16426 -6647
rect 16492 -6673 16522 -6647
rect 16588 -6673 16618 -6647
rect 16684 -6673 16714 -6647
rect 16780 -6673 16810 -6647
rect 16876 -6673 16906 -6647
rect 16972 -6673 17002 -6647
rect 17068 -6673 17098 -6647
rect 7204 -6955 7234 -6929
rect 7300 -6955 7330 -6929
rect 7396 -6955 7426 -6929
rect 7492 -6955 7522 -6929
rect 7588 -6955 7618 -6929
rect 7684 -6955 7714 -6929
rect 7780 -6955 7810 -6929
rect 7876 -6955 7906 -6929
rect 7972 -6955 8002 -6929
rect 8068 -6955 8098 -6929
rect 7204 -7081 7234 -7059
rect 7300 -7081 7330 -7059
rect 7396 -7081 7426 -7059
rect 7492 -7081 7522 -7059
rect 7588 -7081 7618 -7059
rect 7684 -7081 7714 -7059
rect 7780 -7081 7810 -7059
rect 7876 -7081 7906 -7059
rect 7972 -7081 8002 -7059
rect 8068 -7081 8098 -7059
rect 7138 -7101 8164 -7081
rect 7138 -7135 7154 -7101
rect 7188 -7135 7346 -7101
rect 7380 -7135 7538 -7101
rect 7572 -7135 7730 -7101
rect 7764 -7135 7922 -7101
rect 7956 -7135 8114 -7101
rect 8148 -7135 8164 -7101
rect 7138 -7147 8164 -7135
rect 16204 -6955 16234 -6929
rect 16300 -6955 16330 -6929
rect 16396 -6955 16426 -6929
rect 16492 -6955 16522 -6929
rect 16588 -6955 16618 -6929
rect 16684 -6955 16714 -6929
rect 16780 -6955 16810 -6929
rect 16876 -6955 16906 -6929
rect 16972 -6955 17002 -6929
rect 17068 -6955 17098 -6929
rect 16204 -7081 16234 -7059
rect 16300 -7081 16330 -7059
rect 16396 -7081 16426 -7059
rect 16492 -7081 16522 -7059
rect 16588 -7081 16618 -7059
rect 16684 -7081 16714 -7059
rect 16780 -7081 16810 -7059
rect 16876 -7081 16906 -7059
rect 16972 -7081 17002 -7059
rect 17068 -7081 17098 -7059
rect 16138 -7101 17164 -7081
rect 16138 -7135 16154 -7101
rect 16188 -7135 16346 -7101
rect 16380 -7135 16538 -7101
rect 16572 -7135 16730 -7101
rect 16764 -7135 16922 -7101
rect 16956 -7135 17114 -7101
rect 17148 -7135 17164 -7101
rect 16138 -7147 17164 -7135
rect -5560 -7790 -5484 -7774
rect -5560 -7808 -5544 -7790
rect -5582 -7824 -5544 -7808
rect -5500 -7808 -5484 -7790
rect -5382 -7790 -5306 -7774
rect -5382 -7808 -5366 -7790
rect -5500 -7824 -5462 -7808
rect -5582 -7862 -5462 -7824
rect -5404 -7824 -5366 -7808
rect -5322 -7808 -5306 -7790
rect -5204 -7790 -5128 -7774
rect -5204 -7808 -5188 -7790
rect -5322 -7824 -5284 -7808
rect -5404 -7862 -5284 -7824
rect -5226 -7824 -5188 -7808
rect -5144 -7808 -5128 -7790
rect -5026 -7790 -4950 -7774
rect -5026 -7808 -5010 -7790
rect -5144 -7824 -5106 -7808
rect -5226 -7862 -5106 -7824
rect -5048 -7824 -5010 -7808
rect -4966 -7808 -4950 -7790
rect -4848 -7790 -4772 -7774
rect -4848 -7808 -4832 -7790
rect -4966 -7824 -4928 -7808
rect -5048 -7862 -4928 -7824
rect -4870 -7824 -4832 -7808
rect -4788 -7808 -4772 -7790
rect -4670 -7790 -4594 -7774
rect -4670 -7808 -4654 -7790
rect -4788 -7824 -4750 -7808
rect -4870 -7862 -4750 -7824
rect -4692 -7824 -4654 -7808
rect -4610 -7808 -4594 -7790
rect -4492 -7790 -4416 -7774
rect -4492 -7808 -4476 -7790
rect -4610 -7824 -4572 -7808
rect -4692 -7862 -4572 -7824
rect -4514 -7824 -4476 -7808
rect -4432 -7808 -4416 -7790
rect -4314 -7790 -4238 -7774
rect -4314 -7808 -4298 -7790
rect -4432 -7824 -4394 -7808
rect -4514 -7862 -4394 -7824
rect -4336 -7824 -4298 -7808
rect -4254 -7808 -4238 -7790
rect -4136 -7790 -4060 -7774
rect -4136 -7808 -4120 -7790
rect -4254 -7824 -4216 -7808
rect -4336 -7862 -4216 -7824
rect -4158 -7824 -4120 -7808
rect -4076 -7808 -4060 -7790
rect -4076 -7824 -4038 -7808
rect -4158 -7862 -4038 -7824
rect -2105 -8048 -2029 -8032
rect -2105 -8066 -2089 -8048
rect -2127 -8082 -2089 -8066
rect -2045 -8066 -2029 -8048
rect -1927 -8048 -1851 -8032
rect -1927 -8066 -1911 -8048
rect -2045 -8082 -2007 -8066
rect -2127 -8120 -2007 -8082
rect -1949 -8082 -1911 -8066
rect -1867 -8066 -1851 -8048
rect -1749 -8048 -1673 -8032
rect -1749 -8066 -1733 -8048
rect -1867 -8082 -1829 -8066
rect -1949 -8120 -1829 -8082
rect -1771 -8082 -1733 -8066
rect -1689 -8066 -1673 -8048
rect -1571 -8048 -1495 -8032
rect -1571 -8066 -1555 -8048
rect -1689 -8082 -1651 -8066
rect -1771 -8120 -1651 -8082
rect -1593 -8082 -1555 -8066
rect -1511 -8066 -1495 -8048
rect -1393 -8048 -1317 -8032
rect -1393 -8066 -1377 -8048
rect -1511 -8082 -1473 -8066
rect -1593 -8120 -1473 -8082
rect -1415 -8082 -1377 -8066
rect -1333 -8066 -1317 -8048
rect -1215 -8048 -1139 -8032
rect -1215 -8066 -1199 -8048
rect -1333 -8082 -1295 -8066
rect -1415 -8120 -1295 -8082
rect -1237 -8082 -1199 -8066
rect -1155 -8066 -1139 -8048
rect -1037 -8048 -961 -8032
rect -1037 -8066 -1021 -8048
rect -1155 -8082 -1117 -8066
rect -1237 -8120 -1117 -8082
rect -1059 -8082 -1021 -8066
rect -977 -8066 -961 -8048
rect -859 -8048 -783 -8032
rect -859 -8066 -843 -8048
rect -977 -8082 -939 -8066
rect -1059 -8120 -939 -8082
rect -881 -8082 -843 -8066
rect -799 -8066 -783 -8048
rect -681 -8048 -605 -8032
rect -681 -8066 -665 -8048
rect -799 -8082 -761 -8066
rect -881 -8120 -761 -8082
rect -703 -8082 -665 -8066
rect -621 -8066 -605 -8048
rect -503 -8048 -427 -8032
rect -503 -8066 -487 -8048
rect -621 -8082 -583 -8066
rect -703 -8120 -583 -8082
rect -525 -8082 -487 -8066
rect -443 -8066 -427 -8048
rect -325 -8048 -249 -8032
rect -325 -8066 -309 -8048
rect -443 -8082 -405 -8066
rect -525 -8120 -405 -8082
rect -347 -8082 -309 -8066
rect -265 -8066 -249 -8048
rect -147 -8048 -71 -8032
rect -147 -8066 -131 -8048
rect -265 -8082 -227 -8066
rect -347 -8120 -227 -8082
rect -169 -8082 -131 -8066
rect -87 -8066 -71 -8048
rect 31 -8048 107 -8032
rect 31 -8066 47 -8048
rect -87 -8082 -49 -8066
rect -169 -8120 -49 -8082
rect 9 -8082 47 -8066
rect 91 -8066 107 -8048
rect 209 -8048 285 -8032
rect 209 -8066 225 -8048
rect 91 -8082 129 -8066
rect 9 -8120 129 -8082
rect 187 -8082 225 -8066
rect 269 -8066 285 -8048
rect 387 -8048 463 -8032
rect 387 -8066 403 -8048
rect 269 -8082 307 -8066
rect 187 -8120 307 -8082
rect 365 -8082 403 -8066
rect 447 -8066 463 -8048
rect 565 -8048 641 -8032
rect 565 -8066 581 -8048
rect 447 -8082 485 -8066
rect 365 -8120 485 -8082
rect 543 -8082 581 -8066
rect 625 -8066 641 -8048
rect 743 -8048 819 -8032
rect 743 -8066 759 -8048
rect 625 -8082 663 -8066
rect 543 -8120 663 -8082
rect 721 -8082 759 -8066
rect 803 -8066 819 -8048
rect 921 -8048 997 -8032
rect 921 -8066 937 -8048
rect 803 -8082 841 -8066
rect 721 -8120 841 -8082
rect 899 -8082 937 -8066
rect 981 -8066 997 -8048
rect 1099 -8048 1175 -8032
rect 1099 -8066 1115 -8048
rect 981 -8082 1019 -8066
rect 899 -8120 1019 -8082
rect 1077 -8082 1115 -8066
rect 1159 -8066 1175 -8048
rect 1277 -8048 1353 -8032
rect 1277 -8066 1293 -8048
rect 1159 -8082 1197 -8066
rect 1077 -8120 1197 -8082
rect 1255 -8082 1293 -8066
rect 1337 -8066 1353 -8048
rect 1455 -8048 1531 -8032
rect 1455 -8066 1471 -8048
rect 1337 -8082 1375 -8066
rect 1255 -8120 1375 -8082
rect 1433 -8082 1471 -8066
rect 1515 -8066 1531 -8048
rect 1633 -8048 1709 -8032
rect 1633 -8066 1649 -8048
rect 1515 -8082 1553 -8066
rect 1433 -8120 1553 -8082
rect 1611 -8082 1649 -8066
rect 1693 -8066 1709 -8048
rect 1811 -8048 1887 -8032
rect 1811 -8066 1827 -8048
rect 1693 -8082 1731 -8066
rect 1611 -8120 1731 -8082
rect 1789 -8082 1827 -8066
rect 1871 -8066 1887 -8048
rect 1989 -8048 2065 -8032
rect 1989 -8066 2005 -8048
rect 1871 -8082 1909 -8066
rect 1789 -8120 1909 -8082
rect 1967 -8082 2005 -8066
rect 2049 -8066 2065 -8048
rect 2167 -8048 2243 -8032
rect 2167 -8066 2183 -8048
rect 2049 -8082 2087 -8066
rect 1967 -8120 2087 -8082
rect 2145 -8082 2183 -8066
rect 2227 -8066 2243 -8048
rect 2345 -8048 2421 -8032
rect 2345 -8066 2361 -8048
rect 2227 -8082 2265 -8066
rect 2145 -8120 2265 -8082
rect 2323 -8082 2361 -8066
rect 2405 -8066 2421 -8048
rect 2523 -8048 2599 -8032
rect 2523 -8066 2539 -8048
rect 2405 -8082 2443 -8066
rect 2323 -8120 2443 -8082
rect 2501 -8082 2539 -8066
rect 2583 -8066 2599 -8048
rect 2701 -8048 2777 -8032
rect 2701 -8066 2717 -8048
rect 2583 -8082 2621 -8066
rect 2501 -8120 2621 -8082
rect 2679 -8082 2717 -8066
rect 2761 -8066 2777 -8048
rect 2879 -8048 2955 -8032
rect 2879 -8066 2895 -8048
rect 2761 -8082 2799 -8066
rect 2679 -8120 2799 -8082
rect 2857 -8082 2895 -8066
rect 2939 -8066 2955 -8048
rect 3057 -8048 3133 -8032
rect 3057 -8066 3073 -8048
rect 2939 -8082 2977 -8066
rect 2857 -8120 2977 -8082
rect 3035 -8082 3073 -8066
rect 3117 -8066 3133 -8048
rect 3235 -8048 3311 -8032
rect 3235 -8066 3251 -8048
rect 3117 -8082 3155 -8066
rect 3035 -8120 3155 -8082
rect 3213 -8082 3251 -8066
rect 3295 -8066 3311 -8048
rect 3413 -8048 3489 -8032
rect 3413 -8066 3429 -8048
rect 3295 -8082 3333 -8066
rect 3213 -8120 3333 -8082
rect 3391 -8082 3429 -8066
rect 3473 -8066 3489 -8048
rect 3591 -8048 3667 -8032
rect 3591 -8066 3607 -8048
rect 3473 -8082 3511 -8066
rect 3391 -8120 3511 -8082
rect 3569 -8082 3607 -8066
rect 3651 -8066 3667 -8048
rect 3769 -8048 3845 -8032
rect 3769 -8066 3785 -8048
rect 3651 -8082 3689 -8066
rect 3569 -8120 3689 -8082
rect 3747 -8082 3785 -8066
rect 3829 -8066 3845 -8048
rect 3947 -8048 4023 -8032
rect 3947 -8066 3963 -8048
rect 3829 -8082 3867 -8066
rect 3747 -8120 3867 -8082
rect 3925 -8082 3963 -8066
rect 4007 -8066 4023 -8048
rect 4007 -8082 4045 -8066
rect 3925 -8120 4045 -8082
rect -5582 -8180 -5462 -8142
rect -5582 -8196 -5544 -8180
rect -5560 -8214 -5544 -8196
rect -5500 -8196 -5462 -8180
rect -5404 -8180 -5284 -8142
rect -5404 -8196 -5366 -8180
rect -5500 -8214 -5484 -8196
rect -5560 -8230 -5484 -8214
rect -5382 -8214 -5366 -8196
rect -5322 -8196 -5284 -8180
rect -5226 -8180 -5106 -8142
rect -5226 -8196 -5188 -8180
rect -5322 -8214 -5306 -8196
rect -5382 -8230 -5306 -8214
rect -5204 -8214 -5188 -8196
rect -5144 -8196 -5106 -8180
rect -5048 -8180 -4928 -8142
rect -5048 -8196 -5010 -8180
rect -5144 -8214 -5128 -8196
rect -5204 -8230 -5128 -8214
rect -5026 -8214 -5010 -8196
rect -4966 -8196 -4928 -8180
rect -4870 -8180 -4750 -8142
rect -4870 -8196 -4832 -8180
rect -4966 -8214 -4950 -8196
rect -5026 -8230 -4950 -8214
rect -4848 -8214 -4832 -8196
rect -4788 -8196 -4750 -8180
rect -4692 -8180 -4572 -8142
rect -4692 -8196 -4654 -8180
rect -4788 -8214 -4772 -8196
rect -4848 -8230 -4772 -8214
rect -4670 -8214 -4654 -8196
rect -4610 -8196 -4572 -8180
rect -4514 -8180 -4394 -8142
rect -4514 -8196 -4476 -8180
rect -4610 -8214 -4594 -8196
rect -4670 -8230 -4594 -8214
rect -4492 -8214 -4476 -8196
rect -4432 -8196 -4394 -8180
rect -4336 -8180 -4216 -8142
rect -4336 -8196 -4298 -8180
rect -4432 -8214 -4416 -8196
rect -4492 -8230 -4416 -8214
rect -4314 -8214 -4298 -8196
rect -4254 -8196 -4216 -8180
rect -4158 -8180 -4038 -8142
rect -4158 -8196 -4120 -8180
rect -4254 -8214 -4238 -8196
rect -4314 -8230 -4238 -8214
rect -4136 -8214 -4120 -8196
rect -4076 -8196 -4038 -8180
rect -4076 -8214 -4060 -8196
rect -4136 -8230 -4060 -8214
rect -5560 -8340 -5484 -8324
rect -5560 -8358 -5544 -8340
rect -5582 -8374 -5544 -8358
rect -5500 -8358 -5484 -8340
rect -5382 -8340 -5306 -8324
rect -5382 -8358 -5366 -8340
rect -5500 -8374 -5462 -8358
rect -5582 -8412 -5462 -8374
rect -5404 -8374 -5366 -8358
rect -5322 -8358 -5306 -8340
rect -5204 -8340 -5128 -8324
rect -5204 -8358 -5188 -8340
rect -5322 -8374 -5284 -8358
rect -5404 -8412 -5284 -8374
rect -5226 -8374 -5188 -8358
rect -5144 -8358 -5128 -8340
rect -5026 -8340 -4950 -8324
rect -5026 -8358 -5010 -8340
rect -5144 -8374 -5106 -8358
rect -5226 -8412 -5106 -8374
rect -5048 -8374 -5010 -8358
rect -4966 -8358 -4950 -8340
rect -4848 -8340 -4772 -8324
rect -4848 -8358 -4832 -8340
rect -4966 -8374 -4928 -8358
rect -5048 -8412 -4928 -8374
rect -4870 -8374 -4832 -8358
rect -4788 -8358 -4772 -8340
rect -4670 -8340 -4594 -8324
rect -4670 -8358 -4654 -8340
rect -4788 -8374 -4750 -8358
rect -4870 -8412 -4750 -8374
rect -4692 -8374 -4654 -8358
rect -4610 -8358 -4594 -8340
rect -4492 -8340 -4416 -8324
rect -4492 -8358 -4476 -8340
rect -4610 -8374 -4572 -8358
rect -4692 -8412 -4572 -8374
rect -4514 -8374 -4476 -8358
rect -4432 -8358 -4416 -8340
rect -4314 -8340 -4238 -8324
rect -4314 -8358 -4298 -8340
rect -4432 -8374 -4394 -8358
rect -4514 -8412 -4394 -8374
rect -4336 -8374 -4298 -8358
rect -4254 -8358 -4238 -8340
rect -4136 -8340 -4060 -8324
rect -4136 -8358 -4120 -8340
rect -4254 -8374 -4216 -8358
rect -4336 -8412 -4216 -8374
rect -4158 -8374 -4120 -8358
rect -4076 -8358 -4060 -8340
rect -4076 -8374 -4038 -8358
rect -4158 -8412 -4038 -8374
rect -2127 -8438 -2007 -8400
rect -2127 -8454 -2089 -8438
rect -2105 -8472 -2089 -8454
rect -2045 -8454 -2007 -8438
rect -1949 -8438 -1829 -8400
rect -1949 -8454 -1911 -8438
rect -2045 -8472 -2029 -8454
rect -2105 -8488 -2029 -8472
rect -1927 -8472 -1911 -8454
rect -1867 -8454 -1829 -8438
rect -1771 -8438 -1651 -8400
rect -1771 -8454 -1733 -8438
rect -1867 -8472 -1851 -8454
rect -1927 -8488 -1851 -8472
rect -1749 -8472 -1733 -8454
rect -1689 -8454 -1651 -8438
rect -1593 -8438 -1473 -8400
rect -1593 -8454 -1555 -8438
rect -1689 -8472 -1673 -8454
rect -1749 -8488 -1673 -8472
rect -1571 -8472 -1555 -8454
rect -1511 -8454 -1473 -8438
rect -1415 -8438 -1295 -8400
rect -1415 -8454 -1377 -8438
rect -1511 -8472 -1495 -8454
rect -1571 -8488 -1495 -8472
rect -1393 -8472 -1377 -8454
rect -1333 -8454 -1295 -8438
rect -1237 -8438 -1117 -8400
rect -1237 -8454 -1199 -8438
rect -1333 -8472 -1317 -8454
rect -1393 -8488 -1317 -8472
rect -1215 -8472 -1199 -8454
rect -1155 -8454 -1117 -8438
rect -1059 -8438 -939 -8400
rect -1059 -8454 -1021 -8438
rect -1155 -8472 -1139 -8454
rect -1215 -8488 -1139 -8472
rect -1037 -8472 -1021 -8454
rect -977 -8454 -939 -8438
rect -881 -8438 -761 -8400
rect -881 -8454 -843 -8438
rect -977 -8472 -961 -8454
rect -1037 -8488 -961 -8472
rect -859 -8472 -843 -8454
rect -799 -8454 -761 -8438
rect -703 -8438 -583 -8400
rect -703 -8454 -665 -8438
rect -799 -8472 -783 -8454
rect -859 -8488 -783 -8472
rect -681 -8472 -665 -8454
rect -621 -8454 -583 -8438
rect -525 -8438 -405 -8400
rect -525 -8454 -487 -8438
rect -621 -8472 -605 -8454
rect -681 -8488 -605 -8472
rect -503 -8472 -487 -8454
rect -443 -8454 -405 -8438
rect -347 -8438 -227 -8400
rect -347 -8454 -309 -8438
rect -443 -8472 -427 -8454
rect -503 -8488 -427 -8472
rect -325 -8472 -309 -8454
rect -265 -8454 -227 -8438
rect -169 -8438 -49 -8400
rect -169 -8454 -131 -8438
rect -265 -8472 -249 -8454
rect -325 -8488 -249 -8472
rect -147 -8472 -131 -8454
rect -87 -8454 -49 -8438
rect 9 -8438 129 -8400
rect 9 -8454 47 -8438
rect -87 -8472 -71 -8454
rect -147 -8488 -71 -8472
rect 31 -8472 47 -8454
rect 91 -8454 129 -8438
rect 187 -8438 307 -8400
rect 187 -8454 225 -8438
rect 91 -8472 107 -8454
rect 31 -8488 107 -8472
rect 209 -8472 225 -8454
rect 269 -8454 307 -8438
rect 365 -8438 485 -8400
rect 365 -8454 403 -8438
rect 269 -8472 285 -8454
rect 209 -8488 285 -8472
rect 387 -8472 403 -8454
rect 447 -8454 485 -8438
rect 543 -8438 663 -8400
rect 543 -8454 581 -8438
rect 447 -8472 463 -8454
rect 387 -8488 463 -8472
rect 565 -8472 581 -8454
rect 625 -8454 663 -8438
rect 721 -8438 841 -8400
rect 721 -8454 759 -8438
rect 625 -8472 641 -8454
rect 565 -8488 641 -8472
rect 743 -8472 759 -8454
rect 803 -8454 841 -8438
rect 899 -8438 1019 -8400
rect 899 -8454 937 -8438
rect 803 -8472 819 -8454
rect 743 -8488 819 -8472
rect 921 -8472 937 -8454
rect 981 -8454 1019 -8438
rect 1077 -8438 1197 -8400
rect 1077 -8454 1115 -8438
rect 981 -8472 997 -8454
rect 921 -8488 997 -8472
rect 1099 -8472 1115 -8454
rect 1159 -8454 1197 -8438
rect 1255 -8438 1375 -8400
rect 1255 -8454 1293 -8438
rect 1159 -8472 1175 -8454
rect 1099 -8488 1175 -8472
rect 1277 -8472 1293 -8454
rect 1337 -8454 1375 -8438
rect 1433 -8438 1553 -8400
rect 1433 -8454 1471 -8438
rect 1337 -8472 1353 -8454
rect 1277 -8488 1353 -8472
rect 1455 -8472 1471 -8454
rect 1515 -8454 1553 -8438
rect 1611 -8438 1731 -8400
rect 1611 -8454 1649 -8438
rect 1515 -8472 1531 -8454
rect 1455 -8488 1531 -8472
rect 1633 -8472 1649 -8454
rect 1693 -8454 1731 -8438
rect 1789 -8438 1909 -8400
rect 1789 -8454 1827 -8438
rect 1693 -8472 1709 -8454
rect 1633 -8488 1709 -8472
rect 1811 -8472 1827 -8454
rect 1871 -8454 1909 -8438
rect 1967 -8438 2087 -8400
rect 1967 -8454 2005 -8438
rect 1871 -8472 1887 -8454
rect 1811 -8488 1887 -8472
rect 1989 -8472 2005 -8454
rect 2049 -8454 2087 -8438
rect 2145 -8438 2265 -8400
rect 2145 -8454 2183 -8438
rect 2049 -8472 2065 -8454
rect 1989 -8488 2065 -8472
rect 2167 -8472 2183 -8454
rect 2227 -8454 2265 -8438
rect 2323 -8438 2443 -8400
rect 2323 -8454 2361 -8438
rect 2227 -8472 2243 -8454
rect 2167 -8488 2243 -8472
rect 2345 -8472 2361 -8454
rect 2405 -8454 2443 -8438
rect 2501 -8438 2621 -8400
rect 2501 -8454 2539 -8438
rect 2405 -8472 2421 -8454
rect 2345 -8488 2421 -8472
rect 2523 -8472 2539 -8454
rect 2583 -8454 2621 -8438
rect 2679 -8438 2799 -8400
rect 2679 -8454 2717 -8438
rect 2583 -8472 2599 -8454
rect 2523 -8488 2599 -8472
rect 2701 -8472 2717 -8454
rect 2761 -8454 2799 -8438
rect 2857 -8438 2977 -8400
rect 2857 -8454 2895 -8438
rect 2761 -8472 2777 -8454
rect 2701 -8488 2777 -8472
rect 2879 -8472 2895 -8454
rect 2939 -8454 2977 -8438
rect 3035 -8438 3155 -8400
rect 3035 -8454 3073 -8438
rect 2939 -8472 2955 -8454
rect 2879 -8488 2955 -8472
rect 3057 -8472 3073 -8454
rect 3117 -8454 3155 -8438
rect 3213 -8438 3333 -8400
rect 3213 -8454 3251 -8438
rect 3117 -8472 3133 -8454
rect 3057 -8488 3133 -8472
rect 3235 -8472 3251 -8454
rect 3295 -8454 3333 -8438
rect 3391 -8438 3511 -8400
rect 3391 -8454 3429 -8438
rect 3295 -8472 3311 -8454
rect 3235 -8488 3311 -8472
rect 3413 -8472 3429 -8454
rect 3473 -8454 3511 -8438
rect 3569 -8438 3689 -8400
rect 3569 -8454 3607 -8438
rect 3473 -8472 3489 -8454
rect 3413 -8488 3489 -8472
rect 3591 -8472 3607 -8454
rect 3651 -8454 3689 -8438
rect 3747 -8438 3867 -8400
rect 3747 -8454 3785 -8438
rect 3651 -8472 3667 -8454
rect 3591 -8488 3667 -8472
rect 3769 -8472 3785 -8454
rect 3829 -8454 3867 -8438
rect 3925 -8438 4045 -8400
rect 3925 -8454 3963 -8438
rect 3829 -8472 3845 -8454
rect 3769 -8488 3845 -8472
rect 3947 -8472 3963 -8454
rect 4007 -8454 4045 -8438
rect 4007 -8472 4023 -8454
rect 3947 -8488 4023 -8472
rect -5582 -8730 -5462 -8692
rect -5582 -8746 -5544 -8730
rect -5560 -8764 -5544 -8746
rect -5500 -8746 -5462 -8730
rect -5404 -8730 -5284 -8692
rect -5404 -8746 -5366 -8730
rect -5500 -8764 -5484 -8746
rect -5560 -8780 -5484 -8764
rect -5382 -8764 -5366 -8746
rect -5322 -8746 -5284 -8730
rect -5226 -8730 -5106 -8692
rect -5226 -8746 -5188 -8730
rect -5322 -8764 -5306 -8746
rect -5382 -8780 -5306 -8764
rect -5204 -8764 -5188 -8746
rect -5144 -8746 -5106 -8730
rect -5048 -8730 -4928 -8692
rect -5048 -8746 -5010 -8730
rect -5144 -8764 -5128 -8746
rect -5204 -8780 -5128 -8764
rect -5026 -8764 -5010 -8746
rect -4966 -8746 -4928 -8730
rect -4870 -8730 -4750 -8692
rect -4870 -8746 -4832 -8730
rect -4966 -8764 -4950 -8746
rect -5026 -8780 -4950 -8764
rect -4848 -8764 -4832 -8746
rect -4788 -8746 -4750 -8730
rect -4692 -8730 -4572 -8692
rect -4692 -8746 -4654 -8730
rect -4788 -8764 -4772 -8746
rect -4848 -8780 -4772 -8764
rect -4670 -8764 -4654 -8746
rect -4610 -8746 -4572 -8730
rect -4514 -8730 -4394 -8692
rect -4514 -8746 -4476 -8730
rect -4610 -8764 -4594 -8746
rect -4670 -8780 -4594 -8764
rect -4492 -8764 -4476 -8746
rect -4432 -8746 -4394 -8730
rect -4336 -8730 -4216 -8692
rect -4336 -8746 -4298 -8730
rect -4432 -8764 -4416 -8746
rect -4492 -8780 -4416 -8764
rect -4314 -8764 -4298 -8746
rect -4254 -8746 -4216 -8730
rect -4158 -8730 -4038 -8692
rect -4158 -8746 -4120 -8730
rect -4254 -8764 -4238 -8746
rect -4314 -8780 -4238 -8764
rect -4136 -8764 -4120 -8746
rect -4076 -8746 -4038 -8730
rect -4076 -8764 -4060 -8746
rect -4136 -8780 -4060 -8764
rect 6580 -8810 6656 -8794
rect 6580 -8828 6596 -8810
rect 6558 -8844 6596 -8828
rect 6640 -8828 6656 -8810
rect 6758 -8810 6834 -8794
rect 6758 -8828 6774 -8810
rect 6640 -8844 6678 -8828
rect -5560 -8890 -5484 -8874
rect -5560 -8908 -5544 -8890
rect -5582 -8924 -5544 -8908
rect -5500 -8908 -5484 -8890
rect -5382 -8890 -5306 -8874
rect -5382 -8908 -5366 -8890
rect -5500 -8924 -5462 -8908
rect -5582 -8962 -5462 -8924
rect -5404 -8924 -5366 -8908
rect -5322 -8908 -5306 -8890
rect -5204 -8890 -5128 -8874
rect -5204 -8908 -5188 -8890
rect -5322 -8924 -5284 -8908
rect -5404 -8962 -5284 -8924
rect -5226 -8924 -5188 -8908
rect -5144 -8908 -5128 -8890
rect -5026 -8890 -4950 -8874
rect -5026 -8908 -5010 -8890
rect -5144 -8924 -5106 -8908
rect -5226 -8962 -5106 -8924
rect -5048 -8924 -5010 -8908
rect -4966 -8908 -4950 -8890
rect -4848 -8890 -4772 -8874
rect -4848 -8908 -4832 -8890
rect -4966 -8924 -4928 -8908
rect -5048 -8962 -4928 -8924
rect -4870 -8924 -4832 -8908
rect -4788 -8908 -4772 -8890
rect -4670 -8890 -4594 -8874
rect -4670 -8908 -4654 -8890
rect -4788 -8924 -4750 -8908
rect -4870 -8962 -4750 -8924
rect -4692 -8924 -4654 -8908
rect -4610 -8908 -4594 -8890
rect -4492 -8890 -4416 -8874
rect -4492 -8908 -4476 -8890
rect -4610 -8924 -4572 -8908
rect -4692 -8962 -4572 -8924
rect -4514 -8924 -4476 -8908
rect -4432 -8908 -4416 -8890
rect -4314 -8890 -4238 -8874
rect -4314 -8908 -4298 -8890
rect -4432 -8924 -4394 -8908
rect -4514 -8962 -4394 -8924
rect -4336 -8924 -4298 -8908
rect -4254 -8908 -4238 -8890
rect -4136 -8890 -4060 -8874
rect 6558 -8882 6678 -8844
rect 6736 -8844 6774 -8828
rect 6818 -8828 6834 -8810
rect 6936 -8810 7012 -8794
rect 6936 -8828 6952 -8810
rect 6818 -8844 6856 -8828
rect 6736 -8882 6856 -8844
rect 6914 -8844 6952 -8828
rect 6996 -8828 7012 -8810
rect 7114 -8810 7190 -8794
rect 7114 -8828 7130 -8810
rect 6996 -8844 7034 -8828
rect 6914 -8882 7034 -8844
rect 7092 -8844 7130 -8828
rect 7174 -8828 7190 -8810
rect 7292 -8810 7368 -8794
rect 7292 -8828 7308 -8810
rect 7174 -8844 7212 -8828
rect 7092 -8882 7212 -8844
rect 7270 -8844 7308 -8828
rect 7352 -8828 7368 -8810
rect 7470 -8810 7546 -8794
rect 7470 -8828 7486 -8810
rect 7352 -8844 7390 -8828
rect 7270 -8882 7390 -8844
rect 7448 -8844 7486 -8828
rect 7530 -8828 7546 -8810
rect 7648 -8810 7724 -8794
rect 7648 -8828 7664 -8810
rect 7530 -8844 7568 -8828
rect 7448 -8882 7568 -8844
rect 7626 -8844 7664 -8828
rect 7708 -8828 7724 -8810
rect 7826 -8810 7902 -8794
rect 7826 -8828 7842 -8810
rect 7708 -8844 7746 -8828
rect 7626 -8882 7746 -8844
rect 7804 -8844 7842 -8828
rect 7886 -8828 7902 -8810
rect 8004 -8810 8080 -8794
rect 8004 -8828 8020 -8810
rect 7886 -8844 7924 -8828
rect 7804 -8882 7924 -8844
rect 7982 -8844 8020 -8828
rect 8064 -8828 8080 -8810
rect 8182 -8810 8258 -8794
rect 8182 -8828 8198 -8810
rect 8064 -8844 8102 -8828
rect 7982 -8882 8102 -8844
rect 8160 -8844 8198 -8828
rect 8242 -8828 8258 -8810
rect 8360 -8810 8436 -8794
rect 8360 -8828 8376 -8810
rect 8242 -8844 8280 -8828
rect 8160 -8882 8280 -8844
rect 8338 -8844 8376 -8828
rect 8420 -8828 8436 -8810
rect 8538 -8810 8614 -8794
rect 8538 -8828 8554 -8810
rect 8420 -8844 8458 -8828
rect 8338 -8882 8458 -8844
rect 8516 -8844 8554 -8828
rect 8598 -8828 8614 -8810
rect 8716 -8810 8792 -8794
rect 8716 -8828 8732 -8810
rect 8598 -8844 8636 -8828
rect 8516 -8882 8636 -8844
rect 8694 -8844 8732 -8828
rect 8776 -8828 8792 -8810
rect 8894 -8810 8970 -8794
rect 8894 -8828 8910 -8810
rect 8776 -8844 8814 -8828
rect 8694 -8882 8814 -8844
rect 8872 -8844 8910 -8828
rect 8954 -8828 8970 -8810
rect 9072 -8810 9148 -8794
rect 9072 -8828 9088 -8810
rect 8954 -8844 8992 -8828
rect 8872 -8882 8992 -8844
rect 9050 -8844 9088 -8828
rect 9132 -8828 9148 -8810
rect 9250 -8810 9326 -8794
rect 9250 -8828 9266 -8810
rect 9132 -8844 9170 -8828
rect 9050 -8882 9170 -8844
rect 9228 -8844 9266 -8828
rect 9310 -8828 9326 -8810
rect 9310 -8844 9348 -8828
rect 9228 -8882 9348 -8844
rect 10840 -8840 10916 -8824
rect 10840 -8858 10856 -8840
rect 10818 -8874 10856 -8858
rect 10900 -8858 10916 -8840
rect 11132 -8840 11208 -8824
rect 11132 -8858 11148 -8840
rect 10900 -8874 10938 -8858
rect -4136 -8908 -4120 -8890
rect -4254 -8924 -4216 -8908
rect -4336 -8962 -4216 -8924
rect -4158 -8924 -4120 -8908
rect -4076 -8908 -4060 -8890
rect -4076 -8924 -4038 -8908
rect -4158 -8962 -4038 -8924
rect -2105 -9048 -2029 -9032
rect -2105 -9066 -2089 -9048
rect -2127 -9082 -2089 -9066
rect -2045 -9066 -2029 -9048
rect -1927 -9048 -1851 -9032
rect -1927 -9066 -1911 -9048
rect -2045 -9082 -2007 -9066
rect -2127 -9120 -2007 -9082
rect -1949 -9082 -1911 -9066
rect -1867 -9066 -1851 -9048
rect -1749 -9048 -1673 -9032
rect -1749 -9066 -1733 -9048
rect -1867 -9082 -1829 -9066
rect -1949 -9120 -1829 -9082
rect -1771 -9082 -1733 -9066
rect -1689 -9066 -1673 -9048
rect -1571 -9048 -1495 -9032
rect -1571 -9066 -1555 -9048
rect -1689 -9082 -1651 -9066
rect -1771 -9120 -1651 -9082
rect -1593 -9082 -1555 -9066
rect -1511 -9066 -1495 -9048
rect -1393 -9048 -1317 -9032
rect -1393 -9066 -1377 -9048
rect -1511 -9082 -1473 -9066
rect -1593 -9120 -1473 -9082
rect -1415 -9082 -1377 -9066
rect -1333 -9066 -1317 -9048
rect -1215 -9048 -1139 -9032
rect -1215 -9066 -1199 -9048
rect -1333 -9082 -1295 -9066
rect -1415 -9120 -1295 -9082
rect -1237 -9082 -1199 -9066
rect -1155 -9066 -1139 -9048
rect -1037 -9048 -961 -9032
rect -1037 -9066 -1021 -9048
rect -1155 -9082 -1117 -9066
rect -1237 -9120 -1117 -9082
rect -1059 -9082 -1021 -9066
rect -977 -9066 -961 -9048
rect -859 -9048 -783 -9032
rect -859 -9066 -843 -9048
rect -977 -9082 -939 -9066
rect -1059 -9120 -939 -9082
rect -881 -9082 -843 -9066
rect -799 -9066 -783 -9048
rect -681 -9048 -605 -9032
rect -681 -9066 -665 -9048
rect -799 -9082 -761 -9066
rect -881 -9120 -761 -9082
rect -703 -9082 -665 -9066
rect -621 -9066 -605 -9048
rect -503 -9048 -427 -9032
rect -503 -9066 -487 -9048
rect -621 -9082 -583 -9066
rect -703 -9120 -583 -9082
rect -525 -9082 -487 -9066
rect -443 -9066 -427 -9048
rect -325 -9048 -249 -9032
rect -325 -9066 -309 -9048
rect -443 -9082 -405 -9066
rect -525 -9120 -405 -9082
rect -347 -9082 -309 -9066
rect -265 -9066 -249 -9048
rect -147 -9048 -71 -9032
rect -147 -9066 -131 -9048
rect -265 -9082 -227 -9066
rect -347 -9120 -227 -9082
rect -169 -9082 -131 -9066
rect -87 -9066 -71 -9048
rect 31 -9048 107 -9032
rect 31 -9066 47 -9048
rect -87 -9082 -49 -9066
rect -169 -9120 -49 -9082
rect 9 -9082 47 -9066
rect 91 -9066 107 -9048
rect 209 -9048 285 -9032
rect 209 -9066 225 -9048
rect 91 -9082 129 -9066
rect 9 -9120 129 -9082
rect 187 -9082 225 -9066
rect 269 -9066 285 -9048
rect 387 -9048 463 -9032
rect 387 -9066 403 -9048
rect 269 -9082 307 -9066
rect 187 -9120 307 -9082
rect 365 -9082 403 -9066
rect 447 -9066 463 -9048
rect 565 -9048 641 -9032
rect 565 -9066 581 -9048
rect 447 -9082 485 -9066
rect 365 -9120 485 -9082
rect 543 -9082 581 -9066
rect 625 -9066 641 -9048
rect 743 -9048 819 -9032
rect 743 -9066 759 -9048
rect 625 -9082 663 -9066
rect 543 -9120 663 -9082
rect 721 -9082 759 -9066
rect 803 -9066 819 -9048
rect 921 -9048 997 -9032
rect 921 -9066 937 -9048
rect 803 -9082 841 -9066
rect 721 -9120 841 -9082
rect 899 -9082 937 -9066
rect 981 -9066 997 -9048
rect 1099 -9048 1175 -9032
rect 1099 -9066 1115 -9048
rect 981 -9082 1019 -9066
rect 899 -9120 1019 -9082
rect 1077 -9082 1115 -9066
rect 1159 -9066 1175 -9048
rect 1277 -9048 1353 -9032
rect 1277 -9066 1293 -9048
rect 1159 -9082 1197 -9066
rect 1077 -9120 1197 -9082
rect 1255 -9082 1293 -9066
rect 1337 -9066 1353 -9048
rect 1455 -9048 1531 -9032
rect 1455 -9066 1471 -9048
rect 1337 -9082 1375 -9066
rect 1255 -9120 1375 -9082
rect 1433 -9082 1471 -9066
rect 1515 -9066 1531 -9048
rect 1633 -9048 1709 -9032
rect 1633 -9066 1649 -9048
rect 1515 -9082 1553 -9066
rect 1433 -9120 1553 -9082
rect 1611 -9082 1649 -9066
rect 1693 -9066 1709 -9048
rect 1811 -9048 1887 -9032
rect 1811 -9066 1827 -9048
rect 1693 -9082 1731 -9066
rect 1611 -9120 1731 -9082
rect 1789 -9082 1827 -9066
rect 1871 -9066 1887 -9048
rect 1989 -9048 2065 -9032
rect 1989 -9066 2005 -9048
rect 1871 -9082 1909 -9066
rect 1789 -9120 1909 -9082
rect 1967 -9082 2005 -9066
rect 2049 -9066 2065 -9048
rect 2167 -9048 2243 -9032
rect 2167 -9066 2183 -9048
rect 2049 -9082 2087 -9066
rect 1967 -9120 2087 -9082
rect 2145 -9082 2183 -9066
rect 2227 -9066 2243 -9048
rect 2345 -9048 2421 -9032
rect 2345 -9066 2361 -9048
rect 2227 -9082 2265 -9066
rect 2145 -9120 2265 -9082
rect 2323 -9082 2361 -9066
rect 2405 -9066 2421 -9048
rect 2523 -9048 2599 -9032
rect 2523 -9066 2539 -9048
rect 2405 -9082 2443 -9066
rect 2323 -9120 2443 -9082
rect 2501 -9082 2539 -9066
rect 2583 -9066 2599 -9048
rect 2701 -9048 2777 -9032
rect 2701 -9066 2717 -9048
rect 2583 -9082 2621 -9066
rect 2501 -9120 2621 -9082
rect 2679 -9082 2717 -9066
rect 2761 -9066 2777 -9048
rect 2879 -9048 2955 -9032
rect 2879 -9066 2895 -9048
rect 2761 -9082 2799 -9066
rect 2679 -9120 2799 -9082
rect 2857 -9082 2895 -9066
rect 2939 -9066 2955 -9048
rect 3057 -9048 3133 -9032
rect 3057 -9066 3073 -9048
rect 2939 -9082 2977 -9066
rect 2857 -9120 2977 -9082
rect 3035 -9082 3073 -9066
rect 3117 -9066 3133 -9048
rect 3235 -9048 3311 -9032
rect 3235 -9066 3251 -9048
rect 3117 -9082 3155 -9066
rect 3035 -9120 3155 -9082
rect 3213 -9082 3251 -9066
rect 3295 -9066 3311 -9048
rect 3413 -9048 3489 -9032
rect 3413 -9066 3429 -9048
rect 3295 -9082 3333 -9066
rect 3213 -9120 3333 -9082
rect 3391 -9082 3429 -9066
rect 3473 -9066 3489 -9048
rect 3591 -9048 3667 -9032
rect 3591 -9066 3607 -9048
rect 3473 -9082 3511 -9066
rect 3391 -9120 3511 -9082
rect 3569 -9082 3607 -9066
rect 3651 -9066 3667 -9048
rect 3769 -9048 3845 -9032
rect 3769 -9066 3785 -9048
rect 3651 -9082 3689 -9066
rect 3569 -9120 3689 -9082
rect 3747 -9082 3785 -9066
rect 3829 -9066 3845 -9048
rect 3947 -9048 4023 -9032
rect 3947 -9066 3963 -9048
rect 3829 -9082 3867 -9066
rect 3747 -9120 3867 -9082
rect 3925 -9082 3963 -9066
rect 4007 -9066 4023 -9048
rect 4007 -9082 4045 -9066
rect 3925 -9120 4045 -9082
rect -5582 -9280 -5462 -9242
rect -5582 -9296 -5544 -9280
rect -5560 -9314 -5544 -9296
rect -5500 -9296 -5462 -9280
rect -5404 -9280 -5284 -9242
rect -5404 -9296 -5366 -9280
rect -5500 -9314 -5484 -9296
rect -5560 -9330 -5484 -9314
rect -5382 -9314 -5366 -9296
rect -5322 -9296 -5284 -9280
rect -5226 -9280 -5106 -9242
rect -5226 -9296 -5188 -9280
rect -5322 -9314 -5306 -9296
rect -5382 -9330 -5306 -9314
rect -5204 -9314 -5188 -9296
rect -5144 -9296 -5106 -9280
rect -5048 -9280 -4928 -9242
rect -5048 -9296 -5010 -9280
rect -5144 -9314 -5128 -9296
rect -5204 -9330 -5128 -9314
rect -5026 -9314 -5010 -9296
rect -4966 -9296 -4928 -9280
rect -4870 -9280 -4750 -9242
rect -4870 -9296 -4832 -9280
rect -4966 -9314 -4950 -9296
rect -5026 -9330 -4950 -9314
rect -4848 -9314 -4832 -9296
rect -4788 -9296 -4750 -9280
rect -4692 -9280 -4572 -9242
rect -4692 -9296 -4654 -9280
rect -4788 -9314 -4772 -9296
rect -4848 -9330 -4772 -9314
rect -4670 -9314 -4654 -9296
rect -4610 -9296 -4572 -9280
rect -4514 -9280 -4394 -9242
rect -4514 -9296 -4476 -9280
rect -4610 -9314 -4594 -9296
rect -4670 -9330 -4594 -9314
rect -4492 -9314 -4476 -9296
rect -4432 -9296 -4394 -9280
rect -4336 -9280 -4216 -9242
rect -4336 -9296 -4298 -9280
rect -4432 -9314 -4416 -9296
rect -4492 -9330 -4416 -9314
rect -4314 -9314 -4298 -9296
rect -4254 -9296 -4216 -9280
rect -4158 -9280 -4038 -9242
rect -4158 -9296 -4120 -9280
rect -4254 -9314 -4238 -9296
rect -4314 -9330 -4238 -9314
rect -4136 -9314 -4120 -9296
rect -4076 -9296 -4038 -9280
rect -4076 -9314 -4060 -9296
rect -4136 -9330 -4060 -9314
rect -5560 -9440 -5484 -9424
rect -5560 -9458 -5544 -9440
rect -5582 -9474 -5544 -9458
rect -5500 -9458 -5484 -9440
rect -5382 -9440 -5306 -9424
rect -5382 -9458 -5366 -9440
rect -5500 -9474 -5462 -9458
rect -5582 -9512 -5462 -9474
rect -5404 -9474 -5366 -9458
rect -5322 -9458 -5306 -9440
rect -5204 -9440 -5128 -9424
rect -5204 -9458 -5188 -9440
rect -5322 -9474 -5284 -9458
rect -5404 -9512 -5284 -9474
rect -5226 -9474 -5188 -9458
rect -5144 -9458 -5128 -9440
rect -5026 -9440 -4950 -9424
rect -5026 -9458 -5010 -9440
rect -5144 -9474 -5106 -9458
rect -5226 -9512 -5106 -9474
rect -5048 -9474 -5010 -9458
rect -4966 -9458 -4950 -9440
rect -4848 -9440 -4772 -9424
rect -4848 -9458 -4832 -9440
rect -4966 -9474 -4928 -9458
rect -5048 -9512 -4928 -9474
rect -4870 -9474 -4832 -9458
rect -4788 -9458 -4772 -9440
rect -4670 -9440 -4594 -9424
rect -4670 -9458 -4654 -9440
rect -4788 -9474 -4750 -9458
rect -4870 -9512 -4750 -9474
rect -4692 -9474 -4654 -9458
rect -4610 -9458 -4594 -9440
rect -4492 -9440 -4416 -9424
rect -4492 -9458 -4476 -9440
rect -4610 -9474 -4572 -9458
rect -4692 -9512 -4572 -9474
rect -4514 -9474 -4476 -9458
rect -4432 -9458 -4416 -9440
rect -4314 -9440 -4238 -9424
rect -4314 -9458 -4298 -9440
rect -4432 -9474 -4394 -9458
rect -4514 -9512 -4394 -9474
rect -4336 -9474 -4298 -9458
rect -4254 -9458 -4238 -9440
rect -4136 -9440 -4060 -9424
rect -4136 -9458 -4120 -9440
rect -4254 -9474 -4216 -9458
rect -4336 -9512 -4216 -9474
rect -4158 -9474 -4120 -9458
rect -4076 -9458 -4060 -9440
rect 10818 -8912 10938 -8874
rect 11110 -8874 11148 -8858
rect 11192 -8858 11208 -8840
rect 11424 -8840 11500 -8824
rect 11424 -8858 11440 -8840
rect 11192 -8874 11230 -8858
rect 11110 -8912 11230 -8874
rect 11402 -8874 11440 -8858
rect 11484 -8858 11500 -8840
rect 11716 -8840 11792 -8824
rect 11716 -8858 11732 -8840
rect 11484 -8874 11522 -8858
rect 11402 -8912 11522 -8874
rect 11694 -8874 11732 -8858
rect 11776 -8858 11792 -8840
rect 12008 -8840 12084 -8824
rect 12008 -8858 12024 -8840
rect 11776 -8874 11814 -8858
rect 11694 -8912 11814 -8874
rect 11986 -8874 12024 -8858
rect 12068 -8858 12084 -8840
rect 12300 -8840 12376 -8824
rect 12300 -8858 12316 -8840
rect 12068 -8874 12106 -8858
rect 11986 -8912 12106 -8874
rect 12278 -8874 12316 -8858
rect 12360 -8858 12376 -8840
rect 12592 -8840 12668 -8824
rect 12592 -8858 12608 -8840
rect 12360 -8874 12398 -8858
rect 12278 -8912 12398 -8874
rect 12570 -8874 12608 -8858
rect 12652 -8858 12668 -8840
rect 12652 -8874 12690 -8858
rect 12570 -8912 12690 -8874
rect 6558 -9200 6678 -9162
rect 6558 -9216 6596 -9200
rect 6580 -9234 6596 -9216
rect 6640 -9216 6678 -9200
rect 6736 -9200 6856 -9162
rect 6736 -9216 6774 -9200
rect 6640 -9234 6656 -9216
rect 6580 -9250 6656 -9234
rect 6758 -9234 6774 -9216
rect 6818 -9216 6856 -9200
rect 6914 -9200 7034 -9162
rect 6914 -9216 6952 -9200
rect 6818 -9234 6834 -9216
rect 6758 -9250 6834 -9234
rect 6936 -9234 6952 -9216
rect 6996 -9216 7034 -9200
rect 7092 -9200 7212 -9162
rect 7092 -9216 7130 -9200
rect 6996 -9234 7012 -9216
rect 6936 -9250 7012 -9234
rect 7114 -9234 7130 -9216
rect 7174 -9216 7212 -9200
rect 7270 -9200 7390 -9162
rect 7270 -9216 7308 -9200
rect 7174 -9234 7190 -9216
rect 7114 -9250 7190 -9234
rect 7292 -9234 7308 -9216
rect 7352 -9216 7390 -9200
rect 7448 -9200 7568 -9162
rect 7448 -9216 7486 -9200
rect 7352 -9234 7368 -9216
rect 7292 -9250 7368 -9234
rect 7470 -9234 7486 -9216
rect 7530 -9216 7568 -9200
rect 7626 -9200 7746 -9162
rect 7626 -9216 7664 -9200
rect 7530 -9234 7546 -9216
rect 7470 -9250 7546 -9234
rect 7648 -9234 7664 -9216
rect 7708 -9216 7746 -9200
rect 7804 -9200 7924 -9162
rect 7804 -9216 7842 -9200
rect 7708 -9234 7724 -9216
rect 7648 -9250 7724 -9234
rect 7826 -9234 7842 -9216
rect 7886 -9216 7924 -9200
rect 7982 -9200 8102 -9162
rect 7982 -9216 8020 -9200
rect 7886 -9234 7902 -9216
rect 7826 -9250 7902 -9234
rect 8004 -9234 8020 -9216
rect 8064 -9216 8102 -9200
rect 8160 -9200 8280 -9162
rect 8160 -9216 8198 -9200
rect 8064 -9234 8080 -9216
rect 8004 -9250 8080 -9234
rect 8182 -9234 8198 -9216
rect 8242 -9216 8280 -9200
rect 8338 -9200 8458 -9162
rect 8338 -9216 8376 -9200
rect 8242 -9234 8258 -9216
rect 8182 -9250 8258 -9234
rect 8360 -9234 8376 -9216
rect 8420 -9216 8458 -9200
rect 8516 -9200 8636 -9162
rect 8516 -9216 8554 -9200
rect 8420 -9234 8436 -9216
rect 8360 -9250 8436 -9234
rect 8538 -9234 8554 -9216
rect 8598 -9216 8636 -9200
rect 8694 -9200 8814 -9162
rect 8694 -9216 8732 -9200
rect 8598 -9234 8614 -9216
rect 8538 -9250 8614 -9234
rect 8716 -9234 8732 -9216
rect 8776 -9216 8814 -9200
rect 8872 -9200 8992 -9162
rect 8872 -9216 8910 -9200
rect 8776 -9234 8792 -9216
rect 8716 -9250 8792 -9234
rect 8894 -9234 8910 -9216
rect 8954 -9216 8992 -9200
rect 9050 -9200 9170 -9162
rect 9050 -9216 9088 -9200
rect 8954 -9234 8970 -9216
rect 8894 -9250 8970 -9234
rect 9072 -9234 9088 -9216
rect 9132 -9216 9170 -9200
rect 9228 -9200 9348 -9162
rect 9228 -9216 9266 -9200
rect 9132 -9234 9148 -9216
rect 9072 -9250 9148 -9234
rect 9250 -9234 9266 -9216
rect 9310 -9216 9348 -9200
rect 9310 -9234 9326 -9216
rect 9250 -9250 9326 -9234
rect 10818 -9230 10938 -9192
rect 10818 -9246 10856 -9230
rect 10840 -9264 10856 -9246
rect 10900 -9246 10938 -9230
rect 11110 -9230 11230 -9192
rect 11110 -9246 11148 -9230
rect 10900 -9264 10916 -9246
rect 10840 -9280 10916 -9264
rect 11132 -9264 11148 -9246
rect 11192 -9246 11230 -9230
rect 11402 -9230 11522 -9192
rect 11402 -9246 11440 -9230
rect 11192 -9264 11208 -9246
rect 11132 -9280 11208 -9264
rect 11424 -9264 11440 -9246
rect 11484 -9246 11522 -9230
rect 11694 -9230 11814 -9192
rect 11694 -9246 11732 -9230
rect 11484 -9264 11500 -9246
rect 11424 -9280 11500 -9264
rect 11716 -9264 11732 -9246
rect 11776 -9246 11814 -9230
rect 11986 -9230 12106 -9192
rect 11986 -9246 12024 -9230
rect 11776 -9264 11792 -9246
rect 11716 -9280 11792 -9264
rect 12008 -9264 12024 -9246
rect 12068 -9246 12106 -9230
rect 12278 -9230 12398 -9192
rect 12278 -9246 12316 -9230
rect 12068 -9264 12084 -9246
rect 12008 -9280 12084 -9264
rect 12300 -9264 12316 -9246
rect 12360 -9246 12398 -9230
rect 12570 -9230 12690 -9192
rect 12570 -9246 12608 -9230
rect 12360 -9264 12376 -9246
rect 12300 -9280 12376 -9264
rect 12592 -9264 12608 -9246
rect 12652 -9246 12690 -9230
rect 12652 -9264 12668 -9246
rect 12592 -9280 12668 -9264
rect -2127 -9438 -2007 -9400
rect -2127 -9454 -2089 -9438
rect -4076 -9474 -4038 -9458
rect -4158 -9512 -4038 -9474
rect -2105 -9472 -2089 -9454
rect -2045 -9454 -2007 -9438
rect -1949 -9438 -1829 -9400
rect -1949 -9454 -1911 -9438
rect -2045 -9472 -2029 -9454
rect -2105 -9488 -2029 -9472
rect -1927 -9472 -1911 -9454
rect -1867 -9454 -1829 -9438
rect -1771 -9438 -1651 -9400
rect -1771 -9454 -1733 -9438
rect -1867 -9472 -1851 -9454
rect -1927 -9488 -1851 -9472
rect -1749 -9472 -1733 -9454
rect -1689 -9454 -1651 -9438
rect -1593 -9438 -1473 -9400
rect -1593 -9454 -1555 -9438
rect -1689 -9472 -1673 -9454
rect -1749 -9488 -1673 -9472
rect -1571 -9472 -1555 -9454
rect -1511 -9454 -1473 -9438
rect -1415 -9438 -1295 -9400
rect -1415 -9454 -1377 -9438
rect -1511 -9472 -1495 -9454
rect -1571 -9488 -1495 -9472
rect -1393 -9472 -1377 -9454
rect -1333 -9454 -1295 -9438
rect -1237 -9438 -1117 -9400
rect -1237 -9454 -1199 -9438
rect -1333 -9472 -1317 -9454
rect -1393 -9488 -1317 -9472
rect -1215 -9472 -1199 -9454
rect -1155 -9454 -1117 -9438
rect -1059 -9438 -939 -9400
rect -1059 -9454 -1021 -9438
rect -1155 -9472 -1139 -9454
rect -1215 -9488 -1139 -9472
rect -1037 -9472 -1021 -9454
rect -977 -9454 -939 -9438
rect -881 -9438 -761 -9400
rect -881 -9454 -843 -9438
rect -977 -9472 -961 -9454
rect -1037 -9488 -961 -9472
rect -859 -9472 -843 -9454
rect -799 -9454 -761 -9438
rect -703 -9438 -583 -9400
rect -703 -9454 -665 -9438
rect -799 -9472 -783 -9454
rect -859 -9488 -783 -9472
rect -681 -9472 -665 -9454
rect -621 -9454 -583 -9438
rect -525 -9438 -405 -9400
rect -525 -9454 -487 -9438
rect -621 -9472 -605 -9454
rect -681 -9488 -605 -9472
rect -503 -9472 -487 -9454
rect -443 -9454 -405 -9438
rect -347 -9438 -227 -9400
rect -347 -9454 -309 -9438
rect -443 -9472 -427 -9454
rect -503 -9488 -427 -9472
rect -325 -9472 -309 -9454
rect -265 -9454 -227 -9438
rect -169 -9438 -49 -9400
rect -169 -9454 -131 -9438
rect -265 -9472 -249 -9454
rect -325 -9488 -249 -9472
rect -147 -9472 -131 -9454
rect -87 -9454 -49 -9438
rect 9 -9438 129 -9400
rect 9 -9454 47 -9438
rect -87 -9472 -71 -9454
rect -147 -9488 -71 -9472
rect 31 -9472 47 -9454
rect 91 -9454 129 -9438
rect 187 -9438 307 -9400
rect 187 -9454 225 -9438
rect 91 -9472 107 -9454
rect 31 -9488 107 -9472
rect 209 -9472 225 -9454
rect 269 -9454 307 -9438
rect 365 -9438 485 -9400
rect 365 -9454 403 -9438
rect 269 -9472 285 -9454
rect 209 -9488 285 -9472
rect 387 -9472 403 -9454
rect 447 -9454 485 -9438
rect 543 -9438 663 -9400
rect 543 -9454 581 -9438
rect 447 -9472 463 -9454
rect 387 -9488 463 -9472
rect 565 -9472 581 -9454
rect 625 -9454 663 -9438
rect 721 -9438 841 -9400
rect 721 -9454 759 -9438
rect 625 -9472 641 -9454
rect 565 -9488 641 -9472
rect 743 -9472 759 -9454
rect 803 -9454 841 -9438
rect 899 -9438 1019 -9400
rect 899 -9454 937 -9438
rect 803 -9472 819 -9454
rect 743 -9488 819 -9472
rect 921 -9472 937 -9454
rect 981 -9454 1019 -9438
rect 1077 -9438 1197 -9400
rect 1077 -9454 1115 -9438
rect 981 -9472 997 -9454
rect 921 -9488 997 -9472
rect 1099 -9472 1115 -9454
rect 1159 -9454 1197 -9438
rect 1255 -9438 1375 -9400
rect 1255 -9454 1293 -9438
rect 1159 -9472 1175 -9454
rect 1099 -9488 1175 -9472
rect 1277 -9472 1293 -9454
rect 1337 -9454 1375 -9438
rect 1433 -9438 1553 -9400
rect 1433 -9454 1471 -9438
rect 1337 -9472 1353 -9454
rect 1277 -9488 1353 -9472
rect 1455 -9472 1471 -9454
rect 1515 -9454 1553 -9438
rect 1611 -9438 1731 -9400
rect 1611 -9454 1649 -9438
rect 1515 -9472 1531 -9454
rect 1455 -9488 1531 -9472
rect 1633 -9472 1649 -9454
rect 1693 -9454 1731 -9438
rect 1789 -9438 1909 -9400
rect 1789 -9454 1827 -9438
rect 1693 -9472 1709 -9454
rect 1633 -9488 1709 -9472
rect 1811 -9472 1827 -9454
rect 1871 -9454 1909 -9438
rect 1967 -9438 2087 -9400
rect 1967 -9454 2005 -9438
rect 1871 -9472 1887 -9454
rect 1811 -9488 1887 -9472
rect 1989 -9472 2005 -9454
rect 2049 -9454 2087 -9438
rect 2145 -9438 2265 -9400
rect 2145 -9454 2183 -9438
rect 2049 -9472 2065 -9454
rect 1989 -9488 2065 -9472
rect 2167 -9472 2183 -9454
rect 2227 -9454 2265 -9438
rect 2323 -9438 2443 -9400
rect 2323 -9454 2361 -9438
rect 2227 -9472 2243 -9454
rect 2167 -9488 2243 -9472
rect 2345 -9472 2361 -9454
rect 2405 -9454 2443 -9438
rect 2501 -9438 2621 -9400
rect 2501 -9454 2539 -9438
rect 2405 -9472 2421 -9454
rect 2345 -9488 2421 -9472
rect 2523 -9472 2539 -9454
rect 2583 -9454 2621 -9438
rect 2679 -9438 2799 -9400
rect 2679 -9454 2717 -9438
rect 2583 -9472 2599 -9454
rect 2523 -9488 2599 -9472
rect 2701 -9472 2717 -9454
rect 2761 -9454 2799 -9438
rect 2857 -9438 2977 -9400
rect 2857 -9454 2895 -9438
rect 2761 -9472 2777 -9454
rect 2701 -9488 2777 -9472
rect 2879 -9472 2895 -9454
rect 2939 -9454 2977 -9438
rect 3035 -9438 3155 -9400
rect 3035 -9454 3073 -9438
rect 2939 -9472 2955 -9454
rect 2879 -9488 2955 -9472
rect 3057 -9472 3073 -9454
rect 3117 -9454 3155 -9438
rect 3213 -9438 3333 -9400
rect 3213 -9454 3251 -9438
rect 3117 -9472 3133 -9454
rect 3057 -9488 3133 -9472
rect 3235 -9472 3251 -9454
rect 3295 -9454 3333 -9438
rect 3391 -9438 3511 -9400
rect 3391 -9454 3429 -9438
rect 3295 -9472 3311 -9454
rect 3235 -9488 3311 -9472
rect 3413 -9472 3429 -9454
rect 3473 -9454 3511 -9438
rect 3569 -9438 3689 -9400
rect 3569 -9454 3607 -9438
rect 3473 -9472 3489 -9454
rect 3413 -9488 3489 -9472
rect 3591 -9472 3607 -9454
rect 3651 -9454 3689 -9438
rect 3747 -9438 3867 -9400
rect 3747 -9454 3785 -9438
rect 3651 -9472 3667 -9454
rect 3591 -9488 3667 -9472
rect 3769 -9472 3785 -9454
rect 3829 -9454 3867 -9438
rect 3925 -9438 4045 -9400
rect 3925 -9454 3963 -9438
rect 3829 -9472 3845 -9454
rect 3769 -9488 3845 -9472
rect 3947 -9472 3963 -9454
rect 4007 -9454 4045 -9438
rect 4007 -9472 4023 -9454
rect 3947 -9488 4023 -9472
rect 10840 -9610 10916 -9594
rect 10840 -9628 10856 -9610
rect 10818 -9644 10856 -9628
rect 10900 -9628 10916 -9610
rect 11132 -9610 11208 -9594
rect 11132 -9628 11148 -9610
rect 10900 -9644 10938 -9628
rect 10818 -9682 10938 -9644
rect 11110 -9644 11148 -9628
rect 11192 -9628 11208 -9610
rect 11424 -9610 11500 -9594
rect 11424 -9628 11440 -9610
rect 11192 -9644 11230 -9628
rect 11110 -9682 11230 -9644
rect 11402 -9644 11440 -9628
rect 11484 -9628 11500 -9610
rect 11716 -9610 11792 -9594
rect 11716 -9628 11732 -9610
rect 11484 -9644 11522 -9628
rect 11402 -9682 11522 -9644
rect 11694 -9644 11732 -9628
rect 11776 -9628 11792 -9610
rect 12008 -9610 12084 -9594
rect 12008 -9628 12024 -9610
rect 11776 -9644 11814 -9628
rect 11694 -9682 11814 -9644
rect 11986 -9644 12024 -9628
rect 12068 -9628 12084 -9610
rect 12300 -9610 12376 -9594
rect 12300 -9628 12316 -9610
rect 12068 -9644 12106 -9628
rect 11986 -9682 12106 -9644
rect 12278 -9644 12316 -9628
rect 12360 -9628 12376 -9610
rect 12592 -9610 12668 -9594
rect 12592 -9628 12608 -9610
rect 12360 -9644 12398 -9628
rect 12278 -9682 12398 -9644
rect 12570 -9644 12608 -9628
rect 12652 -9628 12668 -9610
rect 12652 -9644 12690 -9628
rect 12570 -9682 12690 -9644
rect 6580 -9710 6656 -9694
rect 6580 -9728 6596 -9710
rect 6558 -9744 6596 -9728
rect 6640 -9728 6656 -9710
rect 6758 -9710 6834 -9694
rect 6758 -9728 6774 -9710
rect 6640 -9744 6678 -9728
rect 6558 -9782 6678 -9744
rect 6736 -9744 6774 -9728
rect 6818 -9728 6834 -9710
rect 6936 -9710 7012 -9694
rect 6936 -9728 6952 -9710
rect 6818 -9744 6856 -9728
rect 6736 -9782 6856 -9744
rect 6914 -9744 6952 -9728
rect 6996 -9728 7012 -9710
rect 7114 -9710 7190 -9694
rect 7114 -9728 7130 -9710
rect 6996 -9744 7034 -9728
rect 6914 -9782 7034 -9744
rect 7092 -9744 7130 -9728
rect 7174 -9728 7190 -9710
rect 7292 -9710 7368 -9694
rect 7292 -9728 7308 -9710
rect 7174 -9744 7212 -9728
rect 7092 -9782 7212 -9744
rect 7270 -9744 7308 -9728
rect 7352 -9728 7368 -9710
rect 7470 -9710 7546 -9694
rect 7470 -9728 7486 -9710
rect 7352 -9744 7390 -9728
rect 7270 -9782 7390 -9744
rect 7448 -9744 7486 -9728
rect 7530 -9728 7546 -9710
rect 7648 -9710 7724 -9694
rect 7648 -9728 7664 -9710
rect 7530 -9744 7568 -9728
rect 7448 -9782 7568 -9744
rect 7626 -9744 7664 -9728
rect 7708 -9728 7724 -9710
rect 7826 -9710 7902 -9694
rect 7826 -9728 7842 -9710
rect 7708 -9744 7746 -9728
rect 7626 -9782 7746 -9744
rect 7804 -9744 7842 -9728
rect 7886 -9728 7902 -9710
rect 8004 -9710 8080 -9694
rect 8004 -9728 8020 -9710
rect 7886 -9744 7924 -9728
rect 7804 -9782 7924 -9744
rect 7982 -9744 8020 -9728
rect 8064 -9728 8080 -9710
rect 8182 -9710 8258 -9694
rect 8182 -9728 8198 -9710
rect 8064 -9744 8102 -9728
rect 7982 -9782 8102 -9744
rect 8160 -9744 8198 -9728
rect 8242 -9728 8258 -9710
rect 8360 -9710 8436 -9694
rect 8360 -9728 8376 -9710
rect 8242 -9744 8280 -9728
rect 8160 -9782 8280 -9744
rect 8338 -9744 8376 -9728
rect 8420 -9728 8436 -9710
rect 8538 -9710 8614 -9694
rect 8538 -9728 8554 -9710
rect 8420 -9744 8458 -9728
rect 8338 -9782 8458 -9744
rect 8516 -9744 8554 -9728
rect 8598 -9728 8614 -9710
rect 8716 -9710 8792 -9694
rect 8716 -9728 8732 -9710
rect 8598 -9744 8636 -9728
rect 8516 -9782 8636 -9744
rect 8694 -9744 8732 -9728
rect 8776 -9728 8792 -9710
rect 8894 -9710 8970 -9694
rect 8894 -9728 8910 -9710
rect 8776 -9744 8814 -9728
rect 8694 -9782 8814 -9744
rect 8872 -9744 8910 -9728
rect 8954 -9728 8970 -9710
rect 9072 -9710 9148 -9694
rect 9072 -9728 9088 -9710
rect 8954 -9744 8992 -9728
rect 8872 -9782 8992 -9744
rect 9050 -9744 9088 -9728
rect 9132 -9728 9148 -9710
rect 9250 -9710 9326 -9694
rect 9250 -9728 9266 -9710
rect 9132 -9744 9170 -9728
rect 9050 -9782 9170 -9744
rect 9228 -9744 9266 -9728
rect 9310 -9728 9326 -9710
rect 9310 -9744 9348 -9728
rect 9228 -9782 9348 -9744
rect -5582 -9830 -5462 -9792
rect -5582 -9846 -5544 -9830
rect -5560 -9864 -5544 -9846
rect -5500 -9846 -5462 -9830
rect -5404 -9830 -5284 -9792
rect -5404 -9846 -5366 -9830
rect -5500 -9864 -5484 -9846
rect -5560 -9880 -5484 -9864
rect -5382 -9864 -5366 -9846
rect -5322 -9846 -5284 -9830
rect -5226 -9830 -5106 -9792
rect -5226 -9846 -5188 -9830
rect -5322 -9864 -5306 -9846
rect -5382 -9880 -5306 -9864
rect -5204 -9864 -5188 -9846
rect -5144 -9846 -5106 -9830
rect -5048 -9830 -4928 -9792
rect -5048 -9846 -5010 -9830
rect -5144 -9864 -5128 -9846
rect -5204 -9880 -5128 -9864
rect -5026 -9864 -5010 -9846
rect -4966 -9846 -4928 -9830
rect -4870 -9830 -4750 -9792
rect -4870 -9846 -4832 -9830
rect -4966 -9864 -4950 -9846
rect -5026 -9880 -4950 -9864
rect -4848 -9864 -4832 -9846
rect -4788 -9846 -4750 -9830
rect -4692 -9830 -4572 -9792
rect -4692 -9846 -4654 -9830
rect -4788 -9864 -4772 -9846
rect -4848 -9880 -4772 -9864
rect -4670 -9864 -4654 -9846
rect -4610 -9846 -4572 -9830
rect -4514 -9830 -4394 -9792
rect -4514 -9846 -4476 -9830
rect -4610 -9864 -4594 -9846
rect -4670 -9880 -4594 -9864
rect -4492 -9864 -4476 -9846
rect -4432 -9846 -4394 -9830
rect -4336 -9830 -4216 -9792
rect -4336 -9846 -4298 -9830
rect -4432 -9864 -4416 -9846
rect -4492 -9880 -4416 -9864
rect -4314 -9864 -4298 -9846
rect -4254 -9846 -4216 -9830
rect -4158 -9830 -4038 -9792
rect -4158 -9846 -4120 -9830
rect -4254 -9864 -4238 -9846
rect -4314 -9880 -4238 -9864
rect -4136 -9864 -4120 -9846
rect -4076 -9846 -4038 -9830
rect -4076 -9864 -4060 -9846
rect -4136 -9880 -4060 -9864
rect -5560 -9990 -5484 -9974
rect -5560 -10008 -5544 -9990
rect -5582 -10024 -5544 -10008
rect -5500 -10008 -5484 -9990
rect -5382 -9990 -5306 -9974
rect -5382 -10008 -5366 -9990
rect -5500 -10024 -5462 -10008
rect -5582 -10062 -5462 -10024
rect -5404 -10024 -5366 -10008
rect -5322 -10008 -5306 -9990
rect -5204 -9990 -5128 -9974
rect -5204 -10008 -5188 -9990
rect -5322 -10024 -5284 -10008
rect -5404 -10062 -5284 -10024
rect -5226 -10024 -5188 -10008
rect -5144 -10008 -5128 -9990
rect -5026 -9990 -4950 -9974
rect -5026 -10008 -5010 -9990
rect -5144 -10024 -5106 -10008
rect -5226 -10062 -5106 -10024
rect -5048 -10024 -5010 -10008
rect -4966 -10008 -4950 -9990
rect -4848 -9990 -4772 -9974
rect -4848 -10008 -4832 -9990
rect -4966 -10024 -4928 -10008
rect -5048 -10062 -4928 -10024
rect -4870 -10024 -4832 -10008
rect -4788 -10008 -4772 -9990
rect -4670 -9990 -4594 -9974
rect -4670 -10008 -4654 -9990
rect -4788 -10024 -4750 -10008
rect -4870 -10062 -4750 -10024
rect -4692 -10024 -4654 -10008
rect -4610 -10008 -4594 -9990
rect -4492 -9990 -4416 -9974
rect -4492 -10008 -4476 -9990
rect -4610 -10024 -4572 -10008
rect -4692 -10062 -4572 -10024
rect -4514 -10024 -4476 -10008
rect -4432 -10008 -4416 -9990
rect -4314 -9990 -4238 -9974
rect -4314 -10008 -4298 -9990
rect -4432 -10024 -4394 -10008
rect -4514 -10062 -4394 -10024
rect -4336 -10024 -4298 -10008
rect -4254 -10008 -4238 -9990
rect -4136 -9990 -4060 -9974
rect -4136 -10008 -4120 -9990
rect -4254 -10024 -4216 -10008
rect -4336 -10062 -4216 -10024
rect -4158 -10024 -4120 -10008
rect -4076 -10008 -4060 -9990
rect -4076 -10024 -4038 -10008
rect -4158 -10062 -4038 -10024
rect -2105 -10048 -2029 -10032
rect -2105 -10066 -2089 -10048
rect -2127 -10082 -2089 -10066
rect -2045 -10066 -2029 -10048
rect -1927 -10048 -1851 -10032
rect -1927 -10066 -1911 -10048
rect -2045 -10082 -2007 -10066
rect -2127 -10120 -2007 -10082
rect -1949 -10082 -1911 -10066
rect -1867 -10066 -1851 -10048
rect -1749 -10048 -1673 -10032
rect -1749 -10066 -1733 -10048
rect -1867 -10082 -1829 -10066
rect -1949 -10120 -1829 -10082
rect -1771 -10082 -1733 -10066
rect -1689 -10066 -1673 -10048
rect -1571 -10048 -1495 -10032
rect -1571 -10066 -1555 -10048
rect -1689 -10082 -1651 -10066
rect -1771 -10120 -1651 -10082
rect -1593 -10082 -1555 -10066
rect -1511 -10066 -1495 -10048
rect -1393 -10048 -1317 -10032
rect -1393 -10066 -1377 -10048
rect -1511 -10082 -1473 -10066
rect -1593 -10120 -1473 -10082
rect -1415 -10082 -1377 -10066
rect -1333 -10066 -1317 -10048
rect -1215 -10048 -1139 -10032
rect -1215 -10066 -1199 -10048
rect -1333 -10082 -1295 -10066
rect -1415 -10120 -1295 -10082
rect -1237 -10082 -1199 -10066
rect -1155 -10066 -1139 -10048
rect -1037 -10048 -961 -10032
rect -1037 -10066 -1021 -10048
rect -1155 -10082 -1117 -10066
rect -1237 -10120 -1117 -10082
rect -1059 -10082 -1021 -10066
rect -977 -10066 -961 -10048
rect -859 -10048 -783 -10032
rect -859 -10066 -843 -10048
rect -977 -10082 -939 -10066
rect -1059 -10120 -939 -10082
rect -881 -10082 -843 -10066
rect -799 -10066 -783 -10048
rect -681 -10048 -605 -10032
rect -681 -10066 -665 -10048
rect -799 -10082 -761 -10066
rect -881 -10120 -761 -10082
rect -703 -10082 -665 -10066
rect -621 -10066 -605 -10048
rect -503 -10048 -427 -10032
rect -503 -10066 -487 -10048
rect -621 -10082 -583 -10066
rect -703 -10120 -583 -10082
rect -525 -10082 -487 -10066
rect -443 -10066 -427 -10048
rect -325 -10048 -249 -10032
rect -325 -10066 -309 -10048
rect -443 -10082 -405 -10066
rect -525 -10120 -405 -10082
rect -347 -10082 -309 -10066
rect -265 -10066 -249 -10048
rect -147 -10048 -71 -10032
rect -147 -10066 -131 -10048
rect -265 -10082 -227 -10066
rect -347 -10120 -227 -10082
rect -169 -10082 -131 -10066
rect -87 -10066 -71 -10048
rect 31 -10048 107 -10032
rect 31 -10066 47 -10048
rect -87 -10082 -49 -10066
rect -169 -10120 -49 -10082
rect 9 -10082 47 -10066
rect 91 -10066 107 -10048
rect 209 -10048 285 -10032
rect 209 -10066 225 -10048
rect 91 -10082 129 -10066
rect 9 -10120 129 -10082
rect 187 -10082 225 -10066
rect 269 -10066 285 -10048
rect 387 -10048 463 -10032
rect 387 -10066 403 -10048
rect 269 -10082 307 -10066
rect 187 -10120 307 -10082
rect 365 -10082 403 -10066
rect 447 -10066 463 -10048
rect 565 -10048 641 -10032
rect 565 -10066 581 -10048
rect 447 -10082 485 -10066
rect 365 -10120 485 -10082
rect 543 -10082 581 -10066
rect 625 -10066 641 -10048
rect 743 -10048 819 -10032
rect 743 -10066 759 -10048
rect 625 -10082 663 -10066
rect 543 -10120 663 -10082
rect 721 -10082 759 -10066
rect 803 -10066 819 -10048
rect 921 -10048 997 -10032
rect 921 -10066 937 -10048
rect 803 -10082 841 -10066
rect 721 -10120 841 -10082
rect 899 -10082 937 -10066
rect 981 -10066 997 -10048
rect 1099 -10048 1175 -10032
rect 1099 -10066 1115 -10048
rect 981 -10082 1019 -10066
rect 899 -10120 1019 -10082
rect 1077 -10082 1115 -10066
rect 1159 -10066 1175 -10048
rect 1277 -10048 1353 -10032
rect 1277 -10066 1293 -10048
rect 1159 -10082 1197 -10066
rect 1077 -10120 1197 -10082
rect 1255 -10082 1293 -10066
rect 1337 -10066 1353 -10048
rect 1455 -10048 1531 -10032
rect 1455 -10066 1471 -10048
rect 1337 -10082 1375 -10066
rect 1255 -10120 1375 -10082
rect 1433 -10082 1471 -10066
rect 1515 -10066 1531 -10048
rect 1633 -10048 1709 -10032
rect 1633 -10066 1649 -10048
rect 1515 -10082 1553 -10066
rect 1433 -10120 1553 -10082
rect 1611 -10082 1649 -10066
rect 1693 -10066 1709 -10048
rect 1811 -10048 1887 -10032
rect 1811 -10066 1827 -10048
rect 1693 -10082 1731 -10066
rect 1611 -10120 1731 -10082
rect 1789 -10082 1827 -10066
rect 1871 -10066 1887 -10048
rect 1989 -10048 2065 -10032
rect 1989 -10066 2005 -10048
rect 1871 -10082 1909 -10066
rect 1789 -10120 1909 -10082
rect 1967 -10082 2005 -10066
rect 2049 -10066 2065 -10048
rect 2167 -10048 2243 -10032
rect 2167 -10066 2183 -10048
rect 2049 -10082 2087 -10066
rect 1967 -10120 2087 -10082
rect 2145 -10082 2183 -10066
rect 2227 -10066 2243 -10048
rect 2345 -10048 2421 -10032
rect 2345 -10066 2361 -10048
rect 2227 -10082 2265 -10066
rect 2145 -10120 2265 -10082
rect 2323 -10082 2361 -10066
rect 2405 -10066 2421 -10048
rect 2523 -10048 2599 -10032
rect 2523 -10066 2539 -10048
rect 2405 -10082 2443 -10066
rect 2323 -10120 2443 -10082
rect 2501 -10082 2539 -10066
rect 2583 -10066 2599 -10048
rect 2701 -10048 2777 -10032
rect 2701 -10066 2717 -10048
rect 2583 -10082 2621 -10066
rect 2501 -10120 2621 -10082
rect 2679 -10082 2717 -10066
rect 2761 -10066 2777 -10048
rect 2879 -10048 2955 -10032
rect 2879 -10066 2895 -10048
rect 2761 -10082 2799 -10066
rect 2679 -10120 2799 -10082
rect 2857 -10082 2895 -10066
rect 2939 -10066 2955 -10048
rect 3057 -10048 3133 -10032
rect 3057 -10066 3073 -10048
rect 2939 -10082 2977 -10066
rect 2857 -10120 2977 -10082
rect 3035 -10082 3073 -10066
rect 3117 -10066 3133 -10048
rect 3235 -10048 3311 -10032
rect 3235 -10066 3251 -10048
rect 3117 -10082 3155 -10066
rect 3035 -10120 3155 -10082
rect 3213 -10082 3251 -10066
rect 3295 -10066 3311 -10048
rect 3413 -10048 3489 -10032
rect 3413 -10066 3429 -10048
rect 3295 -10082 3333 -10066
rect 3213 -10120 3333 -10082
rect 3391 -10082 3429 -10066
rect 3473 -10066 3489 -10048
rect 3591 -10048 3667 -10032
rect 3591 -10066 3607 -10048
rect 3473 -10082 3511 -10066
rect 3391 -10120 3511 -10082
rect 3569 -10082 3607 -10066
rect 3651 -10066 3667 -10048
rect 3769 -10048 3845 -10032
rect 3769 -10066 3785 -10048
rect 3651 -10082 3689 -10066
rect 3569 -10120 3689 -10082
rect 3747 -10082 3785 -10066
rect 3829 -10066 3845 -10048
rect 3947 -10048 4023 -10032
rect 3947 -10066 3963 -10048
rect 3829 -10082 3867 -10066
rect 3747 -10120 3867 -10082
rect 3925 -10082 3963 -10066
rect 4007 -10066 4023 -10048
rect 10818 -10000 10938 -9962
rect 10818 -10016 10856 -10000
rect 10840 -10034 10856 -10016
rect 10900 -10016 10938 -10000
rect 11110 -10000 11230 -9962
rect 11110 -10016 11148 -10000
rect 10900 -10034 10916 -10016
rect 10840 -10050 10916 -10034
rect 11132 -10034 11148 -10016
rect 11192 -10016 11230 -10000
rect 11402 -10000 11522 -9962
rect 11402 -10016 11440 -10000
rect 11192 -10034 11208 -10016
rect 11132 -10050 11208 -10034
rect 11424 -10034 11440 -10016
rect 11484 -10016 11522 -10000
rect 11694 -10000 11814 -9962
rect 11694 -10016 11732 -10000
rect 11484 -10034 11500 -10016
rect 11424 -10050 11500 -10034
rect 11716 -10034 11732 -10016
rect 11776 -10016 11814 -10000
rect 11986 -10000 12106 -9962
rect 11986 -10016 12024 -10000
rect 11776 -10034 11792 -10016
rect 11716 -10050 11792 -10034
rect 12008 -10034 12024 -10016
rect 12068 -10016 12106 -10000
rect 12278 -10000 12398 -9962
rect 12278 -10016 12316 -10000
rect 12068 -10034 12084 -10016
rect 12008 -10050 12084 -10034
rect 12300 -10034 12316 -10016
rect 12360 -10016 12398 -10000
rect 12570 -10000 12690 -9962
rect 12570 -10016 12608 -10000
rect 12360 -10034 12376 -10016
rect 12300 -10050 12376 -10034
rect 12592 -10034 12608 -10016
rect 12652 -10016 12690 -10000
rect 12652 -10034 12668 -10016
rect 12592 -10050 12668 -10034
rect 4007 -10082 4045 -10066
rect 3925 -10120 4045 -10082
rect 6558 -10100 6678 -10062
rect 6558 -10116 6596 -10100
rect -5582 -10380 -5462 -10342
rect -5582 -10396 -5544 -10380
rect -5560 -10414 -5544 -10396
rect -5500 -10396 -5462 -10380
rect -5404 -10380 -5284 -10342
rect -5404 -10396 -5366 -10380
rect -5500 -10414 -5484 -10396
rect -5560 -10430 -5484 -10414
rect -5382 -10414 -5366 -10396
rect -5322 -10396 -5284 -10380
rect -5226 -10380 -5106 -10342
rect -5226 -10396 -5188 -10380
rect -5322 -10414 -5306 -10396
rect -5382 -10430 -5306 -10414
rect -5204 -10414 -5188 -10396
rect -5144 -10396 -5106 -10380
rect -5048 -10380 -4928 -10342
rect -5048 -10396 -5010 -10380
rect -5144 -10414 -5128 -10396
rect -5204 -10430 -5128 -10414
rect -5026 -10414 -5010 -10396
rect -4966 -10396 -4928 -10380
rect -4870 -10380 -4750 -10342
rect -4870 -10396 -4832 -10380
rect -4966 -10414 -4950 -10396
rect -5026 -10430 -4950 -10414
rect -4848 -10414 -4832 -10396
rect -4788 -10396 -4750 -10380
rect -4692 -10380 -4572 -10342
rect -4692 -10396 -4654 -10380
rect -4788 -10414 -4772 -10396
rect -4848 -10430 -4772 -10414
rect -4670 -10414 -4654 -10396
rect -4610 -10396 -4572 -10380
rect -4514 -10380 -4394 -10342
rect -4514 -10396 -4476 -10380
rect -4610 -10414 -4594 -10396
rect -4670 -10430 -4594 -10414
rect -4492 -10414 -4476 -10396
rect -4432 -10396 -4394 -10380
rect -4336 -10380 -4216 -10342
rect -4336 -10396 -4298 -10380
rect -4432 -10414 -4416 -10396
rect -4492 -10430 -4416 -10414
rect -4314 -10414 -4298 -10396
rect -4254 -10396 -4216 -10380
rect -4158 -10380 -4038 -10342
rect -4158 -10396 -4120 -10380
rect -4254 -10414 -4238 -10396
rect -4314 -10430 -4238 -10414
rect -4136 -10414 -4120 -10396
rect -4076 -10396 -4038 -10380
rect -4076 -10414 -4060 -10396
rect 6580 -10134 6596 -10116
rect 6640 -10116 6678 -10100
rect 6736 -10100 6856 -10062
rect 6736 -10116 6774 -10100
rect 6640 -10134 6656 -10116
rect 6580 -10150 6656 -10134
rect 6758 -10134 6774 -10116
rect 6818 -10116 6856 -10100
rect 6914 -10100 7034 -10062
rect 6914 -10116 6952 -10100
rect 6818 -10134 6834 -10116
rect 6758 -10150 6834 -10134
rect 6936 -10134 6952 -10116
rect 6996 -10116 7034 -10100
rect 7092 -10100 7212 -10062
rect 7092 -10116 7130 -10100
rect 6996 -10134 7012 -10116
rect 6936 -10150 7012 -10134
rect 7114 -10134 7130 -10116
rect 7174 -10116 7212 -10100
rect 7270 -10100 7390 -10062
rect 7270 -10116 7308 -10100
rect 7174 -10134 7190 -10116
rect 7114 -10150 7190 -10134
rect 7292 -10134 7308 -10116
rect 7352 -10116 7390 -10100
rect 7448 -10100 7568 -10062
rect 7448 -10116 7486 -10100
rect 7352 -10134 7368 -10116
rect 7292 -10150 7368 -10134
rect 7470 -10134 7486 -10116
rect 7530 -10116 7568 -10100
rect 7626 -10100 7746 -10062
rect 7626 -10116 7664 -10100
rect 7530 -10134 7546 -10116
rect 7470 -10150 7546 -10134
rect 7648 -10134 7664 -10116
rect 7708 -10116 7746 -10100
rect 7804 -10100 7924 -10062
rect 7804 -10116 7842 -10100
rect 7708 -10134 7724 -10116
rect 7648 -10150 7724 -10134
rect 7826 -10134 7842 -10116
rect 7886 -10116 7924 -10100
rect 7982 -10100 8102 -10062
rect 7982 -10116 8020 -10100
rect 7886 -10134 7902 -10116
rect 7826 -10150 7902 -10134
rect 8004 -10134 8020 -10116
rect 8064 -10116 8102 -10100
rect 8160 -10100 8280 -10062
rect 8160 -10116 8198 -10100
rect 8064 -10134 8080 -10116
rect 8004 -10150 8080 -10134
rect 8182 -10134 8198 -10116
rect 8242 -10116 8280 -10100
rect 8338 -10100 8458 -10062
rect 8338 -10116 8376 -10100
rect 8242 -10134 8258 -10116
rect 8182 -10150 8258 -10134
rect 8360 -10134 8376 -10116
rect 8420 -10116 8458 -10100
rect 8516 -10100 8636 -10062
rect 8516 -10116 8554 -10100
rect 8420 -10134 8436 -10116
rect 8360 -10150 8436 -10134
rect 8538 -10134 8554 -10116
rect 8598 -10116 8636 -10100
rect 8694 -10100 8814 -10062
rect 8694 -10116 8732 -10100
rect 8598 -10134 8614 -10116
rect 8538 -10150 8614 -10134
rect 8716 -10134 8732 -10116
rect 8776 -10116 8814 -10100
rect 8872 -10100 8992 -10062
rect 8872 -10116 8910 -10100
rect 8776 -10134 8792 -10116
rect 8716 -10150 8792 -10134
rect 8894 -10134 8910 -10116
rect 8954 -10116 8992 -10100
rect 9050 -10100 9170 -10062
rect 9050 -10116 9088 -10100
rect 8954 -10134 8970 -10116
rect 8894 -10150 8970 -10134
rect 9072 -10134 9088 -10116
rect 9132 -10116 9170 -10100
rect 9228 -10100 9348 -10062
rect 9228 -10116 9266 -10100
rect 9132 -10134 9148 -10116
rect 9072 -10150 9148 -10134
rect 9250 -10134 9266 -10116
rect 9310 -10116 9348 -10100
rect 9310 -10134 9326 -10116
rect 9250 -10150 9326 -10134
rect 10840 -10380 10916 -10364
rect 10840 -10398 10856 -10380
rect -4136 -10430 -4060 -10414
rect -2127 -10438 -2007 -10400
rect -2127 -10454 -2089 -10438
rect -2105 -10472 -2089 -10454
rect -2045 -10454 -2007 -10438
rect -1949 -10438 -1829 -10400
rect -1949 -10454 -1911 -10438
rect -2045 -10472 -2029 -10454
rect -2105 -10488 -2029 -10472
rect -1927 -10472 -1911 -10454
rect -1867 -10454 -1829 -10438
rect -1771 -10438 -1651 -10400
rect -1771 -10454 -1733 -10438
rect -1867 -10472 -1851 -10454
rect -1927 -10488 -1851 -10472
rect -1749 -10472 -1733 -10454
rect -1689 -10454 -1651 -10438
rect -1593 -10438 -1473 -10400
rect -1593 -10454 -1555 -10438
rect -1689 -10472 -1673 -10454
rect -1749 -10488 -1673 -10472
rect -1571 -10472 -1555 -10454
rect -1511 -10454 -1473 -10438
rect -1415 -10438 -1295 -10400
rect -1415 -10454 -1377 -10438
rect -1511 -10472 -1495 -10454
rect -1571 -10488 -1495 -10472
rect -1393 -10472 -1377 -10454
rect -1333 -10454 -1295 -10438
rect -1237 -10438 -1117 -10400
rect -1237 -10454 -1199 -10438
rect -1333 -10472 -1317 -10454
rect -1393 -10488 -1317 -10472
rect -1215 -10472 -1199 -10454
rect -1155 -10454 -1117 -10438
rect -1059 -10438 -939 -10400
rect -1059 -10454 -1021 -10438
rect -1155 -10472 -1139 -10454
rect -1215 -10488 -1139 -10472
rect -1037 -10472 -1021 -10454
rect -977 -10454 -939 -10438
rect -881 -10438 -761 -10400
rect -881 -10454 -843 -10438
rect -977 -10472 -961 -10454
rect -1037 -10488 -961 -10472
rect -859 -10472 -843 -10454
rect -799 -10454 -761 -10438
rect -703 -10438 -583 -10400
rect -703 -10454 -665 -10438
rect -799 -10472 -783 -10454
rect -859 -10488 -783 -10472
rect -681 -10472 -665 -10454
rect -621 -10454 -583 -10438
rect -525 -10438 -405 -10400
rect -525 -10454 -487 -10438
rect -621 -10472 -605 -10454
rect -681 -10488 -605 -10472
rect -503 -10472 -487 -10454
rect -443 -10454 -405 -10438
rect -347 -10438 -227 -10400
rect -347 -10454 -309 -10438
rect -443 -10472 -427 -10454
rect -503 -10488 -427 -10472
rect -325 -10472 -309 -10454
rect -265 -10454 -227 -10438
rect -169 -10438 -49 -10400
rect -169 -10454 -131 -10438
rect -265 -10472 -249 -10454
rect -325 -10488 -249 -10472
rect -147 -10472 -131 -10454
rect -87 -10454 -49 -10438
rect 9 -10438 129 -10400
rect 9 -10454 47 -10438
rect -87 -10472 -71 -10454
rect -147 -10488 -71 -10472
rect 31 -10472 47 -10454
rect 91 -10454 129 -10438
rect 187 -10438 307 -10400
rect 187 -10454 225 -10438
rect 91 -10472 107 -10454
rect 31 -10488 107 -10472
rect 209 -10472 225 -10454
rect 269 -10454 307 -10438
rect 365 -10438 485 -10400
rect 365 -10454 403 -10438
rect 269 -10472 285 -10454
rect 209 -10488 285 -10472
rect 387 -10472 403 -10454
rect 447 -10454 485 -10438
rect 543 -10438 663 -10400
rect 543 -10454 581 -10438
rect 447 -10472 463 -10454
rect 387 -10488 463 -10472
rect 565 -10472 581 -10454
rect 625 -10454 663 -10438
rect 721 -10438 841 -10400
rect 721 -10454 759 -10438
rect 625 -10472 641 -10454
rect 565 -10488 641 -10472
rect 743 -10472 759 -10454
rect 803 -10454 841 -10438
rect 899 -10438 1019 -10400
rect 899 -10454 937 -10438
rect 803 -10472 819 -10454
rect 743 -10488 819 -10472
rect 921 -10472 937 -10454
rect 981 -10454 1019 -10438
rect 1077 -10438 1197 -10400
rect 1077 -10454 1115 -10438
rect 981 -10472 997 -10454
rect 921 -10488 997 -10472
rect 1099 -10472 1115 -10454
rect 1159 -10454 1197 -10438
rect 1255 -10438 1375 -10400
rect 1255 -10454 1293 -10438
rect 1159 -10472 1175 -10454
rect 1099 -10488 1175 -10472
rect 1277 -10472 1293 -10454
rect 1337 -10454 1375 -10438
rect 1433 -10438 1553 -10400
rect 1433 -10454 1471 -10438
rect 1337 -10472 1353 -10454
rect 1277 -10488 1353 -10472
rect 1455 -10472 1471 -10454
rect 1515 -10454 1553 -10438
rect 1611 -10438 1731 -10400
rect 1611 -10454 1649 -10438
rect 1515 -10472 1531 -10454
rect 1455 -10488 1531 -10472
rect 1633 -10472 1649 -10454
rect 1693 -10454 1731 -10438
rect 1789 -10438 1909 -10400
rect 1789 -10454 1827 -10438
rect 1693 -10472 1709 -10454
rect 1633 -10488 1709 -10472
rect 1811 -10472 1827 -10454
rect 1871 -10454 1909 -10438
rect 1967 -10438 2087 -10400
rect 1967 -10454 2005 -10438
rect 1871 -10472 1887 -10454
rect 1811 -10488 1887 -10472
rect 1989 -10472 2005 -10454
rect 2049 -10454 2087 -10438
rect 2145 -10438 2265 -10400
rect 2145 -10454 2183 -10438
rect 2049 -10472 2065 -10454
rect 1989 -10488 2065 -10472
rect 2167 -10472 2183 -10454
rect 2227 -10454 2265 -10438
rect 2323 -10438 2443 -10400
rect 2323 -10454 2361 -10438
rect 2227 -10472 2243 -10454
rect 2167 -10488 2243 -10472
rect 2345 -10472 2361 -10454
rect 2405 -10454 2443 -10438
rect 2501 -10438 2621 -10400
rect 2501 -10454 2539 -10438
rect 2405 -10472 2421 -10454
rect 2345 -10488 2421 -10472
rect 2523 -10472 2539 -10454
rect 2583 -10454 2621 -10438
rect 2679 -10438 2799 -10400
rect 2679 -10454 2717 -10438
rect 2583 -10472 2599 -10454
rect 2523 -10488 2599 -10472
rect 2701 -10472 2717 -10454
rect 2761 -10454 2799 -10438
rect 2857 -10438 2977 -10400
rect 2857 -10454 2895 -10438
rect 2761 -10472 2777 -10454
rect 2701 -10488 2777 -10472
rect 2879 -10472 2895 -10454
rect 2939 -10454 2977 -10438
rect 3035 -10438 3155 -10400
rect 3035 -10454 3073 -10438
rect 2939 -10472 2955 -10454
rect 2879 -10488 2955 -10472
rect 3057 -10472 3073 -10454
rect 3117 -10454 3155 -10438
rect 3213 -10438 3333 -10400
rect 3213 -10454 3251 -10438
rect 3117 -10472 3133 -10454
rect 3057 -10488 3133 -10472
rect 3235 -10472 3251 -10454
rect 3295 -10454 3333 -10438
rect 3391 -10438 3511 -10400
rect 3391 -10454 3429 -10438
rect 3295 -10472 3311 -10454
rect 3235 -10488 3311 -10472
rect 3413 -10472 3429 -10454
rect 3473 -10454 3511 -10438
rect 3569 -10438 3689 -10400
rect 3569 -10454 3607 -10438
rect 3473 -10472 3489 -10454
rect 3413 -10488 3489 -10472
rect 3591 -10472 3607 -10454
rect 3651 -10454 3689 -10438
rect 3747 -10438 3867 -10400
rect 3747 -10454 3785 -10438
rect 3651 -10472 3667 -10454
rect 3591 -10488 3667 -10472
rect 3769 -10472 3785 -10454
rect 3829 -10454 3867 -10438
rect 3925 -10438 4045 -10400
rect 3925 -10454 3963 -10438
rect 3829 -10472 3845 -10454
rect 3769 -10488 3845 -10472
rect 3947 -10472 3963 -10454
rect 4007 -10454 4045 -10438
rect 10818 -10414 10856 -10398
rect 10900 -10398 10916 -10380
rect 11132 -10380 11208 -10364
rect 11132 -10398 11148 -10380
rect 10900 -10414 10938 -10398
rect 10818 -10452 10938 -10414
rect 11110 -10414 11148 -10398
rect 11192 -10398 11208 -10380
rect 11424 -10380 11500 -10364
rect 11424 -10398 11440 -10380
rect 11192 -10414 11230 -10398
rect 11110 -10452 11230 -10414
rect 11402 -10414 11440 -10398
rect 11484 -10398 11500 -10380
rect 11716 -10380 11792 -10364
rect 11716 -10398 11732 -10380
rect 11484 -10414 11522 -10398
rect 11402 -10452 11522 -10414
rect 11694 -10414 11732 -10398
rect 11776 -10398 11792 -10380
rect 12008 -10380 12084 -10364
rect 12008 -10398 12024 -10380
rect 11776 -10414 11814 -10398
rect 11694 -10452 11814 -10414
rect 11986 -10414 12024 -10398
rect 12068 -10398 12084 -10380
rect 12300 -10380 12376 -10364
rect 12300 -10398 12316 -10380
rect 12068 -10414 12106 -10398
rect 11986 -10452 12106 -10414
rect 12278 -10414 12316 -10398
rect 12360 -10398 12376 -10380
rect 12592 -10380 12668 -10364
rect 12592 -10398 12608 -10380
rect 12360 -10414 12398 -10398
rect 12278 -10452 12398 -10414
rect 12570 -10414 12608 -10398
rect 12652 -10398 12668 -10380
rect 12652 -10414 12690 -10398
rect 12570 -10452 12690 -10414
rect 4007 -10472 4023 -10454
rect 3947 -10488 4023 -10472
rect -5560 -10540 -5484 -10524
rect -5560 -10558 -5544 -10540
rect -5582 -10574 -5544 -10558
rect -5500 -10558 -5484 -10540
rect -5382 -10540 -5306 -10524
rect -5382 -10558 -5366 -10540
rect -5500 -10574 -5462 -10558
rect -5582 -10612 -5462 -10574
rect -5404 -10574 -5366 -10558
rect -5322 -10558 -5306 -10540
rect -5204 -10540 -5128 -10524
rect -5204 -10558 -5188 -10540
rect -5322 -10574 -5284 -10558
rect -5404 -10612 -5284 -10574
rect -5226 -10574 -5188 -10558
rect -5144 -10558 -5128 -10540
rect -5026 -10540 -4950 -10524
rect -5026 -10558 -5010 -10540
rect -5144 -10574 -5106 -10558
rect -5226 -10612 -5106 -10574
rect -5048 -10574 -5010 -10558
rect -4966 -10558 -4950 -10540
rect -4848 -10540 -4772 -10524
rect -4848 -10558 -4832 -10540
rect -4966 -10574 -4928 -10558
rect -5048 -10612 -4928 -10574
rect -4870 -10574 -4832 -10558
rect -4788 -10558 -4772 -10540
rect -4670 -10540 -4594 -10524
rect -4670 -10558 -4654 -10540
rect -4788 -10574 -4750 -10558
rect -4870 -10612 -4750 -10574
rect -4692 -10574 -4654 -10558
rect -4610 -10558 -4594 -10540
rect -4492 -10540 -4416 -10524
rect -4492 -10558 -4476 -10540
rect -4610 -10574 -4572 -10558
rect -4692 -10612 -4572 -10574
rect -4514 -10574 -4476 -10558
rect -4432 -10558 -4416 -10540
rect -4314 -10540 -4238 -10524
rect -4314 -10558 -4298 -10540
rect -4432 -10574 -4394 -10558
rect -4514 -10612 -4394 -10574
rect -4336 -10574 -4298 -10558
rect -4254 -10558 -4238 -10540
rect -4136 -10540 -4060 -10524
rect -4136 -10558 -4120 -10540
rect -4254 -10574 -4216 -10558
rect -4336 -10612 -4216 -10574
rect -4158 -10574 -4120 -10558
rect -4076 -10558 -4060 -10540
rect -4076 -10574 -4038 -10558
rect -4158 -10612 -4038 -10574
rect 6580 -10610 6656 -10594
rect 6580 -10628 6596 -10610
rect 6558 -10644 6596 -10628
rect 6640 -10628 6656 -10610
rect 6758 -10610 6834 -10594
rect 6758 -10628 6774 -10610
rect 6640 -10644 6678 -10628
rect 6558 -10682 6678 -10644
rect 6736 -10644 6774 -10628
rect 6818 -10628 6834 -10610
rect 6936 -10610 7012 -10594
rect 6936 -10628 6952 -10610
rect 6818 -10644 6856 -10628
rect 6736 -10682 6856 -10644
rect 6914 -10644 6952 -10628
rect 6996 -10628 7012 -10610
rect 7114 -10610 7190 -10594
rect 7114 -10628 7130 -10610
rect 6996 -10644 7034 -10628
rect 6914 -10682 7034 -10644
rect 7092 -10644 7130 -10628
rect 7174 -10628 7190 -10610
rect 7292 -10610 7368 -10594
rect 7292 -10628 7308 -10610
rect 7174 -10644 7212 -10628
rect 7092 -10682 7212 -10644
rect 7270 -10644 7308 -10628
rect 7352 -10628 7368 -10610
rect 7470 -10610 7546 -10594
rect 7470 -10628 7486 -10610
rect 7352 -10644 7390 -10628
rect 7270 -10682 7390 -10644
rect 7448 -10644 7486 -10628
rect 7530 -10628 7546 -10610
rect 7648 -10610 7724 -10594
rect 7648 -10628 7664 -10610
rect 7530 -10644 7568 -10628
rect 7448 -10682 7568 -10644
rect 7626 -10644 7664 -10628
rect 7708 -10628 7724 -10610
rect 7826 -10610 7902 -10594
rect 7826 -10628 7842 -10610
rect 7708 -10644 7746 -10628
rect 7626 -10682 7746 -10644
rect 7804 -10644 7842 -10628
rect 7886 -10628 7902 -10610
rect 8004 -10610 8080 -10594
rect 8004 -10628 8020 -10610
rect 7886 -10644 7924 -10628
rect 7804 -10682 7924 -10644
rect 7982 -10644 8020 -10628
rect 8064 -10628 8080 -10610
rect 8182 -10610 8258 -10594
rect 8182 -10628 8198 -10610
rect 8064 -10644 8102 -10628
rect 7982 -10682 8102 -10644
rect 8160 -10644 8198 -10628
rect 8242 -10628 8258 -10610
rect 8360 -10610 8436 -10594
rect 8360 -10628 8376 -10610
rect 8242 -10644 8280 -10628
rect 8160 -10682 8280 -10644
rect 8338 -10644 8376 -10628
rect 8420 -10628 8436 -10610
rect 8538 -10610 8614 -10594
rect 8538 -10628 8554 -10610
rect 8420 -10644 8458 -10628
rect 8338 -10682 8458 -10644
rect 8516 -10644 8554 -10628
rect 8598 -10628 8614 -10610
rect 8716 -10610 8792 -10594
rect 8716 -10628 8732 -10610
rect 8598 -10644 8636 -10628
rect 8516 -10682 8636 -10644
rect 8694 -10644 8732 -10628
rect 8776 -10628 8792 -10610
rect 8894 -10610 8970 -10594
rect 8894 -10628 8910 -10610
rect 8776 -10644 8814 -10628
rect 8694 -10682 8814 -10644
rect 8872 -10644 8910 -10628
rect 8954 -10628 8970 -10610
rect 9072 -10610 9148 -10594
rect 9072 -10628 9088 -10610
rect 8954 -10644 8992 -10628
rect 8872 -10682 8992 -10644
rect 9050 -10644 9088 -10628
rect 9132 -10628 9148 -10610
rect 9250 -10610 9326 -10594
rect 9250 -10628 9266 -10610
rect 9132 -10644 9170 -10628
rect 9050 -10682 9170 -10644
rect 9228 -10644 9266 -10628
rect 9310 -10628 9326 -10610
rect 9310 -10644 9348 -10628
rect 9228 -10682 9348 -10644
rect -5582 -10930 -5462 -10892
rect -5582 -10946 -5544 -10930
rect -5560 -10964 -5544 -10946
rect -5500 -10946 -5462 -10930
rect -5404 -10930 -5284 -10892
rect -5404 -10946 -5366 -10930
rect -5500 -10964 -5484 -10946
rect -5560 -10980 -5484 -10964
rect -5382 -10964 -5366 -10946
rect -5322 -10946 -5284 -10930
rect -5226 -10930 -5106 -10892
rect -5226 -10946 -5188 -10930
rect -5322 -10964 -5306 -10946
rect -5382 -10980 -5306 -10964
rect -5204 -10964 -5188 -10946
rect -5144 -10946 -5106 -10930
rect -5048 -10930 -4928 -10892
rect -5048 -10946 -5010 -10930
rect -5144 -10964 -5128 -10946
rect -5204 -10980 -5128 -10964
rect -5026 -10964 -5010 -10946
rect -4966 -10946 -4928 -10930
rect -4870 -10930 -4750 -10892
rect -4870 -10946 -4832 -10930
rect -4966 -10964 -4950 -10946
rect -5026 -10980 -4950 -10964
rect -4848 -10964 -4832 -10946
rect -4788 -10946 -4750 -10930
rect -4692 -10930 -4572 -10892
rect -4692 -10946 -4654 -10930
rect -4788 -10964 -4772 -10946
rect -4848 -10980 -4772 -10964
rect -4670 -10964 -4654 -10946
rect -4610 -10946 -4572 -10930
rect -4514 -10930 -4394 -10892
rect -4514 -10946 -4476 -10930
rect -4610 -10964 -4594 -10946
rect -4670 -10980 -4594 -10964
rect -4492 -10964 -4476 -10946
rect -4432 -10946 -4394 -10930
rect -4336 -10930 -4216 -10892
rect -4336 -10946 -4298 -10930
rect -4432 -10964 -4416 -10946
rect -4492 -10980 -4416 -10964
rect -4314 -10964 -4298 -10946
rect -4254 -10946 -4216 -10930
rect -4158 -10930 -4038 -10892
rect -4158 -10946 -4120 -10930
rect -4254 -10964 -4238 -10946
rect -4314 -10980 -4238 -10964
rect -4136 -10964 -4120 -10946
rect -4076 -10946 -4038 -10930
rect -4076 -10964 -4060 -10946
rect 10818 -10770 10938 -10732
rect 10818 -10786 10856 -10770
rect 10840 -10804 10856 -10786
rect 10900 -10786 10938 -10770
rect 11110 -10770 11230 -10732
rect 11110 -10786 11148 -10770
rect 10900 -10804 10916 -10786
rect 10840 -10820 10916 -10804
rect 11132 -10804 11148 -10786
rect 11192 -10786 11230 -10770
rect 11402 -10770 11522 -10732
rect 11402 -10786 11440 -10770
rect 11192 -10804 11208 -10786
rect 11132 -10820 11208 -10804
rect 11424 -10804 11440 -10786
rect 11484 -10786 11522 -10770
rect 11694 -10770 11814 -10732
rect 11694 -10786 11732 -10770
rect 11484 -10804 11500 -10786
rect 11424 -10820 11500 -10804
rect 11716 -10804 11732 -10786
rect 11776 -10786 11814 -10770
rect 11986 -10770 12106 -10732
rect 11986 -10786 12024 -10770
rect 11776 -10804 11792 -10786
rect 11716 -10820 11792 -10804
rect 12008 -10804 12024 -10786
rect 12068 -10786 12106 -10770
rect 12278 -10770 12398 -10732
rect 12278 -10786 12316 -10770
rect 12068 -10804 12084 -10786
rect 12008 -10820 12084 -10804
rect 12300 -10804 12316 -10786
rect 12360 -10786 12398 -10770
rect 12570 -10770 12690 -10732
rect 12570 -10786 12608 -10770
rect 12360 -10804 12376 -10786
rect 12300 -10820 12376 -10804
rect 12592 -10804 12608 -10786
rect 12652 -10786 12690 -10770
rect 12652 -10804 12668 -10786
rect 12592 -10820 12668 -10804
rect -4136 -10980 -4060 -10964
rect 6558 -11000 6678 -10962
rect 6558 -11016 6596 -11000
rect -2105 -11048 -2029 -11032
rect -2105 -11066 -2089 -11048
rect -5560 -11090 -5484 -11074
rect -5560 -11108 -5544 -11090
rect -5582 -11124 -5544 -11108
rect -5500 -11108 -5484 -11090
rect -5382 -11090 -5306 -11074
rect -5382 -11108 -5366 -11090
rect -5500 -11124 -5462 -11108
rect -5582 -11162 -5462 -11124
rect -5404 -11124 -5366 -11108
rect -5322 -11108 -5306 -11090
rect -5204 -11090 -5128 -11074
rect -5204 -11108 -5188 -11090
rect -5322 -11124 -5284 -11108
rect -5404 -11162 -5284 -11124
rect -5226 -11124 -5188 -11108
rect -5144 -11108 -5128 -11090
rect -5026 -11090 -4950 -11074
rect -5026 -11108 -5010 -11090
rect -5144 -11124 -5106 -11108
rect -5226 -11162 -5106 -11124
rect -5048 -11124 -5010 -11108
rect -4966 -11108 -4950 -11090
rect -4848 -11090 -4772 -11074
rect -4848 -11108 -4832 -11090
rect -4966 -11124 -4928 -11108
rect -5048 -11162 -4928 -11124
rect -4870 -11124 -4832 -11108
rect -4788 -11108 -4772 -11090
rect -4670 -11090 -4594 -11074
rect -4670 -11108 -4654 -11090
rect -4788 -11124 -4750 -11108
rect -4870 -11162 -4750 -11124
rect -4692 -11124 -4654 -11108
rect -4610 -11108 -4594 -11090
rect -4492 -11090 -4416 -11074
rect -4492 -11108 -4476 -11090
rect -4610 -11124 -4572 -11108
rect -4692 -11162 -4572 -11124
rect -4514 -11124 -4476 -11108
rect -4432 -11108 -4416 -11090
rect -4314 -11090 -4238 -11074
rect -4314 -11108 -4298 -11090
rect -4432 -11124 -4394 -11108
rect -4514 -11162 -4394 -11124
rect -4336 -11124 -4298 -11108
rect -4254 -11108 -4238 -11090
rect -4136 -11090 -4060 -11074
rect -4136 -11108 -4120 -11090
rect -4254 -11124 -4216 -11108
rect -4336 -11162 -4216 -11124
rect -4158 -11124 -4120 -11108
rect -4076 -11108 -4060 -11090
rect -2127 -11082 -2089 -11066
rect -2045 -11066 -2029 -11048
rect -1927 -11048 -1851 -11032
rect -1927 -11066 -1911 -11048
rect -2045 -11082 -2007 -11066
rect -4076 -11124 -4038 -11108
rect -2127 -11120 -2007 -11082
rect -1949 -11082 -1911 -11066
rect -1867 -11066 -1851 -11048
rect -1749 -11048 -1673 -11032
rect -1749 -11066 -1733 -11048
rect -1867 -11082 -1829 -11066
rect -1949 -11120 -1829 -11082
rect -1771 -11082 -1733 -11066
rect -1689 -11066 -1673 -11048
rect -1571 -11048 -1495 -11032
rect -1571 -11066 -1555 -11048
rect -1689 -11082 -1651 -11066
rect -1771 -11120 -1651 -11082
rect -1593 -11082 -1555 -11066
rect -1511 -11066 -1495 -11048
rect -1393 -11048 -1317 -11032
rect -1393 -11066 -1377 -11048
rect -1511 -11082 -1473 -11066
rect -1593 -11120 -1473 -11082
rect -1415 -11082 -1377 -11066
rect -1333 -11066 -1317 -11048
rect -1215 -11048 -1139 -11032
rect -1215 -11066 -1199 -11048
rect -1333 -11082 -1295 -11066
rect -1415 -11120 -1295 -11082
rect -1237 -11082 -1199 -11066
rect -1155 -11066 -1139 -11048
rect -1037 -11048 -961 -11032
rect -1037 -11066 -1021 -11048
rect -1155 -11082 -1117 -11066
rect -1237 -11120 -1117 -11082
rect -1059 -11082 -1021 -11066
rect -977 -11066 -961 -11048
rect -859 -11048 -783 -11032
rect -859 -11066 -843 -11048
rect -977 -11082 -939 -11066
rect -1059 -11120 -939 -11082
rect -881 -11082 -843 -11066
rect -799 -11066 -783 -11048
rect -681 -11048 -605 -11032
rect -681 -11066 -665 -11048
rect -799 -11082 -761 -11066
rect -881 -11120 -761 -11082
rect -703 -11082 -665 -11066
rect -621 -11066 -605 -11048
rect -503 -11048 -427 -11032
rect -503 -11066 -487 -11048
rect -621 -11082 -583 -11066
rect -703 -11120 -583 -11082
rect -525 -11082 -487 -11066
rect -443 -11066 -427 -11048
rect -325 -11048 -249 -11032
rect -325 -11066 -309 -11048
rect -443 -11082 -405 -11066
rect -525 -11120 -405 -11082
rect -347 -11082 -309 -11066
rect -265 -11066 -249 -11048
rect -147 -11048 -71 -11032
rect -147 -11066 -131 -11048
rect -265 -11082 -227 -11066
rect -347 -11120 -227 -11082
rect -169 -11082 -131 -11066
rect -87 -11066 -71 -11048
rect 31 -11048 107 -11032
rect 31 -11066 47 -11048
rect -87 -11082 -49 -11066
rect -169 -11120 -49 -11082
rect 9 -11082 47 -11066
rect 91 -11066 107 -11048
rect 209 -11048 285 -11032
rect 209 -11066 225 -11048
rect 91 -11082 129 -11066
rect 9 -11120 129 -11082
rect 187 -11082 225 -11066
rect 269 -11066 285 -11048
rect 387 -11048 463 -11032
rect 387 -11066 403 -11048
rect 269 -11082 307 -11066
rect 187 -11120 307 -11082
rect 365 -11082 403 -11066
rect 447 -11066 463 -11048
rect 565 -11048 641 -11032
rect 565 -11066 581 -11048
rect 447 -11082 485 -11066
rect 365 -11120 485 -11082
rect 543 -11082 581 -11066
rect 625 -11066 641 -11048
rect 743 -11048 819 -11032
rect 743 -11066 759 -11048
rect 625 -11082 663 -11066
rect 543 -11120 663 -11082
rect 721 -11082 759 -11066
rect 803 -11066 819 -11048
rect 921 -11048 997 -11032
rect 921 -11066 937 -11048
rect 803 -11082 841 -11066
rect 721 -11120 841 -11082
rect 899 -11082 937 -11066
rect 981 -11066 997 -11048
rect 1099 -11048 1175 -11032
rect 1099 -11066 1115 -11048
rect 981 -11082 1019 -11066
rect 899 -11120 1019 -11082
rect 1077 -11082 1115 -11066
rect 1159 -11066 1175 -11048
rect 1277 -11048 1353 -11032
rect 1277 -11066 1293 -11048
rect 1159 -11082 1197 -11066
rect 1077 -11120 1197 -11082
rect 1255 -11082 1293 -11066
rect 1337 -11066 1353 -11048
rect 1455 -11048 1531 -11032
rect 1455 -11066 1471 -11048
rect 1337 -11082 1375 -11066
rect 1255 -11120 1375 -11082
rect 1433 -11082 1471 -11066
rect 1515 -11066 1531 -11048
rect 1633 -11048 1709 -11032
rect 1633 -11066 1649 -11048
rect 1515 -11082 1553 -11066
rect 1433 -11120 1553 -11082
rect 1611 -11082 1649 -11066
rect 1693 -11066 1709 -11048
rect 1811 -11048 1887 -11032
rect 1811 -11066 1827 -11048
rect 1693 -11082 1731 -11066
rect 1611 -11120 1731 -11082
rect 1789 -11082 1827 -11066
rect 1871 -11066 1887 -11048
rect 1989 -11048 2065 -11032
rect 1989 -11066 2005 -11048
rect 1871 -11082 1909 -11066
rect 1789 -11120 1909 -11082
rect 1967 -11082 2005 -11066
rect 2049 -11066 2065 -11048
rect 2167 -11048 2243 -11032
rect 2167 -11066 2183 -11048
rect 2049 -11082 2087 -11066
rect 1967 -11120 2087 -11082
rect 2145 -11082 2183 -11066
rect 2227 -11066 2243 -11048
rect 2345 -11048 2421 -11032
rect 2345 -11066 2361 -11048
rect 2227 -11082 2265 -11066
rect 2145 -11120 2265 -11082
rect 2323 -11082 2361 -11066
rect 2405 -11066 2421 -11048
rect 2523 -11048 2599 -11032
rect 2523 -11066 2539 -11048
rect 2405 -11082 2443 -11066
rect 2323 -11120 2443 -11082
rect 2501 -11082 2539 -11066
rect 2583 -11066 2599 -11048
rect 2701 -11048 2777 -11032
rect 2701 -11066 2717 -11048
rect 2583 -11082 2621 -11066
rect 2501 -11120 2621 -11082
rect 2679 -11082 2717 -11066
rect 2761 -11066 2777 -11048
rect 2879 -11048 2955 -11032
rect 2879 -11066 2895 -11048
rect 2761 -11082 2799 -11066
rect 2679 -11120 2799 -11082
rect 2857 -11082 2895 -11066
rect 2939 -11066 2955 -11048
rect 3057 -11048 3133 -11032
rect 3057 -11066 3073 -11048
rect 2939 -11082 2977 -11066
rect 2857 -11120 2977 -11082
rect 3035 -11082 3073 -11066
rect 3117 -11066 3133 -11048
rect 3235 -11048 3311 -11032
rect 3235 -11066 3251 -11048
rect 3117 -11082 3155 -11066
rect 3035 -11120 3155 -11082
rect 3213 -11082 3251 -11066
rect 3295 -11066 3311 -11048
rect 3413 -11048 3489 -11032
rect 3413 -11066 3429 -11048
rect 3295 -11082 3333 -11066
rect 3213 -11120 3333 -11082
rect 3391 -11082 3429 -11066
rect 3473 -11066 3489 -11048
rect 3591 -11048 3667 -11032
rect 3591 -11066 3607 -11048
rect 3473 -11082 3511 -11066
rect 3391 -11120 3511 -11082
rect 3569 -11082 3607 -11066
rect 3651 -11066 3667 -11048
rect 3769 -11048 3845 -11032
rect 3769 -11066 3785 -11048
rect 3651 -11082 3689 -11066
rect 3569 -11120 3689 -11082
rect 3747 -11082 3785 -11066
rect 3829 -11066 3845 -11048
rect 3947 -11048 4023 -11032
rect 3947 -11066 3963 -11048
rect 3829 -11082 3867 -11066
rect 3747 -11120 3867 -11082
rect 3925 -11082 3963 -11066
rect 4007 -11066 4023 -11048
rect 6580 -11034 6596 -11016
rect 6640 -11016 6678 -11000
rect 6736 -11000 6856 -10962
rect 6736 -11016 6774 -11000
rect 6640 -11034 6656 -11016
rect 6580 -11050 6656 -11034
rect 6758 -11034 6774 -11016
rect 6818 -11016 6856 -11000
rect 6914 -11000 7034 -10962
rect 6914 -11016 6952 -11000
rect 6818 -11034 6834 -11016
rect 6758 -11050 6834 -11034
rect 6936 -11034 6952 -11016
rect 6996 -11016 7034 -11000
rect 7092 -11000 7212 -10962
rect 7092 -11016 7130 -11000
rect 6996 -11034 7012 -11016
rect 6936 -11050 7012 -11034
rect 7114 -11034 7130 -11016
rect 7174 -11016 7212 -11000
rect 7270 -11000 7390 -10962
rect 7270 -11016 7308 -11000
rect 7174 -11034 7190 -11016
rect 7114 -11050 7190 -11034
rect 7292 -11034 7308 -11016
rect 7352 -11016 7390 -11000
rect 7448 -11000 7568 -10962
rect 7448 -11016 7486 -11000
rect 7352 -11034 7368 -11016
rect 7292 -11050 7368 -11034
rect 7470 -11034 7486 -11016
rect 7530 -11016 7568 -11000
rect 7626 -11000 7746 -10962
rect 7626 -11016 7664 -11000
rect 7530 -11034 7546 -11016
rect 7470 -11050 7546 -11034
rect 7648 -11034 7664 -11016
rect 7708 -11016 7746 -11000
rect 7804 -11000 7924 -10962
rect 7804 -11016 7842 -11000
rect 7708 -11034 7724 -11016
rect 7648 -11050 7724 -11034
rect 7826 -11034 7842 -11016
rect 7886 -11016 7924 -11000
rect 7982 -11000 8102 -10962
rect 7982 -11016 8020 -11000
rect 7886 -11034 7902 -11016
rect 7826 -11050 7902 -11034
rect 8004 -11034 8020 -11016
rect 8064 -11016 8102 -11000
rect 8160 -11000 8280 -10962
rect 8160 -11016 8198 -11000
rect 8064 -11034 8080 -11016
rect 8004 -11050 8080 -11034
rect 8182 -11034 8198 -11016
rect 8242 -11016 8280 -11000
rect 8338 -11000 8458 -10962
rect 8338 -11016 8376 -11000
rect 8242 -11034 8258 -11016
rect 8182 -11050 8258 -11034
rect 8360 -11034 8376 -11016
rect 8420 -11016 8458 -11000
rect 8516 -11000 8636 -10962
rect 8516 -11016 8554 -11000
rect 8420 -11034 8436 -11016
rect 8360 -11050 8436 -11034
rect 8538 -11034 8554 -11016
rect 8598 -11016 8636 -11000
rect 8694 -11000 8814 -10962
rect 8694 -11016 8732 -11000
rect 8598 -11034 8614 -11016
rect 8538 -11050 8614 -11034
rect 8716 -11034 8732 -11016
rect 8776 -11016 8814 -11000
rect 8872 -11000 8992 -10962
rect 8872 -11016 8910 -11000
rect 8776 -11034 8792 -11016
rect 8716 -11050 8792 -11034
rect 8894 -11034 8910 -11016
rect 8954 -11016 8992 -11000
rect 9050 -11000 9170 -10962
rect 9050 -11016 9088 -11000
rect 8954 -11034 8970 -11016
rect 8894 -11050 8970 -11034
rect 9072 -11034 9088 -11016
rect 9132 -11016 9170 -11000
rect 9228 -11000 9348 -10962
rect 9228 -11016 9266 -11000
rect 9132 -11034 9148 -11016
rect 9072 -11050 9148 -11034
rect 9250 -11034 9266 -11016
rect 9310 -11016 9348 -11000
rect 9310 -11034 9326 -11016
rect 9250 -11050 9326 -11034
rect 4007 -11082 4045 -11066
rect 3925 -11120 4045 -11082
rect -4158 -11162 -4038 -11124
rect -5582 -11480 -5462 -11442
rect -5582 -11496 -5544 -11480
rect -5560 -11514 -5544 -11496
rect -5500 -11496 -5462 -11480
rect -5404 -11480 -5284 -11442
rect -5404 -11496 -5366 -11480
rect -5500 -11514 -5484 -11496
rect -5560 -11530 -5484 -11514
rect -5382 -11514 -5366 -11496
rect -5322 -11496 -5284 -11480
rect -5226 -11480 -5106 -11442
rect -5226 -11496 -5188 -11480
rect -5322 -11514 -5306 -11496
rect -5382 -11530 -5306 -11514
rect -5204 -11514 -5188 -11496
rect -5144 -11496 -5106 -11480
rect -5048 -11480 -4928 -11442
rect -5048 -11496 -5010 -11480
rect -5144 -11514 -5128 -11496
rect -5204 -11530 -5128 -11514
rect -5026 -11514 -5010 -11496
rect -4966 -11496 -4928 -11480
rect -4870 -11480 -4750 -11442
rect -4870 -11496 -4832 -11480
rect -4966 -11514 -4950 -11496
rect -5026 -11530 -4950 -11514
rect -4848 -11514 -4832 -11496
rect -4788 -11496 -4750 -11480
rect -4692 -11480 -4572 -11442
rect -4692 -11496 -4654 -11480
rect -4788 -11514 -4772 -11496
rect -4848 -11530 -4772 -11514
rect -4670 -11514 -4654 -11496
rect -4610 -11496 -4572 -11480
rect -4514 -11480 -4394 -11442
rect -4514 -11496 -4476 -11480
rect -4610 -11514 -4594 -11496
rect -4670 -11530 -4594 -11514
rect -4492 -11514 -4476 -11496
rect -4432 -11496 -4394 -11480
rect -4336 -11480 -4216 -11442
rect -4336 -11496 -4298 -11480
rect -4432 -11514 -4416 -11496
rect -4492 -11530 -4416 -11514
rect -4314 -11514 -4298 -11496
rect -4254 -11496 -4216 -11480
rect -4158 -11480 -4038 -11442
rect 10840 -11150 10916 -11134
rect 10840 -11168 10856 -11150
rect 10818 -11184 10856 -11168
rect 10900 -11168 10916 -11150
rect 11132 -11150 11208 -11134
rect 11132 -11168 11148 -11150
rect 10900 -11184 10938 -11168
rect 10818 -11222 10938 -11184
rect 11110 -11184 11148 -11168
rect 11192 -11168 11208 -11150
rect 11424 -11150 11500 -11134
rect 11424 -11168 11440 -11150
rect 11192 -11184 11230 -11168
rect 11110 -11222 11230 -11184
rect 11402 -11184 11440 -11168
rect 11484 -11168 11500 -11150
rect 11716 -11150 11792 -11134
rect 11716 -11168 11732 -11150
rect 11484 -11184 11522 -11168
rect 11402 -11222 11522 -11184
rect 11694 -11184 11732 -11168
rect 11776 -11168 11792 -11150
rect 12008 -11150 12084 -11134
rect 12008 -11168 12024 -11150
rect 11776 -11184 11814 -11168
rect 11694 -11222 11814 -11184
rect 11986 -11184 12024 -11168
rect 12068 -11168 12084 -11150
rect 12300 -11150 12376 -11134
rect 12300 -11168 12316 -11150
rect 12068 -11184 12106 -11168
rect 11986 -11222 12106 -11184
rect 12278 -11184 12316 -11168
rect 12360 -11168 12376 -11150
rect 12592 -11150 12668 -11134
rect 12592 -11168 12608 -11150
rect 12360 -11184 12398 -11168
rect 12278 -11222 12398 -11184
rect 12570 -11184 12608 -11168
rect 12652 -11168 12668 -11150
rect 12652 -11184 12690 -11168
rect 12570 -11222 12690 -11184
rect -2127 -11438 -2007 -11400
rect -2127 -11454 -2089 -11438
rect -2105 -11472 -2089 -11454
rect -2045 -11454 -2007 -11438
rect -1949 -11438 -1829 -11400
rect -1949 -11454 -1911 -11438
rect -2045 -11472 -2029 -11454
rect -4158 -11496 -4120 -11480
rect -4254 -11514 -4238 -11496
rect -4314 -11530 -4238 -11514
rect -4136 -11514 -4120 -11496
rect -4076 -11496 -4038 -11480
rect -2105 -11488 -2029 -11472
rect -1927 -11472 -1911 -11454
rect -1867 -11454 -1829 -11438
rect -1771 -11438 -1651 -11400
rect -1771 -11454 -1733 -11438
rect -1867 -11472 -1851 -11454
rect -1927 -11488 -1851 -11472
rect -1749 -11472 -1733 -11454
rect -1689 -11454 -1651 -11438
rect -1593 -11438 -1473 -11400
rect -1593 -11454 -1555 -11438
rect -1689 -11472 -1673 -11454
rect -1749 -11488 -1673 -11472
rect -1571 -11472 -1555 -11454
rect -1511 -11454 -1473 -11438
rect -1415 -11438 -1295 -11400
rect -1415 -11454 -1377 -11438
rect -1511 -11472 -1495 -11454
rect -1571 -11488 -1495 -11472
rect -1393 -11472 -1377 -11454
rect -1333 -11454 -1295 -11438
rect -1237 -11438 -1117 -11400
rect -1237 -11454 -1199 -11438
rect -1333 -11472 -1317 -11454
rect -1393 -11488 -1317 -11472
rect -1215 -11472 -1199 -11454
rect -1155 -11454 -1117 -11438
rect -1059 -11438 -939 -11400
rect -1059 -11454 -1021 -11438
rect -1155 -11472 -1139 -11454
rect -1215 -11488 -1139 -11472
rect -1037 -11472 -1021 -11454
rect -977 -11454 -939 -11438
rect -881 -11438 -761 -11400
rect -881 -11454 -843 -11438
rect -977 -11472 -961 -11454
rect -1037 -11488 -961 -11472
rect -859 -11472 -843 -11454
rect -799 -11454 -761 -11438
rect -703 -11438 -583 -11400
rect -703 -11454 -665 -11438
rect -799 -11472 -783 -11454
rect -859 -11488 -783 -11472
rect -681 -11472 -665 -11454
rect -621 -11454 -583 -11438
rect -525 -11438 -405 -11400
rect -525 -11454 -487 -11438
rect -621 -11472 -605 -11454
rect -681 -11488 -605 -11472
rect -503 -11472 -487 -11454
rect -443 -11454 -405 -11438
rect -347 -11438 -227 -11400
rect -347 -11454 -309 -11438
rect -443 -11472 -427 -11454
rect -503 -11488 -427 -11472
rect -325 -11472 -309 -11454
rect -265 -11454 -227 -11438
rect -169 -11438 -49 -11400
rect -169 -11454 -131 -11438
rect -265 -11472 -249 -11454
rect -325 -11488 -249 -11472
rect -147 -11472 -131 -11454
rect -87 -11454 -49 -11438
rect 9 -11438 129 -11400
rect 9 -11454 47 -11438
rect -87 -11472 -71 -11454
rect -147 -11488 -71 -11472
rect 31 -11472 47 -11454
rect 91 -11454 129 -11438
rect 187 -11438 307 -11400
rect 187 -11454 225 -11438
rect 91 -11472 107 -11454
rect 31 -11488 107 -11472
rect 209 -11472 225 -11454
rect 269 -11454 307 -11438
rect 365 -11438 485 -11400
rect 365 -11454 403 -11438
rect 269 -11472 285 -11454
rect 209 -11488 285 -11472
rect 387 -11472 403 -11454
rect 447 -11454 485 -11438
rect 543 -11438 663 -11400
rect 543 -11454 581 -11438
rect 447 -11472 463 -11454
rect 387 -11488 463 -11472
rect 565 -11472 581 -11454
rect 625 -11454 663 -11438
rect 721 -11438 841 -11400
rect 721 -11454 759 -11438
rect 625 -11472 641 -11454
rect 565 -11488 641 -11472
rect 743 -11472 759 -11454
rect 803 -11454 841 -11438
rect 899 -11438 1019 -11400
rect 899 -11454 937 -11438
rect 803 -11472 819 -11454
rect 743 -11488 819 -11472
rect 921 -11472 937 -11454
rect 981 -11454 1019 -11438
rect 1077 -11438 1197 -11400
rect 1077 -11454 1115 -11438
rect 981 -11472 997 -11454
rect 921 -11488 997 -11472
rect 1099 -11472 1115 -11454
rect 1159 -11454 1197 -11438
rect 1255 -11438 1375 -11400
rect 1255 -11454 1293 -11438
rect 1159 -11472 1175 -11454
rect 1099 -11488 1175 -11472
rect 1277 -11472 1293 -11454
rect 1337 -11454 1375 -11438
rect 1433 -11438 1553 -11400
rect 1433 -11454 1471 -11438
rect 1337 -11472 1353 -11454
rect 1277 -11488 1353 -11472
rect 1455 -11472 1471 -11454
rect 1515 -11454 1553 -11438
rect 1611 -11438 1731 -11400
rect 1611 -11454 1649 -11438
rect 1515 -11472 1531 -11454
rect 1455 -11488 1531 -11472
rect 1633 -11472 1649 -11454
rect 1693 -11454 1731 -11438
rect 1789 -11438 1909 -11400
rect 1789 -11454 1827 -11438
rect 1693 -11472 1709 -11454
rect 1633 -11488 1709 -11472
rect 1811 -11472 1827 -11454
rect 1871 -11454 1909 -11438
rect 1967 -11438 2087 -11400
rect 1967 -11454 2005 -11438
rect 1871 -11472 1887 -11454
rect 1811 -11488 1887 -11472
rect 1989 -11472 2005 -11454
rect 2049 -11454 2087 -11438
rect 2145 -11438 2265 -11400
rect 2145 -11454 2183 -11438
rect 2049 -11472 2065 -11454
rect 1989 -11488 2065 -11472
rect 2167 -11472 2183 -11454
rect 2227 -11454 2265 -11438
rect 2323 -11438 2443 -11400
rect 2323 -11454 2361 -11438
rect 2227 -11472 2243 -11454
rect 2167 -11488 2243 -11472
rect 2345 -11472 2361 -11454
rect 2405 -11454 2443 -11438
rect 2501 -11438 2621 -11400
rect 2501 -11454 2539 -11438
rect 2405 -11472 2421 -11454
rect 2345 -11488 2421 -11472
rect 2523 -11472 2539 -11454
rect 2583 -11454 2621 -11438
rect 2679 -11438 2799 -11400
rect 2679 -11454 2717 -11438
rect 2583 -11472 2599 -11454
rect 2523 -11488 2599 -11472
rect 2701 -11472 2717 -11454
rect 2761 -11454 2799 -11438
rect 2857 -11438 2977 -11400
rect 2857 -11454 2895 -11438
rect 2761 -11472 2777 -11454
rect 2701 -11488 2777 -11472
rect 2879 -11472 2895 -11454
rect 2939 -11454 2977 -11438
rect 3035 -11438 3155 -11400
rect 3035 -11454 3073 -11438
rect 2939 -11472 2955 -11454
rect 2879 -11488 2955 -11472
rect 3057 -11472 3073 -11454
rect 3117 -11454 3155 -11438
rect 3213 -11438 3333 -11400
rect 3213 -11454 3251 -11438
rect 3117 -11472 3133 -11454
rect 3057 -11488 3133 -11472
rect 3235 -11472 3251 -11454
rect 3295 -11454 3333 -11438
rect 3391 -11438 3511 -11400
rect 3391 -11454 3429 -11438
rect 3295 -11472 3311 -11454
rect 3235 -11488 3311 -11472
rect 3413 -11472 3429 -11454
rect 3473 -11454 3511 -11438
rect 3569 -11438 3689 -11400
rect 3569 -11454 3607 -11438
rect 3473 -11472 3489 -11454
rect 3413 -11488 3489 -11472
rect 3591 -11472 3607 -11454
rect 3651 -11454 3689 -11438
rect 3747 -11438 3867 -11400
rect 3747 -11454 3785 -11438
rect 3651 -11472 3667 -11454
rect 3591 -11488 3667 -11472
rect 3769 -11472 3785 -11454
rect 3829 -11454 3867 -11438
rect 3925 -11438 4045 -11400
rect 3925 -11454 3963 -11438
rect 3829 -11472 3845 -11454
rect 3769 -11488 3845 -11472
rect 3947 -11472 3963 -11454
rect 4007 -11454 4045 -11438
rect 4007 -11472 4023 -11454
rect 3947 -11488 4023 -11472
rect -4076 -11514 -4060 -11496
rect -4136 -11530 -4060 -11514
rect 6580 -11510 6656 -11494
rect 6580 -11528 6596 -11510
rect 6558 -11544 6596 -11528
rect 6640 -11528 6656 -11510
rect 6758 -11510 6834 -11494
rect 6758 -11528 6774 -11510
rect 6640 -11544 6678 -11528
rect 6558 -11582 6678 -11544
rect 6736 -11544 6774 -11528
rect 6818 -11528 6834 -11510
rect 6936 -11510 7012 -11494
rect 6936 -11528 6952 -11510
rect 6818 -11544 6856 -11528
rect 6736 -11582 6856 -11544
rect 6914 -11544 6952 -11528
rect 6996 -11528 7012 -11510
rect 7114 -11510 7190 -11494
rect 7114 -11528 7130 -11510
rect 6996 -11544 7034 -11528
rect 6914 -11582 7034 -11544
rect 7092 -11544 7130 -11528
rect 7174 -11528 7190 -11510
rect 7292 -11510 7368 -11494
rect 7292 -11528 7308 -11510
rect 7174 -11544 7212 -11528
rect 7092 -11582 7212 -11544
rect 7270 -11544 7308 -11528
rect 7352 -11528 7368 -11510
rect 7470 -11510 7546 -11494
rect 7470 -11528 7486 -11510
rect 7352 -11544 7390 -11528
rect 7270 -11582 7390 -11544
rect 7448 -11544 7486 -11528
rect 7530 -11528 7546 -11510
rect 7648 -11510 7724 -11494
rect 7648 -11528 7664 -11510
rect 7530 -11544 7568 -11528
rect 7448 -11582 7568 -11544
rect 7626 -11544 7664 -11528
rect 7708 -11528 7724 -11510
rect 7826 -11510 7902 -11494
rect 7826 -11528 7842 -11510
rect 7708 -11544 7746 -11528
rect 7626 -11582 7746 -11544
rect 7804 -11544 7842 -11528
rect 7886 -11528 7902 -11510
rect 8004 -11510 8080 -11494
rect 8004 -11528 8020 -11510
rect 7886 -11544 7924 -11528
rect 7804 -11582 7924 -11544
rect 7982 -11544 8020 -11528
rect 8064 -11528 8080 -11510
rect 8182 -11510 8258 -11494
rect 8182 -11528 8198 -11510
rect 8064 -11544 8102 -11528
rect 7982 -11582 8102 -11544
rect 8160 -11544 8198 -11528
rect 8242 -11528 8258 -11510
rect 8360 -11510 8436 -11494
rect 8360 -11528 8376 -11510
rect 8242 -11544 8280 -11528
rect 8160 -11582 8280 -11544
rect 8338 -11544 8376 -11528
rect 8420 -11528 8436 -11510
rect 8538 -11510 8614 -11494
rect 8538 -11528 8554 -11510
rect 8420 -11544 8458 -11528
rect 8338 -11582 8458 -11544
rect 8516 -11544 8554 -11528
rect 8598 -11528 8614 -11510
rect 8716 -11510 8792 -11494
rect 8716 -11528 8732 -11510
rect 8598 -11544 8636 -11528
rect 8516 -11582 8636 -11544
rect 8694 -11544 8732 -11528
rect 8776 -11528 8792 -11510
rect 8894 -11510 8970 -11494
rect 8894 -11528 8910 -11510
rect 8776 -11544 8814 -11528
rect 8694 -11582 8814 -11544
rect 8872 -11544 8910 -11528
rect 8954 -11528 8970 -11510
rect 9072 -11510 9148 -11494
rect 9072 -11528 9088 -11510
rect 8954 -11544 8992 -11528
rect 8872 -11582 8992 -11544
rect 9050 -11544 9088 -11528
rect 9132 -11528 9148 -11510
rect 9250 -11510 9326 -11494
rect 9250 -11528 9266 -11510
rect 9132 -11544 9170 -11528
rect 9050 -11582 9170 -11544
rect 9228 -11544 9266 -11528
rect 9310 -11528 9326 -11510
rect 9310 -11544 9348 -11528
rect 9228 -11582 9348 -11544
rect 10818 -11540 10938 -11502
rect 10818 -11556 10856 -11540
rect 10840 -11574 10856 -11556
rect 10900 -11556 10938 -11540
rect 11110 -11540 11230 -11502
rect 11110 -11556 11148 -11540
rect 10900 -11574 10916 -11556
rect -5560 -11640 -5484 -11624
rect -5560 -11658 -5544 -11640
rect -5582 -11674 -5544 -11658
rect -5500 -11658 -5484 -11640
rect -5382 -11640 -5306 -11624
rect -5382 -11658 -5366 -11640
rect -5500 -11674 -5462 -11658
rect -5582 -11712 -5462 -11674
rect -5404 -11674 -5366 -11658
rect -5322 -11658 -5306 -11640
rect -5204 -11640 -5128 -11624
rect -5204 -11658 -5188 -11640
rect -5322 -11674 -5284 -11658
rect -5404 -11712 -5284 -11674
rect -5226 -11674 -5188 -11658
rect -5144 -11658 -5128 -11640
rect -5026 -11640 -4950 -11624
rect -5026 -11658 -5010 -11640
rect -5144 -11674 -5106 -11658
rect -5226 -11712 -5106 -11674
rect -5048 -11674 -5010 -11658
rect -4966 -11658 -4950 -11640
rect -4848 -11640 -4772 -11624
rect -4848 -11658 -4832 -11640
rect -4966 -11674 -4928 -11658
rect -5048 -11712 -4928 -11674
rect -4870 -11674 -4832 -11658
rect -4788 -11658 -4772 -11640
rect -4670 -11640 -4594 -11624
rect -4670 -11658 -4654 -11640
rect -4788 -11674 -4750 -11658
rect -4870 -11712 -4750 -11674
rect -4692 -11674 -4654 -11658
rect -4610 -11658 -4594 -11640
rect -4492 -11640 -4416 -11624
rect -4492 -11658 -4476 -11640
rect -4610 -11674 -4572 -11658
rect -4692 -11712 -4572 -11674
rect -4514 -11674 -4476 -11658
rect -4432 -11658 -4416 -11640
rect -4314 -11640 -4238 -11624
rect -4314 -11658 -4298 -11640
rect -4432 -11674 -4394 -11658
rect -4514 -11712 -4394 -11674
rect -4336 -11674 -4298 -11658
rect -4254 -11658 -4238 -11640
rect -4136 -11640 -4060 -11624
rect -4136 -11658 -4120 -11640
rect -4254 -11674 -4216 -11658
rect -4336 -11712 -4216 -11674
rect -4158 -11674 -4120 -11658
rect -4076 -11658 -4060 -11640
rect -4076 -11674 -4038 -11658
rect -4158 -11712 -4038 -11674
rect 10840 -11590 10916 -11574
rect 11132 -11574 11148 -11556
rect 11192 -11556 11230 -11540
rect 11402 -11540 11522 -11502
rect 11402 -11556 11440 -11540
rect 11192 -11574 11208 -11556
rect 11132 -11590 11208 -11574
rect 11424 -11574 11440 -11556
rect 11484 -11556 11522 -11540
rect 11694 -11540 11814 -11502
rect 11694 -11556 11732 -11540
rect 11484 -11574 11500 -11556
rect 11424 -11590 11500 -11574
rect 11716 -11574 11732 -11556
rect 11776 -11556 11814 -11540
rect 11986 -11540 12106 -11502
rect 11986 -11556 12024 -11540
rect 11776 -11574 11792 -11556
rect 11716 -11590 11792 -11574
rect 12008 -11574 12024 -11556
rect 12068 -11556 12106 -11540
rect 12278 -11540 12398 -11502
rect 12278 -11556 12316 -11540
rect 12068 -11574 12084 -11556
rect 12008 -11590 12084 -11574
rect 12300 -11574 12316 -11556
rect 12360 -11556 12398 -11540
rect 12570 -11540 12690 -11502
rect 12570 -11556 12608 -11540
rect 12360 -11574 12376 -11556
rect 12300 -11590 12376 -11574
rect 12592 -11574 12608 -11556
rect 12652 -11556 12690 -11540
rect 12652 -11574 12668 -11556
rect 12592 -11590 12668 -11574
rect 6558 -11900 6678 -11862
rect 6558 -11916 6596 -11900
rect 6580 -11934 6596 -11916
rect 6640 -11916 6678 -11900
rect 6736 -11900 6856 -11862
rect 6736 -11916 6774 -11900
rect 6640 -11934 6656 -11916
rect 6580 -11950 6656 -11934
rect 6758 -11934 6774 -11916
rect 6818 -11916 6856 -11900
rect 6914 -11900 7034 -11862
rect 6914 -11916 6952 -11900
rect 6818 -11934 6834 -11916
rect 6758 -11950 6834 -11934
rect 6936 -11934 6952 -11916
rect 6996 -11916 7034 -11900
rect 7092 -11900 7212 -11862
rect 7092 -11916 7130 -11900
rect 6996 -11934 7012 -11916
rect 6936 -11950 7012 -11934
rect 7114 -11934 7130 -11916
rect 7174 -11916 7212 -11900
rect 7270 -11900 7390 -11862
rect 7270 -11916 7308 -11900
rect 7174 -11934 7190 -11916
rect 7114 -11950 7190 -11934
rect 7292 -11934 7308 -11916
rect 7352 -11916 7390 -11900
rect 7448 -11900 7568 -11862
rect 7448 -11916 7486 -11900
rect 7352 -11934 7368 -11916
rect 7292 -11950 7368 -11934
rect 7470 -11934 7486 -11916
rect 7530 -11916 7568 -11900
rect 7626 -11900 7746 -11862
rect 7626 -11916 7664 -11900
rect 7530 -11934 7546 -11916
rect 7470 -11950 7546 -11934
rect 7648 -11934 7664 -11916
rect 7708 -11916 7746 -11900
rect 7804 -11900 7924 -11862
rect 7804 -11916 7842 -11900
rect 7708 -11934 7724 -11916
rect 7648 -11950 7724 -11934
rect 7826 -11934 7842 -11916
rect 7886 -11916 7924 -11900
rect 7982 -11900 8102 -11862
rect 7982 -11916 8020 -11900
rect 7886 -11934 7902 -11916
rect 7826 -11950 7902 -11934
rect 8004 -11934 8020 -11916
rect 8064 -11916 8102 -11900
rect 8160 -11900 8280 -11862
rect 8160 -11916 8198 -11900
rect 8064 -11934 8080 -11916
rect 8004 -11950 8080 -11934
rect 8182 -11934 8198 -11916
rect 8242 -11916 8280 -11900
rect 8338 -11900 8458 -11862
rect 8338 -11916 8376 -11900
rect 8242 -11934 8258 -11916
rect 8182 -11950 8258 -11934
rect 8360 -11934 8376 -11916
rect 8420 -11916 8458 -11900
rect 8516 -11900 8636 -11862
rect 8516 -11916 8554 -11900
rect 8420 -11934 8436 -11916
rect 8360 -11950 8436 -11934
rect 8538 -11934 8554 -11916
rect 8598 -11916 8636 -11900
rect 8694 -11900 8814 -11862
rect 8694 -11916 8732 -11900
rect 8598 -11934 8614 -11916
rect 8538 -11950 8614 -11934
rect 8716 -11934 8732 -11916
rect 8776 -11916 8814 -11900
rect 8872 -11900 8992 -11862
rect 8872 -11916 8910 -11900
rect 8776 -11934 8792 -11916
rect 8716 -11950 8792 -11934
rect 8894 -11934 8910 -11916
rect 8954 -11916 8992 -11900
rect 9050 -11900 9170 -11862
rect 9050 -11916 9088 -11900
rect 8954 -11934 8970 -11916
rect 8894 -11950 8970 -11934
rect 9072 -11934 9088 -11916
rect 9132 -11916 9170 -11900
rect 9228 -11900 9348 -11862
rect 9228 -11916 9266 -11900
rect 9132 -11934 9148 -11916
rect 9072 -11950 9148 -11934
rect 9250 -11934 9266 -11916
rect 9310 -11916 9348 -11900
rect 9310 -11934 9326 -11916
rect 9250 -11950 9326 -11934
rect -5582 -12030 -5462 -11992
rect -5582 -12046 -5544 -12030
rect -5560 -12064 -5544 -12046
rect -5500 -12046 -5462 -12030
rect -5404 -12030 -5284 -11992
rect -5404 -12046 -5366 -12030
rect -5500 -12064 -5484 -12046
rect -5560 -12080 -5484 -12064
rect -5382 -12064 -5366 -12046
rect -5322 -12046 -5284 -12030
rect -5226 -12030 -5106 -11992
rect -5226 -12046 -5188 -12030
rect -5322 -12064 -5306 -12046
rect -5382 -12080 -5306 -12064
rect -5204 -12064 -5188 -12046
rect -5144 -12046 -5106 -12030
rect -5048 -12030 -4928 -11992
rect -5048 -12046 -5010 -12030
rect -5144 -12064 -5128 -12046
rect -5204 -12080 -5128 -12064
rect -5026 -12064 -5010 -12046
rect -4966 -12046 -4928 -12030
rect -4870 -12030 -4750 -11992
rect -4870 -12046 -4832 -12030
rect -4966 -12064 -4950 -12046
rect -5026 -12080 -4950 -12064
rect -4848 -12064 -4832 -12046
rect -4788 -12046 -4750 -12030
rect -4692 -12030 -4572 -11992
rect -4692 -12046 -4654 -12030
rect -4788 -12064 -4772 -12046
rect -4848 -12080 -4772 -12064
rect -4670 -12064 -4654 -12046
rect -4610 -12046 -4572 -12030
rect -4514 -12030 -4394 -11992
rect -4514 -12046 -4476 -12030
rect -4610 -12064 -4594 -12046
rect -4670 -12080 -4594 -12064
rect -4492 -12064 -4476 -12046
rect -4432 -12046 -4394 -12030
rect -4336 -12030 -4216 -11992
rect -4336 -12046 -4298 -12030
rect -4432 -12064 -4416 -12046
rect -4492 -12080 -4416 -12064
rect -4314 -12064 -4298 -12046
rect -4254 -12046 -4216 -12030
rect -4158 -12030 -4038 -11992
rect -4158 -12046 -4120 -12030
rect -4254 -12064 -4238 -12046
rect -4314 -12080 -4238 -12064
rect -4136 -12064 -4120 -12046
rect -4076 -12046 -4038 -12030
rect -4076 -12064 -4060 -12046
rect -4136 -12080 -4060 -12064
rect -2105 -12048 -2029 -12032
rect -2105 -12066 -2089 -12048
rect -2127 -12082 -2089 -12066
rect -2045 -12066 -2029 -12048
rect -1927 -12048 -1851 -12032
rect -1927 -12066 -1911 -12048
rect -2045 -12082 -2007 -12066
rect -2127 -12120 -2007 -12082
rect -1949 -12082 -1911 -12066
rect -1867 -12066 -1851 -12048
rect -1749 -12048 -1673 -12032
rect -1749 -12066 -1733 -12048
rect -1867 -12082 -1829 -12066
rect -1949 -12120 -1829 -12082
rect -1771 -12082 -1733 -12066
rect -1689 -12066 -1673 -12048
rect -1571 -12048 -1495 -12032
rect -1571 -12066 -1555 -12048
rect -1689 -12082 -1651 -12066
rect -1771 -12120 -1651 -12082
rect -1593 -12082 -1555 -12066
rect -1511 -12066 -1495 -12048
rect -1393 -12048 -1317 -12032
rect -1393 -12066 -1377 -12048
rect -1511 -12082 -1473 -12066
rect -1593 -12120 -1473 -12082
rect -1415 -12082 -1377 -12066
rect -1333 -12066 -1317 -12048
rect -1215 -12048 -1139 -12032
rect -1215 -12066 -1199 -12048
rect -1333 -12082 -1295 -12066
rect -1415 -12120 -1295 -12082
rect -1237 -12082 -1199 -12066
rect -1155 -12066 -1139 -12048
rect -1037 -12048 -961 -12032
rect -1037 -12066 -1021 -12048
rect -1155 -12082 -1117 -12066
rect -1237 -12120 -1117 -12082
rect -1059 -12082 -1021 -12066
rect -977 -12066 -961 -12048
rect -859 -12048 -783 -12032
rect -859 -12066 -843 -12048
rect -977 -12082 -939 -12066
rect -1059 -12120 -939 -12082
rect -881 -12082 -843 -12066
rect -799 -12066 -783 -12048
rect -681 -12048 -605 -12032
rect -681 -12066 -665 -12048
rect -799 -12082 -761 -12066
rect -881 -12120 -761 -12082
rect -703 -12082 -665 -12066
rect -621 -12066 -605 -12048
rect -503 -12048 -427 -12032
rect -503 -12066 -487 -12048
rect -621 -12082 -583 -12066
rect -703 -12120 -583 -12082
rect -525 -12082 -487 -12066
rect -443 -12066 -427 -12048
rect -325 -12048 -249 -12032
rect -325 -12066 -309 -12048
rect -443 -12082 -405 -12066
rect -525 -12120 -405 -12082
rect -347 -12082 -309 -12066
rect -265 -12066 -249 -12048
rect -147 -12048 -71 -12032
rect -147 -12066 -131 -12048
rect -265 -12082 -227 -12066
rect -347 -12120 -227 -12082
rect -169 -12082 -131 -12066
rect -87 -12066 -71 -12048
rect 31 -12048 107 -12032
rect 31 -12066 47 -12048
rect -87 -12082 -49 -12066
rect -169 -12120 -49 -12082
rect 9 -12082 47 -12066
rect 91 -12066 107 -12048
rect 209 -12048 285 -12032
rect 209 -12066 225 -12048
rect 91 -12082 129 -12066
rect 9 -12120 129 -12082
rect 187 -12082 225 -12066
rect 269 -12066 285 -12048
rect 387 -12048 463 -12032
rect 387 -12066 403 -12048
rect 269 -12082 307 -12066
rect 187 -12120 307 -12082
rect 365 -12082 403 -12066
rect 447 -12066 463 -12048
rect 565 -12048 641 -12032
rect 565 -12066 581 -12048
rect 447 -12082 485 -12066
rect 365 -12120 485 -12082
rect 543 -12082 581 -12066
rect 625 -12066 641 -12048
rect 743 -12048 819 -12032
rect 743 -12066 759 -12048
rect 625 -12082 663 -12066
rect 543 -12120 663 -12082
rect 721 -12082 759 -12066
rect 803 -12066 819 -12048
rect 921 -12048 997 -12032
rect 921 -12066 937 -12048
rect 803 -12082 841 -12066
rect 721 -12120 841 -12082
rect 899 -12082 937 -12066
rect 981 -12066 997 -12048
rect 1099 -12048 1175 -12032
rect 1099 -12066 1115 -12048
rect 981 -12082 1019 -12066
rect 899 -12120 1019 -12082
rect 1077 -12082 1115 -12066
rect 1159 -12066 1175 -12048
rect 1277 -12048 1353 -12032
rect 1277 -12066 1293 -12048
rect 1159 -12082 1197 -12066
rect 1077 -12120 1197 -12082
rect 1255 -12082 1293 -12066
rect 1337 -12066 1353 -12048
rect 1455 -12048 1531 -12032
rect 1455 -12066 1471 -12048
rect 1337 -12082 1375 -12066
rect 1255 -12120 1375 -12082
rect 1433 -12082 1471 -12066
rect 1515 -12066 1531 -12048
rect 1633 -12048 1709 -12032
rect 1633 -12066 1649 -12048
rect 1515 -12082 1553 -12066
rect 1433 -12120 1553 -12082
rect 1611 -12082 1649 -12066
rect 1693 -12066 1709 -12048
rect 1811 -12048 1887 -12032
rect 1811 -12066 1827 -12048
rect 1693 -12082 1731 -12066
rect 1611 -12120 1731 -12082
rect 1789 -12082 1827 -12066
rect 1871 -12066 1887 -12048
rect 1989 -12048 2065 -12032
rect 1989 -12066 2005 -12048
rect 1871 -12082 1909 -12066
rect 1789 -12120 1909 -12082
rect 1967 -12082 2005 -12066
rect 2049 -12066 2065 -12048
rect 2167 -12048 2243 -12032
rect 2167 -12066 2183 -12048
rect 2049 -12082 2087 -12066
rect 1967 -12120 2087 -12082
rect 2145 -12082 2183 -12066
rect 2227 -12066 2243 -12048
rect 2345 -12048 2421 -12032
rect 2345 -12066 2361 -12048
rect 2227 -12082 2265 -12066
rect 2145 -12120 2265 -12082
rect 2323 -12082 2361 -12066
rect 2405 -12066 2421 -12048
rect 2523 -12048 2599 -12032
rect 2523 -12066 2539 -12048
rect 2405 -12082 2443 -12066
rect 2323 -12120 2443 -12082
rect 2501 -12082 2539 -12066
rect 2583 -12066 2599 -12048
rect 2701 -12048 2777 -12032
rect 2701 -12066 2717 -12048
rect 2583 -12082 2621 -12066
rect 2501 -12120 2621 -12082
rect 2679 -12082 2717 -12066
rect 2761 -12066 2777 -12048
rect 2879 -12048 2955 -12032
rect 2879 -12066 2895 -12048
rect 2761 -12082 2799 -12066
rect 2679 -12120 2799 -12082
rect 2857 -12082 2895 -12066
rect 2939 -12066 2955 -12048
rect 3057 -12048 3133 -12032
rect 3057 -12066 3073 -12048
rect 2939 -12082 2977 -12066
rect 2857 -12120 2977 -12082
rect 3035 -12082 3073 -12066
rect 3117 -12066 3133 -12048
rect 3235 -12048 3311 -12032
rect 3235 -12066 3251 -12048
rect 3117 -12082 3155 -12066
rect 3035 -12120 3155 -12082
rect 3213 -12082 3251 -12066
rect 3295 -12066 3311 -12048
rect 3413 -12048 3489 -12032
rect 3413 -12066 3429 -12048
rect 3295 -12082 3333 -12066
rect 3213 -12120 3333 -12082
rect 3391 -12082 3429 -12066
rect 3473 -12066 3489 -12048
rect 3591 -12048 3667 -12032
rect 3591 -12066 3607 -12048
rect 3473 -12082 3511 -12066
rect 3391 -12120 3511 -12082
rect 3569 -12082 3607 -12066
rect 3651 -12066 3667 -12048
rect 3769 -12048 3845 -12032
rect 3769 -12066 3785 -12048
rect 3651 -12082 3689 -12066
rect 3569 -12120 3689 -12082
rect 3747 -12082 3785 -12066
rect 3829 -12066 3845 -12048
rect 3947 -12048 4023 -12032
rect 3947 -12066 3963 -12048
rect 3829 -12082 3867 -12066
rect 3747 -12120 3867 -12082
rect 3925 -12082 3963 -12066
rect 4007 -12066 4023 -12048
rect 4007 -12082 4045 -12066
rect 3925 -12120 4045 -12082
rect -2127 -12438 -2007 -12400
rect -2127 -12454 -2089 -12438
rect -2105 -12472 -2089 -12454
rect -2045 -12454 -2007 -12438
rect -1949 -12438 -1829 -12400
rect -1949 -12454 -1911 -12438
rect -2045 -12472 -2029 -12454
rect -2105 -12488 -2029 -12472
rect -1927 -12472 -1911 -12454
rect -1867 -12454 -1829 -12438
rect -1771 -12438 -1651 -12400
rect -1771 -12454 -1733 -12438
rect -1867 -12472 -1851 -12454
rect -1927 -12488 -1851 -12472
rect -1749 -12472 -1733 -12454
rect -1689 -12454 -1651 -12438
rect -1593 -12438 -1473 -12400
rect -1593 -12454 -1555 -12438
rect -1689 -12472 -1673 -12454
rect -1749 -12488 -1673 -12472
rect -1571 -12472 -1555 -12454
rect -1511 -12454 -1473 -12438
rect -1415 -12438 -1295 -12400
rect -1415 -12454 -1377 -12438
rect -1511 -12472 -1495 -12454
rect -1571 -12488 -1495 -12472
rect -1393 -12472 -1377 -12454
rect -1333 -12454 -1295 -12438
rect -1237 -12438 -1117 -12400
rect -1237 -12454 -1199 -12438
rect -1333 -12472 -1317 -12454
rect -1393 -12488 -1317 -12472
rect -1215 -12472 -1199 -12454
rect -1155 -12454 -1117 -12438
rect -1059 -12438 -939 -12400
rect -1059 -12454 -1021 -12438
rect -1155 -12472 -1139 -12454
rect -1215 -12488 -1139 -12472
rect -1037 -12472 -1021 -12454
rect -977 -12454 -939 -12438
rect -881 -12438 -761 -12400
rect -881 -12454 -843 -12438
rect -977 -12472 -961 -12454
rect -1037 -12488 -961 -12472
rect -859 -12472 -843 -12454
rect -799 -12454 -761 -12438
rect -703 -12438 -583 -12400
rect -703 -12454 -665 -12438
rect -799 -12472 -783 -12454
rect -859 -12488 -783 -12472
rect -681 -12472 -665 -12454
rect -621 -12454 -583 -12438
rect -525 -12438 -405 -12400
rect -525 -12454 -487 -12438
rect -621 -12472 -605 -12454
rect -681 -12488 -605 -12472
rect -503 -12472 -487 -12454
rect -443 -12454 -405 -12438
rect -347 -12438 -227 -12400
rect -347 -12454 -309 -12438
rect -443 -12472 -427 -12454
rect -503 -12488 -427 -12472
rect -325 -12472 -309 -12454
rect -265 -12454 -227 -12438
rect -169 -12438 -49 -12400
rect -169 -12454 -131 -12438
rect -265 -12472 -249 -12454
rect -325 -12488 -249 -12472
rect -147 -12472 -131 -12454
rect -87 -12454 -49 -12438
rect 9 -12438 129 -12400
rect 9 -12454 47 -12438
rect -87 -12472 -71 -12454
rect -147 -12488 -71 -12472
rect 31 -12472 47 -12454
rect 91 -12454 129 -12438
rect 187 -12438 307 -12400
rect 187 -12454 225 -12438
rect 91 -12472 107 -12454
rect 31 -12488 107 -12472
rect 209 -12472 225 -12454
rect 269 -12454 307 -12438
rect 365 -12438 485 -12400
rect 365 -12454 403 -12438
rect 269 -12472 285 -12454
rect 209 -12488 285 -12472
rect 387 -12472 403 -12454
rect 447 -12454 485 -12438
rect 543 -12438 663 -12400
rect 543 -12454 581 -12438
rect 447 -12472 463 -12454
rect 387 -12488 463 -12472
rect 565 -12472 581 -12454
rect 625 -12454 663 -12438
rect 721 -12438 841 -12400
rect 721 -12454 759 -12438
rect 625 -12472 641 -12454
rect 565 -12488 641 -12472
rect 743 -12472 759 -12454
rect 803 -12454 841 -12438
rect 899 -12438 1019 -12400
rect 899 -12454 937 -12438
rect 803 -12472 819 -12454
rect 743 -12488 819 -12472
rect 921 -12472 937 -12454
rect 981 -12454 1019 -12438
rect 1077 -12438 1197 -12400
rect 1077 -12454 1115 -12438
rect 981 -12472 997 -12454
rect 921 -12488 997 -12472
rect 1099 -12472 1115 -12454
rect 1159 -12454 1197 -12438
rect 1255 -12438 1375 -12400
rect 1255 -12454 1293 -12438
rect 1159 -12472 1175 -12454
rect 1099 -12488 1175 -12472
rect 1277 -12472 1293 -12454
rect 1337 -12454 1375 -12438
rect 1433 -12438 1553 -12400
rect 1433 -12454 1471 -12438
rect 1337 -12472 1353 -12454
rect 1277 -12488 1353 -12472
rect 1455 -12472 1471 -12454
rect 1515 -12454 1553 -12438
rect 1611 -12438 1731 -12400
rect 1611 -12454 1649 -12438
rect 1515 -12472 1531 -12454
rect 1455 -12488 1531 -12472
rect 1633 -12472 1649 -12454
rect 1693 -12454 1731 -12438
rect 1789 -12438 1909 -12400
rect 1789 -12454 1827 -12438
rect 1693 -12472 1709 -12454
rect 1633 -12488 1709 -12472
rect 1811 -12472 1827 -12454
rect 1871 -12454 1909 -12438
rect 1967 -12438 2087 -12400
rect 1967 -12454 2005 -12438
rect 1871 -12472 1887 -12454
rect 1811 -12488 1887 -12472
rect 1989 -12472 2005 -12454
rect 2049 -12454 2087 -12438
rect 2145 -12438 2265 -12400
rect 2145 -12454 2183 -12438
rect 2049 -12472 2065 -12454
rect 1989 -12488 2065 -12472
rect 2167 -12472 2183 -12454
rect 2227 -12454 2265 -12438
rect 2323 -12438 2443 -12400
rect 2323 -12454 2361 -12438
rect 2227 -12472 2243 -12454
rect 2167 -12488 2243 -12472
rect 2345 -12472 2361 -12454
rect 2405 -12454 2443 -12438
rect 2501 -12438 2621 -12400
rect 2501 -12454 2539 -12438
rect 2405 -12472 2421 -12454
rect 2345 -12488 2421 -12472
rect 2523 -12472 2539 -12454
rect 2583 -12454 2621 -12438
rect 2679 -12438 2799 -12400
rect 2679 -12454 2717 -12438
rect 2583 -12472 2599 -12454
rect 2523 -12488 2599 -12472
rect 2701 -12472 2717 -12454
rect 2761 -12454 2799 -12438
rect 2857 -12438 2977 -12400
rect 2857 -12454 2895 -12438
rect 2761 -12472 2777 -12454
rect 2701 -12488 2777 -12472
rect 2879 -12472 2895 -12454
rect 2939 -12454 2977 -12438
rect 3035 -12438 3155 -12400
rect 3035 -12454 3073 -12438
rect 2939 -12472 2955 -12454
rect 2879 -12488 2955 -12472
rect 3057 -12472 3073 -12454
rect 3117 -12454 3155 -12438
rect 3213 -12438 3333 -12400
rect 3213 -12454 3251 -12438
rect 3117 -12472 3133 -12454
rect 3057 -12488 3133 -12472
rect 3235 -12472 3251 -12454
rect 3295 -12454 3333 -12438
rect 3391 -12438 3511 -12400
rect 3391 -12454 3429 -12438
rect 3295 -12472 3311 -12454
rect 3235 -12488 3311 -12472
rect 3413 -12472 3429 -12454
rect 3473 -12454 3511 -12438
rect 3569 -12438 3689 -12400
rect 3569 -12454 3607 -12438
rect 3473 -12472 3489 -12454
rect 3413 -12488 3489 -12472
rect 3591 -12472 3607 -12454
rect 3651 -12454 3689 -12438
rect 3747 -12438 3867 -12400
rect 3747 -12454 3785 -12438
rect 3651 -12472 3667 -12454
rect 3591 -12488 3667 -12472
rect 3769 -12472 3785 -12454
rect 3829 -12454 3867 -12438
rect 3925 -12438 4045 -12400
rect 3925 -12454 3963 -12438
rect 3829 -12472 3845 -12454
rect 3769 -12488 3845 -12472
rect 3947 -12472 3963 -12454
rect 4007 -12454 4045 -12438
rect 4007 -12472 4023 -12454
rect 3947 -12488 4023 -12472
rect -5883 -12628 -5817 -12612
rect -5883 -12662 -5867 -12628
rect -5833 -12662 -5817 -12628
rect -5883 -12678 -5817 -12662
rect -5633 -12628 -5567 -12612
rect -5633 -12662 -5617 -12628
rect -5583 -12662 -5567 -12628
rect -5633 -12678 -5567 -12662
rect -5383 -12628 -5317 -12612
rect -5383 -12662 -5367 -12628
rect -5333 -12662 -5317 -12628
rect -5383 -12678 -5317 -12662
rect -5133 -12628 -5067 -12612
rect -5133 -12662 -5117 -12628
rect -5083 -12662 -5067 -12628
rect -5133 -12678 -5067 -12662
rect -4883 -12628 -4817 -12612
rect -4883 -12662 -4867 -12628
rect -4833 -12662 -4817 -12628
rect -4883 -12678 -4817 -12662
rect -4633 -12628 -4567 -12612
rect -4633 -12662 -4617 -12628
rect -4583 -12662 -4567 -12628
rect -4633 -12678 -4567 -12662
rect -4383 -12628 -4317 -12612
rect -4383 -12662 -4367 -12628
rect -4333 -12662 -4317 -12628
rect -4383 -12678 -4317 -12662
rect -4133 -12628 -4067 -12612
rect -4133 -12662 -4117 -12628
rect -4083 -12662 -4067 -12628
rect -4133 -12678 -4067 -12662
rect -5871 -12700 -5829 -12678
rect -5621 -12700 -5579 -12678
rect -5371 -12700 -5329 -12678
rect -5121 -12700 -5079 -12678
rect -4871 -12700 -4829 -12678
rect -4621 -12700 -4579 -12678
rect -4371 -12700 -4329 -12678
rect -4121 -12700 -4079 -12678
rect -5871 -12962 -5829 -12940
rect -5621 -12962 -5579 -12940
rect -5371 -12962 -5329 -12940
rect -5121 -12962 -5079 -12940
rect -4871 -12962 -4829 -12940
rect -4621 -12962 -4579 -12940
rect -4371 -12962 -4329 -12940
rect -4121 -12962 -4079 -12940
rect -5883 -12978 -5817 -12962
rect -5883 -13012 -5867 -12978
rect -5833 -13012 -5817 -12978
rect -5883 -13028 -5817 -13012
rect -5633 -12978 -5567 -12962
rect -5633 -13012 -5617 -12978
rect -5583 -13012 -5567 -12978
rect -5633 -13028 -5567 -13012
rect -5383 -12978 -5317 -12962
rect -5383 -13012 -5367 -12978
rect -5333 -13012 -5317 -12978
rect -5383 -13028 -5317 -13012
rect -5133 -12978 -5067 -12962
rect -5133 -13012 -5117 -12978
rect -5083 -13012 -5067 -12978
rect -5133 -13028 -5067 -13012
rect -4883 -12978 -4817 -12962
rect -4883 -13012 -4867 -12978
rect -4833 -13012 -4817 -12978
rect -4883 -13028 -4817 -13012
rect -4633 -12978 -4567 -12962
rect -4633 -13012 -4617 -12978
rect -4583 -13012 -4567 -12978
rect -4633 -13028 -4567 -13012
rect -4383 -12978 -4317 -12962
rect -4383 -13012 -4367 -12978
rect -4333 -13012 -4317 -12978
rect -4383 -13028 -4317 -13012
rect -4133 -12978 -4067 -12962
rect -4133 -13012 -4117 -12978
rect -4083 -13012 -4067 -12978
rect -4133 -13028 -4067 -13012
rect -2105 -13048 -2029 -13032
rect -2105 -13066 -2089 -13048
rect -2127 -13082 -2089 -13066
rect -2045 -13066 -2029 -13048
rect -1927 -13048 -1851 -13032
rect -1927 -13066 -1911 -13048
rect -2045 -13082 -2007 -13066
rect -2127 -13120 -2007 -13082
rect -1949 -13082 -1911 -13066
rect -1867 -13066 -1851 -13048
rect -1749 -13048 -1673 -13032
rect -1749 -13066 -1733 -13048
rect -1867 -13082 -1829 -13066
rect -1949 -13120 -1829 -13082
rect -1771 -13082 -1733 -13066
rect -1689 -13066 -1673 -13048
rect -1571 -13048 -1495 -13032
rect -1571 -13066 -1555 -13048
rect -1689 -13082 -1651 -13066
rect -1771 -13120 -1651 -13082
rect -1593 -13082 -1555 -13066
rect -1511 -13066 -1495 -13048
rect -1393 -13048 -1317 -13032
rect -1393 -13066 -1377 -13048
rect -1511 -13082 -1473 -13066
rect -1593 -13120 -1473 -13082
rect -1415 -13082 -1377 -13066
rect -1333 -13066 -1317 -13048
rect -1215 -13048 -1139 -13032
rect -1215 -13066 -1199 -13048
rect -1333 -13082 -1295 -13066
rect -1415 -13120 -1295 -13082
rect -1237 -13082 -1199 -13066
rect -1155 -13066 -1139 -13048
rect -1037 -13048 -961 -13032
rect -1037 -13066 -1021 -13048
rect -1155 -13082 -1117 -13066
rect -1237 -13120 -1117 -13082
rect -1059 -13082 -1021 -13066
rect -977 -13066 -961 -13048
rect -859 -13048 -783 -13032
rect -859 -13066 -843 -13048
rect -977 -13082 -939 -13066
rect -1059 -13120 -939 -13082
rect -881 -13082 -843 -13066
rect -799 -13066 -783 -13048
rect -681 -13048 -605 -13032
rect -681 -13066 -665 -13048
rect -799 -13082 -761 -13066
rect -881 -13120 -761 -13082
rect -703 -13082 -665 -13066
rect -621 -13066 -605 -13048
rect -503 -13048 -427 -13032
rect -503 -13066 -487 -13048
rect -621 -13082 -583 -13066
rect -703 -13120 -583 -13082
rect -525 -13082 -487 -13066
rect -443 -13066 -427 -13048
rect -325 -13048 -249 -13032
rect -325 -13066 -309 -13048
rect -443 -13082 -405 -13066
rect -525 -13120 -405 -13082
rect -347 -13082 -309 -13066
rect -265 -13066 -249 -13048
rect -147 -13048 -71 -13032
rect -147 -13066 -131 -13048
rect -265 -13082 -227 -13066
rect -347 -13120 -227 -13082
rect -169 -13082 -131 -13066
rect -87 -13066 -71 -13048
rect 31 -13048 107 -13032
rect 31 -13066 47 -13048
rect -87 -13082 -49 -13066
rect -169 -13120 -49 -13082
rect 9 -13082 47 -13066
rect 91 -13066 107 -13048
rect 209 -13048 285 -13032
rect 209 -13066 225 -13048
rect 91 -13082 129 -13066
rect 9 -13120 129 -13082
rect 187 -13082 225 -13066
rect 269 -13066 285 -13048
rect 387 -13048 463 -13032
rect 387 -13066 403 -13048
rect 269 -13082 307 -13066
rect 187 -13120 307 -13082
rect 365 -13082 403 -13066
rect 447 -13066 463 -13048
rect 565 -13048 641 -13032
rect 565 -13066 581 -13048
rect 447 -13082 485 -13066
rect 365 -13120 485 -13082
rect 543 -13082 581 -13066
rect 625 -13066 641 -13048
rect 743 -13048 819 -13032
rect 743 -13066 759 -13048
rect 625 -13082 663 -13066
rect 543 -13120 663 -13082
rect 721 -13082 759 -13066
rect 803 -13066 819 -13048
rect 921 -13048 997 -13032
rect 921 -13066 937 -13048
rect 803 -13082 841 -13066
rect 721 -13120 841 -13082
rect 899 -13082 937 -13066
rect 981 -13066 997 -13048
rect 1099 -13048 1175 -13032
rect 1099 -13066 1115 -13048
rect 981 -13082 1019 -13066
rect 899 -13120 1019 -13082
rect 1077 -13082 1115 -13066
rect 1159 -13066 1175 -13048
rect 1277 -13048 1353 -13032
rect 1277 -13066 1293 -13048
rect 1159 -13082 1197 -13066
rect 1077 -13120 1197 -13082
rect 1255 -13082 1293 -13066
rect 1337 -13066 1353 -13048
rect 1455 -13048 1531 -13032
rect 1455 -13066 1471 -13048
rect 1337 -13082 1375 -13066
rect 1255 -13120 1375 -13082
rect 1433 -13082 1471 -13066
rect 1515 -13066 1531 -13048
rect 1633 -13048 1709 -13032
rect 1633 -13066 1649 -13048
rect 1515 -13082 1553 -13066
rect 1433 -13120 1553 -13082
rect 1611 -13082 1649 -13066
rect 1693 -13066 1709 -13048
rect 1811 -13048 1887 -13032
rect 1811 -13066 1827 -13048
rect 1693 -13082 1731 -13066
rect 1611 -13120 1731 -13082
rect 1789 -13082 1827 -13066
rect 1871 -13066 1887 -13048
rect 1989 -13048 2065 -13032
rect 1989 -13066 2005 -13048
rect 1871 -13082 1909 -13066
rect 1789 -13120 1909 -13082
rect 1967 -13082 2005 -13066
rect 2049 -13066 2065 -13048
rect 2167 -13048 2243 -13032
rect 2167 -13066 2183 -13048
rect 2049 -13082 2087 -13066
rect 1967 -13120 2087 -13082
rect 2145 -13082 2183 -13066
rect 2227 -13066 2243 -13048
rect 2345 -13048 2421 -13032
rect 2345 -13066 2361 -13048
rect 2227 -13082 2265 -13066
rect 2145 -13120 2265 -13082
rect 2323 -13082 2361 -13066
rect 2405 -13066 2421 -13048
rect 2523 -13048 2599 -13032
rect 2523 -13066 2539 -13048
rect 2405 -13082 2443 -13066
rect 2323 -13120 2443 -13082
rect 2501 -13082 2539 -13066
rect 2583 -13066 2599 -13048
rect 2701 -13048 2777 -13032
rect 2701 -13066 2717 -13048
rect 2583 -13082 2621 -13066
rect 2501 -13120 2621 -13082
rect 2679 -13082 2717 -13066
rect 2761 -13066 2777 -13048
rect 2879 -13048 2955 -13032
rect 2879 -13066 2895 -13048
rect 2761 -13082 2799 -13066
rect 2679 -13120 2799 -13082
rect 2857 -13082 2895 -13066
rect 2939 -13066 2955 -13048
rect 3057 -13048 3133 -13032
rect 3057 -13066 3073 -13048
rect 2939 -13082 2977 -13066
rect 2857 -13120 2977 -13082
rect 3035 -13082 3073 -13066
rect 3117 -13066 3133 -13048
rect 3235 -13048 3311 -13032
rect 3235 -13066 3251 -13048
rect 3117 -13082 3155 -13066
rect 3035 -13120 3155 -13082
rect 3213 -13082 3251 -13066
rect 3295 -13066 3311 -13048
rect 3413 -13048 3489 -13032
rect 3413 -13066 3429 -13048
rect 3295 -13082 3333 -13066
rect 3213 -13120 3333 -13082
rect 3391 -13082 3429 -13066
rect 3473 -13066 3489 -13048
rect 3591 -13048 3667 -13032
rect 3591 -13066 3607 -13048
rect 3473 -13082 3511 -13066
rect 3391 -13120 3511 -13082
rect 3569 -13082 3607 -13066
rect 3651 -13066 3667 -13048
rect 3769 -13048 3845 -13032
rect 3769 -13066 3785 -13048
rect 3651 -13082 3689 -13066
rect 3569 -13120 3689 -13082
rect 3747 -13082 3785 -13066
rect 3829 -13066 3845 -13048
rect 3947 -13048 4023 -13032
rect 3947 -13066 3963 -13048
rect 3829 -13082 3867 -13066
rect 3747 -13120 3867 -13082
rect 3925 -13082 3963 -13066
rect 4007 -13066 4023 -13048
rect 4007 -13082 4045 -13066
rect 3925 -13120 4045 -13082
rect -5883 -13308 -5817 -13292
rect -5883 -13342 -5867 -13308
rect -5833 -13342 -5817 -13308
rect -5883 -13358 -5817 -13342
rect -5633 -13308 -5567 -13292
rect -5633 -13342 -5617 -13308
rect -5583 -13342 -5567 -13308
rect -5633 -13358 -5567 -13342
rect -5383 -13308 -5317 -13292
rect -5383 -13342 -5367 -13308
rect -5333 -13342 -5317 -13308
rect -5383 -13358 -5317 -13342
rect -5133 -13308 -5067 -13292
rect -5133 -13342 -5117 -13308
rect -5083 -13342 -5067 -13308
rect -5133 -13358 -5067 -13342
rect -4883 -13308 -4817 -13292
rect -4883 -13342 -4867 -13308
rect -4833 -13342 -4817 -13308
rect -4883 -13358 -4817 -13342
rect -4633 -13308 -4567 -13292
rect -4633 -13342 -4617 -13308
rect -4583 -13342 -4567 -13308
rect -4633 -13358 -4567 -13342
rect -4383 -13308 -4317 -13292
rect -4383 -13342 -4367 -13308
rect -4333 -13342 -4317 -13308
rect -4383 -13358 -4317 -13342
rect -4133 -13308 -4067 -13292
rect -4133 -13342 -4117 -13308
rect -4083 -13342 -4067 -13308
rect -4133 -13358 -4067 -13342
rect -5871 -13380 -5829 -13358
rect -5621 -13380 -5579 -13358
rect -5371 -13380 -5329 -13358
rect -5121 -13380 -5079 -13358
rect -4871 -13380 -4829 -13358
rect -4621 -13380 -4579 -13358
rect -4371 -13380 -4329 -13358
rect -4121 -13380 -4079 -13358
rect -2127 -13438 -2007 -13400
rect -2127 -13454 -2089 -13438
rect -2105 -13472 -2089 -13454
rect -2045 -13454 -2007 -13438
rect -1949 -13438 -1829 -13400
rect -1949 -13454 -1911 -13438
rect -2045 -13472 -2029 -13454
rect -2105 -13488 -2029 -13472
rect -1927 -13472 -1911 -13454
rect -1867 -13454 -1829 -13438
rect -1771 -13438 -1651 -13400
rect -1771 -13454 -1733 -13438
rect -1867 -13472 -1851 -13454
rect -1927 -13488 -1851 -13472
rect -1749 -13472 -1733 -13454
rect -1689 -13454 -1651 -13438
rect -1593 -13438 -1473 -13400
rect -1593 -13454 -1555 -13438
rect -1689 -13472 -1673 -13454
rect -1749 -13488 -1673 -13472
rect -1571 -13472 -1555 -13454
rect -1511 -13454 -1473 -13438
rect -1415 -13438 -1295 -13400
rect -1415 -13454 -1377 -13438
rect -1511 -13472 -1495 -13454
rect -1571 -13488 -1495 -13472
rect -1393 -13472 -1377 -13454
rect -1333 -13454 -1295 -13438
rect -1237 -13438 -1117 -13400
rect -1237 -13454 -1199 -13438
rect -1333 -13472 -1317 -13454
rect -1393 -13488 -1317 -13472
rect -1215 -13472 -1199 -13454
rect -1155 -13454 -1117 -13438
rect -1059 -13438 -939 -13400
rect -1059 -13454 -1021 -13438
rect -1155 -13472 -1139 -13454
rect -1215 -13488 -1139 -13472
rect -1037 -13472 -1021 -13454
rect -977 -13454 -939 -13438
rect -881 -13438 -761 -13400
rect -881 -13454 -843 -13438
rect -977 -13472 -961 -13454
rect -1037 -13488 -961 -13472
rect -859 -13472 -843 -13454
rect -799 -13454 -761 -13438
rect -703 -13438 -583 -13400
rect -703 -13454 -665 -13438
rect -799 -13472 -783 -13454
rect -859 -13488 -783 -13472
rect -681 -13472 -665 -13454
rect -621 -13454 -583 -13438
rect -525 -13438 -405 -13400
rect -525 -13454 -487 -13438
rect -621 -13472 -605 -13454
rect -681 -13488 -605 -13472
rect -503 -13472 -487 -13454
rect -443 -13454 -405 -13438
rect -347 -13438 -227 -13400
rect -347 -13454 -309 -13438
rect -443 -13472 -427 -13454
rect -503 -13488 -427 -13472
rect -325 -13472 -309 -13454
rect -265 -13454 -227 -13438
rect -169 -13438 -49 -13400
rect -169 -13454 -131 -13438
rect -265 -13472 -249 -13454
rect -325 -13488 -249 -13472
rect -147 -13472 -131 -13454
rect -87 -13454 -49 -13438
rect 9 -13438 129 -13400
rect 9 -13454 47 -13438
rect -87 -13472 -71 -13454
rect -147 -13488 -71 -13472
rect 31 -13472 47 -13454
rect 91 -13454 129 -13438
rect 187 -13438 307 -13400
rect 187 -13454 225 -13438
rect 91 -13472 107 -13454
rect 31 -13488 107 -13472
rect 209 -13472 225 -13454
rect 269 -13454 307 -13438
rect 365 -13438 485 -13400
rect 365 -13454 403 -13438
rect 269 -13472 285 -13454
rect 209 -13488 285 -13472
rect 387 -13472 403 -13454
rect 447 -13454 485 -13438
rect 543 -13438 663 -13400
rect 543 -13454 581 -13438
rect 447 -13472 463 -13454
rect 387 -13488 463 -13472
rect 565 -13472 581 -13454
rect 625 -13454 663 -13438
rect 721 -13438 841 -13400
rect 721 -13454 759 -13438
rect 625 -13472 641 -13454
rect 565 -13488 641 -13472
rect 743 -13472 759 -13454
rect 803 -13454 841 -13438
rect 899 -13438 1019 -13400
rect 899 -13454 937 -13438
rect 803 -13472 819 -13454
rect 743 -13488 819 -13472
rect 921 -13472 937 -13454
rect 981 -13454 1019 -13438
rect 1077 -13438 1197 -13400
rect 1077 -13454 1115 -13438
rect 981 -13472 997 -13454
rect 921 -13488 997 -13472
rect 1099 -13472 1115 -13454
rect 1159 -13454 1197 -13438
rect 1255 -13438 1375 -13400
rect 1255 -13454 1293 -13438
rect 1159 -13472 1175 -13454
rect 1099 -13488 1175 -13472
rect 1277 -13472 1293 -13454
rect 1337 -13454 1375 -13438
rect 1433 -13438 1553 -13400
rect 1433 -13454 1471 -13438
rect 1337 -13472 1353 -13454
rect 1277 -13488 1353 -13472
rect 1455 -13472 1471 -13454
rect 1515 -13454 1553 -13438
rect 1611 -13438 1731 -13400
rect 1611 -13454 1649 -13438
rect 1515 -13472 1531 -13454
rect 1455 -13488 1531 -13472
rect 1633 -13472 1649 -13454
rect 1693 -13454 1731 -13438
rect 1789 -13438 1909 -13400
rect 1789 -13454 1827 -13438
rect 1693 -13472 1709 -13454
rect 1633 -13488 1709 -13472
rect 1811 -13472 1827 -13454
rect 1871 -13454 1909 -13438
rect 1967 -13438 2087 -13400
rect 1967 -13454 2005 -13438
rect 1871 -13472 1887 -13454
rect 1811 -13488 1887 -13472
rect 1989 -13472 2005 -13454
rect 2049 -13454 2087 -13438
rect 2145 -13438 2265 -13400
rect 2145 -13454 2183 -13438
rect 2049 -13472 2065 -13454
rect 1989 -13488 2065 -13472
rect 2167 -13472 2183 -13454
rect 2227 -13454 2265 -13438
rect 2323 -13438 2443 -13400
rect 2323 -13454 2361 -13438
rect 2227 -13472 2243 -13454
rect 2167 -13488 2243 -13472
rect 2345 -13472 2361 -13454
rect 2405 -13454 2443 -13438
rect 2501 -13438 2621 -13400
rect 2501 -13454 2539 -13438
rect 2405 -13472 2421 -13454
rect 2345 -13488 2421 -13472
rect 2523 -13472 2539 -13454
rect 2583 -13454 2621 -13438
rect 2679 -13438 2799 -13400
rect 2679 -13454 2717 -13438
rect 2583 -13472 2599 -13454
rect 2523 -13488 2599 -13472
rect 2701 -13472 2717 -13454
rect 2761 -13454 2799 -13438
rect 2857 -13438 2977 -13400
rect 2857 -13454 2895 -13438
rect 2761 -13472 2777 -13454
rect 2701 -13488 2777 -13472
rect 2879 -13472 2895 -13454
rect 2939 -13454 2977 -13438
rect 3035 -13438 3155 -13400
rect 3035 -13454 3073 -13438
rect 2939 -13472 2955 -13454
rect 2879 -13488 2955 -13472
rect 3057 -13472 3073 -13454
rect 3117 -13454 3155 -13438
rect 3213 -13438 3333 -13400
rect 3213 -13454 3251 -13438
rect 3117 -13472 3133 -13454
rect 3057 -13488 3133 -13472
rect 3235 -13472 3251 -13454
rect 3295 -13454 3333 -13438
rect 3391 -13438 3511 -13400
rect 3391 -13454 3429 -13438
rect 3295 -13472 3311 -13454
rect 3235 -13488 3311 -13472
rect 3413 -13472 3429 -13454
rect 3473 -13454 3511 -13438
rect 3569 -13438 3689 -13400
rect 3569 -13454 3607 -13438
rect 3473 -13472 3489 -13454
rect 3413 -13488 3489 -13472
rect 3591 -13472 3607 -13454
rect 3651 -13454 3689 -13438
rect 3747 -13438 3867 -13400
rect 3747 -13454 3785 -13438
rect 3651 -13472 3667 -13454
rect 3591 -13488 3667 -13472
rect 3769 -13472 3785 -13454
rect 3829 -13454 3867 -13438
rect 3925 -13438 4045 -13400
rect 3925 -13454 3963 -13438
rect 3829 -13472 3845 -13454
rect 3769 -13488 3845 -13472
rect 3947 -13472 3963 -13454
rect 4007 -13454 4045 -13438
rect 4007 -13472 4023 -13454
rect 3947 -13488 4023 -13472
rect -5871 -13642 -5829 -13620
rect -5621 -13642 -5579 -13620
rect -5371 -13642 -5329 -13620
rect -5121 -13642 -5079 -13620
rect -4871 -13642 -4829 -13620
rect -4621 -13642 -4579 -13620
rect -4371 -13642 -4329 -13620
rect -4121 -13642 -4079 -13620
rect -5883 -13658 -5817 -13642
rect -5883 -13692 -5867 -13658
rect -5833 -13692 -5817 -13658
rect -5883 -13708 -5817 -13692
rect -5633 -13658 -5567 -13642
rect -5633 -13692 -5617 -13658
rect -5583 -13692 -5567 -13658
rect -5633 -13708 -5567 -13692
rect -5383 -13658 -5317 -13642
rect -5383 -13692 -5367 -13658
rect -5333 -13692 -5317 -13658
rect -5383 -13708 -5317 -13692
rect -5133 -13658 -5067 -13642
rect -5133 -13692 -5117 -13658
rect -5083 -13692 -5067 -13658
rect -5133 -13708 -5067 -13692
rect -4883 -13658 -4817 -13642
rect -4883 -13692 -4867 -13658
rect -4833 -13692 -4817 -13658
rect -4883 -13708 -4817 -13692
rect -4633 -13658 -4567 -13642
rect -4633 -13692 -4617 -13658
rect -4583 -13692 -4567 -13658
rect -4633 -13708 -4567 -13692
rect -4383 -13658 -4317 -13642
rect -4383 -13692 -4367 -13658
rect -4333 -13692 -4317 -13658
rect -4383 -13708 -4317 -13692
rect -4133 -13658 -4067 -13642
rect -4133 -13692 -4117 -13658
rect -4083 -13692 -4067 -13658
rect -4133 -13708 -4067 -13692
rect -2105 -14048 -2029 -14032
rect -2105 -14066 -2089 -14048
rect -2127 -14082 -2089 -14066
rect -2045 -14066 -2029 -14048
rect -1927 -14048 -1851 -14032
rect -1927 -14066 -1911 -14048
rect -2045 -14082 -2007 -14066
rect -2127 -14120 -2007 -14082
rect -1949 -14082 -1911 -14066
rect -1867 -14066 -1851 -14048
rect -1749 -14048 -1673 -14032
rect -1749 -14066 -1733 -14048
rect -1867 -14082 -1829 -14066
rect -1949 -14120 -1829 -14082
rect -1771 -14082 -1733 -14066
rect -1689 -14066 -1673 -14048
rect -1571 -14048 -1495 -14032
rect -1571 -14066 -1555 -14048
rect -1689 -14082 -1651 -14066
rect -1771 -14120 -1651 -14082
rect -1593 -14082 -1555 -14066
rect -1511 -14066 -1495 -14048
rect -1393 -14048 -1317 -14032
rect -1393 -14066 -1377 -14048
rect -1511 -14082 -1473 -14066
rect -1593 -14120 -1473 -14082
rect -1415 -14082 -1377 -14066
rect -1333 -14066 -1317 -14048
rect -1215 -14048 -1139 -14032
rect -1215 -14066 -1199 -14048
rect -1333 -14082 -1295 -14066
rect -1415 -14120 -1295 -14082
rect -1237 -14082 -1199 -14066
rect -1155 -14066 -1139 -14048
rect -1037 -14048 -961 -14032
rect -1037 -14066 -1021 -14048
rect -1155 -14082 -1117 -14066
rect -1237 -14120 -1117 -14082
rect -1059 -14082 -1021 -14066
rect -977 -14066 -961 -14048
rect -859 -14048 -783 -14032
rect -859 -14066 -843 -14048
rect -977 -14082 -939 -14066
rect -1059 -14120 -939 -14082
rect -881 -14082 -843 -14066
rect -799 -14066 -783 -14048
rect -681 -14048 -605 -14032
rect -681 -14066 -665 -14048
rect -799 -14082 -761 -14066
rect -881 -14120 -761 -14082
rect -703 -14082 -665 -14066
rect -621 -14066 -605 -14048
rect -503 -14048 -427 -14032
rect -503 -14066 -487 -14048
rect -621 -14082 -583 -14066
rect -703 -14120 -583 -14082
rect -525 -14082 -487 -14066
rect -443 -14066 -427 -14048
rect -325 -14048 -249 -14032
rect -325 -14066 -309 -14048
rect -443 -14082 -405 -14066
rect -525 -14120 -405 -14082
rect -347 -14082 -309 -14066
rect -265 -14066 -249 -14048
rect -147 -14048 -71 -14032
rect -147 -14066 -131 -14048
rect -265 -14082 -227 -14066
rect -347 -14120 -227 -14082
rect -169 -14082 -131 -14066
rect -87 -14066 -71 -14048
rect 31 -14048 107 -14032
rect 31 -14066 47 -14048
rect -87 -14082 -49 -14066
rect -169 -14120 -49 -14082
rect 9 -14082 47 -14066
rect 91 -14066 107 -14048
rect 209 -14048 285 -14032
rect 209 -14066 225 -14048
rect 91 -14082 129 -14066
rect 9 -14120 129 -14082
rect 187 -14082 225 -14066
rect 269 -14066 285 -14048
rect 387 -14048 463 -14032
rect 387 -14066 403 -14048
rect 269 -14082 307 -14066
rect 187 -14120 307 -14082
rect 365 -14082 403 -14066
rect 447 -14066 463 -14048
rect 565 -14048 641 -14032
rect 565 -14066 581 -14048
rect 447 -14082 485 -14066
rect 365 -14120 485 -14082
rect 543 -14082 581 -14066
rect 625 -14066 641 -14048
rect 743 -14048 819 -14032
rect 743 -14066 759 -14048
rect 625 -14082 663 -14066
rect 543 -14120 663 -14082
rect 721 -14082 759 -14066
rect 803 -14066 819 -14048
rect 921 -14048 997 -14032
rect 921 -14066 937 -14048
rect 803 -14082 841 -14066
rect 721 -14120 841 -14082
rect 899 -14082 937 -14066
rect 981 -14066 997 -14048
rect 1099 -14048 1175 -14032
rect 1099 -14066 1115 -14048
rect 981 -14082 1019 -14066
rect 899 -14120 1019 -14082
rect 1077 -14082 1115 -14066
rect 1159 -14066 1175 -14048
rect 1277 -14048 1353 -14032
rect 1277 -14066 1293 -14048
rect 1159 -14082 1197 -14066
rect 1077 -14120 1197 -14082
rect 1255 -14082 1293 -14066
rect 1337 -14066 1353 -14048
rect 1455 -14048 1531 -14032
rect 1455 -14066 1471 -14048
rect 1337 -14082 1375 -14066
rect 1255 -14120 1375 -14082
rect 1433 -14082 1471 -14066
rect 1515 -14066 1531 -14048
rect 1633 -14048 1709 -14032
rect 1633 -14066 1649 -14048
rect 1515 -14082 1553 -14066
rect 1433 -14120 1553 -14082
rect 1611 -14082 1649 -14066
rect 1693 -14066 1709 -14048
rect 1811 -14048 1887 -14032
rect 1811 -14066 1827 -14048
rect 1693 -14082 1731 -14066
rect 1611 -14120 1731 -14082
rect 1789 -14082 1827 -14066
rect 1871 -14066 1887 -14048
rect 1989 -14048 2065 -14032
rect 1989 -14066 2005 -14048
rect 1871 -14082 1909 -14066
rect 1789 -14120 1909 -14082
rect 1967 -14082 2005 -14066
rect 2049 -14066 2065 -14048
rect 2167 -14048 2243 -14032
rect 2167 -14066 2183 -14048
rect 2049 -14082 2087 -14066
rect 1967 -14120 2087 -14082
rect 2145 -14082 2183 -14066
rect 2227 -14066 2243 -14048
rect 2345 -14048 2421 -14032
rect 2345 -14066 2361 -14048
rect 2227 -14082 2265 -14066
rect 2145 -14120 2265 -14082
rect 2323 -14082 2361 -14066
rect 2405 -14066 2421 -14048
rect 2523 -14048 2599 -14032
rect 2523 -14066 2539 -14048
rect 2405 -14082 2443 -14066
rect 2323 -14120 2443 -14082
rect 2501 -14082 2539 -14066
rect 2583 -14066 2599 -14048
rect 2701 -14048 2777 -14032
rect 2701 -14066 2717 -14048
rect 2583 -14082 2621 -14066
rect 2501 -14120 2621 -14082
rect 2679 -14082 2717 -14066
rect 2761 -14066 2777 -14048
rect 2879 -14048 2955 -14032
rect 2879 -14066 2895 -14048
rect 2761 -14082 2799 -14066
rect 2679 -14120 2799 -14082
rect 2857 -14082 2895 -14066
rect 2939 -14066 2955 -14048
rect 3057 -14048 3133 -14032
rect 3057 -14066 3073 -14048
rect 2939 -14082 2977 -14066
rect 2857 -14120 2977 -14082
rect 3035 -14082 3073 -14066
rect 3117 -14066 3133 -14048
rect 3235 -14048 3311 -14032
rect 3235 -14066 3251 -14048
rect 3117 -14082 3155 -14066
rect 3035 -14120 3155 -14082
rect 3213 -14082 3251 -14066
rect 3295 -14066 3311 -14048
rect 3413 -14048 3489 -14032
rect 3413 -14066 3429 -14048
rect 3295 -14082 3333 -14066
rect 3213 -14120 3333 -14082
rect 3391 -14082 3429 -14066
rect 3473 -14066 3489 -14048
rect 3591 -14048 3667 -14032
rect 3591 -14066 3607 -14048
rect 3473 -14082 3511 -14066
rect 3391 -14120 3511 -14082
rect 3569 -14082 3607 -14066
rect 3651 -14066 3667 -14048
rect 3769 -14048 3845 -14032
rect 3769 -14066 3785 -14048
rect 3651 -14082 3689 -14066
rect 3569 -14120 3689 -14082
rect 3747 -14082 3785 -14066
rect 3829 -14066 3845 -14048
rect 3947 -14048 4023 -14032
rect 3947 -14066 3963 -14048
rect 3829 -14082 3867 -14066
rect 3747 -14120 3867 -14082
rect 3925 -14082 3963 -14066
rect 4007 -14066 4023 -14048
rect 5645 -14048 5721 -14032
rect 5645 -14066 5661 -14048
rect 4007 -14082 4045 -14066
rect 3925 -14120 4045 -14082
rect 5623 -14082 5661 -14066
rect 5705 -14066 5721 -14048
rect 5823 -14048 5899 -14032
rect 5823 -14066 5839 -14048
rect 5705 -14082 5743 -14066
rect 5623 -14120 5743 -14082
rect 5801 -14082 5839 -14066
rect 5883 -14066 5899 -14048
rect 6001 -14048 6077 -14032
rect 6001 -14066 6017 -14048
rect 5883 -14082 5921 -14066
rect 5801 -14120 5921 -14082
rect 5979 -14082 6017 -14066
rect 6061 -14066 6077 -14048
rect 6179 -14048 6255 -14032
rect 6179 -14066 6195 -14048
rect 6061 -14082 6099 -14066
rect 5979 -14120 6099 -14082
rect 6157 -14082 6195 -14066
rect 6239 -14066 6255 -14048
rect 6357 -14048 6433 -14032
rect 6357 -14066 6373 -14048
rect 6239 -14082 6277 -14066
rect 6157 -14120 6277 -14082
rect 6335 -14082 6373 -14066
rect 6417 -14066 6433 -14048
rect 6535 -14048 6611 -14032
rect 6535 -14066 6551 -14048
rect 6417 -14082 6455 -14066
rect 6335 -14120 6455 -14082
rect 6513 -14082 6551 -14066
rect 6595 -14066 6611 -14048
rect 6713 -14048 6789 -14032
rect 6713 -14066 6729 -14048
rect 6595 -14082 6633 -14066
rect 6513 -14120 6633 -14082
rect 6691 -14082 6729 -14066
rect 6773 -14066 6789 -14048
rect 6891 -14048 6967 -14032
rect 6891 -14066 6907 -14048
rect 6773 -14082 6811 -14066
rect 6691 -14120 6811 -14082
rect 6869 -14082 6907 -14066
rect 6951 -14066 6967 -14048
rect 7069 -14048 7145 -14032
rect 7069 -14066 7085 -14048
rect 6951 -14082 6989 -14066
rect 6869 -14120 6989 -14082
rect 7047 -14082 7085 -14066
rect 7129 -14066 7145 -14048
rect 7247 -14048 7323 -14032
rect 7247 -14066 7263 -14048
rect 7129 -14082 7167 -14066
rect 7047 -14120 7167 -14082
rect 7225 -14082 7263 -14066
rect 7307 -14066 7323 -14048
rect 7425 -14048 7501 -14032
rect 7425 -14066 7441 -14048
rect 7307 -14082 7345 -14066
rect 7225 -14120 7345 -14082
rect 7403 -14082 7441 -14066
rect 7485 -14066 7501 -14048
rect 7603 -14048 7679 -14032
rect 7603 -14066 7619 -14048
rect 7485 -14082 7523 -14066
rect 7403 -14120 7523 -14082
rect 7581 -14082 7619 -14066
rect 7663 -14066 7679 -14048
rect 7781 -14048 7857 -14032
rect 7781 -14066 7797 -14048
rect 7663 -14082 7701 -14066
rect 7581 -14120 7701 -14082
rect 7759 -14082 7797 -14066
rect 7841 -14066 7857 -14048
rect 7959 -14048 8035 -14032
rect 7959 -14066 7975 -14048
rect 7841 -14082 7879 -14066
rect 7759 -14120 7879 -14082
rect 7937 -14082 7975 -14066
rect 8019 -14066 8035 -14048
rect 8137 -14048 8213 -14032
rect 8137 -14066 8153 -14048
rect 8019 -14082 8057 -14066
rect 7937 -14120 8057 -14082
rect 8115 -14082 8153 -14066
rect 8197 -14066 8213 -14048
rect 8315 -14048 8391 -14032
rect 8315 -14066 8331 -14048
rect 8197 -14082 8235 -14066
rect 8115 -14120 8235 -14082
rect 8293 -14082 8331 -14066
rect 8375 -14066 8391 -14048
rect 8493 -14048 8569 -14032
rect 8493 -14066 8509 -14048
rect 8375 -14082 8413 -14066
rect 8293 -14120 8413 -14082
rect 8471 -14082 8509 -14066
rect 8553 -14066 8569 -14048
rect 8671 -14048 8747 -14032
rect 8671 -14066 8687 -14048
rect 8553 -14082 8591 -14066
rect 8471 -14120 8591 -14082
rect 8649 -14082 8687 -14066
rect 8731 -14066 8747 -14048
rect 8849 -14048 8925 -14032
rect 8849 -14066 8865 -14048
rect 8731 -14082 8769 -14066
rect 8649 -14120 8769 -14082
rect 8827 -14082 8865 -14066
rect 8909 -14066 8925 -14048
rect 9027 -14048 9103 -14032
rect 9027 -14066 9043 -14048
rect 8909 -14082 8947 -14066
rect 8827 -14120 8947 -14082
rect 9005 -14082 9043 -14066
rect 9087 -14066 9103 -14048
rect 9205 -14048 9281 -14032
rect 9205 -14066 9221 -14048
rect 9087 -14082 9125 -14066
rect 9005 -14120 9125 -14082
rect 9183 -14082 9221 -14066
rect 9265 -14066 9281 -14048
rect 9383 -14048 9459 -14032
rect 9383 -14066 9399 -14048
rect 9265 -14082 9303 -14066
rect 9183 -14120 9303 -14082
rect 9361 -14082 9399 -14066
rect 9443 -14066 9459 -14048
rect 9561 -14048 9637 -14032
rect 9561 -14066 9577 -14048
rect 9443 -14082 9481 -14066
rect 9361 -14120 9481 -14082
rect 9539 -14082 9577 -14066
rect 9621 -14066 9637 -14048
rect 9739 -14048 9815 -14032
rect 9739 -14066 9755 -14048
rect 9621 -14082 9659 -14066
rect 9539 -14120 9659 -14082
rect 9717 -14082 9755 -14066
rect 9799 -14066 9815 -14048
rect 9917 -14048 9993 -14032
rect 9917 -14066 9933 -14048
rect 9799 -14082 9837 -14066
rect 9717 -14120 9837 -14082
rect 9895 -14082 9933 -14066
rect 9977 -14066 9993 -14048
rect 10095 -14048 10171 -14032
rect 10095 -14066 10111 -14048
rect 9977 -14082 10015 -14066
rect 9895 -14120 10015 -14082
rect 10073 -14082 10111 -14066
rect 10155 -14066 10171 -14048
rect 10273 -14048 10349 -14032
rect 10273 -14066 10289 -14048
rect 10155 -14082 10193 -14066
rect 10073 -14120 10193 -14082
rect 10251 -14082 10289 -14066
rect 10333 -14066 10349 -14048
rect 10451 -14048 10527 -14032
rect 10451 -14066 10467 -14048
rect 10333 -14082 10371 -14066
rect 10251 -14120 10371 -14082
rect 10429 -14082 10467 -14066
rect 10511 -14066 10527 -14048
rect 10629 -14048 10705 -14032
rect 10629 -14066 10645 -14048
rect 10511 -14082 10549 -14066
rect 10429 -14120 10549 -14082
rect 10607 -14082 10645 -14066
rect 10689 -14066 10705 -14048
rect 10807 -14048 10883 -14032
rect 10807 -14066 10823 -14048
rect 10689 -14082 10727 -14066
rect 10607 -14120 10727 -14082
rect 10785 -14082 10823 -14066
rect 10867 -14066 10883 -14048
rect 10985 -14048 11061 -14032
rect 10985 -14066 11001 -14048
rect 10867 -14082 10905 -14066
rect 10785 -14120 10905 -14082
rect 10963 -14082 11001 -14066
rect 11045 -14066 11061 -14048
rect 11163 -14048 11239 -14032
rect 11163 -14066 11179 -14048
rect 11045 -14082 11083 -14066
rect 10963 -14120 11083 -14082
rect 11141 -14082 11179 -14066
rect 11223 -14066 11239 -14048
rect 11341 -14048 11417 -14032
rect 11341 -14066 11357 -14048
rect 11223 -14082 11261 -14066
rect 11141 -14120 11261 -14082
rect 11319 -14082 11357 -14066
rect 11401 -14066 11417 -14048
rect 11519 -14048 11595 -14032
rect 11519 -14066 11535 -14048
rect 11401 -14082 11439 -14066
rect 11319 -14120 11439 -14082
rect 11497 -14082 11535 -14066
rect 11579 -14066 11595 -14048
rect 11697 -14048 11773 -14032
rect 11697 -14066 11713 -14048
rect 11579 -14082 11617 -14066
rect 11497 -14120 11617 -14082
rect 11675 -14082 11713 -14066
rect 11757 -14066 11773 -14048
rect 11875 -14048 11951 -14032
rect 11875 -14066 11891 -14048
rect 11757 -14082 11795 -14066
rect 11675 -14120 11795 -14082
rect 11853 -14082 11891 -14066
rect 11935 -14066 11951 -14048
rect 12053 -14048 12129 -14032
rect 12053 -14066 12069 -14048
rect 11935 -14082 11973 -14066
rect 11853 -14120 11973 -14082
rect 12031 -14082 12069 -14066
rect 12113 -14066 12129 -14048
rect 12231 -14048 12307 -14032
rect 12231 -14066 12247 -14048
rect 12113 -14082 12151 -14066
rect 12031 -14120 12151 -14082
rect 12209 -14082 12247 -14066
rect 12291 -14066 12307 -14048
rect 12409 -14048 12485 -14032
rect 12409 -14066 12425 -14048
rect 12291 -14082 12329 -14066
rect 12209 -14120 12329 -14082
rect 12387 -14082 12425 -14066
rect 12469 -14066 12485 -14048
rect 12587 -14048 12663 -14032
rect 12587 -14066 12603 -14048
rect 12469 -14082 12507 -14066
rect 12387 -14120 12507 -14082
rect 12565 -14082 12603 -14066
rect 12647 -14066 12663 -14048
rect 12647 -14082 12685 -14066
rect 12565 -14120 12685 -14082
rect -5960 -14310 -5884 -14294
rect -5960 -14328 -5944 -14310
rect -5982 -14344 -5944 -14328
rect -5900 -14328 -5884 -14310
rect -5782 -14310 -5706 -14294
rect -5782 -14328 -5766 -14310
rect -5900 -14344 -5862 -14328
rect -5982 -14382 -5862 -14344
rect -5804 -14344 -5766 -14328
rect -5722 -14328 -5706 -14310
rect -5604 -14310 -5528 -14294
rect -5604 -14328 -5588 -14310
rect -5722 -14344 -5684 -14328
rect -5804 -14382 -5684 -14344
rect -5626 -14344 -5588 -14328
rect -5544 -14328 -5528 -14310
rect -5426 -14310 -5350 -14294
rect -5426 -14328 -5410 -14310
rect -5544 -14344 -5506 -14328
rect -5626 -14382 -5506 -14344
rect -5448 -14344 -5410 -14328
rect -5366 -14328 -5350 -14310
rect -5248 -14310 -5172 -14294
rect -5248 -14328 -5232 -14310
rect -5366 -14344 -5328 -14328
rect -5448 -14382 -5328 -14344
rect -5270 -14344 -5232 -14328
rect -5188 -14328 -5172 -14310
rect -5070 -14310 -4994 -14294
rect -5070 -14328 -5054 -14310
rect -5188 -14344 -5150 -14328
rect -5270 -14382 -5150 -14344
rect -5092 -14344 -5054 -14328
rect -5010 -14328 -4994 -14310
rect -4892 -14310 -4816 -14294
rect -4892 -14328 -4876 -14310
rect -5010 -14344 -4972 -14328
rect -5092 -14382 -4972 -14344
rect -4914 -14344 -4876 -14328
rect -4832 -14328 -4816 -14310
rect -4714 -14310 -4638 -14294
rect -4714 -14328 -4698 -14310
rect -4832 -14344 -4794 -14328
rect -4914 -14382 -4794 -14344
rect -4736 -14344 -4698 -14328
rect -4654 -14328 -4638 -14310
rect -4536 -14310 -4460 -14294
rect -4536 -14328 -4520 -14310
rect -4654 -14344 -4616 -14328
rect -4736 -14382 -4616 -14344
rect -4558 -14344 -4520 -14328
rect -4476 -14328 -4460 -14310
rect -4358 -14310 -4282 -14294
rect -4358 -14328 -4342 -14310
rect -4476 -14344 -4438 -14328
rect -4558 -14382 -4438 -14344
rect -4380 -14344 -4342 -14328
rect -4298 -14328 -4282 -14310
rect -4180 -14310 -4104 -14294
rect -4180 -14328 -4164 -14310
rect -4298 -14344 -4260 -14328
rect -4380 -14382 -4260 -14344
rect -4202 -14344 -4164 -14328
rect -4120 -14328 -4104 -14310
rect -4120 -14344 -4082 -14328
rect -4202 -14382 -4082 -14344
rect -2127 -14438 -2007 -14400
rect -2127 -14454 -2089 -14438
rect -2105 -14472 -2089 -14454
rect -2045 -14454 -2007 -14438
rect -1949 -14438 -1829 -14400
rect -1949 -14454 -1911 -14438
rect -2045 -14472 -2029 -14454
rect -2105 -14488 -2029 -14472
rect -1927 -14472 -1911 -14454
rect -1867 -14454 -1829 -14438
rect -1771 -14438 -1651 -14400
rect -1771 -14454 -1733 -14438
rect -1867 -14472 -1851 -14454
rect -1927 -14488 -1851 -14472
rect -1749 -14472 -1733 -14454
rect -1689 -14454 -1651 -14438
rect -1593 -14438 -1473 -14400
rect -1593 -14454 -1555 -14438
rect -1689 -14472 -1673 -14454
rect -1749 -14488 -1673 -14472
rect -1571 -14472 -1555 -14454
rect -1511 -14454 -1473 -14438
rect -1415 -14438 -1295 -14400
rect -1415 -14454 -1377 -14438
rect -1511 -14472 -1495 -14454
rect -1571 -14488 -1495 -14472
rect -1393 -14472 -1377 -14454
rect -1333 -14454 -1295 -14438
rect -1237 -14438 -1117 -14400
rect -1237 -14454 -1199 -14438
rect -1333 -14472 -1317 -14454
rect -1393 -14488 -1317 -14472
rect -1215 -14472 -1199 -14454
rect -1155 -14454 -1117 -14438
rect -1059 -14438 -939 -14400
rect -1059 -14454 -1021 -14438
rect -1155 -14472 -1139 -14454
rect -1215 -14488 -1139 -14472
rect -1037 -14472 -1021 -14454
rect -977 -14454 -939 -14438
rect -881 -14438 -761 -14400
rect -881 -14454 -843 -14438
rect -977 -14472 -961 -14454
rect -1037 -14488 -961 -14472
rect -859 -14472 -843 -14454
rect -799 -14454 -761 -14438
rect -703 -14438 -583 -14400
rect -703 -14454 -665 -14438
rect -799 -14472 -783 -14454
rect -859 -14488 -783 -14472
rect -681 -14472 -665 -14454
rect -621 -14454 -583 -14438
rect -525 -14438 -405 -14400
rect -525 -14454 -487 -14438
rect -621 -14472 -605 -14454
rect -681 -14488 -605 -14472
rect -503 -14472 -487 -14454
rect -443 -14454 -405 -14438
rect -347 -14438 -227 -14400
rect -347 -14454 -309 -14438
rect -443 -14472 -427 -14454
rect -503 -14488 -427 -14472
rect -325 -14472 -309 -14454
rect -265 -14454 -227 -14438
rect -169 -14438 -49 -14400
rect -169 -14454 -131 -14438
rect -265 -14472 -249 -14454
rect -325 -14488 -249 -14472
rect -147 -14472 -131 -14454
rect -87 -14454 -49 -14438
rect 9 -14438 129 -14400
rect 9 -14454 47 -14438
rect -87 -14472 -71 -14454
rect -147 -14488 -71 -14472
rect 31 -14472 47 -14454
rect 91 -14454 129 -14438
rect 187 -14438 307 -14400
rect 187 -14454 225 -14438
rect 91 -14472 107 -14454
rect 31 -14488 107 -14472
rect 209 -14472 225 -14454
rect 269 -14454 307 -14438
rect 365 -14438 485 -14400
rect 365 -14454 403 -14438
rect 269 -14472 285 -14454
rect 209 -14488 285 -14472
rect 387 -14472 403 -14454
rect 447 -14454 485 -14438
rect 543 -14438 663 -14400
rect 543 -14454 581 -14438
rect 447 -14472 463 -14454
rect 387 -14488 463 -14472
rect 565 -14472 581 -14454
rect 625 -14454 663 -14438
rect 721 -14438 841 -14400
rect 721 -14454 759 -14438
rect 625 -14472 641 -14454
rect 565 -14488 641 -14472
rect 743 -14472 759 -14454
rect 803 -14454 841 -14438
rect 899 -14438 1019 -14400
rect 899 -14454 937 -14438
rect 803 -14472 819 -14454
rect 743 -14488 819 -14472
rect 921 -14472 937 -14454
rect 981 -14454 1019 -14438
rect 1077 -14438 1197 -14400
rect 1077 -14454 1115 -14438
rect 981 -14472 997 -14454
rect 921 -14488 997 -14472
rect 1099 -14472 1115 -14454
rect 1159 -14454 1197 -14438
rect 1255 -14438 1375 -14400
rect 1255 -14454 1293 -14438
rect 1159 -14472 1175 -14454
rect 1099 -14488 1175 -14472
rect 1277 -14472 1293 -14454
rect 1337 -14454 1375 -14438
rect 1433 -14438 1553 -14400
rect 1433 -14454 1471 -14438
rect 1337 -14472 1353 -14454
rect 1277 -14488 1353 -14472
rect 1455 -14472 1471 -14454
rect 1515 -14454 1553 -14438
rect 1611 -14438 1731 -14400
rect 1611 -14454 1649 -14438
rect 1515 -14472 1531 -14454
rect 1455 -14488 1531 -14472
rect 1633 -14472 1649 -14454
rect 1693 -14454 1731 -14438
rect 1789 -14438 1909 -14400
rect 1789 -14454 1827 -14438
rect 1693 -14472 1709 -14454
rect 1633 -14488 1709 -14472
rect 1811 -14472 1827 -14454
rect 1871 -14454 1909 -14438
rect 1967 -14438 2087 -14400
rect 1967 -14454 2005 -14438
rect 1871 -14472 1887 -14454
rect 1811 -14488 1887 -14472
rect 1989 -14472 2005 -14454
rect 2049 -14454 2087 -14438
rect 2145 -14438 2265 -14400
rect 2145 -14454 2183 -14438
rect 2049 -14472 2065 -14454
rect 1989 -14488 2065 -14472
rect 2167 -14472 2183 -14454
rect 2227 -14454 2265 -14438
rect 2323 -14438 2443 -14400
rect 2323 -14454 2361 -14438
rect 2227 -14472 2243 -14454
rect 2167 -14488 2243 -14472
rect 2345 -14472 2361 -14454
rect 2405 -14454 2443 -14438
rect 2501 -14438 2621 -14400
rect 2501 -14454 2539 -14438
rect 2405 -14472 2421 -14454
rect 2345 -14488 2421 -14472
rect 2523 -14472 2539 -14454
rect 2583 -14454 2621 -14438
rect 2679 -14438 2799 -14400
rect 2679 -14454 2717 -14438
rect 2583 -14472 2599 -14454
rect 2523 -14488 2599 -14472
rect 2701 -14472 2717 -14454
rect 2761 -14454 2799 -14438
rect 2857 -14438 2977 -14400
rect 2857 -14454 2895 -14438
rect 2761 -14472 2777 -14454
rect 2701 -14488 2777 -14472
rect 2879 -14472 2895 -14454
rect 2939 -14454 2977 -14438
rect 3035 -14438 3155 -14400
rect 3035 -14454 3073 -14438
rect 2939 -14472 2955 -14454
rect 2879 -14488 2955 -14472
rect 3057 -14472 3073 -14454
rect 3117 -14454 3155 -14438
rect 3213 -14438 3333 -14400
rect 3213 -14454 3251 -14438
rect 3117 -14472 3133 -14454
rect 3057 -14488 3133 -14472
rect 3235 -14472 3251 -14454
rect 3295 -14454 3333 -14438
rect 3391 -14438 3511 -14400
rect 3391 -14454 3429 -14438
rect 3295 -14472 3311 -14454
rect 3235 -14488 3311 -14472
rect 3413 -14472 3429 -14454
rect 3473 -14454 3511 -14438
rect 3569 -14438 3689 -14400
rect 3569 -14454 3607 -14438
rect 3473 -14472 3489 -14454
rect 3413 -14488 3489 -14472
rect 3591 -14472 3607 -14454
rect 3651 -14454 3689 -14438
rect 3747 -14438 3867 -14400
rect 3747 -14454 3785 -14438
rect 3651 -14472 3667 -14454
rect 3591 -14488 3667 -14472
rect 3769 -14472 3785 -14454
rect 3829 -14454 3867 -14438
rect 3925 -14438 4045 -14400
rect 3925 -14454 3963 -14438
rect 3829 -14472 3845 -14454
rect 3769 -14488 3845 -14472
rect 3947 -14472 3963 -14454
rect 4007 -14454 4045 -14438
rect 5623 -14438 5743 -14400
rect 5623 -14454 5661 -14438
rect 4007 -14472 4023 -14454
rect 3947 -14488 4023 -14472
rect 5645 -14472 5661 -14454
rect 5705 -14454 5743 -14438
rect 5801 -14438 5921 -14400
rect 5801 -14454 5839 -14438
rect 5705 -14472 5721 -14454
rect 5645 -14488 5721 -14472
rect 5823 -14472 5839 -14454
rect 5883 -14454 5921 -14438
rect 5979 -14438 6099 -14400
rect 5979 -14454 6017 -14438
rect 5883 -14472 5899 -14454
rect 5823 -14488 5899 -14472
rect 6001 -14472 6017 -14454
rect 6061 -14454 6099 -14438
rect 6157 -14438 6277 -14400
rect 6157 -14454 6195 -14438
rect 6061 -14472 6077 -14454
rect 6001 -14488 6077 -14472
rect 6179 -14472 6195 -14454
rect 6239 -14454 6277 -14438
rect 6335 -14438 6455 -14400
rect 6335 -14454 6373 -14438
rect 6239 -14472 6255 -14454
rect 6179 -14488 6255 -14472
rect 6357 -14472 6373 -14454
rect 6417 -14454 6455 -14438
rect 6513 -14438 6633 -14400
rect 6513 -14454 6551 -14438
rect 6417 -14472 6433 -14454
rect 6357 -14488 6433 -14472
rect 6535 -14472 6551 -14454
rect 6595 -14454 6633 -14438
rect 6691 -14438 6811 -14400
rect 6691 -14454 6729 -14438
rect 6595 -14472 6611 -14454
rect 6535 -14488 6611 -14472
rect 6713 -14472 6729 -14454
rect 6773 -14454 6811 -14438
rect 6869 -14438 6989 -14400
rect 6869 -14454 6907 -14438
rect 6773 -14472 6789 -14454
rect 6713 -14488 6789 -14472
rect 6891 -14472 6907 -14454
rect 6951 -14454 6989 -14438
rect 7047 -14438 7167 -14400
rect 7047 -14454 7085 -14438
rect 6951 -14472 6967 -14454
rect 6891 -14488 6967 -14472
rect 7069 -14472 7085 -14454
rect 7129 -14454 7167 -14438
rect 7225 -14438 7345 -14400
rect 7225 -14454 7263 -14438
rect 7129 -14472 7145 -14454
rect 7069 -14488 7145 -14472
rect 7247 -14472 7263 -14454
rect 7307 -14454 7345 -14438
rect 7403 -14438 7523 -14400
rect 7403 -14454 7441 -14438
rect 7307 -14472 7323 -14454
rect 7247 -14488 7323 -14472
rect 7425 -14472 7441 -14454
rect 7485 -14454 7523 -14438
rect 7581 -14438 7701 -14400
rect 7581 -14454 7619 -14438
rect 7485 -14472 7501 -14454
rect 7425 -14488 7501 -14472
rect 7603 -14472 7619 -14454
rect 7663 -14454 7701 -14438
rect 7759 -14438 7879 -14400
rect 7759 -14454 7797 -14438
rect 7663 -14472 7679 -14454
rect 7603 -14488 7679 -14472
rect 7781 -14472 7797 -14454
rect 7841 -14454 7879 -14438
rect 7937 -14438 8057 -14400
rect 7937 -14454 7975 -14438
rect 7841 -14472 7857 -14454
rect 7781 -14488 7857 -14472
rect 7959 -14472 7975 -14454
rect 8019 -14454 8057 -14438
rect 8115 -14438 8235 -14400
rect 8115 -14454 8153 -14438
rect 8019 -14472 8035 -14454
rect 7959 -14488 8035 -14472
rect 8137 -14472 8153 -14454
rect 8197 -14454 8235 -14438
rect 8293 -14438 8413 -14400
rect 8293 -14454 8331 -14438
rect 8197 -14472 8213 -14454
rect 8137 -14488 8213 -14472
rect 8315 -14472 8331 -14454
rect 8375 -14454 8413 -14438
rect 8471 -14438 8591 -14400
rect 8471 -14454 8509 -14438
rect 8375 -14472 8391 -14454
rect 8315 -14488 8391 -14472
rect 8493 -14472 8509 -14454
rect 8553 -14454 8591 -14438
rect 8649 -14438 8769 -14400
rect 8649 -14454 8687 -14438
rect 8553 -14472 8569 -14454
rect 8493 -14488 8569 -14472
rect 8671 -14472 8687 -14454
rect 8731 -14454 8769 -14438
rect 8827 -14438 8947 -14400
rect 8827 -14454 8865 -14438
rect 8731 -14472 8747 -14454
rect 8671 -14488 8747 -14472
rect 8849 -14472 8865 -14454
rect 8909 -14454 8947 -14438
rect 9005 -14438 9125 -14400
rect 9005 -14454 9043 -14438
rect 8909 -14472 8925 -14454
rect 8849 -14488 8925 -14472
rect 9027 -14472 9043 -14454
rect 9087 -14454 9125 -14438
rect 9183 -14438 9303 -14400
rect 9183 -14454 9221 -14438
rect 9087 -14472 9103 -14454
rect 9027 -14488 9103 -14472
rect 9205 -14472 9221 -14454
rect 9265 -14454 9303 -14438
rect 9361 -14438 9481 -14400
rect 9361 -14454 9399 -14438
rect 9265 -14472 9281 -14454
rect 9205 -14488 9281 -14472
rect 9383 -14472 9399 -14454
rect 9443 -14454 9481 -14438
rect 9539 -14438 9659 -14400
rect 9539 -14454 9577 -14438
rect 9443 -14472 9459 -14454
rect 9383 -14488 9459 -14472
rect 9561 -14472 9577 -14454
rect 9621 -14454 9659 -14438
rect 9717 -14438 9837 -14400
rect 9717 -14454 9755 -14438
rect 9621 -14472 9637 -14454
rect 9561 -14488 9637 -14472
rect 9739 -14472 9755 -14454
rect 9799 -14454 9837 -14438
rect 9895 -14438 10015 -14400
rect 9895 -14454 9933 -14438
rect 9799 -14472 9815 -14454
rect 9739 -14488 9815 -14472
rect 9917 -14472 9933 -14454
rect 9977 -14454 10015 -14438
rect 10073 -14438 10193 -14400
rect 10073 -14454 10111 -14438
rect 9977 -14472 9993 -14454
rect 9917 -14488 9993 -14472
rect 10095 -14472 10111 -14454
rect 10155 -14454 10193 -14438
rect 10251 -14438 10371 -14400
rect 10251 -14454 10289 -14438
rect 10155 -14472 10171 -14454
rect 10095 -14488 10171 -14472
rect 10273 -14472 10289 -14454
rect 10333 -14454 10371 -14438
rect 10429 -14438 10549 -14400
rect 10429 -14454 10467 -14438
rect 10333 -14472 10349 -14454
rect 10273 -14488 10349 -14472
rect 10451 -14472 10467 -14454
rect 10511 -14454 10549 -14438
rect 10607 -14438 10727 -14400
rect 10607 -14454 10645 -14438
rect 10511 -14472 10527 -14454
rect 10451 -14488 10527 -14472
rect 10629 -14472 10645 -14454
rect 10689 -14454 10727 -14438
rect 10785 -14438 10905 -14400
rect 10785 -14454 10823 -14438
rect 10689 -14472 10705 -14454
rect 10629 -14488 10705 -14472
rect 10807 -14472 10823 -14454
rect 10867 -14454 10905 -14438
rect 10963 -14438 11083 -14400
rect 10963 -14454 11001 -14438
rect 10867 -14472 10883 -14454
rect 10807 -14488 10883 -14472
rect 10985 -14472 11001 -14454
rect 11045 -14454 11083 -14438
rect 11141 -14438 11261 -14400
rect 11141 -14454 11179 -14438
rect 11045 -14472 11061 -14454
rect 10985 -14488 11061 -14472
rect 11163 -14472 11179 -14454
rect 11223 -14454 11261 -14438
rect 11319 -14438 11439 -14400
rect 11319 -14454 11357 -14438
rect 11223 -14472 11239 -14454
rect 11163 -14488 11239 -14472
rect 11341 -14472 11357 -14454
rect 11401 -14454 11439 -14438
rect 11497 -14438 11617 -14400
rect 11497 -14454 11535 -14438
rect 11401 -14472 11417 -14454
rect 11341 -14488 11417 -14472
rect 11519 -14472 11535 -14454
rect 11579 -14454 11617 -14438
rect 11675 -14438 11795 -14400
rect 11675 -14454 11713 -14438
rect 11579 -14472 11595 -14454
rect 11519 -14488 11595 -14472
rect 11697 -14472 11713 -14454
rect 11757 -14454 11795 -14438
rect 11853 -14438 11973 -14400
rect 11853 -14454 11891 -14438
rect 11757 -14472 11773 -14454
rect 11697 -14488 11773 -14472
rect 11875 -14472 11891 -14454
rect 11935 -14454 11973 -14438
rect 12031 -14438 12151 -14400
rect 12031 -14454 12069 -14438
rect 11935 -14472 11951 -14454
rect 11875 -14488 11951 -14472
rect 12053 -14472 12069 -14454
rect 12113 -14454 12151 -14438
rect 12209 -14438 12329 -14400
rect 12209 -14454 12247 -14438
rect 12113 -14472 12129 -14454
rect 12053 -14488 12129 -14472
rect 12231 -14472 12247 -14454
rect 12291 -14454 12329 -14438
rect 12387 -14438 12507 -14400
rect 12387 -14454 12425 -14438
rect 12291 -14472 12307 -14454
rect 12231 -14488 12307 -14472
rect 12409 -14472 12425 -14454
rect 12469 -14454 12507 -14438
rect 12565 -14438 12685 -14400
rect 12565 -14454 12603 -14438
rect 12469 -14472 12485 -14454
rect 12409 -14488 12485 -14472
rect 12587 -14472 12603 -14454
rect 12647 -14454 12685 -14438
rect 12647 -14472 12663 -14454
rect 12587 -14488 12663 -14472
rect -5982 -14700 -5862 -14662
rect -5982 -14716 -5944 -14700
rect -5960 -14734 -5944 -14716
rect -5900 -14716 -5862 -14700
rect -5804 -14700 -5684 -14662
rect -5804 -14716 -5766 -14700
rect -5900 -14734 -5884 -14716
rect -5960 -14750 -5884 -14734
rect -5782 -14734 -5766 -14716
rect -5722 -14716 -5684 -14700
rect -5626 -14700 -5506 -14662
rect -5626 -14716 -5588 -14700
rect -5722 -14734 -5706 -14716
rect -5782 -14750 -5706 -14734
rect -5604 -14734 -5588 -14716
rect -5544 -14716 -5506 -14700
rect -5448 -14700 -5328 -14662
rect -5448 -14716 -5410 -14700
rect -5544 -14734 -5528 -14716
rect -5604 -14750 -5528 -14734
rect -5426 -14734 -5410 -14716
rect -5366 -14716 -5328 -14700
rect -5270 -14700 -5150 -14662
rect -5270 -14716 -5232 -14700
rect -5366 -14734 -5350 -14716
rect -5426 -14750 -5350 -14734
rect -5248 -14734 -5232 -14716
rect -5188 -14716 -5150 -14700
rect -5092 -14700 -4972 -14662
rect -5092 -14716 -5054 -14700
rect -5188 -14734 -5172 -14716
rect -5248 -14750 -5172 -14734
rect -5070 -14734 -5054 -14716
rect -5010 -14716 -4972 -14700
rect -4914 -14700 -4794 -14662
rect -4914 -14716 -4876 -14700
rect -5010 -14734 -4994 -14716
rect -5070 -14750 -4994 -14734
rect -4892 -14734 -4876 -14716
rect -4832 -14716 -4794 -14700
rect -4736 -14700 -4616 -14662
rect -4736 -14716 -4698 -14700
rect -4832 -14734 -4816 -14716
rect -4892 -14750 -4816 -14734
rect -4714 -14734 -4698 -14716
rect -4654 -14716 -4616 -14700
rect -4558 -14700 -4438 -14662
rect -4558 -14716 -4520 -14700
rect -4654 -14734 -4638 -14716
rect -4714 -14750 -4638 -14734
rect -4536 -14734 -4520 -14716
rect -4476 -14716 -4438 -14700
rect -4380 -14700 -4260 -14662
rect -4380 -14716 -4342 -14700
rect -4476 -14734 -4460 -14716
rect -4536 -14750 -4460 -14734
rect -4358 -14734 -4342 -14716
rect -4298 -14716 -4260 -14700
rect -4202 -14700 -4082 -14662
rect -4202 -14716 -4164 -14700
rect -4298 -14734 -4282 -14716
rect -4358 -14750 -4282 -14734
rect -4180 -14734 -4164 -14716
rect -4120 -14716 -4082 -14700
rect -4120 -14734 -4104 -14716
rect -4180 -14750 -4104 -14734
rect -5960 -15010 -5884 -14994
rect -5960 -15028 -5944 -15010
rect -5982 -15044 -5944 -15028
rect -5900 -15028 -5884 -15010
rect -5782 -15010 -5706 -14994
rect -5782 -15028 -5766 -15010
rect -5900 -15044 -5862 -15028
rect -5982 -15082 -5862 -15044
rect -5804 -15044 -5766 -15028
rect -5722 -15028 -5706 -15010
rect -5604 -15010 -5528 -14994
rect -5604 -15028 -5588 -15010
rect -5722 -15044 -5684 -15028
rect -5804 -15082 -5684 -15044
rect -5626 -15044 -5588 -15028
rect -5544 -15028 -5528 -15010
rect -5426 -15010 -5350 -14994
rect -5426 -15028 -5410 -15010
rect -5544 -15044 -5506 -15028
rect -5626 -15082 -5506 -15044
rect -5448 -15044 -5410 -15028
rect -5366 -15028 -5350 -15010
rect -5248 -15010 -5172 -14994
rect -5248 -15028 -5232 -15010
rect -5366 -15044 -5328 -15028
rect -5448 -15082 -5328 -15044
rect -5270 -15044 -5232 -15028
rect -5188 -15028 -5172 -15010
rect -5070 -15010 -4994 -14994
rect -5070 -15028 -5054 -15010
rect -5188 -15044 -5150 -15028
rect -5270 -15082 -5150 -15044
rect -5092 -15044 -5054 -15028
rect -5010 -15028 -4994 -15010
rect -4892 -15010 -4816 -14994
rect -4892 -15028 -4876 -15010
rect -5010 -15044 -4972 -15028
rect -5092 -15082 -4972 -15044
rect -4914 -15044 -4876 -15028
rect -4832 -15028 -4816 -15010
rect -4714 -15010 -4638 -14994
rect -4714 -15028 -4698 -15010
rect -4832 -15044 -4794 -15028
rect -4914 -15082 -4794 -15044
rect -4736 -15044 -4698 -15028
rect -4654 -15028 -4638 -15010
rect -4536 -15010 -4460 -14994
rect -4536 -15028 -4520 -15010
rect -4654 -15044 -4616 -15028
rect -4736 -15082 -4616 -15044
rect -4558 -15044 -4520 -15028
rect -4476 -15028 -4460 -15010
rect -4358 -15010 -4282 -14994
rect -4358 -15028 -4342 -15010
rect -4476 -15044 -4438 -15028
rect -4558 -15082 -4438 -15044
rect -4380 -15044 -4342 -15028
rect -4298 -15028 -4282 -15010
rect -4180 -15010 -4104 -14994
rect -4180 -15028 -4164 -15010
rect -4298 -15044 -4260 -15028
rect -4380 -15082 -4260 -15044
rect -4202 -15044 -4164 -15028
rect -4120 -15028 -4104 -15010
rect -4120 -15044 -4082 -15028
rect -4202 -15082 -4082 -15044
rect -2105 -15048 -2029 -15032
rect -2105 -15066 -2089 -15048
rect -2127 -15082 -2089 -15066
rect -2045 -15066 -2029 -15048
rect -1927 -15048 -1851 -15032
rect -1927 -15066 -1911 -15048
rect -2045 -15082 -2007 -15066
rect -2127 -15120 -2007 -15082
rect -1949 -15082 -1911 -15066
rect -1867 -15066 -1851 -15048
rect -1749 -15048 -1673 -15032
rect -1749 -15066 -1733 -15048
rect -1867 -15082 -1829 -15066
rect -1949 -15120 -1829 -15082
rect -1771 -15082 -1733 -15066
rect -1689 -15066 -1673 -15048
rect -1571 -15048 -1495 -15032
rect -1571 -15066 -1555 -15048
rect -1689 -15082 -1651 -15066
rect -1771 -15120 -1651 -15082
rect -1593 -15082 -1555 -15066
rect -1511 -15066 -1495 -15048
rect -1393 -15048 -1317 -15032
rect -1393 -15066 -1377 -15048
rect -1511 -15082 -1473 -15066
rect -1593 -15120 -1473 -15082
rect -1415 -15082 -1377 -15066
rect -1333 -15066 -1317 -15048
rect -1215 -15048 -1139 -15032
rect -1215 -15066 -1199 -15048
rect -1333 -15082 -1295 -15066
rect -1415 -15120 -1295 -15082
rect -1237 -15082 -1199 -15066
rect -1155 -15066 -1139 -15048
rect -1037 -15048 -961 -15032
rect -1037 -15066 -1021 -15048
rect -1155 -15082 -1117 -15066
rect -1237 -15120 -1117 -15082
rect -1059 -15082 -1021 -15066
rect -977 -15066 -961 -15048
rect -859 -15048 -783 -15032
rect -859 -15066 -843 -15048
rect -977 -15082 -939 -15066
rect -1059 -15120 -939 -15082
rect -881 -15082 -843 -15066
rect -799 -15066 -783 -15048
rect -681 -15048 -605 -15032
rect -681 -15066 -665 -15048
rect -799 -15082 -761 -15066
rect -881 -15120 -761 -15082
rect -703 -15082 -665 -15066
rect -621 -15066 -605 -15048
rect -503 -15048 -427 -15032
rect -503 -15066 -487 -15048
rect -621 -15082 -583 -15066
rect -703 -15120 -583 -15082
rect -525 -15082 -487 -15066
rect -443 -15066 -427 -15048
rect -325 -15048 -249 -15032
rect -325 -15066 -309 -15048
rect -443 -15082 -405 -15066
rect -525 -15120 -405 -15082
rect -347 -15082 -309 -15066
rect -265 -15066 -249 -15048
rect -147 -15048 -71 -15032
rect -147 -15066 -131 -15048
rect -265 -15082 -227 -15066
rect -347 -15120 -227 -15082
rect -169 -15082 -131 -15066
rect -87 -15066 -71 -15048
rect 31 -15048 107 -15032
rect 31 -15066 47 -15048
rect -87 -15082 -49 -15066
rect -169 -15120 -49 -15082
rect 9 -15082 47 -15066
rect 91 -15066 107 -15048
rect 209 -15048 285 -15032
rect 209 -15066 225 -15048
rect 91 -15082 129 -15066
rect 9 -15120 129 -15082
rect 187 -15082 225 -15066
rect 269 -15066 285 -15048
rect 387 -15048 463 -15032
rect 387 -15066 403 -15048
rect 269 -15082 307 -15066
rect 187 -15120 307 -15082
rect 365 -15082 403 -15066
rect 447 -15066 463 -15048
rect 565 -15048 641 -15032
rect 565 -15066 581 -15048
rect 447 -15082 485 -15066
rect 365 -15120 485 -15082
rect 543 -15082 581 -15066
rect 625 -15066 641 -15048
rect 743 -15048 819 -15032
rect 743 -15066 759 -15048
rect 625 -15082 663 -15066
rect 543 -15120 663 -15082
rect 721 -15082 759 -15066
rect 803 -15066 819 -15048
rect 921 -15048 997 -15032
rect 921 -15066 937 -15048
rect 803 -15082 841 -15066
rect 721 -15120 841 -15082
rect 899 -15082 937 -15066
rect 981 -15066 997 -15048
rect 1099 -15048 1175 -15032
rect 1099 -15066 1115 -15048
rect 981 -15082 1019 -15066
rect 899 -15120 1019 -15082
rect 1077 -15082 1115 -15066
rect 1159 -15066 1175 -15048
rect 1277 -15048 1353 -15032
rect 1277 -15066 1293 -15048
rect 1159 -15082 1197 -15066
rect 1077 -15120 1197 -15082
rect 1255 -15082 1293 -15066
rect 1337 -15066 1353 -15048
rect 1455 -15048 1531 -15032
rect 1455 -15066 1471 -15048
rect 1337 -15082 1375 -15066
rect 1255 -15120 1375 -15082
rect 1433 -15082 1471 -15066
rect 1515 -15066 1531 -15048
rect 1633 -15048 1709 -15032
rect 1633 -15066 1649 -15048
rect 1515 -15082 1553 -15066
rect 1433 -15120 1553 -15082
rect 1611 -15082 1649 -15066
rect 1693 -15066 1709 -15048
rect 1811 -15048 1887 -15032
rect 1811 -15066 1827 -15048
rect 1693 -15082 1731 -15066
rect 1611 -15120 1731 -15082
rect 1789 -15082 1827 -15066
rect 1871 -15066 1887 -15048
rect 1989 -15048 2065 -15032
rect 1989 -15066 2005 -15048
rect 1871 -15082 1909 -15066
rect 1789 -15120 1909 -15082
rect 1967 -15082 2005 -15066
rect 2049 -15066 2065 -15048
rect 2167 -15048 2243 -15032
rect 2167 -15066 2183 -15048
rect 2049 -15082 2087 -15066
rect 1967 -15120 2087 -15082
rect 2145 -15082 2183 -15066
rect 2227 -15066 2243 -15048
rect 2345 -15048 2421 -15032
rect 2345 -15066 2361 -15048
rect 2227 -15082 2265 -15066
rect 2145 -15120 2265 -15082
rect 2323 -15082 2361 -15066
rect 2405 -15066 2421 -15048
rect 2523 -15048 2599 -15032
rect 2523 -15066 2539 -15048
rect 2405 -15082 2443 -15066
rect 2323 -15120 2443 -15082
rect 2501 -15082 2539 -15066
rect 2583 -15066 2599 -15048
rect 2701 -15048 2777 -15032
rect 2701 -15066 2717 -15048
rect 2583 -15082 2621 -15066
rect 2501 -15120 2621 -15082
rect 2679 -15082 2717 -15066
rect 2761 -15066 2777 -15048
rect 2879 -15048 2955 -15032
rect 2879 -15066 2895 -15048
rect 2761 -15082 2799 -15066
rect 2679 -15120 2799 -15082
rect 2857 -15082 2895 -15066
rect 2939 -15066 2955 -15048
rect 3057 -15048 3133 -15032
rect 3057 -15066 3073 -15048
rect 2939 -15082 2977 -15066
rect 2857 -15120 2977 -15082
rect 3035 -15082 3073 -15066
rect 3117 -15066 3133 -15048
rect 3235 -15048 3311 -15032
rect 3235 -15066 3251 -15048
rect 3117 -15082 3155 -15066
rect 3035 -15120 3155 -15082
rect 3213 -15082 3251 -15066
rect 3295 -15066 3311 -15048
rect 3413 -15048 3489 -15032
rect 3413 -15066 3429 -15048
rect 3295 -15082 3333 -15066
rect 3213 -15120 3333 -15082
rect 3391 -15082 3429 -15066
rect 3473 -15066 3489 -15048
rect 3591 -15048 3667 -15032
rect 3591 -15066 3607 -15048
rect 3473 -15082 3511 -15066
rect 3391 -15120 3511 -15082
rect 3569 -15082 3607 -15066
rect 3651 -15066 3667 -15048
rect 3769 -15048 3845 -15032
rect 3769 -15066 3785 -15048
rect 3651 -15082 3689 -15066
rect 3569 -15120 3689 -15082
rect 3747 -15082 3785 -15066
rect 3829 -15066 3845 -15048
rect 3947 -15048 4023 -15032
rect 3947 -15066 3963 -15048
rect 3829 -15082 3867 -15066
rect 3747 -15120 3867 -15082
rect 3925 -15082 3963 -15066
rect 4007 -15066 4023 -15048
rect 4007 -15082 4045 -15066
rect 5645 -15048 5721 -15032
rect 5645 -15066 5661 -15048
rect 3925 -15120 4045 -15082
rect 5623 -15082 5661 -15066
rect 5705 -15066 5721 -15048
rect 5823 -15048 5899 -15032
rect 5823 -15066 5839 -15048
rect 5705 -15082 5743 -15066
rect 5623 -15120 5743 -15082
rect 5801 -15082 5839 -15066
rect 5883 -15066 5899 -15048
rect 6001 -15048 6077 -15032
rect 6001 -15066 6017 -15048
rect 5883 -15082 5921 -15066
rect 5801 -15120 5921 -15082
rect 5979 -15082 6017 -15066
rect 6061 -15066 6077 -15048
rect 6179 -15048 6255 -15032
rect 6179 -15066 6195 -15048
rect 6061 -15082 6099 -15066
rect 5979 -15120 6099 -15082
rect 6157 -15082 6195 -15066
rect 6239 -15066 6255 -15048
rect 6357 -15048 6433 -15032
rect 6357 -15066 6373 -15048
rect 6239 -15082 6277 -15066
rect 6157 -15120 6277 -15082
rect 6335 -15082 6373 -15066
rect 6417 -15066 6433 -15048
rect 6535 -15048 6611 -15032
rect 6535 -15066 6551 -15048
rect 6417 -15082 6455 -15066
rect 6335 -15120 6455 -15082
rect 6513 -15082 6551 -15066
rect 6595 -15066 6611 -15048
rect 6713 -15048 6789 -15032
rect 6713 -15066 6729 -15048
rect 6595 -15082 6633 -15066
rect 6513 -15120 6633 -15082
rect 6691 -15082 6729 -15066
rect 6773 -15066 6789 -15048
rect 6891 -15048 6967 -15032
rect 6891 -15066 6907 -15048
rect 6773 -15082 6811 -15066
rect 6691 -15120 6811 -15082
rect 6869 -15082 6907 -15066
rect 6951 -15066 6967 -15048
rect 7069 -15048 7145 -15032
rect 7069 -15066 7085 -15048
rect 6951 -15082 6989 -15066
rect 6869 -15120 6989 -15082
rect 7047 -15082 7085 -15066
rect 7129 -15066 7145 -15048
rect 7247 -15048 7323 -15032
rect 7247 -15066 7263 -15048
rect 7129 -15082 7167 -15066
rect 7047 -15120 7167 -15082
rect 7225 -15082 7263 -15066
rect 7307 -15066 7323 -15048
rect 7425 -15048 7501 -15032
rect 7425 -15066 7441 -15048
rect 7307 -15082 7345 -15066
rect 7225 -15120 7345 -15082
rect 7403 -15082 7441 -15066
rect 7485 -15066 7501 -15048
rect 7603 -15048 7679 -15032
rect 7603 -15066 7619 -15048
rect 7485 -15082 7523 -15066
rect 7403 -15120 7523 -15082
rect 7581 -15082 7619 -15066
rect 7663 -15066 7679 -15048
rect 7781 -15048 7857 -15032
rect 7781 -15066 7797 -15048
rect 7663 -15082 7701 -15066
rect 7581 -15120 7701 -15082
rect 7759 -15082 7797 -15066
rect 7841 -15066 7857 -15048
rect 7959 -15048 8035 -15032
rect 7959 -15066 7975 -15048
rect 7841 -15082 7879 -15066
rect 7759 -15120 7879 -15082
rect 7937 -15082 7975 -15066
rect 8019 -15066 8035 -15048
rect 8137 -15048 8213 -15032
rect 8137 -15066 8153 -15048
rect 8019 -15082 8057 -15066
rect 7937 -15120 8057 -15082
rect 8115 -15082 8153 -15066
rect 8197 -15066 8213 -15048
rect 8315 -15048 8391 -15032
rect 8315 -15066 8331 -15048
rect 8197 -15082 8235 -15066
rect 8115 -15120 8235 -15082
rect 8293 -15082 8331 -15066
rect 8375 -15066 8391 -15048
rect 8493 -15048 8569 -15032
rect 8493 -15066 8509 -15048
rect 8375 -15082 8413 -15066
rect 8293 -15120 8413 -15082
rect 8471 -15082 8509 -15066
rect 8553 -15066 8569 -15048
rect 8671 -15048 8747 -15032
rect 8671 -15066 8687 -15048
rect 8553 -15082 8591 -15066
rect 8471 -15120 8591 -15082
rect 8649 -15082 8687 -15066
rect 8731 -15066 8747 -15048
rect 8849 -15048 8925 -15032
rect 8849 -15066 8865 -15048
rect 8731 -15082 8769 -15066
rect 8649 -15120 8769 -15082
rect 8827 -15082 8865 -15066
rect 8909 -15066 8925 -15048
rect 9027 -15048 9103 -15032
rect 9027 -15066 9043 -15048
rect 8909 -15082 8947 -15066
rect 8827 -15120 8947 -15082
rect 9005 -15082 9043 -15066
rect 9087 -15066 9103 -15048
rect 9205 -15048 9281 -15032
rect 9205 -15066 9221 -15048
rect 9087 -15082 9125 -15066
rect 9005 -15120 9125 -15082
rect 9183 -15082 9221 -15066
rect 9265 -15066 9281 -15048
rect 9383 -15048 9459 -15032
rect 9383 -15066 9399 -15048
rect 9265 -15082 9303 -15066
rect 9183 -15120 9303 -15082
rect 9361 -15082 9399 -15066
rect 9443 -15066 9459 -15048
rect 9561 -15048 9637 -15032
rect 9561 -15066 9577 -15048
rect 9443 -15082 9481 -15066
rect 9361 -15120 9481 -15082
rect 9539 -15082 9577 -15066
rect 9621 -15066 9637 -15048
rect 9739 -15048 9815 -15032
rect 9739 -15066 9755 -15048
rect 9621 -15082 9659 -15066
rect 9539 -15120 9659 -15082
rect 9717 -15082 9755 -15066
rect 9799 -15066 9815 -15048
rect 9917 -15048 9993 -15032
rect 9917 -15066 9933 -15048
rect 9799 -15082 9837 -15066
rect 9717 -15120 9837 -15082
rect 9895 -15082 9933 -15066
rect 9977 -15066 9993 -15048
rect 10095 -15048 10171 -15032
rect 10095 -15066 10111 -15048
rect 9977 -15082 10015 -15066
rect 9895 -15120 10015 -15082
rect 10073 -15082 10111 -15066
rect 10155 -15066 10171 -15048
rect 10273 -15048 10349 -15032
rect 10273 -15066 10289 -15048
rect 10155 -15082 10193 -15066
rect 10073 -15120 10193 -15082
rect 10251 -15082 10289 -15066
rect 10333 -15066 10349 -15048
rect 10451 -15048 10527 -15032
rect 10451 -15066 10467 -15048
rect 10333 -15082 10371 -15066
rect 10251 -15120 10371 -15082
rect 10429 -15082 10467 -15066
rect 10511 -15066 10527 -15048
rect 10629 -15048 10705 -15032
rect 10629 -15066 10645 -15048
rect 10511 -15082 10549 -15066
rect 10429 -15120 10549 -15082
rect 10607 -15082 10645 -15066
rect 10689 -15066 10705 -15048
rect 10807 -15048 10883 -15032
rect 10807 -15066 10823 -15048
rect 10689 -15082 10727 -15066
rect 10607 -15120 10727 -15082
rect 10785 -15082 10823 -15066
rect 10867 -15066 10883 -15048
rect 10985 -15048 11061 -15032
rect 10985 -15066 11001 -15048
rect 10867 -15082 10905 -15066
rect 10785 -15120 10905 -15082
rect 10963 -15082 11001 -15066
rect 11045 -15066 11061 -15048
rect 11163 -15048 11239 -15032
rect 11163 -15066 11179 -15048
rect 11045 -15082 11083 -15066
rect 10963 -15120 11083 -15082
rect 11141 -15082 11179 -15066
rect 11223 -15066 11239 -15048
rect 11341 -15048 11417 -15032
rect 11341 -15066 11357 -15048
rect 11223 -15082 11261 -15066
rect 11141 -15120 11261 -15082
rect 11319 -15082 11357 -15066
rect 11401 -15066 11417 -15048
rect 11519 -15048 11595 -15032
rect 11519 -15066 11535 -15048
rect 11401 -15082 11439 -15066
rect 11319 -15120 11439 -15082
rect 11497 -15082 11535 -15066
rect 11579 -15066 11595 -15048
rect 11697 -15048 11773 -15032
rect 11697 -15066 11713 -15048
rect 11579 -15082 11617 -15066
rect 11497 -15120 11617 -15082
rect 11675 -15082 11713 -15066
rect 11757 -15066 11773 -15048
rect 11875 -15048 11951 -15032
rect 11875 -15066 11891 -15048
rect 11757 -15082 11795 -15066
rect 11675 -15120 11795 -15082
rect 11853 -15082 11891 -15066
rect 11935 -15066 11951 -15048
rect 12053 -15048 12129 -15032
rect 12053 -15066 12069 -15048
rect 11935 -15082 11973 -15066
rect 11853 -15120 11973 -15082
rect 12031 -15082 12069 -15066
rect 12113 -15066 12129 -15048
rect 12231 -15048 12307 -15032
rect 12231 -15066 12247 -15048
rect 12113 -15082 12151 -15066
rect 12031 -15120 12151 -15082
rect 12209 -15082 12247 -15066
rect 12291 -15066 12307 -15048
rect 12409 -15048 12485 -15032
rect 12409 -15066 12425 -15048
rect 12291 -15082 12329 -15066
rect 12209 -15120 12329 -15082
rect 12387 -15082 12425 -15066
rect 12469 -15066 12485 -15048
rect 12587 -15048 12663 -15032
rect 12587 -15066 12603 -15048
rect 12469 -15082 12507 -15066
rect 12387 -15120 12507 -15082
rect 12565 -15082 12603 -15066
rect 12647 -15066 12663 -15048
rect 12647 -15082 12685 -15066
rect 12565 -15120 12685 -15082
rect -5982 -15400 -5862 -15362
rect -5982 -15416 -5944 -15400
rect -5960 -15434 -5944 -15416
rect -5900 -15416 -5862 -15400
rect -5804 -15400 -5684 -15362
rect -5804 -15416 -5766 -15400
rect -5900 -15434 -5884 -15416
rect -5960 -15450 -5884 -15434
rect -5782 -15434 -5766 -15416
rect -5722 -15416 -5684 -15400
rect -5626 -15400 -5506 -15362
rect -5626 -15416 -5588 -15400
rect -5722 -15434 -5706 -15416
rect -5782 -15450 -5706 -15434
rect -5604 -15434 -5588 -15416
rect -5544 -15416 -5506 -15400
rect -5448 -15400 -5328 -15362
rect -5448 -15416 -5410 -15400
rect -5544 -15434 -5528 -15416
rect -5604 -15450 -5528 -15434
rect -5426 -15434 -5410 -15416
rect -5366 -15416 -5328 -15400
rect -5270 -15400 -5150 -15362
rect -5270 -15416 -5232 -15400
rect -5366 -15434 -5350 -15416
rect -5426 -15450 -5350 -15434
rect -5248 -15434 -5232 -15416
rect -5188 -15416 -5150 -15400
rect -5092 -15400 -4972 -15362
rect -5092 -15416 -5054 -15400
rect -5188 -15434 -5172 -15416
rect -5248 -15450 -5172 -15434
rect -5070 -15434 -5054 -15416
rect -5010 -15416 -4972 -15400
rect -4914 -15400 -4794 -15362
rect -4914 -15416 -4876 -15400
rect -5010 -15434 -4994 -15416
rect -5070 -15450 -4994 -15434
rect -4892 -15434 -4876 -15416
rect -4832 -15416 -4794 -15400
rect -4736 -15400 -4616 -15362
rect -4736 -15416 -4698 -15400
rect -4832 -15434 -4816 -15416
rect -4892 -15450 -4816 -15434
rect -4714 -15434 -4698 -15416
rect -4654 -15416 -4616 -15400
rect -4558 -15400 -4438 -15362
rect -4558 -15416 -4520 -15400
rect -4654 -15434 -4638 -15416
rect -4714 -15450 -4638 -15434
rect -4536 -15434 -4520 -15416
rect -4476 -15416 -4438 -15400
rect -4380 -15400 -4260 -15362
rect -4380 -15416 -4342 -15400
rect -4476 -15434 -4460 -15416
rect -4536 -15450 -4460 -15434
rect -4358 -15434 -4342 -15416
rect -4298 -15416 -4260 -15400
rect -4202 -15400 -4082 -15362
rect -4202 -15416 -4164 -15400
rect -4298 -15434 -4282 -15416
rect -4358 -15450 -4282 -15434
rect -4180 -15434 -4164 -15416
rect -4120 -15416 -4082 -15400
rect -4120 -15434 -4104 -15416
rect -4180 -15450 -4104 -15434
rect -2127 -15438 -2007 -15400
rect -2127 -15454 -2089 -15438
rect -2105 -15472 -2089 -15454
rect -2045 -15454 -2007 -15438
rect -1949 -15438 -1829 -15400
rect -1949 -15454 -1911 -15438
rect -2045 -15472 -2029 -15454
rect -2105 -15488 -2029 -15472
rect -1927 -15472 -1911 -15454
rect -1867 -15454 -1829 -15438
rect -1771 -15438 -1651 -15400
rect -1771 -15454 -1733 -15438
rect -1867 -15472 -1851 -15454
rect -1927 -15488 -1851 -15472
rect -1749 -15472 -1733 -15454
rect -1689 -15454 -1651 -15438
rect -1593 -15438 -1473 -15400
rect -1593 -15454 -1555 -15438
rect -1689 -15472 -1673 -15454
rect -1749 -15488 -1673 -15472
rect -1571 -15472 -1555 -15454
rect -1511 -15454 -1473 -15438
rect -1415 -15438 -1295 -15400
rect -1415 -15454 -1377 -15438
rect -1511 -15472 -1495 -15454
rect -1571 -15488 -1495 -15472
rect -1393 -15472 -1377 -15454
rect -1333 -15454 -1295 -15438
rect -1237 -15438 -1117 -15400
rect -1237 -15454 -1199 -15438
rect -1333 -15472 -1317 -15454
rect -1393 -15488 -1317 -15472
rect -1215 -15472 -1199 -15454
rect -1155 -15454 -1117 -15438
rect -1059 -15438 -939 -15400
rect -1059 -15454 -1021 -15438
rect -1155 -15472 -1139 -15454
rect -1215 -15488 -1139 -15472
rect -1037 -15472 -1021 -15454
rect -977 -15454 -939 -15438
rect -881 -15438 -761 -15400
rect -881 -15454 -843 -15438
rect -977 -15472 -961 -15454
rect -1037 -15488 -961 -15472
rect -859 -15472 -843 -15454
rect -799 -15454 -761 -15438
rect -703 -15438 -583 -15400
rect -703 -15454 -665 -15438
rect -799 -15472 -783 -15454
rect -859 -15488 -783 -15472
rect -681 -15472 -665 -15454
rect -621 -15454 -583 -15438
rect -525 -15438 -405 -15400
rect -525 -15454 -487 -15438
rect -621 -15472 -605 -15454
rect -681 -15488 -605 -15472
rect -503 -15472 -487 -15454
rect -443 -15454 -405 -15438
rect -347 -15438 -227 -15400
rect -347 -15454 -309 -15438
rect -443 -15472 -427 -15454
rect -503 -15488 -427 -15472
rect -325 -15472 -309 -15454
rect -265 -15454 -227 -15438
rect -169 -15438 -49 -15400
rect -169 -15454 -131 -15438
rect -265 -15472 -249 -15454
rect -325 -15488 -249 -15472
rect -147 -15472 -131 -15454
rect -87 -15454 -49 -15438
rect 9 -15438 129 -15400
rect 9 -15454 47 -15438
rect -87 -15472 -71 -15454
rect -147 -15488 -71 -15472
rect 31 -15472 47 -15454
rect 91 -15454 129 -15438
rect 187 -15438 307 -15400
rect 187 -15454 225 -15438
rect 91 -15472 107 -15454
rect 31 -15488 107 -15472
rect 209 -15472 225 -15454
rect 269 -15454 307 -15438
rect 365 -15438 485 -15400
rect 365 -15454 403 -15438
rect 269 -15472 285 -15454
rect 209 -15488 285 -15472
rect 387 -15472 403 -15454
rect 447 -15454 485 -15438
rect 543 -15438 663 -15400
rect 543 -15454 581 -15438
rect 447 -15472 463 -15454
rect 387 -15488 463 -15472
rect 565 -15472 581 -15454
rect 625 -15454 663 -15438
rect 721 -15438 841 -15400
rect 721 -15454 759 -15438
rect 625 -15472 641 -15454
rect 565 -15488 641 -15472
rect 743 -15472 759 -15454
rect 803 -15454 841 -15438
rect 899 -15438 1019 -15400
rect 899 -15454 937 -15438
rect 803 -15472 819 -15454
rect 743 -15488 819 -15472
rect 921 -15472 937 -15454
rect 981 -15454 1019 -15438
rect 1077 -15438 1197 -15400
rect 1077 -15454 1115 -15438
rect 981 -15472 997 -15454
rect 921 -15488 997 -15472
rect 1099 -15472 1115 -15454
rect 1159 -15454 1197 -15438
rect 1255 -15438 1375 -15400
rect 1255 -15454 1293 -15438
rect 1159 -15472 1175 -15454
rect 1099 -15488 1175 -15472
rect 1277 -15472 1293 -15454
rect 1337 -15454 1375 -15438
rect 1433 -15438 1553 -15400
rect 1433 -15454 1471 -15438
rect 1337 -15472 1353 -15454
rect 1277 -15488 1353 -15472
rect 1455 -15472 1471 -15454
rect 1515 -15454 1553 -15438
rect 1611 -15438 1731 -15400
rect 1611 -15454 1649 -15438
rect 1515 -15472 1531 -15454
rect 1455 -15488 1531 -15472
rect 1633 -15472 1649 -15454
rect 1693 -15454 1731 -15438
rect 1789 -15438 1909 -15400
rect 1789 -15454 1827 -15438
rect 1693 -15472 1709 -15454
rect 1633 -15488 1709 -15472
rect 1811 -15472 1827 -15454
rect 1871 -15454 1909 -15438
rect 1967 -15438 2087 -15400
rect 1967 -15454 2005 -15438
rect 1871 -15472 1887 -15454
rect 1811 -15488 1887 -15472
rect 1989 -15472 2005 -15454
rect 2049 -15454 2087 -15438
rect 2145 -15438 2265 -15400
rect 2145 -15454 2183 -15438
rect 2049 -15472 2065 -15454
rect 1989 -15488 2065 -15472
rect 2167 -15472 2183 -15454
rect 2227 -15454 2265 -15438
rect 2323 -15438 2443 -15400
rect 2323 -15454 2361 -15438
rect 2227 -15472 2243 -15454
rect 2167 -15488 2243 -15472
rect 2345 -15472 2361 -15454
rect 2405 -15454 2443 -15438
rect 2501 -15438 2621 -15400
rect 2501 -15454 2539 -15438
rect 2405 -15472 2421 -15454
rect 2345 -15488 2421 -15472
rect 2523 -15472 2539 -15454
rect 2583 -15454 2621 -15438
rect 2679 -15438 2799 -15400
rect 2679 -15454 2717 -15438
rect 2583 -15472 2599 -15454
rect 2523 -15488 2599 -15472
rect 2701 -15472 2717 -15454
rect 2761 -15454 2799 -15438
rect 2857 -15438 2977 -15400
rect 2857 -15454 2895 -15438
rect 2761 -15472 2777 -15454
rect 2701 -15488 2777 -15472
rect 2879 -15472 2895 -15454
rect 2939 -15454 2977 -15438
rect 3035 -15438 3155 -15400
rect 3035 -15454 3073 -15438
rect 2939 -15472 2955 -15454
rect 2879 -15488 2955 -15472
rect 3057 -15472 3073 -15454
rect 3117 -15454 3155 -15438
rect 3213 -15438 3333 -15400
rect 3213 -15454 3251 -15438
rect 3117 -15472 3133 -15454
rect 3057 -15488 3133 -15472
rect 3235 -15472 3251 -15454
rect 3295 -15454 3333 -15438
rect 3391 -15438 3511 -15400
rect 3391 -15454 3429 -15438
rect 3295 -15472 3311 -15454
rect 3235 -15488 3311 -15472
rect 3413 -15472 3429 -15454
rect 3473 -15454 3511 -15438
rect 3569 -15438 3689 -15400
rect 3569 -15454 3607 -15438
rect 3473 -15472 3489 -15454
rect 3413 -15488 3489 -15472
rect 3591 -15472 3607 -15454
rect 3651 -15454 3689 -15438
rect 3747 -15438 3867 -15400
rect 3747 -15454 3785 -15438
rect 3651 -15472 3667 -15454
rect 3591 -15488 3667 -15472
rect 3769 -15472 3785 -15454
rect 3829 -15454 3867 -15438
rect 3925 -15438 4045 -15400
rect 3925 -15454 3963 -15438
rect 3829 -15472 3845 -15454
rect 3769 -15488 3845 -15472
rect 3947 -15472 3963 -15454
rect 4007 -15454 4045 -15438
rect 5623 -15438 5743 -15400
rect 5623 -15454 5661 -15438
rect 4007 -15472 4023 -15454
rect 3947 -15488 4023 -15472
rect 5645 -15472 5661 -15454
rect 5705 -15454 5743 -15438
rect 5801 -15438 5921 -15400
rect 5801 -15454 5839 -15438
rect 5705 -15472 5721 -15454
rect 5645 -15488 5721 -15472
rect 5823 -15472 5839 -15454
rect 5883 -15454 5921 -15438
rect 5979 -15438 6099 -15400
rect 5979 -15454 6017 -15438
rect 5883 -15472 5899 -15454
rect 5823 -15488 5899 -15472
rect 6001 -15472 6017 -15454
rect 6061 -15454 6099 -15438
rect 6157 -15438 6277 -15400
rect 6157 -15454 6195 -15438
rect 6061 -15472 6077 -15454
rect 6001 -15488 6077 -15472
rect 6179 -15472 6195 -15454
rect 6239 -15454 6277 -15438
rect 6335 -15438 6455 -15400
rect 6335 -15454 6373 -15438
rect 6239 -15472 6255 -15454
rect 6179 -15488 6255 -15472
rect 6357 -15472 6373 -15454
rect 6417 -15454 6455 -15438
rect 6513 -15438 6633 -15400
rect 6513 -15454 6551 -15438
rect 6417 -15472 6433 -15454
rect 6357 -15488 6433 -15472
rect 6535 -15472 6551 -15454
rect 6595 -15454 6633 -15438
rect 6691 -15438 6811 -15400
rect 6691 -15454 6729 -15438
rect 6595 -15472 6611 -15454
rect 6535 -15488 6611 -15472
rect 6713 -15472 6729 -15454
rect 6773 -15454 6811 -15438
rect 6869 -15438 6989 -15400
rect 6869 -15454 6907 -15438
rect 6773 -15472 6789 -15454
rect 6713 -15488 6789 -15472
rect 6891 -15472 6907 -15454
rect 6951 -15454 6989 -15438
rect 7047 -15438 7167 -15400
rect 7047 -15454 7085 -15438
rect 6951 -15472 6967 -15454
rect 6891 -15488 6967 -15472
rect 7069 -15472 7085 -15454
rect 7129 -15454 7167 -15438
rect 7225 -15438 7345 -15400
rect 7225 -15454 7263 -15438
rect 7129 -15472 7145 -15454
rect 7069 -15488 7145 -15472
rect 7247 -15472 7263 -15454
rect 7307 -15454 7345 -15438
rect 7403 -15438 7523 -15400
rect 7403 -15454 7441 -15438
rect 7307 -15472 7323 -15454
rect 7247 -15488 7323 -15472
rect 7425 -15472 7441 -15454
rect 7485 -15454 7523 -15438
rect 7581 -15438 7701 -15400
rect 7581 -15454 7619 -15438
rect 7485 -15472 7501 -15454
rect 7425 -15488 7501 -15472
rect 7603 -15472 7619 -15454
rect 7663 -15454 7701 -15438
rect 7759 -15438 7879 -15400
rect 7759 -15454 7797 -15438
rect 7663 -15472 7679 -15454
rect 7603 -15488 7679 -15472
rect 7781 -15472 7797 -15454
rect 7841 -15454 7879 -15438
rect 7937 -15438 8057 -15400
rect 7937 -15454 7975 -15438
rect 7841 -15472 7857 -15454
rect 7781 -15488 7857 -15472
rect 7959 -15472 7975 -15454
rect 8019 -15454 8057 -15438
rect 8115 -15438 8235 -15400
rect 8115 -15454 8153 -15438
rect 8019 -15472 8035 -15454
rect 7959 -15488 8035 -15472
rect 8137 -15472 8153 -15454
rect 8197 -15454 8235 -15438
rect 8293 -15438 8413 -15400
rect 8293 -15454 8331 -15438
rect 8197 -15472 8213 -15454
rect 8137 -15488 8213 -15472
rect 8315 -15472 8331 -15454
rect 8375 -15454 8413 -15438
rect 8471 -15438 8591 -15400
rect 8471 -15454 8509 -15438
rect 8375 -15472 8391 -15454
rect 8315 -15488 8391 -15472
rect 8493 -15472 8509 -15454
rect 8553 -15454 8591 -15438
rect 8649 -15438 8769 -15400
rect 8649 -15454 8687 -15438
rect 8553 -15472 8569 -15454
rect 8493 -15488 8569 -15472
rect 8671 -15472 8687 -15454
rect 8731 -15454 8769 -15438
rect 8827 -15438 8947 -15400
rect 8827 -15454 8865 -15438
rect 8731 -15472 8747 -15454
rect 8671 -15488 8747 -15472
rect 8849 -15472 8865 -15454
rect 8909 -15454 8947 -15438
rect 9005 -15438 9125 -15400
rect 9005 -15454 9043 -15438
rect 8909 -15472 8925 -15454
rect 8849 -15488 8925 -15472
rect 9027 -15472 9043 -15454
rect 9087 -15454 9125 -15438
rect 9183 -15438 9303 -15400
rect 9183 -15454 9221 -15438
rect 9087 -15472 9103 -15454
rect 9027 -15488 9103 -15472
rect 9205 -15472 9221 -15454
rect 9265 -15454 9303 -15438
rect 9361 -15438 9481 -15400
rect 9361 -15454 9399 -15438
rect 9265 -15472 9281 -15454
rect 9205 -15488 9281 -15472
rect 9383 -15472 9399 -15454
rect 9443 -15454 9481 -15438
rect 9539 -15438 9659 -15400
rect 9539 -15454 9577 -15438
rect 9443 -15472 9459 -15454
rect 9383 -15488 9459 -15472
rect 9561 -15472 9577 -15454
rect 9621 -15454 9659 -15438
rect 9717 -15438 9837 -15400
rect 9717 -15454 9755 -15438
rect 9621 -15472 9637 -15454
rect 9561 -15488 9637 -15472
rect 9739 -15472 9755 -15454
rect 9799 -15454 9837 -15438
rect 9895 -15438 10015 -15400
rect 9895 -15454 9933 -15438
rect 9799 -15472 9815 -15454
rect 9739 -15488 9815 -15472
rect 9917 -15472 9933 -15454
rect 9977 -15454 10015 -15438
rect 10073 -15438 10193 -15400
rect 10073 -15454 10111 -15438
rect 9977 -15472 9993 -15454
rect 9917 -15488 9993 -15472
rect 10095 -15472 10111 -15454
rect 10155 -15454 10193 -15438
rect 10251 -15438 10371 -15400
rect 10251 -15454 10289 -15438
rect 10155 -15472 10171 -15454
rect 10095 -15488 10171 -15472
rect 10273 -15472 10289 -15454
rect 10333 -15454 10371 -15438
rect 10429 -15438 10549 -15400
rect 10429 -15454 10467 -15438
rect 10333 -15472 10349 -15454
rect 10273 -15488 10349 -15472
rect 10451 -15472 10467 -15454
rect 10511 -15454 10549 -15438
rect 10607 -15438 10727 -15400
rect 10607 -15454 10645 -15438
rect 10511 -15472 10527 -15454
rect 10451 -15488 10527 -15472
rect 10629 -15472 10645 -15454
rect 10689 -15454 10727 -15438
rect 10785 -15438 10905 -15400
rect 10785 -15454 10823 -15438
rect 10689 -15472 10705 -15454
rect 10629 -15488 10705 -15472
rect 10807 -15472 10823 -15454
rect 10867 -15454 10905 -15438
rect 10963 -15438 11083 -15400
rect 10963 -15454 11001 -15438
rect 10867 -15472 10883 -15454
rect 10807 -15488 10883 -15472
rect 10985 -15472 11001 -15454
rect 11045 -15454 11083 -15438
rect 11141 -15438 11261 -15400
rect 11141 -15454 11179 -15438
rect 11045 -15472 11061 -15454
rect 10985 -15488 11061 -15472
rect 11163 -15472 11179 -15454
rect 11223 -15454 11261 -15438
rect 11319 -15438 11439 -15400
rect 11319 -15454 11357 -15438
rect 11223 -15472 11239 -15454
rect 11163 -15488 11239 -15472
rect 11341 -15472 11357 -15454
rect 11401 -15454 11439 -15438
rect 11497 -15438 11617 -15400
rect 11497 -15454 11535 -15438
rect 11401 -15472 11417 -15454
rect 11341 -15488 11417 -15472
rect 11519 -15472 11535 -15454
rect 11579 -15454 11617 -15438
rect 11675 -15438 11795 -15400
rect 11675 -15454 11713 -15438
rect 11579 -15472 11595 -15454
rect 11519 -15488 11595 -15472
rect 11697 -15472 11713 -15454
rect 11757 -15454 11795 -15438
rect 11853 -15438 11973 -15400
rect 11853 -15454 11891 -15438
rect 11757 -15472 11773 -15454
rect 11697 -15488 11773 -15472
rect 11875 -15472 11891 -15454
rect 11935 -15454 11973 -15438
rect 12031 -15438 12151 -15400
rect 12031 -15454 12069 -15438
rect 11935 -15472 11951 -15454
rect 11875 -15488 11951 -15472
rect 12053 -15472 12069 -15454
rect 12113 -15454 12151 -15438
rect 12209 -15438 12329 -15400
rect 12209 -15454 12247 -15438
rect 12113 -15472 12129 -15454
rect 12053 -15488 12129 -15472
rect 12231 -15472 12247 -15454
rect 12291 -15454 12329 -15438
rect 12387 -15438 12507 -15400
rect 12387 -15454 12425 -15438
rect 12291 -15472 12307 -15454
rect 12231 -15488 12307 -15472
rect 12409 -15472 12425 -15454
rect 12469 -15454 12507 -15438
rect 12565 -15438 12685 -15400
rect 12565 -15454 12603 -15438
rect 12469 -15472 12485 -15454
rect 12409 -15488 12485 -15472
rect 12587 -15472 12603 -15454
rect 12647 -15454 12685 -15438
rect 12647 -15472 12663 -15454
rect 12587 -15488 12663 -15472
rect -5960 -15710 -5884 -15694
rect -5960 -15728 -5944 -15710
rect -5982 -15744 -5944 -15728
rect -5900 -15728 -5884 -15710
rect -5782 -15710 -5706 -15694
rect -5782 -15728 -5766 -15710
rect -5900 -15744 -5862 -15728
rect -5982 -15782 -5862 -15744
rect -5804 -15744 -5766 -15728
rect -5722 -15728 -5706 -15710
rect -5604 -15710 -5528 -15694
rect -5604 -15728 -5588 -15710
rect -5722 -15744 -5684 -15728
rect -5804 -15782 -5684 -15744
rect -5626 -15744 -5588 -15728
rect -5544 -15728 -5528 -15710
rect -5426 -15710 -5350 -15694
rect -5426 -15728 -5410 -15710
rect -5544 -15744 -5506 -15728
rect -5626 -15782 -5506 -15744
rect -5448 -15744 -5410 -15728
rect -5366 -15728 -5350 -15710
rect -5248 -15710 -5172 -15694
rect -5248 -15728 -5232 -15710
rect -5366 -15744 -5328 -15728
rect -5448 -15782 -5328 -15744
rect -5270 -15744 -5232 -15728
rect -5188 -15728 -5172 -15710
rect -5070 -15710 -4994 -15694
rect -5070 -15728 -5054 -15710
rect -5188 -15744 -5150 -15728
rect -5270 -15782 -5150 -15744
rect -5092 -15744 -5054 -15728
rect -5010 -15728 -4994 -15710
rect -4892 -15710 -4816 -15694
rect -4892 -15728 -4876 -15710
rect -5010 -15744 -4972 -15728
rect -5092 -15782 -4972 -15744
rect -4914 -15744 -4876 -15728
rect -4832 -15728 -4816 -15710
rect -4714 -15710 -4638 -15694
rect -4714 -15728 -4698 -15710
rect -4832 -15744 -4794 -15728
rect -4914 -15782 -4794 -15744
rect -4736 -15744 -4698 -15728
rect -4654 -15728 -4638 -15710
rect -4536 -15710 -4460 -15694
rect -4536 -15728 -4520 -15710
rect -4654 -15744 -4616 -15728
rect -4736 -15782 -4616 -15744
rect -4558 -15744 -4520 -15728
rect -4476 -15728 -4460 -15710
rect -4358 -15710 -4282 -15694
rect -4358 -15728 -4342 -15710
rect -4476 -15744 -4438 -15728
rect -4558 -15782 -4438 -15744
rect -4380 -15744 -4342 -15728
rect -4298 -15728 -4282 -15710
rect -4180 -15710 -4104 -15694
rect -4180 -15728 -4164 -15710
rect -4298 -15744 -4260 -15728
rect -4380 -15782 -4260 -15744
rect -4202 -15744 -4164 -15728
rect -4120 -15728 -4104 -15710
rect -4120 -15744 -4082 -15728
rect -4202 -15782 -4082 -15744
rect -2105 -16048 -2029 -16032
rect -5982 -16100 -5862 -16062
rect -5982 -16116 -5944 -16100
rect -5960 -16134 -5944 -16116
rect -5900 -16116 -5862 -16100
rect -5804 -16100 -5684 -16062
rect -5804 -16116 -5766 -16100
rect -5900 -16134 -5884 -16116
rect -5960 -16150 -5884 -16134
rect -5782 -16134 -5766 -16116
rect -5722 -16116 -5684 -16100
rect -5626 -16100 -5506 -16062
rect -5626 -16116 -5588 -16100
rect -5722 -16134 -5706 -16116
rect -5782 -16150 -5706 -16134
rect -5604 -16134 -5588 -16116
rect -5544 -16116 -5506 -16100
rect -5448 -16100 -5328 -16062
rect -5448 -16116 -5410 -16100
rect -5544 -16134 -5528 -16116
rect -5604 -16150 -5528 -16134
rect -5426 -16134 -5410 -16116
rect -5366 -16116 -5328 -16100
rect -5270 -16100 -5150 -16062
rect -5270 -16116 -5232 -16100
rect -5366 -16134 -5350 -16116
rect -5426 -16150 -5350 -16134
rect -5248 -16134 -5232 -16116
rect -5188 -16116 -5150 -16100
rect -5092 -16100 -4972 -16062
rect -5092 -16116 -5054 -16100
rect -5188 -16134 -5172 -16116
rect -5248 -16150 -5172 -16134
rect -5070 -16134 -5054 -16116
rect -5010 -16116 -4972 -16100
rect -4914 -16100 -4794 -16062
rect -4914 -16116 -4876 -16100
rect -5010 -16134 -4994 -16116
rect -5070 -16150 -4994 -16134
rect -4892 -16134 -4876 -16116
rect -4832 -16116 -4794 -16100
rect -4736 -16100 -4616 -16062
rect -4736 -16116 -4698 -16100
rect -4832 -16134 -4816 -16116
rect -4892 -16150 -4816 -16134
rect -4714 -16134 -4698 -16116
rect -4654 -16116 -4616 -16100
rect -4558 -16100 -4438 -16062
rect -4558 -16116 -4520 -16100
rect -4654 -16134 -4638 -16116
rect -4714 -16150 -4638 -16134
rect -4536 -16134 -4520 -16116
rect -4476 -16116 -4438 -16100
rect -4380 -16100 -4260 -16062
rect -4380 -16116 -4342 -16100
rect -4476 -16134 -4460 -16116
rect -4536 -16150 -4460 -16134
rect -4358 -16134 -4342 -16116
rect -4298 -16116 -4260 -16100
rect -4202 -16100 -4082 -16062
rect -2105 -16066 -2089 -16048
rect -4202 -16116 -4164 -16100
rect -4298 -16134 -4282 -16116
rect -4358 -16150 -4282 -16134
rect -4180 -16134 -4164 -16116
rect -4120 -16116 -4082 -16100
rect -2127 -16082 -2089 -16066
rect -2045 -16066 -2029 -16048
rect -1927 -16048 -1851 -16032
rect -1927 -16066 -1911 -16048
rect -2045 -16082 -2007 -16066
rect -4120 -16134 -4104 -16116
rect -2127 -16120 -2007 -16082
rect -1949 -16082 -1911 -16066
rect -1867 -16066 -1851 -16048
rect -1749 -16048 -1673 -16032
rect -1749 -16066 -1733 -16048
rect -1867 -16082 -1829 -16066
rect -1949 -16120 -1829 -16082
rect -1771 -16082 -1733 -16066
rect -1689 -16066 -1673 -16048
rect -1571 -16048 -1495 -16032
rect -1571 -16066 -1555 -16048
rect -1689 -16082 -1651 -16066
rect -1771 -16120 -1651 -16082
rect -1593 -16082 -1555 -16066
rect -1511 -16066 -1495 -16048
rect -1393 -16048 -1317 -16032
rect -1393 -16066 -1377 -16048
rect -1511 -16082 -1473 -16066
rect -1593 -16120 -1473 -16082
rect -1415 -16082 -1377 -16066
rect -1333 -16066 -1317 -16048
rect -1215 -16048 -1139 -16032
rect -1215 -16066 -1199 -16048
rect -1333 -16082 -1295 -16066
rect -1415 -16120 -1295 -16082
rect -1237 -16082 -1199 -16066
rect -1155 -16066 -1139 -16048
rect -1037 -16048 -961 -16032
rect -1037 -16066 -1021 -16048
rect -1155 -16082 -1117 -16066
rect -1237 -16120 -1117 -16082
rect -1059 -16082 -1021 -16066
rect -977 -16066 -961 -16048
rect -859 -16048 -783 -16032
rect -859 -16066 -843 -16048
rect -977 -16082 -939 -16066
rect -1059 -16120 -939 -16082
rect -881 -16082 -843 -16066
rect -799 -16066 -783 -16048
rect -681 -16048 -605 -16032
rect -681 -16066 -665 -16048
rect -799 -16082 -761 -16066
rect -881 -16120 -761 -16082
rect -703 -16082 -665 -16066
rect -621 -16066 -605 -16048
rect -503 -16048 -427 -16032
rect -503 -16066 -487 -16048
rect -621 -16082 -583 -16066
rect -703 -16120 -583 -16082
rect -525 -16082 -487 -16066
rect -443 -16066 -427 -16048
rect -325 -16048 -249 -16032
rect -325 -16066 -309 -16048
rect -443 -16082 -405 -16066
rect -525 -16120 -405 -16082
rect -347 -16082 -309 -16066
rect -265 -16066 -249 -16048
rect -147 -16048 -71 -16032
rect -147 -16066 -131 -16048
rect -265 -16082 -227 -16066
rect -347 -16120 -227 -16082
rect -169 -16082 -131 -16066
rect -87 -16066 -71 -16048
rect 31 -16048 107 -16032
rect 31 -16066 47 -16048
rect -87 -16082 -49 -16066
rect -169 -16120 -49 -16082
rect 9 -16082 47 -16066
rect 91 -16066 107 -16048
rect 209 -16048 285 -16032
rect 209 -16066 225 -16048
rect 91 -16082 129 -16066
rect 9 -16120 129 -16082
rect 187 -16082 225 -16066
rect 269 -16066 285 -16048
rect 387 -16048 463 -16032
rect 387 -16066 403 -16048
rect 269 -16082 307 -16066
rect 187 -16120 307 -16082
rect 365 -16082 403 -16066
rect 447 -16066 463 -16048
rect 565 -16048 641 -16032
rect 565 -16066 581 -16048
rect 447 -16082 485 -16066
rect 365 -16120 485 -16082
rect 543 -16082 581 -16066
rect 625 -16066 641 -16048
rect 743 -16048 819 -16032
rect 743 -16066 759 -16048
rect 625 -16082 663 -16066
rect 543 -16120 663 -16082
rect 721 -16082 759 -16066
rect 803 -16066 819 -16048
rect 921 -16048 997 -16032
rect 921 -16066 937 -16048
rect 803 -16082 841 -16066
rect 721 -16120 841 -16082
rect 899 -16082 937 -16066
rect 981 -16066 997 -16048
rect 1099 -16048 1175 -16032
rect 1099 -16066 1115 -16048
rect 981 -16082 1019 -16066
rect 899 -16120 1019 -16082
rect 1077 -16082 1115 -16066
rect 1159 -16066 1175 -16048
rect 1277 -16048 1353 -16032
rect 1277 -16066 1293 -16048
rect 1159 -16082 1197 -16066
rect 1077 -16120 1197 -16082
rect 1255 -16082 1293 -16066
rect 1337 -16066 1353 -16048
rect 1455 -16048 1531 -16032
rect 1455 -16066 1471 -16048
rect 1337 -16082 1375 -16066
rect 1255 -16120 1375 -16082
rect 1433 -16082 1471 -16066
rect 1515 -16066 1531 -16048
rect 1633 -16048 1709 -16032
rect 1633 -16066 1649 -16048
rect 1515 -16082 1553 -16066
rect 1433 -16120 1553 -16082
rect 1611 -16082 1649 -16066
rect 1693 -16066 1709 -16048
rect 1811 -16048 1887 -16032
rect 1811 -16066 1827 -16048
rect 1693 -16082 1731 -16066
rect 1611 -16120 1731 -16082
rect 1789 -16082 1827 -16066
rect 1871 -16066 1887 -16048
rect 1989 -16048 2065 -16032
rect 1989 -16066 2005 -16048
rect 1871 -16082 1909 -16066
rect 1789 -16120 1909 -16082
rect 1967 -16082 2005 -16066
rect 2049 -16066 2065 -16048
rect 2167 -16048 2243 -16032
rect 2167 -16066 2183 -16048
rect 2049 -16082 2087 -16066
rect 1967 -16120 2087 -16082
rect 2145 -16082 2183 -16066
rect 2227 -16066 2243 -16048
rect 2345 -16048 2421 -16032
rect 2345 -16066 2361 -16048
rect 2227 -16082 2265 -16066
rect 2145 -16120 2265 -16082
rect 2323 -16082 2361 -16066
rect 2405 -16066 2421 -16048
rect 2523 -16048 2599 -16032
rect 2523 -16066 2539 -16048
rect 2405 -16082 2443 -16066
rect 2323 -16120 2443 -16082
rect 2501 -16082 2539 -16066
rect 2583 -16066 2599 -16048
rect 2701 -16048 2777 -16032
rect 2701 -16066 2717 -16048
rect 2583 -16082 2621 -16066
rect 2501 -16120 2621 -16082
rect 2679 -16082 2717 -16066
rect 2761 -16066 2777 -16048
rect 2879 -16048 2955 -16032
rect 2879 -16066 2895 -16048
rect 2761 -16082 2799 -16066
rect 2679 -16120 2799 -16082
rect 2857 -16082 2895 -16066
rect 2939 -16066 2955 -16048
rect 3057 -16048 3133 -16032
rect 3057 -16066 3073 -16048
rect 2939 -16082 2977 -16066
rect 2857 -16120 2977 -16082
rect 3035 -16082 3073 -16066
rect 3117 -16066 3133 -16048
rect 3235 -16048 3311 -16032
rect 3235 -16066 3251 -16048
rect 3117 -16082 3155 -16066
rect 3035 -16120 3155 -16082
rect 3213 -16082 3251 -16066
rect 3295 -16066 3311 -16048
rect 3413 -16048 3489 -16032
rect 3413 -16066 3429 -16048
rect 3295 -16082 3333 -16066
rect 3213 -16120 3333 -16082
rect 3391 -16082 3429 -16066
rect 3473 -16066 3489 -16048
rect 3591 -16048 3667 -16032
rect 3591 -16066 3607 -16048
rect 3473 -16082 3511 -16066
rect 3391 -16120 3511 -16082
rect 3569 -16082 3607 -16066
rect 3651 -16066 3667 -16048
rect 3769 -16048 3845 -16032
rect 3769 -16066 3785 -16048
rect 3651 -16082 3689 -16066
rect 3569 -16120 3689 -16082
rect 3747 -16082 3785 -16066
rect 3829 -16066 3845 -16048
rect 3947 -16048 4023 -16032
rect 3947 -16066 3963 -16048
rect 3829 -16082 3867 -16066
rect 3747 -16120 3867 -16082
rect 3925 -16082 3963 -16066
rect 4007 -16066 4023 -16048
rect 5645 -16048 5721 -16032
rect 5645 -16066 5661 -16048
rect 4007 -16082 4045 -16066
rect 3925 -16120 4045 -16082
rect 5623 -16082 5661 -16066
rect 5705 -16066 5721 -16048
rect 5823 -16048 5899 -16032
rect 5823 -16066 5839 -16048
rect 5705 -16082 5743 -16066
rect 5623 -16120 5743 -16082
rect 5801 -16082 5839 -16066
rect 5883 -16066 5899 -16048
rect 6001 -16048 6077 -16032
rect 6001 -16066 6017 -16048
rect 5883 -16082 5921 -16066
rect 5801 -16120 5921 -16082
rect 5979 -16082 6017 -16066
rect 6061 -16066 6077 -16048
rect 6179 -16048 6255 -16032
rect 6179 -16066 6195 -16048
rect 6061 -16082 6099 -16066
rect 5979 -16120 6099 -16082
rect 6157 -16082 6195 -16066
rect 6239 -16066 6255 -16048
rect 6357 -16048 6433 -16032
rect 6357 -16066 6373 -16048
rect 6239 -16082 6277 -16066
rect 6157 -16120 6277 -16082
rect 6335 -16082 6373 -16066
rect 6417 -16066 6433 -16048
rect 6535 -16048 6611 -16032
rect 6535 -16066 6551 -16048
rect 6417 -16082 6455 -16066
rect 6335 -16120 6455 -16082
rect 6513 -16082 6551 -16066
rect 6595 -16066 6611 -16048
rect 6713 -16048 6789 -16032
rect 6713 -16066 6729 -16048
rect 6595 -16082 6633 -16066
rect 6513 -16120 6633 -16082
rect 6691 -16082 6729 -16066
rect 6773 -16066 6789 -16048
rect 6891 -16048 6967 -16032
rect 6891 -16066 6907 -16048
rect 6773 -16082 6811 -16066
rect 6691 -16120 6811 -16082
rect 6869 -16082 6907 -16066
rect 6951 -16066 6967 -16048
rect 7069 -16048 7145 -16032
rect 7069 -16066 7085 -16048
rect 6951 -16082 6989 -16066
rect 6869 -16120 6989 -16082
rect 7047 -16082 7085 -16066
rect 7129 -16066 7145 -16048
rect 7247 -16048 7323 -16032
rect 7247 -16066 7263 -16048
rect 7129 -16082 7167 -16066
rect 7047 -16120 7167 -16082
rect 7225 -16082 7263 -16066
rect 7307 -16066 7323 -16048
rect 7425 -16048 7501 -16032
rect 7425 -16066 7441 -16048
rect 7307 -16082 7345 -16066
rect 7225 -16120 7345 -16082
rect 7403 -16082 7441 -16066
rect 7485 -16066 7501 -16048
rect 7603 -16048 7679 -16032
rect 7603 -16066 7619 -16048
rect 7485 -16082 7523 -16066
rect 7403 -16120 7523 -16082
rect 7581 -16082 7619 -16066
rect 7663 -16066 7679 -16048
rect 7781 -16048 7857 -16032
rect 7781 -16066 7797 -16048
rect 7663 -16082 7701 -16066
rect 7581 -16120 7701 -16082
rect 7759 -16082 7797 -16066
rect 7841 -16066 7857 -16048
rect 7959 -16048 8035 -16032
rect 7959 -16066 7975 -16048
rect 7841 -16082 7879 -16066
rect 7759 -16120 7879 -16082
rect 7937 -16082 7975 -16066
rect 8019 -16066 8035 -16048
rect 8137 -16048 8213 -16032
rect 8137 -16066 8153 -16048
rect 8019 -16082 8057 -16066
rect 7937 -16120 8057 -16082
rect 8115 -16082 8153 -16066
rect 8197 -16066 8213 -16048
rect 8315 -16048 8391 -16032
rect 8315 -16066 8331 -16048
rect 8197 -16082 8235 -16066
rect 8115 -16120 8235 -16082
rect 8293 -16082 8331 -16066
rect 8375 -16066 8391 -16048
rect 8493 -16048 8569 -16032
rect 8493 -16066 8509 -16048
rect 8375 -16082 8413 -16066
rect 8293 -16120 8413 -16082
rect 8471 -16082 8509 -16066
rect 8553 -16066 8569 -16048
rect 8671 -16048 8747 -16032
rect 8671 -16066 8687 -16048
rect 8553 -16082 8591 -16066
rect 8471 -16120 8591 -16082
rect 8649 -16082 8687 -16066
rect 8731 -16066 8747 -16048
rect 8849 -16048 8925 -16032
rect 8849 -16066 8865 -16048
rect 8731 -16082 8769 -16066
rect 8649 -16120 8769 -16082
rect 8827 -16082 8865 -16066
rect 8909 -16066 8925 -16048
rect 9027 -16048 9103 -16032
rect 9027 -16066 9043 -16048
rect 8909 -16082 8947 -16066
rect 8827 -16120 8947 -16082
rect 9005 -16082 9043 -16066
rect 9087 -16066 9103 -16048
rect 9205 -16048 9281 -16032
rect 9205 -16066 9221 -16048
rect 9087 -16082 9125 -16066
rect 9005 -16120 9125 -16082
rect 9183 -16082 9221 -16066
rect 9265 -16066 9281 -16048
rect 9383 -16048 9459 -16032
rect 9383 -16066 9399 -16048
rect 9265 -16082 9303 -16066
rect 9183 -16120 9303 -16082
rect 9361 -16082 9399 -16066
rect 9443 -16066 9459 -16048
rect 9561 -16048 9637 -16032
rect 9561 -16066 9577 -16048
rect 9443 -16082 9481 -16066
rect 9361 -16120 9481 -16082
rect 9539 -16082 9577 -16066
rect 9621 -16066 9637 -16048
rect 9739 -16048 9815 -16032
rect 9739 -16066 9755 -16048
rect 9621 -16082 9659 -16066
rect 9539 -16120 9659 -16082
rect 9717 -16082 9755 -16066
rect 9799 -16066 9815 -16048
rect 9917 -16048 9993 -16032
rect 9917 -16066 9933 -16048
rect 9799 -16082 9837 -16066
rect 9717 -16120 9837 -16082
rect 9895 -16082 9933 -16066
rect 9977 -16066 9993 -16048
rect 10095 -16048 10171 -16032
rect 10095 -16066 10111 -16048
rect 9977 -16082 10015 -16066
rect 9895 -16120 10015 -16082
rect 10073 -16082 10111 -16066
rect 10155 -16066 10171 -16048
rect 10273 -16048 10349 -16032
rect 10273 -16066 10289 -16048
rect 10155 -16082 10193 -16066
rect 10073 -16120 10193 -16082
rect 10251 -16082 10289 -16066
rect 10333 -16066 10349 -16048
rect 10451 -16048 10527 -16032
rect 10451 -16066 10467 -16048
rect 10333 -16082 10371 -16066
rect 10251 -16120 10371 -16082
rect 10429 -16082 10467 -16066
rect 10511 -16066 10527 -16048
rect 10629 -16048 10705 -16032
rect 10629 -16066 10645 -16048
rect 10511 -16082 10549 -16066
rect 10429 -16120 10549 -16082
rect 10607 -16082 10645 -16066
rect 10689 -16066 10705 -16048
rect 10807 -16048 10883 -16032
rect 10807 -16066 10823 -16048
rect 10689 -16082 10727 -16066
rect 10607 -16120 10727 -16082
rect 10785 -16082 10823 -16066
rect 10867 -16066 10883 -16048
rect 10985 -16048 11061 -16032
rect 10985 -16066 11001 -16048
rect 10867 -16082 10905 -16066
rect 10785 -16120 10905 -16082
rect 10963 -16082 11001 -16066
rect 11045 -16066 11061 -16048
rect 11163 -16048 11239 -16032
rect 11163 -16066 11179 -16048
rect 11045 -16082 11083 -16066
rect 10963 -16120 11083 -16082
rect 11141 -16082 11179 -16066
rect 11223 -16066 11239 -16048
rect 11341 -16048 11417 -16032
rect 11341 -16066 11357 -16048
rect 11223 -16082 11261 -16066
rect 11141 -16120 11261 -16082
rect 11319 -16082 11357 -16066
rect 11401 -16066 11417 -16048
rect 11519 -16048 11595 -16032
rect 11519 -16066 11535 -16048
rect 11401 -16082 11439 -16066
rect 11319 -16120 11439 -16082
rect 11497 -16082 11535 -16066
rect 11579 -16066 11595 -16048
rect 11697 -16048 11773 -16032
rect 11697 -16066 11713 -16048
rect 11579 -16082 11617 -16066
rect 11497 -16120 11617 -16082
rect 11675 -16082 11713 -16066
rect 11757 -16066 11773 -16048
rect 11875 -16048 11951 -16032
rect 11875 -16066 11891 -16048
rect 11757 -16082 11795 -16066
rect 11675 -16120 11795 -16082
rect 11853 -16082 11891 -16066
rect 11935 -16066 11951 -16048
rect 12053 -16048 12129 -16032
rect 12053 -16066 12069 -16048
rect 11935 -16082 11973 -16066
rect 11853 -16120 11973 -16082
rect 12031 -16082 12069 -16066
rect 12113 -16066 12129 -16048
rect 12231 -16048 12307 -16032
rect 12231 -16066 12247 -16048
rect 12113 -16082 12151 -16066
rect 12031 -16120 12151 -16082
rect 12209 -16082 12247 -16066
rect 12291 -16066 12307 -16048
rect 12409 -16048 12485 -16032
rect 12409 -16066 12425 -16048
rect 12291 -16082 12329 -16066
rect 12209 -16120 12329 -16082
rect 12387 -16082 12425 -16066
rect 12469 -16066 12485 -16048
rect 12587 -16048 12663 -16032
rect 12587 -16066 12603 -16048
rect 12469 -16082 12507 -16066
rect 12387 -16120 12507 -16082
rect 12565 -16082 12603 -16066
rect 12647 -16066 12663 -16048
rect 12647 -16082 12685 -16066
rect 12565 -16120 12685 -16082
rect -4180 -16150 -4104 -16134
rect -5960 -16410 -5884 -16394
rect -5960 -16428 -5944 -16410
rect -5982 -16444 -5944 -16428
rect -5900 -16428 -5884 -16410
rect -5782 -16410 -5706 -16394
rect -5782 -16428 -5766 -16410
rect -5900 -16444 -5862 -16428
rect -5982 -16482 -5862 -16444
rect -5804 -16444 -5766 -16428
rect -5722 -16428 -5706 -16410
rect -5604 -16410 -5528 -16394
rect -5604 -16428 -5588 -16410
rect -5722 -16444 -5684 -16428
rect -5804 -16482 -5684 -16444
rect -5626 -16444 -5588 -16428
rect -5544 -16428 -5528 -16410
rect -5426 -16410 -5350 -16394
rect -5426 -16428 -5410 -16410
rect -5544 -16444 -5506 -16428
rect -5626 -16482 -5506 -16444
rect -5448 -16444 -5410 -16428
rect -5366 -16428 -5350 -16410
rect -5248 -16410 -5172 -16394
rect -5248 -16428 -5232 -16410
rect -5366 -16444 -5328 -16428
rect -5448 -16482 -5328 -16444
rect -5270 -16444 -5232 -16428
rect -5188 -16428 -5172 -16410
rect -5070 -16410 -4994 -16394
rect -5070 -16428 -5054 -16410
rect -5188 -16444 -5150 -16428
rect -5270 -16482 -5150 -16444
rect -5092 -16444 -5054 -16428
rect -5010 -16428 -4994 -16410
rect -4892 -16410 -4816 -16394
rect -4892 -16428 -4876 -16410
rect -5010 -16444 -4972 -16428
rect -5092 -16482 -4972 -16444
rect -4914 -16444 -4876 -16428
rect -4832 -16428 -4816 -16410
rect -4714 -16410 -4638 -16394
rect -4714 -16428 -4698 -16410
rect -4832 -16444 -4794 -16428
rect -4914 -16482 -4794 -16444
rect -4736 -16444 -4698 -16428
rect -4654 -16428 -4638 -16410
rect -4536 -16410 -4460 -16394
rect -4536 -16428 -4520 -16410
rect -4654 -16444 -4616 -16428
rect -4736 -16482 -4616 -16444
rect -4558 -16444 -4520 -16428
rect -4476 -16428 -4460 -16410
rect -4358 -16410 -4282 -16394
rect -4358 -16428 -4342 -16410
rect -4476 -16444 -4438 -16428
rect -4558 -16482 -4438 -16444
rect -4380 -16444 -4342 -16428
rect -4298 -16428 -4282 -16410
rect -4180 -16410 -4104 -16394
rect -4180 -16428 -4164 -16410
rect -4298 -16444 -4260 -16428
rect -4380 -16482 -4260 -16444
rect -4202 -16444 -4164 -16428
rect -4120 -16428 -4104 -16410
rect -4120 -16444 -4082 -16428
rect -4202 -16482 -4082 -16444
rect -2127 -16438 -2007 -16400
rect -2127 -16454 -2089 -16438
rect -2105 -16472 -2089 -16454
rect -2045 -16454 -2007 -16438
rect -1949 -16438 -1829 -16400
rect -1949 -16454 -1911 -16438
rect -2045 -16472 -2029 -16454
rect -2105 -16488 -2029 -16472
rect -1927 -16472 -1911 -16454
rect -1867 -16454 -1829 -16438
rect -1771 -16438 -1651 -16400
rect -1771 -16454 -1733 -16438
rect -1867 -16472 -1851 -16454
rect -1927 -16488 -1851 -16472
rect -1749 -16472 -1733 -16454
rect -1689 -16454 -1651 -16438
rect -1593 -16438 -1473 -16400
rect -1593 -16454 -1555 -16438
rect -1689 -16472 -1673 -16454
rect -1749 -16488 -1673 -16472
rect -1571 -16472 -1555 -16454
rect -1511 -16454 -1473 -16438
rect -1415 -16438 -1295 -16400
rect -1415 -16454 -1377 -16438
rect -1511 -16472 -1495 -16454
rect -1571 -16488 -1495 -16472
rect -1393 -16472 -1377 -16454
rect -1333 -16454 -1295 -16438
rect -1237 -16438 -1117 -16400
rect -1237 -16454 -1199 -16438
rect -1333 -16472 -1317 -16454
rect -1393 -16488 -1317 -16472
rect -1215 -16472 -1199 -16454
rect -1155 -16454 -1117 -16438
rect -1059 -16438 -939 -16400
rect -1059 -16454 -1021 -16438
rect -1155 -16472 -1139 -16454
rect -1215 -16488 -1139 -16472
rect -1037 -16472 -1021 -16454
rect -977 -16454 -939 -16438
rect -881 -16438 -761 -16400
rect -881 -16454 -843 -16438
rect -977 -16472 -961 -16454
rect -1037 -16488 -961 -16472
rect -859 -16472 -843 -16454
rect -799 -16454 -761 -16438
rect -703 -16438 -583 -16400
rect -703 -16454 -665 -16438
rect -799 -16472 -783 -16454
rect -859 -16488 -783 -16472
rect -681 -16472 -665 -16454
rect -621 -16454 -583 -16438
rect -525 -16438 -405 -16400
rect -525 -16454 -487 -16438
rect -621 -16472 -605 -16454
rect -681 -16488 -605 -16472
rect -503 -16472 -487 -16454
rect -443 -16454 -405 -16438
rect -347 -16438 -227 -16400
rect -347 -16454 -309 -16438
rect -443 -16472 -427 -16454
rect -503 -16488 -427 -16472
rect -325 -16472 -309 -16454
rect -265 -16454 -227 -16438
rect -169 -16438 -49 -16400
rect -169 -16454 -131 -16438
rect -265 -16472 -249 -16454
rect -325 -16488 -249 -16472
rect -147 -16472 -131 -16454
rect -87 -16454 -49 -16438
rect 9 -16438 129 -16400
rect 9 -16454 47 -16438
rect -87 -16472 -71 -16454
rect -147 -16488 -71 -16472
rect 31 -16472 47 -16454
rect 91 -16454 129 -16438
rect 187 -16438 307 -16400
rect 187 -16454 225 -16438
rect 91 -16472 107 -16454
rect 31 -16488 107 -16472
rect 209 -16472 225 -16454
rect 269 -16454 307 -16438
rect 365 -16438 485 -16400
rect 365 -16454 403 -16438
rect 269 -16472 285 -16454
rect 209 -16488 285 -16472
rect 387 -16472 403 -16454
rect 447 -16454 485 -16438
rect 543 -16438 663 -16400
rect 543 -16454 581 -16438
rect 447 -16472 463 -16454
rect 387 -16488 463 -16472
rect 565 -16472 581 -16454
rect 625 -16454 663 -16438
rect 721 -16438 841 -16400
rect 721 -16454 759 -16438
rect 625 -16472 641 -16454
rect 565 -16488 641 -16472
rect 743 -16472 759 -16454
rect 803 -16454 841 -16438
rect 899 -16438 1019 -16400
rect 899 -16454 937 -16438
rect 803 -16472 819 -16454
rect 743 -16488 819 -16472
rect 921 -16472 937 -16454
rect 981 -16454 1019 -16438
rect 1077 -16438 1197 -16400
rect 1077 -16454 1115 -16438
rect 981 -16472 997 -16454
rect 921 -16488 997 -16472
rect 1099 -16472 1115 -16454
rect 1159 -16454 1197 -16438
rect 1255 -16438 1375 -16400
rect 1255 -16454 1293 -16438
rect 1159 -16472 1175 -16454
rect 1099 -16488 1175 -16472
rect 1277 -16472 1293 -16454
rect 1337 -16454 1375 -16438
rect 1433 -16438 1553 -16400
rect 1433 -16454 1471 -16438
rect 1337 -16472 1353 -16454
rect 1277 -16488 1353 -16472
rect 1455 -16472 1471 -16454
rect 1515 -16454 1553 -16438
rect 1611 -16438 1731 -16400
rect 1611 -16454 1649 -16438
rect 1515 -16472 1531 -16454
rect 1455 -16488 1531 -16472
rect 1633 -16472 1649 -16454
rect 1693 -16454 1731 -16438
rect 1789 -16438 1909 -16400
rect 1789 -16454 1827 -16438
rect 1693 -16472 1709 -16454
rect 1633 -16488 1709 -16472
rect 1811 -16472 1827 -16454
rect 1871 -16454 1909 -16438
rect 1967 -16438 2087 -16400
rect 1967 -16454 2005 -16438
rect 1871 -16472 1887 -16454
rect 1811 -16488 1887 -16472
rect 1989 -16472 2005 -16454
rect 2049 -16454 2087 -16438
rect 2145 -16438 2265 -16400
rect 2145 -16454 2183 -16438
rect 2049 -16472 2065 -16454
rect 1989 -16488 2065 -16472
rect 2167 -16472 2183 -16454
rect 2227 -16454 2265 -16438
rect 2323 -16438 2443 -16400
rect 2323 -16454 2361 -16438
rect 2227 -16472 2243 -16454
rect 2167 -16488 2243 -16472
rect 2345 -16472 2361 -16454
rect 2405 -16454 2443 -16438
rect 2501 -16438 2621 -16400
rect 2501 -16454 2539 -16438
rect 2405 -16472 2421 -16454
rect 2345 -16488 2421 -16472
rect 2523 -16472 2539 -16454
rect 2583 -16454 2621 -16438
rect 2679 -16438 2799 -16400
rect 2679 -16454 2717 -16438
rect 2583 -16472 2599 -16454
rect 2523 -16488 2599 -16472
rect 2701 -16472 2717 -16454
rect 2761 -16454 2799 -16438
rect 2857 -16438 2977 -16400
rect 2857 -16454 2895 -16438
rect 2761 -16472 2777 -16454
rect 2701 -16488 2777 -16472
rect 2879 -16472 2895 -16454
rect 2939 -16454 2977 -16438
rect 3035 -16438 3155 -16400
rect 3035 -16454 3073 -16438
rect 2939 -16472 2955 -16454
rect 2879 -16488 2955 -16472
rect 3057 -16472 3073 -16454
rect 3117 -16454 3155 -16438
rect 3213 -16438 3333 -16400
rect 3213 -16454 3251 -16438
rect 3117 -16472 3133 -16454
rect 3057 -16488 3133 -16472
rect 3235 -16472 3251 -16454
rect 3295 -16454 3333 -16438
rect 3391 -16438 3511 -16400
rect 3391 -16454 3429 -16438
rect 3295 -16472 3311 -16454
rect 3235 -16488 3311 -16472
rect 3413 -16472 3429 -16454
rect 3473 -16454 3511 -16438
rect 3569 -16438 3689 -16400
rect 3569 -16454 3607 -16438
rect 3473 -16472 3489 -16454
rect 3413 -16488 3489 -16472
rect 3591 -16472 3607 -16454
rect 3651 -16454 3689 -16438
rect 3747 -16438 3867 -16400
rect 3747 -16454 3785 -16438
rect 3651 -16472 3667 -16454
rect 3591 -16488 3667 -16472
rect 3769 -16472 3785 -16454
rect 3829 -16454 3867 -16438
rect 3925 -16438 4045 -16400
rect 3925 -16454 3963 -16438
rect 3829 -16472 3845 -16454
rect 3769 -16488 3845 -16472
rect 3947 -16472 3963 -16454
rect 4007 -16454 4045 -16438
rect 5623 -16438 5743 -16400
rect 5623 -16454 5661 -16438
rect 4007 -16472 4023 -16454
rect 3947 -16488 4023 -16472
rect 5645 -16472 5661 -16454
rect 5705 -16454 5743 -16438
rect 5801 -16438 5921 -16400
rect 5801 -16454 5839 -16438
rect 5705 -16472 5721 -16454
rect 5645 -16488 5721 -16472
rect 5823 -16472 5839 -16454
rect 5883 -16454 5921 -16438
rect 5979 -16438 6099 -16400
rect 5979 -16454 6017 -16438
rect 5883 -16472 5899 -16454
rect 5823 -16488 5899 -16472
rect 6001 -16472 6017 -16454
rect 6061 -16454 6099 -16438
rect 6157 -16438 6277 -16400
rect 6157 -16454 6195 -16438
rect 6061 -16472 6077 -16454
rect 6001 -16488 6077 -16472
rect 6179 -16472 6195 -16454
rect 6239 -16454 6277 -16438
rect 6335 -16438 6455 -16400
rect 6335 -16454 6373 -16438
rect 6239 -16472 6255 -16454
rect 6179 -16488 6255 -16472
rect 6357 -16472 6373 -16454
rect 6417 -16454 6455 -16438
rect 6513 -16438 6633 -16400
rect 6513 -16454 6551 -16438
rect 6417 -16472 6433 -16454
rect 6357 -16488 6433 -16472
rect 6535 -16472 6551 -16454
rect 6595 -16454 6633 -16438
rect 6691 -16438 6811 -16400
rect 6691 -16454 6729 -16438
rect 6595 -16472 6611 -16454
rect 6535 -16488 6611 -16472
rect 6713 -16472 6729 -16454
rect 6773 -16454 6811 -16438
rect 6869 -16438 6989 -16400
rect 6869 -16454 6907 -16438
rect 6773 -16472 6789 -16454
rect 6713 -16488 6789 -16472
rect 6891 -16472 6907 -16454
rect 6951 -16454 6989 -16438
rect 7047 -16438 7167 -16400
rect 7047 -16454 7085 -16438
rect 6951 -16472 6967 -16454
rect 6891 -16488 6967 -16472
rect 7069 -16472 7085 -16454
rect 7129 -16454 7167 -16438
rect 7225 -16438 7345 -16400
rect 7225 -16454 7263 -16438
rect 7129 -16472 7145 -16454
rect 7069 -16488 7145 -16472
rect 7247 -16472 7263 -16454
rect 7307 -16454 7345 -16438
rect 7403 -16438 7523 -16400
rect 7403 -16454 7441 -16438
rect 7307 -16472 7323 -16454
rect 7247 -16488 7323 -16472
rect 7425 -16472 7441 -16454
rect 7485 -16454 7523 -16438
rect 7581 -16438 7701 -16400
rect 7581 -16454 7619 -16438
rect 7485 -16472 7501 -16454
rect 7425 -16488 7501 -16472
rect 7603 -16472 7619 -16454
rect 7663 -16454 7701 -16438
rect 7759 -16438 7879 -16400
rect 7759 -16454 7797 -16438
rect 7663 -16472 7679 -16454
rect 7603 -16488 7679 -16472
rect 7781 -16472 7797 -16454
rect 7841 -16454 7879 -16438
rect 7937 -16438 8057 -16400
rect 7937 -16454 7975 -16438
rect 7841 -16472 7857 -16454
rect 7781 -16488 7857 -16472
rect 7959 -16472 7975 -16454
rect 8019 -16454 8057 -16438
rect 8115 -16438 8235 -16400
rect 8115 -16454 8153 -16438
rect 8019 -16472 8035 -16454
rect 7959 -16488 8035 -16472
rect 8137 -16472 8153 -16454
rect 8197 -16454 8235 -16438
rect 8293 -16438 8413 -16400
rect 8293 -16454 8331 -16438
rect 8197 -16472 8213 -16454
rect 8137 -16488 8213 -16472
rect 8315 -16472 8331 -16454
rect 8375 -16454 8413 -16438
rect 8471 -16438 8591 -16400
rect 8471 -16454 8509 -16438
rect 8375 -16472 8391 -16454
rect 8315 -16488 8391 -16472
rect 8493 -16472 8509 -16454
rect 8553 -16454 8591 -16438
rect 8649 -16438 8769 -16400
rect 8649 -16454 8687 -16438
rect 8553 -16472 8569 -16454
rect 8493 -16488 8569 -16472
rect 8671 -16472 8687 -16454
rect 8731 -16454 8769 -16438
rect 8827 -16438 8947 -16400
rect 8827 -16454 8865 -16438
rect 8731 -16472 8747 -16454
rect 8671 -16488 8747 -16472
rect 8849 -16472 8865 -16454
rect 8909 -16454 8947 -16438
rect 9005 -16438 9125 -16400
rect 9005 -16454 9043 -16438
rect 8909 -16472 8925 -16454
rect 8849 -16488 8925 -16472
rect 9027 -16472 9043 -16454
rect 9087 -16454 9125 -16438
rect 9183 -16438 9303 -16400
rect 9183 -16454 9221 -16438
rect 9087 -16472 9103 -16454
rect 9027 -16488 9103 -16472
rect 9205 -16472 9221 -16454
rect 9265 -16454 9303 -16438
rect 9361 -16438 9481 -16400
rect 9361 -16454 9399 -16438
rect 9265 -16472 9281 -16454
rect 9205 -16488 9281 -16472
rect 9383 -16472 9399 -16454
rect 9443 -16454 9481 -16438
rect 9539 -16438 9659 -16400
rect 9539 -16454 9577 -16438
rect 9443 -16472 9459 -16454
rect 9383 -16488 9459 -16472
rect 9561 -16472 9577 -16454
rect 9621 -16454 9659 -16438
rect 9717 -16438 9837 -16400
rect 9717 -16454 9755 -16438
rect 9621 -16472 9637 -16454
rect 9561 -16488 9637 -16472
rect 9739 -16472 9755 -16454
rect 9799 -16454 9837 -16438
rect 9895 -16438 10015 -16400
rect 9895 -16454 9933 -16438
rect 9799 -16472 9815 -16454
rect 9739 -16488 9815 -16472
rect 9917 -16472 9933 -16454
rect 9977 -16454 10015 -16438
rect 10073 -16438 10193 -16400
rect 10073 -16454 10111 -16438
rect 9977 -16472 9993 -16454
rect 9917 -16488 9993 -16472
rect 10095 -16472 10111 -16454
rect 10155 -16454 10193 -16438
rect 10251 -16438 10371 -16400
rect 10251 -16454 10289 -16438
rect 10155 -16472 10171 -16454
rect 10095 -16488 10171 -16472
rect 10273 -16472 10289 -16454
rect 10333 -16454 10371 -16438
rect 10429 -16438 10549 -16400
rect 10429 -16454 10467 -16438
rect 10333 -16472 10349 -16454
rect 10273 -16488 10349 -16472
rect 10451 -16472 10467 -16454
rect 10511 -16454 10549 -16438
rect 10607 -16438 10727 -16400
rect 10607 -16454 10645 -16438
rect 10511 -16472 10527 -16454
rect 10451 -16488 10527 -16472
rect 10629 -16472 10645 -16454
rect 10689 -16454 10727 -16438
rect 10785 -16438 10905 -16400
rect 10785 -16454 10823 -16438
rect 10689 -16472 10705 -16454
rect 10629 -16488 10705 -16472
rect 10807 -16472 10823 -16454
rect 10867 -16454 10905 -16438
rect 10963 -16438 11083 -16400
rect 10963 -16454 11001 -16438
rect 10867 -16472 10883 -16454
rect 10807 -16488 10883 -16472
rect 10985 -16472 11001 -16454
rect 11045 -16454 11083 -16438
rect 11141 -16438 11261 -16400
rect 11141 -16454 11179 -16438
rect 11045 -16472 11061 -16454
rect 10985 -16488 11061 -16472
rect 11163 -16472 11179 -16454
rect 11223 -16454 11261 -16438
rect 11319 -16438 11439 -16400
rect 11319 -16454 11357 -16438
rect 11223 -16472 11239 -16454
rect 11163 -16488 11239 -16472
rect 11341 -16472 11357 -16454
rect 11401 -16454 11439 -16438
rect 11497 -16438 11617 -16400
rect 11497 -16454 11535 -16438
rect 11401 -16472 11417 -16454
rect 11341 -16488 11417 -16472
rect 11519 -16472 11535 -16454
rect 11579 -16454 11617 -16438
rect 11675 -16438 11795 -16400
rect 11675 -16454 11713 -16438
rect 11579 -16472 11595 -16454
rect 11519 -16488 11595 -16472
rect 11697 -16472 11713 -16454
rect 11757 -16454 11795 -16438
rect 11853 -16438 11973 -16400
rect 11853 -16454 11891 -16438
rect 11757 -16472 11773 -16454
rect 11697 -16488 11773 -16472
rect 11875 -16472 11891 -16454
rect 11935 -16454 11973 -16438
rect 12031 -16438 12151 -16400
rect 12031 -16454 12069 -16438
rect 11935 -16472 11951 -16454
rect 11875 -16488 11951 -16472
rect 12053 -16472 12069 -16454
rect 12113 -16454 12151 -16438
rect 12209 -16438 12329 -16400
rect 12209 -16454 12247 -16438
rect 12113 -16472 12129 -16454
rect 12053 -16488 12129 -16472
rect 12231 -16472 12247 -16454
rect 12291 -16454 12329 -16438
rect 12387 -16438 12507 -16400
rect 12387 -16454 12425 -16438
rect 12291 -16472 12307 -16454
rect 12231 -16488 12307 -16472
rect 12409 -16472 12425 -16454
rect 12469 -16454 12507 -16438
rect 12565 -16438 12685 -16400
rect 12565 -16454 12603 -16438
rect 12469 -16472 12485 -16454
rect 12409 -16488 12485 -16472
rect 12587 -16472 12603 -16454
rect 12647 -16454 12685 -16438
rect 12647 -16472 12663 -16454
rect 12587 -16488 12663 -16472
rect -5982 -16800 -5862 -16762
rect -5982 -16816 -5944 -16800
rect -5960 -16834 -5944 -16816
rect -5900 -16816 -5862 -16800
rect -5804 -16800 -5684 -16762
rect -5804 -16816 -5766 -16800
rect -5900 -16834 -5884 -16816
rect -5960 -16850 -5884 -16834
rect -5782 -16834 -5766 -16816
rect -5722 -16816 -5684 -16800
rect -5626 -16800 -5506 -16762
rect -5626 -16816 -5588 -16800
rect -5722 -16834 -5706 -16816
rect -5782 -16850 -5706 -16834
rect -5604 -16834 -5588 -16816
rect -5544 -16816 -5506 -16800
rect -5448 -16800 -5328 -16762
rect -5448 -16816 -5410 -16800
rect -5544 -16834 -5528 -16816
rect -5604 -16850 -5528 -16834
rect -5426 -16834 -5410 -16816
rect -5366 -16816 -5328 -16800
rect -5270 -16800 -5150 -16762
rect -5270 -16816 -5232 -16800
rect -5366 -16834 -5350 -16816
rect -5426 -16850 -5350 -16834
rect -5248 -16834 -5232 -16816
rect -5188 -16816 -5150 -16800
rect -5092 -16800 -4972 -16762
rect -5092 -16816 -5054 -16800
rect -5188 -16834 -5172 -16816
rect -5248 -16850 -5172 -16834
rect -5070 -16834 -5054 -16816
rect -5010 -16816 -4972 -16800
rect -4914 -16800 -4794 -16762
rect -4914 -16816 -4876 -16800
rect -5010 -16834 -4994 -16816
rect -5070 -16850 -4994 -16834
rect -4892 -16834 -4876 -16816
rect -4832 -16816 -4794 -16800
rect -4736 -16800 -4616 -16762
rect -4736 -16816 -4698 -16800
rect -4832 -16834 -4816 -16816
rect -4892 -16850 -4816 -16834
rect -4714 -16834 -4698 -16816
rect -4654 -16816 -4616 -16800
rect -4558 -16800 -4438 -16762
rect -4558 -16816 -4520 -16800
rect -4654 -16834 -4638 -16816
rect -4714 -16850 -4638 -16834
rect -4536 -16834 -4520 -16816
rect -4476 -16816 -4438 -16800
rect -4380 -16800 -4260 -16762
rect -4380 -16816 -4342 -16800
rect -4476 -16834 -4460 -16816
rect -4536 -16850 -4460 -16834
rect -4358 -16834 -4342 -16816
rect -4298 -16816 -4260 -16800
rect -4202 -16800 -4082 -16762
rect -4202 -16816 -4164 -16800
rect -4298 -16834 -4282 -16816
rect -4358 -16850 -4282 -16834
rect -4180 -16834 -4164 -16816
rect -4120 -16816 -4082 -16800
rect -4120 -16834 -4104 -16816
rect -4180 -16850 -4104 -16834
<< polycont >>
rect 7154 2673 7188 2707
rect 7346 2673 7380 2707
rect 7538 2673 7572 2707
rect 7730 2673 7764 2707
rect 7922 2673 7956 2707
rect 8114 2673 8148 2707
rect 16154 2673 16188 2707
rect 16346 2673 16380 2707
rect 16538 2673 16572 2707
rect 16730 2673 16764 2707
rect 16922 2673 16956 2707
rect 17114 2673 17148 2707
rect 7154 1865 7188 1899
rect 7346 1865 7380 1899
rect 7538 1865 7572 1899
rect 7730 1865 7764 1899
rect 7922 1865 7956 1899
rect 8114 1865 8148 1899
rect 16154 1865 16188 1899
rect 16346 1865 16380 1899
rect 16538 1865 16572 1899
rect 16730 1865 16764 1899
rect 16922 1865 16956 1899
rect 17114 1865 17148 1899
rect 7154 873 7188 907
rect 7346 873 7380 907
rect 7538 873 7572 907
rect 7730 873 7764 907
rect 7922 873 7956 907
rect 8114 873 8148 907
rect 16154 873 16188 907
rect 16346 873 16380 907
rect 16538 873 16572 907
rect 16730 873 16764 907
rect 16922 873 16956 907
rect 17114 873 17148 907
rect 7154 65 7188 99
rect 7346 65 7380 99
rect 7538 65 7572 99
rect 7730 65 7764 99
rect 7922 65 7956 99
rect 8114 65 8148 99
rect 16154 65 16188 99
rect 16346 65 16380 99
rect 16538 65 16572 99
rect 16730 65 16764 99
rect 16922 65 16956 99
rect 17114 65 17148 99
rect 7154 -927 7188 -893
rect 7346 -927 7380 -893
rect 7538 -927 7572 -893
rect 7730 -927 7764 -893
rect 7922 -927 7956 -893
rect 8114 -927 8148 -893
rect 16154 -927 16188 -893
rect 16346 -927 16380 -893
rect 16538 -927 16572 -893
rect 16730 -927 16764 -893
rect 16922 -927 16956 -893
rect 17114 -927 17148 -893
rect -6218 -2073 -6174 -2039
rect -6040 -2073 -5996 -2039
rect -5862 -2073 -5818 -2039
rect -5684 -2073 -5640 -2039
rect -5506 -2073 -5462 -2039
rect -5328 -2073 -5284 -2039
rect -5150 -2073 -5106 -2039
rect -4972 -2073 -4928 -2039
rect -4794 -2073 -4750 -2039
rect -4616 -2073 -4572 -2039
rect -4438 -2073 -4394 -2039
rect -4260 -2073 -4216 -2039
rect -4082 -2073 -4038 -2039
rect -3904 -2073 -3860 -2039
rect -3726 -2073 -3682 -2039
rect -3548 -2073 -3504 -2039
rect -6218 -2481 -6174 -2447
rect -6040 -2481 -5996 -2447
rect -5862 -2481 -5818 -2447
rect -5684 -2481 -5640 -2447
rect -5506 -2481 -5462 -2447
rect -5328 -2481 -5284 -2447
rect -5150 -2481 -5106 -2447
rect -4972 -2481 -4928 -2447
rect -4794 -2481 -4750 -2447
rect -4616 -2481 -4572 -2447
rect -4438 -2481 -4394 -2447
rect -4260 -2481 -4216 -2447
rect -4082 -2481 -4038 -2447
rect -3904 -2481 -3860 -2447
rect -3726 -2481 -3682 -2447
rect -3548 -2481 -3504 -2447
rect -1370 -2825 -1326 -2791
rect -1192 -2825 -1148 -2791
rect -1014 -2825 -970 -2791
rect -836 -2825 -792 -2791
rect -658 -2825 -614 -2791
rect -480 -2825 -436 -2791
rect -302 -2825 -258 -2791
rect -124 -2825 -80 -2791
rect 54 -2825 98 -2791
rect 232 -2825 276 -2791
rect 410 -2825 454 -2791
rect 588 -2825 632 -2791
rect 766 -2825 810 -2791
rect 944 -2825 988 -2791
rect 1122 -2825 1166 -2791
rect 1300 -2825 1344 -2791
rect 1478 -2825 1522 -2791
rect 1656 -2825 1700 -2791
rect 1834 -2825 1878 -2791
rect 2012 -2825 2056 -2791
rect 2190 -2825 2234 -2791
rect 2368 -2825 2412 -2791
rect 2546 -2825 2590 -2791
rect -6218 -2943 -6174 -2909
rect -6040 -2943 -5996 -2909
rect -5862 -2943 -5818 -2909
rect -5684 -2943 -5640 -2909
rect -5506 -2943 -5462 -2909
rect -5328 -2943 -5284 -2909
rect -5150 -2943 -5106 -2909
rect -4972 -2943 -4928 -2909
rect -4794 -2943 -4750 -2909
rect -4616 -2943 -4572 -2909
rect -4438 -2943 -4394 -2909
rect -4260 -2943 -4216 -2909
rect -4082 -2943 -4038 -2909
rect -3904 -2943 -3860 -2909
rect -3726 -2943 -3682 -2909
rect -3548 -2943 -3504 -2909
rect -1370 -3233 -1326 -3199
rect -1192 -3233 -1148 -3199
rect -1014 -3233 -970 -3199
rect -836 -3233 -792 -3199
rect -658 -3233 -614 -3199
rect -480 -3233 -436 -3199
rect -302 -3233 -258 -3199
rect -124 -3233 -80 -3199
rect 54 -3233 98 -3199
rect 232 -3233 276 -3199
rect 410 -3233 454 -3199
rect 588 -3233 632 -3199
rect 766 -3233 810 -3199
rect 944 -3233 988 -3199
rect 1122 -3233 1166 -3199
rect 1300 -3233 1344 -3199
rect 1478 -3233 1522 -3199
rect 1656 -3233 1700 -3199
rect 1834 -3233 1878 -3199
rect 2012 -3233 2056 -3199
rect 2190 -3233 2234 -3199
rect 2368 -3233 2412 -3199
rect 2546 -3233 2590 -3199
rect -6218 -3351 -6174 -3317
rect -6040 -3351 -5996 -3317
rect -5862 -3351 -5818 -3317
rect -5684 -3351 -5640 -3317
rect -5506 -3351 -5462 -3317
rect -5328 -3351 -5284 -3317
rect -5150 -3351 -5106 -3317
rect -4972 -3351 -4928 -3317
rect -4794 -3351 -4750 -3317
rect -4616 -3351 -4572 -3317
rect -4438 -3351 -4394 -3317
rect -4260 -3351 -4216 -3317
rect -4082 -3351 -4038 -3317
rect -3904 -3351 -3860 -3317
rect -3726 -3351 -3682 -3317
rect -3548 -3351 -3504 -3317
rect -1370 -3725 -1326 -3691
rect -6218 -3813 -6174 -3779
rect -6040 -3813 -5996 -3779
rect -5862 -3813 -5818 -3779
rect -5684 -3813 -5640 -3779
rect -5506 -3813 -5462 -3779
rect -5328 -3813 -5284 -3779
rect -5150 -3813 -5106 -3779
rect -4972 -3813 -4928 -3779
rect -4794 -3813 -4750 -3779
rect -4616 -3813 -4572 -3779
rect -4438 -3813 -4394 -3779
rect -4260 -3813 -4216 -3779
rect -4082 -3813 -4038 -3779
rect -3904 -3813 -3860 -3779
rect -3726 -3813 -3682 -3779
rect -1192 -3725 -1148 -3691
rect -1014 -3725 -970 -3691
rect -836 -3725 -792 -3691
rect -658 -3725 -614 -3691
rect -480 -3725 -436 -3691
rect -302 -3725 -258 -3691
rect -124 -3725 -80 -3691
rect 54 -3725 98 -3691
rect 232 -3725 276 -3691
rect 410 -3725 454 -3691
rect 588 -3725 632 -3691
rect 766 -3725 810 -3691
rect 944 -3725 988 -3691
rect 1122 -3725 1166 -3691
rect 1300 -3725 1344 -3691
rect 1478 -3725 1522 -3691
rect 1656 -3725 1700 -3691
rect 1834 -3725 1878 -3691
rect 2012 -3725 2056 -3691
rect 2190 -3725 2234 -3691
rect 2368 -3725 2412 -3691
rect 2546 -3725 2590 -3691
rect -3548 -3813 -3504 -3779
rect -1370 -4133 -1326 -4099
rect -6218 -4221 -6174 -4187
rect -6040 -4221 -5996 -4187
rect -5862 -4221 -5818 -4187
rect -5684 -4221 -5640 -4187
rect -5506 -4221 -5462 -4187
rect -5328 -4221 -5284 -4187
rect -5150 -4221 -5106 -4187
rect -4972 -4221 -4928 -4187
rect -4794 -4221 -4750 -4187
rect -4616 -4221 -4572 -4187
rect -4438 -4221 -4394 -4187
rect -4260 -4221 -4216 -4187
rect -4082 -4221 -4038 -4187
rect -3904 -4221 -3860 -4187
rect -3726 -4221 -3682 -4187
rect -1192 -4133 -1148 -4099
rect -1014 -4133 -970 -4099
rect -836 -4133 -792 -4099
rect -658 -4133 -614 -4099
rect -480 -4133 -436 -4099
rect -302 -4133 -258 -4099
rect -124 -4133 -80 -4099
rect 54 -4133 98 -4099
rect 232 -4133 276 -4099
rect 410 -4133 454 -4099
rect 588 -4133 632 -4099
rect 766 -4133 810 -4099
rect 944 -4133 988 -4099
rect 1122 -4133 1166 -4099
rect 1300 -4133 1344 -4099
rect 1478 -4133 1522 -4099
rect 1656 -4133 1700 -4099
rect 1834 -4133 1878 -4099
rect 2012 -4133 2056 -4099
rect 2190 -4133 2234 -4099
rect 2368 -4133 2412 -4099
rect 2546 -4133 2590 -4099
rect -3548 -4221 -3504 -4187
rect -1370 -4625 -1326 -4591
rect -6218 -4683 -6174 -4649
rect -6040 -4683 -5996 -4649
rect -5862 -4683 -5818 -4649
rect -5684 -4683 -5640 -4649
rect -5506 -4683 -5462 -4649
rect -5328 -4683 -5284 -4649
rect -5150 -4683 -5106 -4649
rect -4972 -4683 -4928 -4649
rect -4794 -4683 -4750 -4649
rect -4616 -4683 -4572 -4649
rect -4438 -4683 -4394 -4649
rect -4260 -4683 -4216 -4649
rect -4082 -4683 -4038 -4649
rect -3904 -4683 -3860 -4649
rect -3726 -4683 -3682 -4649
rect -3548 -4683 -3504 -4649
rect -1192 -4625 -1148 -4591
rect -1014 -4625 -970 -4591
rect -836 -4625 -792 -4591
rect -658 -4625 -614 -4591
rect -480 -4625 -436 -4591
rect -302 -4625 -258 -4591
rect -124 -4625 -80 -4591
rect 54 -4625 98 -4591
rect 232 -4625 276 -4591
rect 410 -4625 454 -4591
rect 588 -4625 632 -4591
rect 766 -4625 810 -4591
rect 944 -4625 988 -4591
rect 1122 -4625 1166 -4591
rect 1300 -4625 1344 -4591
rect 1478 -4625 1522 -4591
rect 1656 -4625 1700 -4591
rect 1834 -4625 1878 -4591
rect 2012 -4625 2056 -4591
rect 2190 -4625 2234 -4591
rect 2368 -4625 2412 -4591
rect 2546 -4625 2590 -4591
rect -6218 -5091 -6174 -5057
rect -6040 -5091 -5996 -5057
rect -5862 -5091 -5818 -5057
rect -5684 -5091 -5640 -5057
rect -5506 -5091 -5462 -5057
rect -5328 -5091 -5284 -5057
rect -5150 -5091 -5106 -5057
rect -4972 -5091 -4928 -5057
rect -4794 -5091 -4750 -5057
rect -4616 -5091 -4572 -5057
rect -4438 -5091 -4394 -5057
rect -4260 -5091 -4216 -5057
rect -4082 -5091 -4038 -5057
rect -3904 -5091 -3860 -5057
rect -3726 -5091 -3682 -5057
rect -1370 -5033 -1326 -4999
rect -1192 -5033 -1148 -4999
rect -1014 -5033 -970 -4999
rect -836 -5033 -792 -4999
rect -658 -5033 -614 -4999
rect -480 -5033 -436 -4999
rect -302 -5033 -258 -4999
rect -124 -5033 -80 -4999
rect 54 -5033 98 -4999
rect 232 -5033 276 -4999
rect 410 -5033 454 -4999
rect 588 -5033 632 -4999
rect 766 -5033 810 -4999
rect 944 -5033 988 -4999
rect 1122 -5033 1166 -4999
rect 1300 -5033 1344 -4999
rect 1478 -5033 1522 -4999
rect 1656 -5033 1700 -4999
rect 1834 -5033 1878 -4999
rect 2012 -5033 2056 -4999
rect 2190 -5033 2234 -4999
rect 2368 -5033 2412 -4999
rect 2546 -5033 2590 -4999
rect -3548 -5091 -3504 -5057
rect -6218 -5553 -6174 -5519
rect -6040 -5553 -5996 -5519
rect -5862 -5553 -5818 -5519
rect -5684 -5553 -5640 -5519
rect -5506 -5553 -5462 -5519
rect -5328 -5553 -5284 -5519
rect -5150 -5553 -5106 -5519
rect -4972 -5553 -4928 -5519
rect -4794 -5553 -4750 -5519
rect -4616 -5553 -4572 -5519
rect -4438 -5553 -4394 -5519
rect -4260 -5553 -4216 -5519
rect -4082 -5553 -4038 -5519
rect -3904 -5553 -3860 -5519
rect -3726 -5553 -3682 -5519
rect -3548 -5553 -3504 -5519
rect -1370 -5525 -1326 -5491
rect -1192 -5525 -1148 -5491
rect -1014 -5525 -970 -5491
rect -836 -5525 -792 -5491
rect -658 -5525 -614 -5491
rect -480 -5525 -436 -5491
rect -302 -5525 -258 -5491
rect -124 -5525 -80 -5491
rect 54 -5525 98 -5491
rect 232 -5525 276 -5491
rect 410 -5525 454 -5491
rect 588 -5525 632 -5491
rect 766 -5525 810 -5491
rect 944 -5525 988 -5491
rect 1122 -5525 1166 -5491
rect 1300 -5525 1344 -5491
rect 1478 -5525 1522 -5491
rect 1656 -5525 1700 -5491
rect 1834 -5525 1878 -5491
rect 2012 -5525 2056 -5491
rect 2190 -5525 2234 -5491
rect 2368 -5525 2412 -5491
rect 2546 -5525 2590 -5491
rect -6218 -5961 -6174 -5927
rect -6040 -5961 -5996 -5927
rect -5862 -5961 -5818 -5927
rect -5684 -5961 -5640 -5927
rect -5506 -5961 -5462 -5927
rect -5328 -5961 -5284 -5927
rect -5150 -5961 -5106 -5927
rect -4972 -5961 -4928 -5927
rect -4794 -5961 -4750 -5927
rect -4616 -5961 -4572 -5927
rect -4438 -5961 -4394 -5927
rect -4260 -5961 -4216 -5927
rect -4082 -5961 -4038 -5927
rect -3904 -5961 -3860 -5927
rect -3726 -5961 -3682 -5927
rect -3548 -5961 -3504 -5927
rect -1370 -5933 -1326 -5899
rect -1192 -5933 -1148 -5899
rect -1014 -5933 -970 -5899
rect -836 -5933 -792 -5899
rect -658 -5933 -614 -5899
rect -480 -5933 -436 -5899
rect -302 -5933 -258 -5899
rect -124 -5933 -80 -5899
rect 54 -5933 98 -5899
rect 232 -5933 276 -5899
rect 410 -5933 454 -5899
rect 588 -5933 632 -5899
rect 766 -5933 810 -5899
rect 944 -5933 988 -5899
rect 1122 -5933 1166 -5899
rect 1300 -5933 1344 -5899
rect 1478 -5933 1522 -5899
rect 1656 -5933 1700 -5899
rect 1834 -5933 1878 -5899
rect 2012 -5933 2056 -5899
rect 2190 -5933 2234 -5899
rect 2368 -5933 2412 -5899
rect 2546 -5933 2590 -5899
rect 7154 -1735 7188 -1701
rect 7346 -1735 7380 -1701
rect 7538 -1735 7572 -1701
rect 7730 -1735 7764 -1701
rect 7922 -1735 7956 -1701
rect 8114 -1735 8148 -1701
rect 16154 -1735 16188 -1701
rect 16346 -1735 16380 -1701
rect 16538 -1735 16572 -1701
rect 16730 -1735 16764 -1701
rect 16922 -1735 16956 -1701
rect 17114 -1735 17148 -1701
rect 7154 -2727 7188 -2693
rect 7346 -2727 7380 -2693
rect 7538 -2727 7572 -2693
rect 7730 -2727 7764 -2693
rect 7922 -2727 7956 -2693
rect 8114 -2727 8148 -2693
rect 16154 -2727 16188 -2693
rect 16346 -2727 16380 -2693
rect 16538 -2727 16572 -2693
rect 16730 -2727 16764 -2693
rect 16922 -2727 16956 -2693
rect 17114 -2727 17148 -2693
rect 7154 -3535 7188 -3501
rect 7346 -3535 7380 -3501
rect 7538 -3535 7572 -3501
rect 7730 -3535 7764 -3501
rect 7922 -3535 7956 -3501
rect 8114 -3535 8148 -3501
rect 16154 -3535 16188 -3501
rect 16346 -3535 16380 -3501
rect 16538 -3535 16572 -3501
rect 16730 -3535 16764 -3501
rect 16922 -3535 16956 -3501
rect 17114 -3535 17148 -3501
rect 7154 -4527 7188 -4493
rect 7346 -4527 7380 -4493
rect 7538 -4527 7572 -4493
rect 7730 -4527 7764 -4493
rect 7922 -4527 7956 -4493
rect 8114 -4527 8148 -4493
rect 16154 -4527 16188 -4493
rect 16346 -4527 16380 -4493
rect 16538 -4527 16572 -4493
rect 16730 -4527 16764 -4493
rect 16922 -4527 16956 -4493
rect 17114 -4527 17148 -4493
rect 7154 -5335 7188 -5301
rect 7346 -5335 7380 -5301
rect 7538 -5335 7572 -5301
rect 7730 -5335 7764 -5301
rect 7922 -5335 7956 -5301
rect 8114 -5335 8148 -5301
rect 16154 -5335 16188 -5301
rect 16346 -5335 16380 -5301
rect 16538 -5335 16572 -5301
rect 16730 -5335 16764 -5301
rect 16922 -5335 16956 -5301
rect 17114 -5335 17148 -5301
rect 7154 -6327 7188 -6293
rect 7346 -6327 7380 -6293
rect 7538 -6327 7572 -6293
rect 7730 -6327 7764 -6293
rect 7922 -6327 7956 -6293
rect 8114 -6327 8148 -6293
rect 16154 -6327 16188 -6293
rect 16346 -6327 16380 -6293
rect 16538 -6327 16572 -6293
rect 16730 -6327 16764 -6293
rect 16922 -6327 16956 -6293
rect 17114 -6327 17148 -6293
rect 7154 -7135 7188 -7101
rect 7346 -7135 7380 -7101
rect 7538 -7135 7572 -7101
rect 7730 -7135 7764 -7101
rect 7922 -7135 7956 -7101
rect 8114 -7135 8148 -7101
rect 16154 -7135 16188 -7101
rect 16346 -7135 16380 -7101
rect 16538 -7135 16572 -7101
rect 16730 -7135 16764 -7101
rect 16922 -7135 16956 -7101
rect 17114 -7135 17148 -7101
rect -5544 -7824 -5500 -7790
rect -5366 -7824 -5322 -7790
rect -5188 -7824 -5144 -7790
rect -5010 -7824 -4966 -7790
rect -4832 -7824 -4788 -7790
rect -4654 -7824 -4610 -7790
rect -4476 -7824 -4432 -7790
rect -4298 -7824 -4254 -7790
rect -4120 -7824 -4076 -7790
rect -2089 -8082 -2045 -8048
rect -1911 -8082 -1867 -8048
rect -1733 -8082 -1689 -8048
rect -1555 -8082 -1511 -8048
rect -1377 -8082 -1333 -8048
rect -1199 -8082 -1155 -8048
rect -1021 -8082 -977 -8048
rect -843 -8082 -799 -8048
rect -665 -8082 -621 -8048
rect -487 -8082 -443 -8048
rect -309 -8082 -265 -8048
rect -131 -8082 -87 -8048
rect 47 -8082 91 -8048
rect 225 -8082 269 -8048
rect 403 -8082 447 -8048
rect 581 -8082 625 -8048
rect 759 -8082 803 -8048
rect 937 -8082 981 -8048
rect 1115 -8082 1159 -8048
rect 1293 -8082 1337 -8048
rect 1471 -8082 1515 -8048
rect 1649 -8082 1693 -8048
rect 1827 -8082 1871 -8048
rect 2005 -8082 2049 -8048
rect 2183 -8082 2227 -8048
rect 2361 -8082 2405 -8048
rect 2539 -8082 2583 -8048
rect 2717 -8082 2761 -8048
rect 2895 -8082 2939 -8048
rect 3073 -8082 3117 -8048
rect 3251 -8082 3295 -8048
rect 3429 -8082 3473 -8048
rect 3607 -8082 3651 -8048
rect 3785 -8082 3829 -8048
rect 3963 -8082 4007 -8048
rect -5544 -8214 -5500 -8180
rect -5366 -8214 -5322 -8180
rect -5188 -8214 -5144 -8180
rect -5010 -8214 -4966 -8180
rect -4832 -8214 -4788 -8180
rect -4654 -8214 -4610 -8180
rect -4476 -8214 -4432 -8180
rect -4298 -8214 -4254 -8180
rect -4120 -8214 -4076 -8180
rect -5544 -8374 -5500 -8340
rect -5366 -8374 -5322 -8340
rect -5188 -8374 -5144 -8340
rect -5010 -8374 -4966 -8340
rect -4832 -8374 -4788 -8340
rect -4654 -8374 -4610 -8340
rect -4476 -8374 -4432 -8340
rect -4298 -8374 -4254 -8340
rect -4120 -8374 -4076 -8340
rect -2089 -8472 -2045 -8438
rect -1911 -8472 -1867 -8438
rect -1733 -8472 -1689 -8438
rect -1555 -8472 -1511 -8438
rect -1377 -8472 -1333 -8438
rect -1199 -8472 -1155 -8438
rect -1021 -8472 -977 -8438
rect -843 -8472 -799 -8438
rect -665 -8472 -621 -8438
rect -487 -8472 -443 -8438
rect -309 -8472 -265 -8438
rect -131 -8472 -87 -8438
rect 47 -8472 91 -8438
rect 225 -8472 269 -8438
rect 403 -8472 447 -8438
rect 581 -8472 625 -8438
rect 759 -8472 803 -8438
rect 937 -8472 981 -8438
rect 1115 -8472 1159 -8438
rect 1293 -8472 1337 -8438
rect 1471 -8472 1515 -8438
rect 1649 -8472 1693 -8438
rect 1827 -8472 1871 -8438
rect 2005 -8472 2049 -8438
rect 2183 -8472 2227 -8438
rect 2361 -8472 2405 -8438
rect 2539 -8472 2583 -8438
rect 2717 -8472 2761 -8438
rect 2895 -8472 2939 -8438
rect 3073 -8472 3117 -8438
rect 3251 -8472 3295 -8438
rect 3429 -8472 3473 -8438
rect 3607 -8472 3651 -8438
rect 3785 -8472 3829 -8438
rect 3963 -8472 4007 -8438
rect -5544 -8764 -5500 -8730
rect -5366 -8764 -5322 -8730
rect -5188 -8764 -5144 -8730
rect -5010 -8764 -4966 -8730
rect -4832 -8764 -4788 -8730
rect -4654 -8764 -4610 -8730
rect -4476 -8764 -4432 -8730
rect -4298 -8764 -4254 -8730
rect -4120 -8764 -4076 -8730
rect 6596 -8844 6640 -8810
rect -5544 -8924 -5500 -8890
rect -5366 -8924 -5322 -8890
rect -5188 -8924 -5144 -8890
rect -5010 -8924 -4966 -8890
rect -4832 -8924 -4788 -8890
rect -4654 -8924 -4610 -8890
rect -4476 -8924 -4432 -8890
rect -4298 -8924 -4254 -8890
rect 6774 -8844 6818 -8810
rect 6952 -8844 6996 -8810
rect 7130 -8844 7174 -8810
rect 7308 -8844 7352 -8810
rect 7486 -8844 7530 -8810
rect 7664 -8844 7708 -8810
rect 7842 -8844 7886 -8810
rect 8020 -8844 8064 -8810
rect 8198 -8844 8242 -8810
rect 8376 -8844 8420 -8810
rect 8554 -8844 8598 -8810
rect 8732 -8844 8776 -8810
rect 8910 -8844 8954 -8810
rect 9088 -8844 9132 -8810
rect 9266 -8844 9310 -8810
rect 10856 -8874 10900 -8840
rect -4120 -8924 -4076 -8890
rect -2089 -9082 -2045 -9048
rect -1911 -9082 -1867 -9048
rect -1733 -9082 -1689 -9048
rect -1555 -9082 -1511 -9048
rect -1377 -9082 -1333 -9048
rect -1199 -9082 -1155 -9048
rect -1021 -9082 -977 -9048
rect -843 -9082 -799 -9048
rect -665 -9082 -621 -9048
rect -487 -9082 -443 -9048
rect -309 -9082 -265 -9048
rect -131 -9082 -87 -9048
rect 47 -9082 91 -9048
rect 225 -9082 269 -9048
rect 403 -9082 447 -9048
rect 581 -9082 625 -9048
rect 759 -9082 803 -9048
rect 937 -9082 981 -9048
rect 1115 -9082 1159 -9048
rect 1293 -9082 1337 -9048
rect 1471 -9082 1515 -9048
rect 1649 -9082 1693 -9048
rect 1827 -9082 1871 -9048
rect 2005 -9082 2049 -9048
rect 2183 -9082 2227 -9048
rect 2361 -9082 2405 -9048
rect 2539 -9082 2583 -9048
rect 2717 -9082 2761 -9048
rect 2895 -9082 2939 -9048
rect 3073 -9082 3117 -9048
rect 3251 -9082 3295 -9048
rect 3429 -9082 3473 -9048
rect 3607 -9082 3651 -9048
rect 3785 -9082 3829 -9048
rect 3963 -9082 4007 -9048
rect -5544 -9314 -5500 -9280
rect -5366 -9314 -5322 -9280
rect -5188 -9314 -5144 -9280
rect -5010 -9314 -4966 -9280
rect -4832 -9314 -4788 -9280
rect -4654 -9314 -4610 -9280
rect -4476 -9314 -4432 -9280
rect -4298 -9314 -4254 -9280
rect -4120 -9314 -4076 -9280
rect -5544 -9474 -5500 -9440
rect -5366 -9474 -5322 -9440
rect -5188 -9474 -5144 -9440
rect -5010 -9474 -4966 -9440
rect -4832 -9474 -4788 -9440
rect -4654 -9474 -4610 -9440
rect -4476 -9474 -4432 -9440
rect -4298 -9474 -4254 -9440
rect -4120 -9474 -4076 -9440
rect 11148 -8874 11192 -8840
rect 11440 -8874 11484 -8840
rect 11732 -8874 11776 -8840
rect 12024 -8874 12068 -8840
rect 12316 -8874 12360 -8840
rect 12608 -8874 12652 -8840
rect 6596 -9234 6640 -9200
rect 6774 -9234 6818 -9200
rect 6952 -9234 6996 -9200
rect 7130 -9234 7174 -9200
rect 7308 -9234 7352 -9200
rect 7486 -9234 7530 -9200
rect 7664 -9234 7708 -9200
rect 7842 -9234 7886 -9200
rect 8020 -9234 8064 -9200
rect 8198 -9234 8242 -9200
rect 8376 -9234 8420 -9200
rect 8554 -9234 8598 -9200
rect 8732 -9234 8776 -9200
rect 8910 -9234 8954 -9200
rect 9088 -9234 9132 -9200
rect 9266 -9234 9310 -9200
rect 10856 -9264 10900 -9230
rect 11148 -9264 11192 -9230
rect 11440 -9264 11484 -9230
rect 11732 -9264 11776 -9230
rect 12024 -9264 12068 -9230
rect 12316 -9264 12360 -9230
rect 12608 -9264 12652 -9230
rect -2089 -9472 -2045 -9438
rect -1911 -9472 -1867 -9438
rect -1733 -9472 -1689 -9438
rect -1555 -9472 -1511 -9438
rect -1377 -9472 -1333 -9438
rect -1199 -9472 -1155 -9438
rect -1021 -9472 -977 -9438
rect -843 -9472 -799 -9438
rect -665 -9472 -621 -9438
rect -487 -9472 -443 -9438
rect -309 -9472 -265 -9438
rect -131 -9472 -87 -9438
rect 47 -9472 91 -9438
rect 225 -9472 269 -9438
rect 403 -9472 447 -9438
rect 581 -9472 625 -9438
rect 759 -9472 803 -9438
rect 937 -9472 981 -9438
rect 1115 -9472 1159 -9438
rect 1293 -9472 1337 -9438
rect 1471 -9472 1515 -9438
rect 1649 -9472 1693 -9438
rect 1827 -9472 1871 -9438
rect 2005 -9472 2049 -9438
rect 2183 -9472 2227 -9438
rect 2361 -9472 2405 -9438
rect 2539 -9472 2583 -9438
rect 2717 -9472 2761 -9438
rect 2895 -9472 2939 -9438
rect 3073 -9472 3117 -9438
rect 3251 -9472 3295 -9438
rect 3429 -9472 3473 -9438
rect 3607 -9472 3651 -9438
rect 3785 -9472 3829 -9438
rect 3963 -9472 4007 -9438
rect 10856 -9644 10900 -9610
rect 11148 -9644 11192 -9610
rect 11440 -9644 11484 -9610
rect 11732 -9644 11776 -9610
rect 12024 -9644 12068 -9610
rect 12316 -9644 12360 -9610
rect 12608 -9644 12652 -9610
rect 6596 -9744 6640 -9710
rect 6774 -9744 6818 -9710
rect 6952 -9744 6996 -9710
rect 7130 -9744 7174 -9710
rect 7308 -9744 7352 -9710
rect 7486 -9744 7530 -9710
rect 7664 -9744 7708 -9710
rect 7842 -9744 7886 -9710
rect 8020 -9744 8064 -9710
rect 8198 -9744 8242 -9710
rect 8376 -9744 8420 -9710
rect 8554 -9744 8598 -9710
rect 8732 -9744 8776 -9710
rect 8910 -9744 8954 -9710
rect 9088 -9744 9132 -9710
rect 9266 -9744 9310 -9710
rect -5544 -9864 -5500 -9830
rect -5366 -9864 -5322 -9830
rect -5188 -9864 -5144 -9830
rect -5010 -9864 -4966 -9830
rect -4832 -9864 -4788 -9830
rect -4654 -9864 -4610 -9830
rect -4476 -9864 -4432 -9830
rect -4298 -9864 -4254 -9830
rect -4120 -9864 -4076 -9830
rect -5544 -10024 -5500 -9990
rect -5366 -10024 -5322 -9990
rect -5188 -10024 -5144 -9990
rect -5010 -10024 -4966 -9990
rect -4832 -10024 -4788 -9990
rect -4654 -10024 -4610 -9990
rect -4476 -10024 -4432 -9990
rect -4298 -10024 -4254 -9990
rect -4120 -10024 -4076 -9990
rect -2089 -10082 -2045 -10048
rect -1911 -10082 -1867 -10048
rect -1733 -10082 -1689 -10048
rect -1555 -10082 -1511 -10048
rect -1377 -10082 -1333 -10048
rect -1199 -10082 -1155 -10048
rect -1021 -10082 -977 -10048
rect -843 -10082 -799 -10048
rect -665 -10082 -621 -10048
rect -487 -10082 -443 -10048
rect -309 -10082 -265 -10048
rect -131 -10082 -87 -10048
rect 47 -10082 91 -10048
rect 225 -10082 269 -10048
rect 403 -10082 447 -10048
rect 581 -10082 625 -10048
rect 759 -10082 803 -10048
rect 937 -10082 981 -10048
rect 1115 -10082 1159 -10048
rect 1293 -10082 1337 -10048
rect 1471 -10082 1515 -10048
rect 1649 -10082 1693 -10048
rect 1827 -10082 1871 -10048
rect 2005 -10082 2049 -10048
rect 2183 -10082 2227 -10048
rect 2361 -10082 2405 -10048
rect 2539 -10082 2583 -10048
rect 2717 -10082 2761 -10048
rect 2895 -10082 2939 -10048
rect 3073 -10082 3117 -10048
rect 3251 -10082 3295 -10048
rect 3429 -10082 3473 -10048
rect 3607 -10082 3651 -10048
rect 3785 -10082 3829 -10048
rect 3963 -10082 4007 -10048
rect 10856 -10034 10900 -10000
rect 11148 -10034 11192 -10000
rect 11440 -10034 11484 -10000
rect 11732 -10034 11776 -10000
rect 12024 -10034 12068 -10000
rect 12316 -10034 12360 -10000
rect 12608 -10034 12652 -10000
rect -5544 -10414 -5500 -10380
rect -5366 -10414 -5322 -10380
rect -5188 -10414 -5144 -10380
rect -5010 -10414 -4966 -10380
rect -4832 -10414 -4788 -10380
rect -4654 -10414 -4610 -10380
rect -4476 -10414 -4432 -10380
rect -4298 -10414 -4254 -10380
rect -4120 -10414 -4076 -10380
rect 6596 -10134 6640 -10100
rect 6774 -10134 6818 -10100
rect 6952 -10134 6996 -10100
rect 7130 -10134 7174 -10100
rect 7308 -10134 7352 -10100
rect 7486 -10134 7530 -10100
rect 7664 -10134 7708 -10100
rect 7842 -10134 7886 -10100
rect 8020 -10134 8064 -10100
rect 8198 -10134 8242 -10100
rect 8376 -10134 8420 -10100
rect 8554 -10134 8598 -10100
rect 8732 -10134 8776 -10100
rect 8910 -10134 8954 -10100
rect 9088 -10134 9132 -10100
rect 9266 -10134 9310 -10100
rect -2089 -10472 -2045 -10438
rect -1911 -10472 -1867 -10438
rect -1733 -10472 -1689 -10438
rect -1555 -10472 -1511 -10438
rect -1377 -10472 -1333 -10438
rect -1199 -10472 -1155 -10438
rect -1021 -10472 -977 -10438
rect -843 -10472 -799 -10438
rect -665 -10472 -621 -10438
rect -487 -10472 -443 -10438
rect -309 -10472 -265 -10438
rect -131 -10472 -87 -10438
rect 47 -10472 91 -10438
rect 225 -10472 269 -10438
rect 403 -10472 447 -10438
rect 581 -10472 625 -10438
rect 759 -10472 803 -10438
rect 937 -10472 981 -10438
rect 1115 -10472 1159 -10438
rect 1293 -10472 1337 -10438
rect 1471 -10472 1515 -10438
rect 1649 -10472 1693 -10438
rect 1827 -10472 1871 -10438
rect 2005 -10472 2049 -10438
rect 2183 -10472 2227 -10438
rect 2361 -10472 2405 -10438
rect 2539 -10472 2583 -10438
rect 2717 -10472 2761 -10438
rect 2895 -10472 2939 -10438
rect 3073 -10472 3117 -10438
rect 3251 -10472 3295 -10438
rect 3429 -10472 3473 -10438
rect 3607 -10472 3651 -10438
rect 3785 -10472 3829 -10438
rect 3963 -10472 4007 -10438
rect 10856 -10414 10900 -10380
rect 11148 -10414 11192 -10380
rect 11440 -10414 11484 -10380
rect 11732 -10414 11776 -10380
rect 12024 -10414 12068 -10380
rect 12316 -10414 12360 -10380
rect 12608 -10414 12652 -10380
rect -5544 -10574 -5500 -10540
rect -5366 -10574 -5322 -10540
rect -5188 -10574 -5144 -10540
rect -5010 -10574 -4966 -10540
rect -4832 -10574 -4788 -10540
rect -4654 -10574 -4610 -10540
rect -4476 -10574 -4432 -10540
rect -4298 -10574 -4254 -10540
rect -4120 -10574 -4076 -10540
rect 6596 -10644 6640 -10610
rect 6774 -10644 6818 -10610
rect 6952 -10644 6996 -10610
rect 7130 -10644 7174 -10610
rect 7308 -10644 7352 -10610
rect 7486 -10644 7530 -10610
rect 7664 -10644 7708 -10610
rect 7842 -10644 7886 -10610
rect 8020 -10644 8064 -10610
rect 8198 -10644 8242 -10610
rect 8376 -10644 8420 -10610
rect 8554 -10644 8598 -10610
rect 8732 -10644 8776 -10610
rect 8910 -10644 8954 -10610
rect 9088 -10644 9132 -10610
rect 9266 -10644 9310 -10610
rect -5544 -10964 -5500 -10930
rect -5366 -10964 -5322 -10930
rect -5188 -10964 -5144 -10930
rect -5010 -10964 -4966 -10930
rect -4832 -10964 -4788 -10930
rect -4654 -10964 -4610 -10930
rect -4476 -10964 -4432 -10930
rect -4298 -10964 -4254 -10930
rect -4120 -10964 -4076 -10930
rect 10856 -10804 10900 -10770
rect 11148 -10804 11192 -10770
rect 11440 -10804 11484 -10770
rect 11732 -10804 11776 -10770
rect 12024 -10804 12068 -10770
rect 12316 -10804 12360 -10770
rect 12608 -10804 12652 -10770
rect -5544 -11124 -5500 -11090
rect -5366 -11124 -5322 -11090
rect -5188 -11124 -5144 -11090
rect -5010 -11124 -4966 -11090
rect -4832 -11124 -4788 -11090
rect -4654 -11124 -4610 -11090
rect -4476 -11124 -4432 -11090
rect -4298 -11124 -4254 -11090
rect -4120 -11124 -4076 -11090
rect -2089 -11082 -2045 -11048
rect -1911 -11082 -1867 -11048
rect -1733 -11082 -1689 -11048
rect -1555 -11082 -1511 -11048
rect -1377 -11082 -1333 -11048
rect -1199 -11082 -1155 -11048
rect -1021 -11082 -977 -11048
rect -843 -11082 -799 -11048
rect -665 -11082 -621 -11048
rect -487 -11082 -443 -11048
rect -309 -11082 -265 -11048
rect -131 -11082 -87 -11048
rect 47 -11082 91 -11048
rect 225 -11082 269 -11048
rect 403 -11082 447 -11048
rect 581 -11082 625 -11048
rect 759 -11082 803 -11048
rect 937 -11082 981 -11048
rect 1115 -11082 1159 -11048
rect 1293 -11082 1337 -11048
rect 1471 -11082 1515 -11048
rect 1649 -11082 1693 -11048
rect 1827 -11082 1871 -11048
rect 2005 -11082 2049 -11048
rect 2183 -11082 2227 -11048
rect 2361 -11082 2405 -11048
rect 2539 -11082 2583 -11048
rect 2717 -11082 2761 -11048
rect 2895 -11082 2939 -11048
rect 3073 -11082 3117 -11048
rect 3251 -11082 3295 -11048
rect 3429 -11082 3473 -11048
rect 3607 -11082 3651 -11048
rect 3785 -11082 3829 -11048
rect 3963 -11082 4007 -11048
rect 6596 -11034 6640 -11000
rect 6774 -11034 6818 -11000
rect 6952 -11034 6996 -11000
rect 7130 -11034 7174 -11000
rect 7308 -11034 7352 -11000
rect 7486 -11034 7530 -11000
rect 7664 -11034 7708 -11000
rect 7842 -11034 7886 -11000
rect 8020 -11034 8064 -11000
rect 8198 -11034 8242 -11000
rect 8376 -11034 8420 -11000
rect 8554 -11034 8598 -11000
rect 8732 -11034 8776 -11000
rect 8910 -11034 8954 -11000
rect 9088 -11034 9132 -11000
rect 9266 -11034 9310 -11000
rect -5544 -11514 -5500 -11480
rect -5366 -11514 -5322 -11480
rect -5188 -11514 -5144 -11480
rect -5010 -11514 -4966 -11480
rect -4832 -11514 -4788 -11480
rect -4654 -11514 -4610 -11480
rect -4476 -11514 -4432 -11480
rect -4298 -11514 -4254 -11480
rect 10856 -11184 10900 -11150
rect 11148 -11184 11192 -11150
rect 11440 -11184 11484 -11150
rect 11732 -11184 11776 -11150
rect 12024 -11184 12068 -11150
rect 12316 -11184 12360 -11150
rect 12608 -11184 12652 -11150
rect -2089 -11472 -2045 -11438
rect -4120 -11514 -4076 -11480
rect -1911 -11472 -1867 -11438
rect -1733 -11472 -1689 -11438
rect -1555 -11472 -1511 -11438
rect -1377 -11472 -1333 -11438
rect -1199 -11472 -1155 -11438
rect -1021 -11472 -977 -11438
rect -843 -11472 -799 -11438
rect -665 -11472 -621 -11438
rect -487 -11472 -443 -11438
rect -309 -11472 -265 -11438
rect -131 -11472 -87 -11438
rect 47 -11472 91 -11438
rect 225 -11472 269 -11438
rect 403 -11472 447 -11438
rect 581 -11472 625 -11438
rect 759 -11472 803 -11438
rect 937 -11472 981 -11438
rect 1115 -11472 1159 -11438
rect 1293 -11472 1337 -11438
rect 1471 -11472 1515 -11438
rect 1649 -11472 1693 -11438
rect 1827 -11472 1871 -11438
rect 2005 -11472 2049 -11438
rect 2183 -11472 2227 -11438
rect 2361 -11472 2405 -11438
rect 2539 -11472 2583 -11438
rect 2717 -11472 2761 -11438
rect 2895 -11472 2939 -11438
rect 3073 -11472 3117 -11438
rect 3251 -11472 3295 -11438
rect 3429 -11472 3473 -11438
rect 3607 -11472 3651 -11438
rect 3785 -11472 3829 -11438
rect 3963 -11472 4007 -11438
rect 6596 -11544 6640 -11510
rect 6774 -11544 6818 -11510
rect 6952 -11544 6996 -11510
rect 7130 -11544 7174 -11510
rect 7308 -11544 7352 -11510
rect 7486 -11544 7530 -11510
rect 7664 -11544 7708 -11510
rect 7842 -11544 7886 -11510
rect 8020 -11544 8064 -11510
rect 8198 -11544 8242 -11510
rect 8376 -11544 8420 -11510
rect 8554 -11544 8598 -11510
rect 8732 -11544 8776 -11510
rect 8910 -11544 8954 -11510
rect 9088 -11544 9132 -11510
rect 9266 -11544 9310 -11510
rect 10856 -11574 10900 -11540
rect -5544 -11674 -5500 -11640
rect -5366 -11674 -5322 -11640
rect -5188 -11674 -5144 -11640
rect -5010 -11674 -4966 -11640
rect -4832 -11674 -4788 -11640
rect -4654 -11674 -4610 -11640
rect -4476 -11674 -4432 -11640
rect -4298 -11674 -4254 -11640
rect -4120 -11674 -4076 -11640
rect 11148 -11574 11192 -11540
rect 11440 -11574 11484 -11540
rect 11732 -11574 11776 -11540
rect 12024 -11574 12068 -11540
rect 12316 -11574 12360 -11540
rect 12608 -11574 12652 -11540
rect 6596 -11934 6640 -11900
rect 6774 -11934 6818 -11900
rect 6952 -11934 6996 -11900
rect 7130 -11934 7174 -11900
rect 7308 -11934 7352 -11900
rect 7486 -11934 7530 -11900
rect 7664 -11934 7708 -11900
rect 7842 -11934 7886 -11900
rect 8020 -11934 8064 -11900
rect 8198 -11934 8242 -11900
rect 8376 -11934 8420 -11900
rect 8554 -11934 8598 -11900
rect 8732 -11934 8776 -11900
rect 8910 -11934 8954 -11900
rect 9088 -11934 9132 -11900
rect 9266 -11934 9310 -11900
rect -5544 -12064 -5500 -12030
rect -5366 -12064 -5322 -12030
rect -5188 -12064 -5144 -12030
rect -5010 -12064 -4966 -12030
rect -4832 -12064 -4788 -12030
rect -4654 -12064 -4610 -12030
rect -4476 -12064 -4432 -12030
rect -4298 -12064 -4254 -12030
rect -4120 -12064 -4076 -12030
rect -2089 -12082 -2045 -12048
rect -1911 -12082 -1867 -12048
rect -1733 -12082 -1689 -12048
rect -1555 -12082 -1511 -12048
rect -1377 -12082 -1333 -12048
rect -1199 -12082 -1155 -12048
rect -1021 -12082 -977 -12048
rect -843 -12082 -799 -12048
rect -665 -12082 -621 -12048
rect -487 -12082 -443 -12048
rect -309 -12082 -265 -12048
rect -131 -12082 -87 -12048
rect 47 -12082 91 -12048
rect 225 -12082 269 -12048
rect 403 -12082 447 -12048
rect 581 -12082 625 -12048
rect 759 -12082 803 -12048
rect 937 -12082 981 -12048
rect 1115 -12082 1159 -12048
rect 1293 -12082 1337 -12048
rect 1471 -12082 1515 -12048
rect 1649 -12082 1693 -12048
rect 1827 -12082 1871 -12048
rect 2005 -12082 2049 -12048
rect 2183 -12082 2227 -12048
rect 2361 -12082 2405 -12048
rect 2539 -12082 2583 -12048
rect 2717 -12082 2761 -12048
rect 2895 -12082 2939 -12048
rect 3073 -12082 3117 -12048
rect 3251 -12082 3295 -12048
rect 3429 -12082 3473 -12048
rect 3607 -12082 3651 -12048
rect 3785 -12082 3829 -12048
rect 3963 -12082 4007 -12048
rect -2089 -12472 -2045 -12438
rect -1911 -12472 -1867 -12438
rect -1733 -12472 -1689 -12438
rect -1555 -12472 -1511 -12438
rect -1377 -12472 -1333 -12438
rect -1199 -12472 -1155 -12438
rect -1021 -12472 -977 -12438
rect -843 -12472 -799 -12438
rect -665 -12472 -621 -12438
rect -487 -12472 -443 -12438
rect -309 -12472 -265 -12438
rect -131 -12472 -87 -12438
rect 47 -12472 91 -12438
rect 225 -12472 269 -12438
rect 403 -12472 447 -12438
rect 581 -12472 625 -12438
rect 759 -12472 803 -12438
rect 937 -12472 981 -12438
rect 1115 -12472 1159 -12438
rect 1293 -12472 1337 -12438
rect 1471 -12472 1515 -12438
rect 1649 -12472 1693 -12438
rect 1827 -12472 1871 -12438
rect 2005 -12472 2049 -12438
rect 2183 -12472 2227 -12438
rect 2361 -12472 2405 -12438
rect 2539 -12472 2583 -12438
rect 2717 -12472 2761 -12438
rect 2895 -12472 2939 -12438
rect 3073 -12472 3117 -12438
rect 3251 -12472 3295 -12438
rect 3429 -12472 3473 -12438
rect 3607 -12472 3651 -12438
rect 3785 -12472 3829 -12438
rect 3963 -12472 4007 -12438
rect -5867 -12662 -5833 -12628
rect -5617 -12662 -5583 -12628
rect -5367 -12662 -5333 -12628
rect -5117 -12662 -5083 -12628
rect -4867 -12662 -4833 -12628
rect -4617 -12662 -4583 -12628
rect -4367 -12662 -4333 -12628
rect -4117 -12662 -4083 -12628
rect -5867 -13012 -5833 -12978
rect -5617 -13012 -5583 -12978
rect -5367 -13012 -5333 -12978
rect -5117 -13012 -5083 -12978
rect -4867 -13012 -4833 -12978
rect -4617 -13012 -4583 -12978
rect -4367 -13012 -4333 -12978
rect -4117 -13012 -4083 -12978
rect -2089 -13082 -2045 -13048
rect -1911 -13082 -1867 -13048
rect -1733 -13082 -1689 -13048
rect -1555 -13082 -1511 -13048
rect -1377 -13082 -1333 -13048
rect -1199 -13082 -1155 -13048
rect -1021 -13082 -977 -13048
rect -843 -13082 -799 -13048
rect -665 -13082 -621 -13048
rect -487 -13082 -443 -13048
rect -309 -13082 -265 -13048
rect -131 -13082 -87 -13048
rect 47 -13082 91 -13048
rect 225 -13082 269 -13048
rect 403 -13082 447 -13048
rect 581 -13082 625 -13048
rect 759 -13082 803 -13048
rect 937 -13082 981 -13048
rect 1115 -13082 1159 -13048
rect 1293 -13082 1337 -13048
rect 1471 -13082 1515 -13048
rect 1649 -13082 1693 -13048
rect 1827 -13082 1871 -13048
rect 2005 -13082 2049 -13048
rect 2183 -13082 2227 -13048
rect 2361 -13082 2405 -13048
rect 2539 -13082 2583 -13048
rect 2717 -13082 2761 -13048
rect 2895 -13082 2939 -13048
rect 3073 -13082 3117 -13048
rect 3251 -13082 3295 -13048
rect 3429 -13082 3473 -13048
rect 3607 -13082 3651 -13048
rect 3785 -13082 3829 -13048
rect 3963 -13082 4007 -13048
rect -5867 -13342 -5833 -13308
rect -5617 -13342 -5583 -13308
rect -5367 -13342 -5333 -13308
rect -5117 -13342 -5083 -13308
rect -4867 -13342 -4833 -13308
rect -4617 -13342 -4583 -13308
rect -4367 -13342 -4333 -13308
rect -4117 -13342 -4083 -13308
rect -2089 -13472 -2045 -13438
rect -1911 -13472 -1867 -13438
rect -1733 -13472 -1689 -13438
rect -1555 -13472 -1511 -13438
rect -1377 -13472 -1333 -13438
rect -1199 -13472 -1155 -13438
rect -1021 -13472 -977 -13438
rect -843 -13472 -799 -13438
rect -665 -13472 -621 -13438
rect -487 -13472 -443 -13438
rect -309 -13472 -265 -13438
rect -131 -13472 -87 -13438
rect 47 -13472 91 -13438
rect 225 -13472 269 -13438
rect 403 -13472 447 -13438
rect 581 -13472 625 -13438
rect 759 -13472 803 -13438
rect 937 -13472 981 -13438
rect 1115 -13472 1159 -13438
rect 1293 -13472 1337 -13438
rect 1471 -13472 1515 -13438
rect 1649 -13472 1693 -13438
rect 1827 -13472 1871 -13438
rect 2005 -13472 2049 -13438
rect 2183 -13472 2227 -13438
rect 2361 -13472 2405 -13438
rect 2539 -13472 2583 -13438
rect 2717 -13472 2761 -13438
rect 2895 -13472 2939 -13438
rect 3073 -13472 3117 -13438
rect 3251 -13472 3295 -13438
rect 3429 -13472 3473 -13438
rect 3607 -13472 3651 -13438
rect 3785 -13472 3829 -13438
rect 3963 -13472 4007 -13438
rect -5867 -13692 -5833 -13658
rect -5617 -13692 -5583 -13658
rect -5367 -13692 -5333 -13658
rect -5117 -13692 -5083 -13658
rect -4867 -13692 -4833 -13658
rect -4617 -13692 -4583 -13658
rect -4367 -13692 -4333 -13658
rect -4117 -13692 -4083 -13658
rect -2089 -14082 -2045 -14048
rect -1911 -14082 -1867 -14048
rect -1733 -14082 -1689 -14048
rect -1555 -14082 -1511 -14048
rect -1377 -14082 -1333 -14048
rect -1199 -14082 -1155 -14048
rect -1021 -14082 -977 -14048
rect -843 -14082 -799 -14048
rect -665 -14082 -621 -14048
rect -487 -14082 -443 -14048
rect -309 -14082 -265 -14048
rect -131 -14082 -87 -14048
rect 47 -14082 91 -14048
rect 225 -14082 269 -14048
rect 403 -14082 447 -14048
rect 581 -14082 625 -14048
rect 759 -14082 803 -14048
rect 937 -14082 981 -14048
rect 1115 -14082 1159 -14048
rect 1293 -14082 1337 -14048
rect 1471 -14082 1515 -14048
rect 1649 -14082 1693 -14048
rect 1827 -14082 1871 -14048
rect 2005 -14082 2049 -14048
rect 2183 -14082 2227 -14048
rect 2361 -14082 2405 -14048
rect 2539 -14082 2583 -14048
rect 2717 -14082 2761 -14048
rect 2895 -14082 2939 -14048
rect 3073 -14082 3117 -14048
rect 3251 -14082 3295 -14048
rect 3429 -14082 3473 -14048
rect 3607 -14082 3651 -14048
rect 3785 -14082 3829 -14048
rect 3963 -14082 4007 -14048
rect 5661 -14082 5705 -14048
rect 5839 -14082 5883 -14048
rect 6017 -14082 6061 -14048
rect 6195 -14082 6239 -14048
rect 6373 -14082 6417 -14048
rect 6551 -14082 6595 -14048
rect 6729 -14082 6773 -14048
rect 6907 -14082 6951 -14048
rect 7085 -14082 7129 -14048
rect 7263 -14082 7307 -14048
rect 7441 -14082 7485 -14048
rect 7619 -14082 7663 -14048
rect 7797 -14082 7841 -14048
rect 7975 -14082 8019 -14048
rect 8153 -14082 8197 -14048
rect 8331 -14082 8375 -14048
rect 8509 -14082 8553 -14048
rect 8687 -14082 8731 -14048
rect 8865 -14082 8909 -14048
rect 9043 -14082 9087 -14048
rect 9221 -14082 9265 -14048
rect 9399 -14082 9443 -14048
rect 9577 -14082 9621 -14048
rect 9755 -14082 9799 -14048
rect 9933 -14082 9977 -14048
rect 10111 -14082 10155 -14048
rect 10289 -14082 10333 -14048
rect 10467 -14082 10511 -14048
rect 10645 -14082 10689 -14048
rect 10823 -14082 10867 -14048
rect 11001 -14082 11045 -14048
rect 11179 -14082 11223 -14048
rect 11357 -14082 11401 -14048
rect 11535 -14082 11579 -14048
rect 11713 -14082 11757 -14048
rect 11891 -14082 11935 -14048
rect 12069 -14082 12113 -14048
rect 12247 -14082 12291 -14048
rect 12425 -14082 12469 -14048
rect 12603 -14082 12647 -14048
rect -5944 -14344 -5900 -14310
rect -5766 -14344 -5722 -14310
rect -5588 -14344 -5544 -14310
rect -5410 -14344 -5366 -14310
rect -5232 -14344 -5188 -14310
rect -5054 -14344 -5010 -14310
rect -4876 -14344 -4832 -14310
rect -4698 -14344 -4654 -14310
rect -4520 -14344 -4476 -14310
rect -4342 -14344 -4298 -14310
rect -4164 -14344 -4120 -14310
rect -2089 -14472 -2045 -14438
rect -1911 -14472 -1867 -14438
rect -1733 -14472 -1689 -14438
rect -1555 -14472 -1511 -14438
rect -1377 -14472 -1333 -14438
rect -1199 -14472 -1155 -14438
rect -1021 -14472 -977 -14438
rect -843 -14472 -799 -14438
rect -665 -14472 -621 -14438
rect -487 -14472 -443 -14438
rect -309 -14472 -265 -14438
rect -131 -14472 -87 -14438
rect 47 -14472 91 -14438
rect 225 -14472 269 -14438
rect 403 -14472 447 -14438
rect 581 -14472 625 -14438
rect 759 -14472 803 -14438
rect 937 -14472 981 -14438
rect 1115 -14472 1159 -14438
rect 1293 -14472 1337 -14438
rect 1471 -14472 1515 -14438
rect 1649 -14472 1693 -14438
rect 1827 -14472 1871 -14438
rect 2005 -14472 2049 -14438
rect 2183 -14472 2227 -14438
rect 2361 -14472 2405 -14438
rect 2539 -14472 2583 -14438
rect 2717 -14472 2761 -14438
rect 2895 -14472 2939 -14438
rect 3073 -14472 3117 -14438
rect 3251 -14472 3295 -14438
rect 3429 -14472 3473 -14438
rect 3607 -14472 3651 -14438
rect 3785 -14472 3829 -14438
rect 3963 -14472 4007 -14438
rect 5661 -14472 5705 -14438
rect 5839 -14472 5883 -14438
rect 6017 -14472 6061 -14438
rect 6195 -14472 6239 -14438
rect 6373 -14472 6417 -14438
rect 6551 -14472 6595 -14438
rect 6729 -14472 6773 -14438
rect 6907 -14472 6951 -14438
rect 7085 -14472 7129 -14438
rect 7263 -14472 7307 -14438
rect 7441 -14472 7485 -14438
rect 7619 -14472 7663 -14438
rect 7797 -14472 7841 -14438
rect 7975 -14472 8019 -14438
rect 8153 -14472 8197 -14438
rect 8331 -14472 8375 -14438
rect 8509 -14472 8553 -14438
rect 8687 -14472 8731 -14438
rect 8865 -14472 8909 -14438
rect 9043 -14472 9087 -14438
rect 9221 -14472 9265 -14438
rect 9399 -14472 9443 -14438
rect 9577 -14472 9621 -14438
rect 9755 -14472 9799 -14438
rect 9933 -14472 9977 -14438
rect 10111 -14472 10155 -14438
rect 10289 -14472 10333 -14438
rect 10467 -14472 10511 -14438
rect 10645 -14472 10689 -14438
rect 10823 -14472 10867 -14438
rect 11001 -14472 11045 -14438
rect 11179 -14472 11223 -14438
rect 11357 -14472 11401 -14438
rect 11535 -14472 11579 -14438
rect 11713 -14472 11757 -14438
rect 11891 -14472 11935 -14438
rect 12069 -14472 12113 -14438
rect 12247 -14472 12291 -14438
rect 12425 -14472 12469 -14438
rect 12603 -14472 12647 -14438
rect -5944 -14734 -5900 -14700
rect -5766 -14734 -5722 -14700
rect -5588 -14734 -5544 -14700
rect -5410 -14734 -5366 -14700
rect -5232 -14734 -5188 -14700
rect -5054 -14734 -5010 -14700
rect -4876 -14734 -4832 -14700
rect -4698 -14734 -4654 -14700
rect -4520 -14734 -4476 -14700
rect -4342 -14734 -4298 -14700
rect -4164 -14734 -4120 -14700
rect -5944 -15044 -5900 -15010
rect -5766 -15044 -5722 -15010
rect -5588 -15044 -5544 -15010
rect -5410 -15044 -5366 -15010
rect -5232 -15044 -5188 -15010
rect -5054 -15044 -5010 -15010
rect -4876 -15044 -4832 -15010
rect -4698 -15044 -4654 -15010
rect -4520 -15044 -4476 -15010
rect -4342 -15044 -4298 -15010
rect -4164 -15044 -4120 -15010
rect -2089 -15082 -2045 -15048
rect -1911 -15082 -1867 -15048
rect -1733 -15082 -1689 -15048
rect -1555 -15082 -1511 -15048
rect -1377 -15082 -1333 -15048
rect -1199 -15082 -1155 -15048
rect -1021 -15082 -977 -15048
rect -843 -15082 -799 -15048
rect -665 -15082 -621 -15048
rect -487 -15082 -443 -15048
rect -309 -15082 -265 -15048
rect -131 -15082 -87 -15048
rect 47 -15082 91 -15048
rect 225 -15082 269 -15048
rect 403 -15082 447 -15048
rect 581 -15082 625 -15048
rect 759 -15082 803 -15048
rect 937 -15082 981 -15048
rect 1115 -15082 1159 -15048
rect 1293 -15082 1337 -15048
rect 1471 -15082 1515 -15048
rect 1649 -15082 1693 -15048
rect 1827 -15082 1871 -15048
rect 2005 -15082 2049 -15048
rect 2183 -15082 2227 -15048
rect 2361 -15082 2405 -15048
rect 2539 -15082 2583 -15048
rect 2717 -15082 2761 -15048
rect 2895 -15082 2939 -15048
rect 3073 -15082 3117 -15048
rect 3251 -15082 3295 -15048
rect 3429 -15082 3473 -15048
rect 3607 -15082 3651 -15048
rect 3785 -15082 3829 -15048
rect 3963 -15082 4007 -15048
rect 5661 -15082 5705 -15048
rect 5839 -15082 5883 -15048
rect 6017 -15082 6061 -15048
rect 6195 -15082 6239 -15048
rect 6373 -15082 6417 -15048
rect 6551 -15082 6595 -15048
rect 6729 -15082 6773 -15048
rect 6907 -15082 6951 -15048
rect 7085 -15082 7129 -15048
rect 7263 -15082 7307 -15048
rect 7441 -15082 7485 -15048
rect 7619 -15082 7663 -15048
rect 7797 -15082 7841 -15048
rect 7975 -15082 8019 -15048
rect 8153 -15082 8197 -15048
rect 8331 -15082 8375 -15048
rect 8509 -15082 8553 -15048
rect 8687 -15082 8731 -15048
rect 8865 -15082 8909 -15048
rect 9043 -15082 9087 -15048
rect 9221 -15082 9265 -15048
rect 9399 -15082 9443 -15048
rect 9577 -15082 9621 -15048
rect 9755 -15082 9799 -15048
rect 9933 -15082 9977 -15048
rect 10111 -15082 10155 -15048
rect 10289 -15082 10333 -15048
rect 10467 -15082 10511 -15048
rect 10645 -15082 10689 -15048
rect 10823 -15082 10867 -15048
rect 11001 -15082 11045 -15048
rect 11179 -15082 11223 -15048
rect 11357 -15082 11401 -15048
rect 11535 -15082 11579 -15048
rect 11713 -15082 11757 -15048
rect 11891 -15082 11935 -15048
rect 12069 -15082 12113 -15048
rect 12247 -15082 12291 -15048
rect 12425 -15082 12469 -15048
rect 12603 -15082 12647 -15048
rect -5944 -15434 -5900 -15400
rect -5766 -15434 -5722 -15400
rect -5588 -15434 -5544 -15400
rect -5410 -15434 -5366 -15400
rect -5232 -15434 -5188 -15400
rect -5054 -15434 -5010 -15400
rect -4876 -15434 -4832 -15400
rect -4698 -15434 -4654 -15400
rect -4520 -15434 -4476 -15400
rect -4342 -15434 -4298 -15400
rect -4164 -15434 -4120 -15400
rect -2089 -15472 -2045 -15438
rect -1911 -15472 -1867 -15438
rect -1733 -15472 -1689 -15438
rect -1555 -15472 -1511 -15438
rect -1377 -15472 -1333 -15438
rect -1199 -15472 -1155 -15438
rect -1021 -15472 -977 -15438
rect -843 -15472 -799 -15438
rect -665 -15472 -621 -15438
rect -487 -15472 -443 -15438
rect -309 -15472 -265 -15438
rect -131 -15472 -87 -15438
rect 47 -15472 91 -15438
rect 225 -15472 269 -15438
rect 403 -15472 447 -15438
rect 581 -15472 625 -15438
rect 759 -15472 803 -15438
rect 937 -15472 981 -15438
rect 1115 -15472 1159 -15438
rect 1293 -15472 1337 -15438
rect 1471 -15472 1515 -15438
rect 1649 -15472 1693 -15438
rect 1827 -15472 1871 -15438
rect 2005 -15472 2049 -15438
rect 2183 -15472 2227 -15438
rect 2361 -15472 2405 -15438
rect 2539 -15472 2583 -15438
rect 2717 -15472 2761 -15438
rect 2895 -15472 2939 -15438
rect 3073 -15472 3117 -15438
rect 3251 -15472 3295 -15438
rect 3429 -15472 3473 -15438
rect 3607 -15472 3651 -15438
rect 3785 -15472 3829 -15438
rect 3963 -15472 4007 -15438
rect 5661 -15472 5705 -15438
rect 5839 -15472 5883 -15438
rect 6017 -15472 6061 -15438
rect 6195 -15472 6239 -15438
rect 6373 -15472 6417 -15438
rect 6551 -15472 6595 -15438
rect 6729 -15472 6773 -15438
rect 6907 -15472 6951 -15438
rect 7085 -15472 7129 -15438
rect 7263 -15472 7307 -15438
rect 7441 -15472 7485 -15438
rect 7619 -15472 7663 -15438
rect 7797 -15472 7841 -15438
rect 7975 -15472 8019 -15438
rect 8153 -15472 8197 -15438
rect 8331 -15472 8375 -15438
rect 8509 -15472 8553 -15438
rect 8687 -15472 8731 -15438
rect 8865 -15472 8909 -15438
rect 9043 -15472 9087 -15438
rect 9221 -15472 9265 -15438
rect 9399 -15472 9443 -15438
rect 9577 -15472 9621 -15438
rect 9755 -15472 9799 -15438
rect 9933 -15472 9977 -15438
rect 10111 -15472 10155 -15438
rect 10289 -15472 10333 -15438
rect 10467 -15472 10511 -15438
rect 10645 -15472 10689 -15438
rect 10823 -15472 10867 -15438
rect 11001 -15472 11045 -15438
rect 11179 -15472 11223 -15438
rect 11357 -15472 11401 -15438
rect 11535 -15472 11579 -15438
rect 11713 -15472 11757 -15438
rect 11891 -15472 11935 -15438
rect 12069 -15472 12113 -15438
rect 12247 -15472 12291 -15438
rect 12425 -15472 12469 -15438
rect 12603 -15472 12647 -15438
rect -5944 -15744 -5900 -15710
rect -5766 -15744 -5722 -15710
rect -5588 -15744 -5544 -15710
rect -5410 -15744 -5366 -15710
rect -5232 -15744 -5188 -15710
rect -5054 -15744 -5010 -15710
rect -4876 -15744 -4832 -15710
rect -4698 -15744 -4654 -15710
rect -4520 -15744 -4476 -15710
rect -4342 -15744 -4298 -15710
rect -4164 -15744 -4120 -15710
rect -5944 -16134 -5900 -16100
rect -5766 -16134 -5722 -16100
rect -5588 -16134 -5544 -16100
rect -5410 -16134 -5366 -16100
rect -5232 -16134 -5188 -16100
rect -5054 -16134 -5010 -16100
rect -4876 -16134 -4832 -16100
rect -4698 -16134 -4654 -16100
rect -4520 -16134 -4476 -16100
rect -4342 -16134 -4298 -16100
rect -4164 -16134 -4120 -16100
rect -2089 -16082 -2045 -16048
rect -1911 -16082 -1867 -16048
rect -1733 -16082 -1689 -16048
rect -1555 -16082 -1511 -16048
rect -1377 -16082 -1333 -16048
rect -1199 -16082 -1155 -16048
rect -1021 -16082 -977 -16048
rect -843 -16082 -799 -16048
rect -665 -16082 -621 -16048
rect -487 -16082 -443 -16048
rect -309 -16082 -265 -16048
rect -131 -16082 -87 -16048
rect 47 -16082 91 -16048
rect 225 -16082 269 -16048
rect 403 -16082 447 -16048
rect 581 -16082 625 -16048
rect 759 -16082 803 -16048
rect 937 -16082 981 -16048
rect 1115 -16082 1159 -16048
rect 1293 -16082 1337 -16048
rect 1471 -16082 1515 -16048
rect 1649 -16082 1693 -16048
rect 1827 -16082 1871 -16048
rect 2005 -16082 2049 -16048
rect 2183 -16082 2227 -16048
rect 2361 -16082 2405 -16048
rect 2539 -16082 2583 -16048
rect 2717 -16082 2761 -16048
rect 2895 -16082 2939 -16048
rect 3073 -16082 3117 -16048
rect 3251 -16082 3295 -16048
rect 3429 -16082 3473 -16048
rect 3607 -16082 3651 -16048
rect 3785 -16082 3829 -16048
rect 3963 -16082 4007 -16048
rect 5661 -16082 5705 -16048
rect 5839 -16082 5883 -16048
rect 6017 -16082 6061 -16048
rect 6195 -16082 6239 -16048
rect 6373 -16082 6417 -16048
rect 6551 -16082 6595 -16048
rect 6729 -16082 6773 -16048
rect 6907 -16082 6951 -16048
rect 7085 -16082 7129 -16048
rect 7263 -16082 7307 -16048
rect 7441 -16082 7485 -16048
rect 7619 -16082 7663 -16048
rect 7797 -16082 7841 -16048
rect 7975 -16082 8019 -16048
rect 8153 -16082 8197 -16048
rect 8331 -16082 8375 -16048
rect 8509 -16082 8553 -16048
rect 8687 -16082 8731 -16048
rect 8865 -16082 8909 -16048
rect 9043 -16082 9087 -16048
rect 9221 -16082 9265 -16048
rect 9399 -16082 9443 -16048
rect 9577 -16082 9621 -16048
rect 9755 -16082 9799 -16048
rect 9933 -16082 9977 -16048
rect 10111 -16082 10155 -16048
rect 10289 -16082 10333 -16048
rect 10467 -16082 10511 -16048
rect 10645 -16082 10689 -16048
rect 10823 -16082 10867 -16048
rect 11001 -16082 11045 -16048
rect 11179 -16082 11223 -16048
rect 11357 -16082 11401 -16048
rect 11535 -16082 11579 -16048
rect 11713 -16082 11757 -16048
rect 11891 -16082 11935 -16048
rect 12069 -16082 12113 -16048
rect 12247 -16082 12291 -16048
rect 12425 -16082 12469 -16048
rect 12603 -16082 12647 -16048
rect -5944 -16444 -5900 -16410
rect -5766 -16444 -5722 -16410
rect -5588 -16444 -5544 -16410
rect -5410 -16444 -5366 -16410
rect -5232 -16444 -5188 -16410
rect -5054 -16444 -5010 -16410
rect -4876 -16444 -4832 -16410
rect -4698 -16444 -4654 -16410
rect -4520 -16444 -4476 -16410
rect -4342 -16444 -4298 -16410
rect -4164 -16444 -4120 -16410
rect -2089 -16472 -2045 -16438
rect -1911 -16472 -1867 -16438
rect -1733 -16472 -1689 -16438
rect -1555 -16472 -1511 -16438
rect -1377 -16472 -1333 -16438
rect -1199 -16472 -1155 -16438
rect -1021 -16472 -977 -16438
rect -843 -16472 -799 -16438
rect -665 -16472 -621 -16438
rect -487 -16472 -443 -16438
rect -309 -16472 -265 -16438
rect -131 -16472 -87 -16438
rect 47 -16472 91 -16438
rect 225 -16472 269 -16438
rect 403 -16472 447 -16438
rect 581 -16472 625 -16438
rect 759 -16472 803 -16438
rect 937 -16472 981 -16438
rect 1115 -16472 1159 -16438
rect 1293 -16472 1337 -16438
rect 1471 -16472 1515 -16438
rect 1649 -16472 1693 -16438
rect 1827 -16472 1871 -16438
rect 2005 -16472 2049 -16438
rect 2183 -16472 2227 -16438
rect 2361 -16472 2405 -16438
rect 2539 -16472 2583 -16438
rect 2717 -16472 2761 -16438
rect 2895 -16472 2939 -16438
rect 3073 -16472 3117 -16438
rect 3251 -16472 3295 -16438
rect 3429 -16472 3473 -16438
rect 3607 -16472 3651 -16438
rect 3785 -16472 3829 -16438
rect 3963 -16472 4007 -16438
rect 5661 -16472 5705 -16438
rect 5839 -16472 5883 -16438
rect 6017 -16472 6061 -16438
rect 6195 -16472 6239 -16438
rect 6373 -16472 6417 -16438
rect 6551 -16472 6595 -16438
rect 6729 -16472 6773 -16438
rect 6907 -16472 6951 -16438
rect 7085 -16472 7129 -16438
rect 7263 -16472 7307 -16438
rect 7441 -16472 7485 -16438
rect 7619 -16472 7663 -16438
rect 7797 -16472 7841 -16438
rect 7975 -16472 8019 -16438
rect 8153 -16472 8197 -16438
rect 8331 -16472 8375 -16438
rect 8509 -16472 8553 -16438
rect 8687 -16472 8731 -16438
rect 8865 -16472 8909 -16438
rect 9043 -16472 9087 -16438
rect 9221 -16472 9265 -16438
rect 9399 -16472 9443 -16438
rect 9577 -16472 9621 -16438
rect 9755 -16472 9799 -16438
rect 9933 -16472 9977 -16438
rect 10111 -16472 10155 -16438
rect 10289 -16472 10333 -16438
rect 10467 -16472 10511 -16438
rect 10645 -16472 10689 -16438
rect 10823 -16472 10867 -16438
rect 11001 -16472 11045 -16438
rect 11179 -16472 11223 -16438
rect 11357 -16472 11401 -16438
rect 11535 -16472 11579 -16438
rect 11713 -16472 11757 -16438
rect 11891 -16472 11935 -16438
rect 12069 -16472 12113 -16438
rect 12247 -16472 12291 -16438
rect 12425 -16472 12469 -16438
rect 12603 -16472 12647 -16438
rect -5944 -16834 -5900 -16800
rect -5766 -16834 -5722 -16800
rect -5588 -16834 -5544 -16800
rect -5410 -16834 -5366 -16800
rect -5232 -16834 -5188 -16800
rect -5054 -16834 -5010 -16800
rect -4876 -16834 -4832 -16800
rect -4698 -16834 -4654 -16800
rect -4520 -16834 -4476 -16800
rect -4342 -16834 -4298 -16800
rect -4164 -16834 -4120 -16800
<< locali >>
rect 7040 2775 7136 2809
rect 8166 2775 8262 2809
rect 7040 2713 7074 2775
rect 8228 2713 8262 2775
rect 7138 2673 7154 2707
rect 7188 2673 7204 2707
rect 7330 2673 7346 2707
rect 7380 2673 7396 2707
rect 7522 2673 7538 2707
rect 7572 2673 7588 2707
rect 7714 2673 7730 2707
rect 7764 2673 7780 2707
rect 7906 2673 7922 2707
rect 7956 2673 7972 2707
rect 8098 2673 8114 2707
rect 8148 2673 8164 2707
rect 7154 2613 7188 2629
rect 7154 2349 7188 2365
rect 7250 2613 7284 2629
rect 7250 2349 7284 2365
rect 7346 2613 7380 2629
rect 7346 2349 7380 2365
rect 7442 2613 7476 2629
rect 7442 2349 7476 2365
rect 7538 2613 7572 2629
rect 7538 2349 7572 2365
rect 7634 2613 7668 2629
rect 7634 2349 7668 2365
rect 7730 2613 7764 2629
rect 7730 2349 7764 2365
rect 7826 2613 7860 2629
rect 7826 2349 7860 2365
rect 7922 2613 7956 2629
rect 7922 2349 7956 2365
rect 8018 2613 8052 2629
rect 8018 2349 8052 2365
rect 8114 2613 8148 2629
rect 8114 2349 8148 2365
rect 7040 2265 7074 2327
rect 8228 2265 8262 2327
rect 7040 2231 7136 2265
rect 8166 2231 8262 2265
rect 16040 2775 16136 2809
rect 17166 2775 17262 2809
rect 16040 2713 16074 2775
rect 17228 2713 17262 2775
rect 16138 2673 16154 2707
rect 16188 2673 16204 2707
rect 16330 2673 16346 2707
rect 16380 2673 16396 2707
rect 16522 2673 16538 2707
rect 16572 2673 16588 2707
rect 16714 2673 16730 2707
rect 16764 2673 16780 2707
rect 16906 2673 16922 2707
rect 16956 2673 16972 2707
rect 17098 2673 17114 2707
rect 17148 2673 17164 2707
rect 16154 2613 16188 2629
rect 16154 2349 16188 2365
rect 16250 2613 16284 2629
rect 16250 2349 16284 2365
rect 16346 2613 16380 2629
rect 16346 2349 16380 2365
rect 16442 2613 16476 2629
rect 16442 2349 16476 2365
rect 16538 2613 16572 2629
rect 16538 2349 16572 2365
rect 16634 2613 16668 2629
rect 16634 2349 16668 2365
rect 16730 2613 16764 2629
rect 16730 2349 16764 2365
rect 16826 2613 16860 2629
rect 16826 2349 16860 2365
rect 16922 2613 16956 2629
rect 16922 2349 16956 2365
rect 17018 2613 17052 2629
rect 17018 2349 17052 2365
rect 17114 2613 17148 2629
rect 17114 2349 17148 2365
rect 16040 2265 16074 2327
rect 17228 2265 17262 2327
rect 16040 2231 16136 2265
rect 17166 2231 17262 2265
rect 7040 2123 7136 2157
rect 8166 2123 8262 2157
rect 7040 2063 7074 2123
rect 8228 2061 8262 2123
rect 7154 2033 7188 2049
rect 7154 1937 7188 1953
rect 7250 2033 7284 2049
rect 7250 1937 7284 1953
rect 7346 2033 7380 2049
rect 7346 1937 7380 1953
rect 7442 2033 7476 2049
rect 7442 1937 7476 1953
rect 7538 2033 7572 2049
rect 7538 1937 7572 1953
rect 7634 2033 7668 2049
rect 7634 1937 7668 1953
rect 7730 2033 7764 2049
rect 7730 1937 7764 1953
rect 7826 2033 7860 2049
rect 7826 1937 7860 1953
rect 7922 2033 7956 2049
rect 7922 1937 7956 1953
rect 8018 2033 8052 2049
rect 8018 1937 8052 1953
rect 8114 2033 8148 2049
rect 8114 1937 8148 1953
rect 7138 1865 7154 1899
rect 7188 1865 7204 1899
rect 7330 1865 7346 1899
rect 7380 1865 7396 1899
rect 7522 1865 7538 1899
rect 7572 1865 7588 1899
rect 7714 1865 7730 1899
rect 7764 1865 7780 1899
rect 7906 1865 7922 1899
rect 7956 1865 7972 1899
rect 8098 1865 8114 1899
rect 8148 1865 8164 1899
rect 7040 1801 7074 1863
rect 8228 1801 8262 1863
rect 7040 1767 7136 1801
rect 8166 1767 8262 1801
rect 16040 2123 16136 2157
rect 17166 2123 17262 2157
rect 16040 2063 16074 2123
rect 17228 2061 17262 2123
rect 16154 2033 16188 2049
rect 16154 1937 16188 1953
rect 16250 2033 16284 2049
rect 16250 1937 16284 1953
rect 16346 2033 16380 2049
rect 16346 1937 16380 1953
rect 16442 2033 16476 2049
rect 16442 1937 16476 1953
rect 16538 2033 16572 2049
rect 16538 1937 16572 1953
rect 16634 2033 16668 2049
rect 16634 1937 16668 1953
rect 16730 2033 16764 2049
rect 16730 1937 16764 1953
rect 16826 2033 16860 2049
rect 16826 1937 16860 1953
rect 16922 2033 16956 2049
rect 16922 1937 16956 1953
rect 17018 2033 17052 2049
rect 17018 1937 17052 1953
rect 17114 2033 17148 2049
rect 17114 1937 17148 1953
rect 16138 1865 16154 1899
rect 16188 1865 16204 1899
rect 16330 1865 16346 1899
rect 16380 1865 16396 1899
rect 16522 1865 16538 1899
rect 16572 1865 16588 1899
rect 16714 1865 16730 1899
rect 16764 1865 16780 1899
rect 16906 1865 16922 1899
rect 16956 1865 16972 1899
rect 17098 1865 17114 1899
rect 17148 1865 17164 1899
rect 16040 1801 16074 1863
rect 17228 1801 17262 1863
rect 16040 1767 16136 1801
rect 17166 1767 17262 1801
rect 7040 975 7136 1009
rect 8166 975 8262 1009
rect 7040 913 7074 975
rect 8228 913 8262 975
rect 7138 873 7154 907
rect 7188 873 7204 907
rect 7330 873 7346 907
rect 7380 873 7396 907
rect 7522 873 7538 907
rect 7572 873 7588 907
rect 7714 873 7730 907
rect 7764 873 7780 907
rect 7906 873 7922 907
rect 7956 873 7972 907
rect 8098 873 8114 907
rect 8148 873 8164 907
rect 7154 813 7188 829
rect 7154 549 7188 565
rect 7250 813 7284 829
rect 7250 549 7284 565
rect 7346 813 7380 829
rect 7346 549 7380 565
rect 7442 813 7476 829
rect 7442 549 7476 565
rect 7538 813 7572 829
rect 7538 549 7572 565
rect 7634 813 7668 829
rect 7634 549 7668 565
rect 7730 813 7764 829
rect 7730 549 7764 565
rect 7826 813 7860 829
rect 7826 549 7860 565
rect 7922 813 7956 829
rect 7922 549 7956 565
rect 8018 813 8052 829
rect 8018 549 8052 565
rect 8114 813 8148 829
rect 8114 549 8148 565
rect 7040 465 7074 527
rect 8228 465 8262 527
rect 7040 431 7136 465
rect 8166 431 8262 465
rect 16040 975 16136 1009
rect 17166 975 17262 1009
rect 16040 913 16074 975
rect 17228 913 17262 975
rect 16138 873 16154 907
rect 16188 873 16204 907
rect 16330 873 16346 907
rect 16380 873 16396 907
rect 16522 873 16538 907
rect 16572 873 16588 907
rect 16714 873 16730 907
rect 16764 873 16780 907
rect 16906 873 16922 907
rect 16956 873 16972 907
rect 17098 873 17114 907
rect 17148 873 17164 907
rect 16154 813 16188 829
rect 16154 549 16188 565
rect 16250 813 16284 829
rect 16250 549 16284 565
rect 16346 813 16380 829
rect 16346 549 16380 565
rect 16442 813 16476 829
rect 16442 549 16476 565
rect 16538 813 16572 829
rect 16538 549 16572 565
rect 16634 813 16668 829
rect 16634 549 16668 565
rect 16730 813 16764 829
rect 16730 549 16764 565
rect 16826 813 16860 829
rect 16826 549 16860 565
rect 16922 813 16956 829
rect 16922 549 16956 565
rect 17018 813 17052 829
rect 17018 549 17052 565
rect 17114 813 17148 829
rect 17114 549 17148 565
rect 16040 465 16074 527
rect 17228 465 17262 527
rect 16040 431 16136 465
rect 17166 431 17262 465
rect 7040 323 7136 357
rect 8166 323 8262 357
rect 7040 263 7074 323
rect 8228 261 8262 323
rect 7154 233 7188 249
rect 7154 137 7188 153
rect 7250 233 7284 249
rect 7250 137 7284 153
rect 7346 233 7380 249
rect 7346 137 7380 153
rect 7442 233 7476 249
rect 7442 137 7476 153
rect 7538 233 7572 249
rect 7538 137 7572 153
rect 7634 233 7668 249
rect 7634 137 7668 153
rect 7730 233 7764 249
rect 7730 137 7764 153
rect 7826 233 7860 249
rect 7826 137 7860 153
rect 7922 233 7956 249
rect 7922 137 7956 153
rect 8018 233 8052 249
rect 8018 137 8052 153
rect 8114 233 8148 249
rect 8114 137 8148 153
rect 7138 65 7154 99
rect 7188 65 7204 99
rect 7330 65 7346 99
rect 7380 65 7396 99
rect 7522 65 7538 99
rect 7572 65 7588 99
rect 7714 65 7730 99
rect 7764 65 7780 99
rect 7906 65 7922 99
rect 7956 65 7972 99
rect 8098 65 8114 99
rect 8148 65 8164 99
rect 7040 1 7074 63
rect 8228 1 8262 63
rect 7040 -33 7136 1
rect 8166 -33 8262 1
rect 16040 323 16136 357
rect 17166 323 17262 357
rect 16040 263 16074 323
rect 17228 261 17262 323
rect 16154 233 16188 249
rect 16154 137 16188 153
rect 16250 233 16284 249
rect 16250 137 16284 153
rect 16346 233 16380 249
rect 16346 137 16380 153
rect 16442 233 16476 249
rect 16442 137 16476 153
rect 16538 233 16572 249
rect 16538 137 16572 153
rect 16634 233 16668 249
rect 16634 137 16668 153
rect 16730 233 16764 249
rect 16730 137 16764 153
rect 16826 233 16860 249
rect 16826 137 16860 153
rect 16922 233 16956 249
rect 16922 137 16956 153
rect 17018 233 17052 249
rect 17018 137 17052 153
rect 17114 233 17148 249
rect 17114 137 17148 153
rect 16138 65 16154 99
rect 16188 65 16204 99
rect 16330 65 16346 99
rect 16380 65 16396 99
rect 16522 65 16538 99
rect 16572 65 16588 99
rect 16714 65 16730 99
rect 16764 65 16780 99
rect 16906 65 16922 99
rect 16956 65 16972 99
rect 17098 65 17114 99
rect 17148 65 17164 99
rect 16040 1 16074 63
rect 17228 1 17262 63
rect 16040 -33 16136 1
rect 17166 -33 17262 1
rect 7040 -825 7136 -791
rect 8166 -825 8262 -791
rect 7040 -887 7074 -825
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect 3610 -1520 3703 -1353
rect 8228 -887 8262 -825
rect 7138 -927 7154 -893
rect 7188 -927 7204 -893
rect 7330 -927 7346 -893
rect 7380 -927 7396 -893
rect 7522 -927 7538 -893
rect 7572 -927 7588 -893
rect 7714 -927 7730 -893
rect 7764 -927 7780 -893
rect 7906 -927 7922 -893
rect 7956 -927 7972 -893
rect 8098 -927 8114 -893
rect 8148 -927 8164 -893
rect 7154 -987 7188 -971
rect 7154 -1251 7188 -1235
rect 7250 -987 7284 -971
rect 7250 -1251 7284 -1235
rect 7346 -987 7380 -971
rect 7346 -1251 7380 -1235
rect 7442 -987 7476 -971
rect 7442 -1251 7476 -1235
rect 7538 -987 7572 -971
rect 7538 -1251 7572 -1235
rect 7634 -987 7668 -971
rect 7634 -1251 7668 -1235
rect 7730 -987 7764 -971
rect 7730 -1251 7764 -1235
rect 7826 -987 7860 -971
rect 7826 -1251 7860 -1235
rect 7922 -987 7956 -971
rect 7922 -1251 7956 -1235
rect 8018 -987 8052 -971
rect 8018 -1251 8052 -1235
rect 8114 -987 8148 -971
rect 8114 -1251 8148 -1235
rect 7040 -1335 7074 -1273
rect 8228 -1335 8262 -1273
rect 7040 -1369 7136 -1335
rect 8166 -1369 8262 -1335
rect 16040 -825 16136 -791
rect 17166 -825 17262 -791
rect 16040 -887 16074 -825
rect 17228 -887 17262 -825
rect 16138 -927 16154 -893
rect 16188 -927 16204 -893
rect 16330 -927 16346 -893
rect 16380 -927 16396 -893
rect 16522 -927 16538 -893
rect 16572 -927 16588 -893
rect 16714 -927 16730 -893
rect 16764 -927 16780 -893
rect 16906 -927 16922 -893
rect 16956 -927 16972 -893
rect 17098 -927 17114 -893
rect 17148 -927 17164 -893
rect 16154 -987 16188 -971
rect 16154 -1251 16188 -1235
rect 16250 -987 16284 -971
rect 16250 -1251 16284 -1235
rect 16346 -987 16380 -971
rect 16346 -1251 16380 -1235
rect 16442 -987 16476 -971
rect 16442 -1251 16476 -1235
rect 16538 -987 16572 -971
rect 16538 -1251 16572 -1235
rect 16634 -987 16668 -971
rect 16634 -1251 16668 -1235
rect 16730 -987 16764 -971
rect 16730 -1251 16764 -1235
rect 16826 -987 16860 -971
rect 16826 -1251 16860 -1235
rect 16922 -987 16956 -971
rect 16922 -1251 16956 -1235
rect 17018 -987 17052 -971
rect 17018 -1251 17052 -1235
rect 17114 -987 17148 -971
rect 17114 -1251 17148 -1235
rect 16040 -1335 16074 -1273
rect 17228 -1335 17262 -1273
rect 16040 -1369 16136 -1335
rect 17166 -1369 17262 -1335
rect -6234 -2073 -6218 -2039
rect -6174 -2073 -6158 -2039
rect -6056 -2073 -6040 -2039
rect -5996 -2073 -5980 -2039
rect -5878 -2073 -5862 -2039
rect -5818 -2073 -5802 -2039
rect -5700 -2073 -5684 -2039
rect -5640 -2073 -5624 -2039
rect -5522 -2073 -5506 -2039
rect -5462 -2073 -5446 -2039
rect -5344 -2073 -5328 -2039
rect -5284 -2073 -5268 -2039
rect -5166 -2073 -5150 -2039
rect -5106 -2073 -5090 -2039
rect -4988 -2073 -4972 -2039
rect -4928 -2073 -4912 -2039
rect -4810 -2073 -4794 -2039
rect -4750 -2073 -4734 -2039
rect -4632 -2073 -4616 -2039
rect -4572 -2073 -4556 -2039
rect -4454 -2073 -4438 -2039
rect -4394 -2073 -4378 -2039
rect -4276 -2073 -4260 -2039
rect -4216 -2073 -4200 -2039
rect -4098 -2073 -4082 -2039
rect -4038 -2073 -4022 -2039
rect -3920 -2073 -3904 -2039
rect -3860 -2073 -3844 -2039
rect -3742 -2073 -3726 -2039
rect -3682 -2073 -3666 -2039
rect -3564 -2073 -3548 -2039
rect -3504 -2073 -3488 -2039
rect -6302 -2132 -6268 -2116
rect -6302 -2404 -6268 -2388
rect -6124 -2132 -6090 -2116
rect -6124 -2404 -6090 -2388
rect -5946 -2132 -5912 -2116
rect -5946 -2404 -5912 -2388
rect -5768 -2132 -5734 -2116
rect -5768 -2404 -5734 -2388
rect -5590 -2132 -5556 -2116
rect -5590 -2404 -5556 -2388
rect -5412 -2132 -5378 -2116
rect -5412 -2404 -5378 -2388
rect -5234 -2132 -5200 -2116
rect -5234 -2404 -5200 -2388
rect -5056 -2132 -5022 -2116
rect -5056 -2404 -5022 -2388
rect -4878 -2132 -4844 -2116
rect -4878 -2404 -4844 -2388
rect -4700 -2132 -4666 -2116
rect -4700 -2404 -4666 -2388
rect -4522 -2132 -4488 -2116
rect -4522 -2404 -4488 -2388
rect -4344 -2132 -4310 -2116
rect -4344 -2404 -4310 -2388
rect -4166 -2132 -4132 -2116
rect -4166 -2404 -4132 -2388
rect -3988 -2132 -3954 -2116
rect -3988 -2404 -3954 -2388
rect -3810 -2132 -3776 -2116
rect -3810 -2404 -3776 -2388
rect -3632 -2132 -3598 -2116
rect -3632 -2404 -3598 -2388
rect -3454 -2132 -3420 -2116
rect -3454 -2404 -3420 -2388
rect -6234 -2481 -6218 -2447
rect -6174 -2481 -6158 -2447
rect -6056 -2481 -6040 -2447
rect -5996 -2481 -5980 -2447
rect -5878 -2481 -5862 -2447
rect -5818 -2481 -5802 -2447
rect -5700 -2481 -5684 -2447
rect -5640 -2481 -5624 -2447
rect -5522 -2481 -5506 -2447
rect -5462 -2481 -5446 -2447
rect -5344 -2481 -5328 -2447
rect -5284 -2481 -5268 -2447
rect -5166 -2481 -5150 -2447
rect -5106 -2481 -5090 -2447
rect -4988 -2481 -4972 -2447
rect -4928 -2481 -4912 -2447
rect -4810 -2481 -4794 -2447
rect -4750 -2481 -4734 -2447
rect -4632 -2481 -4616 -2447
rect -4572 -2481 -4556 -2447
rect -4454 -2481 -4438 -2447
rect -4394 -2481 -4378 -2447
rect -4276 -2481 -4260 -2447
rect -4216 -2481 -4200 -2447
rect -4098 -2481 -4082 -2447
rect -4038 -2481 -4022 -2447
rect -3920 -2481 -3904 -2447
rect -3860 -2481 -3844 -2447
rect -3742 -2481 -3726 -2447
rect -3682 -2481 -3666 -2447
rect -3564 -2481 -3548 -2447
rect -3504 -2481 -3488 -2447
rect -1386 -2825 -1370 -2791
rect -1326 -2825 -1310 -2791
rect -1208 -2825 -1192 -2791
rect -1148 -2825 -1132 -2791
rect -1030 -2825 -1014 -2791
rect -970 -2825 -954 -2791
rect -852 -2825 -836 -2791
rect -792 -2825 -776 -2791
rect -674 -2825 -658 -2791
rect -614 -2825 -598 -2791
rect -496 -2825 -480 -2791
rect -436 -2825 -420 -2791
rect -318 -2825 -302 -2791
rect -258 -2825 -242 -2791
rect -140 -2825 -124 -2791
rect -80 -2825 -64 -2791
rect 38 -2825 54 -2791
rect 98 -2825 114 -2791
rect 216 -2825 232 -2791
rect 276 -2825 292 -2791
rect 394 -2825 410 -2791
rect 454 -2825 470 -2791
rect 572 -2825 588 -2791
rect 632 -2825 648 -2791
rect 750 -2825 766 -2791
rect 810 -2825 826 -2791
rect 928 -2825 944 -2791
rect 988 -2825 1004 -2791
rect 1106 -2825 1122 -2791
rect 1166 -2825 1182 -2791
rect 1284 -2825 1300 -2791
rect 1344 -2825 1360 -2791
rect 1462 -2825 1478 -2791
rect 1522 -2825 1538 -2791
rect 1640 -2825 1656 -2791
rect 1700 -2825 1716 -2791
rect 1818 -2825 1834 -2791
rect 1878 -2825 1894 -2791
rect 1996 -2825 2012 -2791
rect 2056 -2825 2072 -2791
rect 2174 -2825 2190 -2791
rect 2234 -2825 2250 -2791
rect 2352 -2825 2368 -2791
rect 2412 -2825 2428 -2791
rect 2530 -2825 2546 -2791
rect 2590 -2825 2606 -2791
rect -1454 -2884 -1420 -2868
rect -6234 -2943 -6218 -2909
rect -6174 -2943 -6158 -2909
rect -6056 -2943 -6040 -2909
rect -5996 -2943 -5980 -2909
rect -5878 -2943 -5862 -2909
rect -5818 -2943 -5802 -2909
rect -5700 -2943 -5684 -2909
rect -5640 -2943 -5624 -2909
rect -5522 -2943 -5506 -2909
rect -5462 -2943 -5446 -2909
rect -5344 -2943 -5328 -2909
rect -5284 -2943 -5268 -2909
rect -5166 -2943 -5150 -2909
rect -5106 -2943 -5090 -2909
rect -4988 -2943 -4972 -2909
rect -4928 -2943 -4912 -2909
rect -4810 -2943 -4794 -2909
rect -4750 -2943 -4734 -2909
rect -4632 -2943 -4616 -2909
rect -4572 -2943 -4556 -2909
rect -4454 -2943 -4438 -2909
rect -4394 -2943 -4378 -2909
rect -4276 -2943 -4260 -2909
rect -4216 -2943 -4200 -2909
rect -4098 -2943 -4082 -2909
rect -4038 -2943 -4022 -2909
rect -3920 -2943 -3904 -2909
rect -3860 -2943 -3844 -2909
rect -3742 -2943 -3726 -2909
rect -3682 -2943 -3666 -2909
rect -3564 -2943 -3548 -2909
rect -3504 -2943 -3488 -2909
rect -6302 -3002 -6268 -2986
rect -6302 -3274 -6268 -3258
rect -6124 -3002 -6090 -2986
rect -6124 -3274 -6090 -3258
rect -5946 -3002 -5912 -2986
rect -5946 -3274 -5912 -3258
rect -5768 -3002 -5734 -2986
rect -5768 -3274 -5734 -3258
rect -5590 -3002 -5556 -2986
rect -5590 -3274 -5556 -3258
rect -5412 -3002 -5378 -2986
rect -5412 -3274 -5378 -3258
rect -5234 -3002 -5200 -2986
rect -5234 -3274 -5200 -3258
rect -5056 -3002 -5022 -2986
rect -5056 -3274 -5022 -3258
rect -4878 -3002 -4844 -2986
rect -4878 -3274 -4844 -3258
rect -4700 -3002 -4666 -2986
rect -4700 -3274 -4666 -3258
rect -4522 -3002 -4488 -2986
rect -4522 -3274 -4488 -3258
rect -4344 -3002 -4310 -2986
rect -4344 -3274 -4310 -3258
rect -4166 -3002 -4132 -2986
rect -4166 -3274 -4132 -3258
rect -3988 -3002 -3954 -2986
rect -3988 -3274 -3954 -3258
rect -3810 -3002 -3776 -2986
rect -3810 -3274 -3776 -3258
rect -3632 -3002 -3598 -2986
rect -3632 -3274 -3598 -3258
rect -3454 -3002 -3420 -2986
rect -2210 -3043 -1984 -3019
rect -2210 -3221 -2186 -3043
rect -2008 -3221 -1984 -3043
rect -1454 -3156 -1420 -3140
rect -1276 -2884 -1242 -2868
rect -1276 -3156 -1242 -3140
rect -1098 -2884 -1064 -2868
rect -1098 -3156 -1064 -3140
rect -920 -2884 -886 -2868
rect -920 -3156 -886 -3140
rect -742 -2884 -708 -2868
rect -742 -3156 -708 -3140
rect -564 -2884 -530 -2868
rect -564 -3156 -530 -3140
rect -386 -2884 -352 -2868
rect -386 -3156 -352 -3140
rect -208 -2884 -174 -2868
rect -208 -3156 -174 -3140
rect -30 -2884 4 -2868
rect -30 -3156 4 -3140
rect 148 -2884 182 -2868
rect 148 -3156 182 -3140
rect 326 -2884 360 -2868
rect 326 -3156 360 -3140
rect 504 -2884 538 -2868
rect 504 -3156 538 -3140
rect 682 -2884 716 -2868
rect 682 -3156 716 -3140
rect 860 -2884 894 -2868
rect 860 -3156 894 -3140
rect 1038 -2884 1072 -2868
rect 1038 -3156 1072 -3140
rect 1216 -2884 1250 -2868
rect 1216 -3156 1250 -3140
rect 1394 -2884 1428 -2868
rect 1394 -3156 1428 -3140
rect 1572 -2884 1606 -2868
rect 1572 -3156 1606 -3140
rect 1750 -2884 1784 -2868
rect 1750 -3156 1784 -3140
rect 1928 -2884 1962 -2868
rect 1928 -3156 1962 -3140
rect 2106 -2884 2140 -2868
rect 2106 -3156 2140 -3140
rect 2284 -2884 2318 -2868
rect 2284 -3156 2318 -3140
rect 2462 -2884 2496 -2868
rect 2462 -3156 2496 -3140
rect 2640 -2884 2674 -2868
rect 2640 -3156 2674 -3140
rect -2210 -3245 -1984 -3221
rect -1386 -3233 -1370 -3199
rect -1326 -3233 -1310 -3199
rect -1208 -3233 -1192 -3199
rect -1148 -3233 -1132 -3199
rect -1030 -3233 -1014 -3199
rect -970 -3233 -954 -3199
rect -852 -3233 -836 -3199
rect -792 -3233 -776 -3199
rect -674 -3233 -658 -3199
rect -614 -3233 -598 -3199
rect -496 -3233 -480 -3199
rect -436 -3233 -420 -3199
rect -318 -3233 -302 -3199
rect -258 -3233 -242 -3199
rect -140 -3233 -124 -3199
rect -80 -3233 -64 -3199
rect 38 -3233 54 -3199
rect 98 -3233 114 -3199
rect 216 -3233 232 -3199
rect 276 -3233 292 -3199
rect 394 -3233 410 -3199
rect 454 -3233 470 -3199
rect 572 -3233 588 -3199
rect 632 -3233 648 -3199
rect 750 -3233 766 -3199
rect 810 -3233 826 -3199
rect 928 -3233 944 -3199
rect 988 -3233 1004 -3199
rect 1106 -3233 1122 -3199
rect 1166 -3233 1182 -3199
rect 1284 -3233 1300 -3199
rect 1344 -3233 1360 -3199
rect 1462 -3233 1478 -3199
rect 1522 -3233 1538 -3199
rect 1640 -3233 1656 -3199
rect 1700 -3233 1716 -3199
rect 1818 -3233 1834 -3199
rect 1878 -3233 1894 -3199
rect 1996 -3233 2012 -3199
rect 2056 -3233 2072 -3199
rect 2174 -3233 2190 -3199
rect 2234 -3233 2250 -3199
rect 2352 -3233 2368 -3199
rect 2412 -3233 2428 -3199
rect 2530 -3233 2546 -3199
rect 2590 -3233 2606 -3199
rect -3454 -3274 -3420 -3258
rect -6234 -3351 -6218 -3317
rect -6174 -3351 -6158 -3317
rect -6056 -3351 -6040 -3317
rect -5996 -3351 -5980 -3317
rect -5878 -3351 -5862 -3317
rect -5818 -3351 -5802 -3317
rect -5700 -3351 -5684 -3317
rect -5640 -3351 -5624 -3317
rect -5522 -3351 -5506 -3317
rect -5462 -3351 -5446 -3317
rect -5344 -3351 -5328 -3317
rect -5284 -3351 -5268 -3317
rect -5166 -3351 -5150 -3317
rect -5106 -3351 -5090 -3317
rect -4988 -3351 -4972 -3317
rect -4928 -3351 -4912 -3317
rect -4810 -3351 -4794 -3317
rect -4750 -3351 -4734 -3317
rect -4632 -3351 -4616 -3317
rect -4572 -3351 -4556 -3317
rect -4454 -3351 -4438 -3317
rect -4394 -3351 -4378 -3317
rect -4276 -3351 -4260 -3317
rect -4216 -3351 -4200 -3317
rect -4098 -3351 -4082 -3317
rect -4038 -3351 -4022 -3317
rect -3920 -3351 -3904 -3317
rect -3860 -3351 -3844 -3317
rect -3742 -3351 -3726 -3317
rect -3682 -3351 -3666 -3317
rect -3564 -3351 -3548 -3317
rect -3504 -3351 -3488 -3317
rect -1386 -3725 -1370 -3691
rect -1326 -3725 -1310 -3691
rect -1208 -3725 -1192 -3691
rect -1148 -3725 -1132 -3691
rect -1030 -3725 -1014 -3691
rect -970 -3725 -954 -3691
rect -852 -3725 -836 -3691
rect -792 -3725 -776 -3691
rect -674 -3725 -658 -3691
rect -614 -3725 -598 -3691
rect -496 -3725 -480 -3691
rect -436 -3725 -420 -3691
rect -318 -3725 -302 -3691
rect -258 -3725 -242 -3691
rect -140 -3725 -124 -3691
rect -80 -3725 -64 -3691
rect 38 -3725 54 -3691
rect 98 -3725 114 -3691
rect 216 -3725 232 -3691
rect 276 -3725 292 -3691
rect 394 -3725 410 -3691
rect 454 -3725 470 -3691
rect 572 -3725 588 -3691
rect 632 -3725 648 -3691
rect 750 -3725 766 -3691
rect 810 -3725 826 -3691
rect 928 -3725 944 -3691
rect 988 -3725 1004 -3691
rect 1106 -3725 1122 -3691
rect 1166 -3725 1182 -3691
rect 1284 -3725 1300 -3691
rect 1344 -3725 1360 -3691
rect 1462 -3725 1478 -3691
rect 1522 -3725 1538 -3691
rect 1640 -3725 1656 -3691
rect 1700 -3725 1716 -3691
rect 1818 -3725 1834 -3691
rect 1878 -3725 1894 -3691
rect 1996 -3725 2012 -3691
rect 2056 -3725 2072 -3691
rect 2174 -3725 2190 -3691
rect 2234 -3725 2250 -3691
rect 2352 -3725 2368 -3691
rect 2412 -3725 2428 -3691
rect 2530 -3725 2546 -3691
rect 2590 -3725 2606 -3691
rect -6234 -3813 -6218 -3779
rect -6174 -3813 -6158 -3779
rect -6056 -3813 -6040 -3779
rect -5996 -3813 -5980 -3779
rect -5878 -3813 -5862 -3779
rect -5818 -3813 -5802 -3779
rect -5700 -3813 -5684 -3779
rect -5640 -3813 -5624 -3779
rect -5522 -3813 -5506 -3779
rect -5462 -3813 -5446 -3779
rect -5344 -3813 -5328 -3779
rect -5284 -3813 -5268 -3779
rect -5166 -3813 -5150 -3779
rect -5106 -3813 -5090 -3779
rect -4988 -3813 -4972 -3779
rect -4928 -3813 -4912 -3779
rect -4810 -3813 -4794 -3779
rect -4750 -3813 -4734 -3779
rect -4632 -3813 -4616 -3779
rect -4572 -3813 -4556 -3779
rect -4454 -3813 -4438 -3779
rect -4394 -3813 -4378 -3779
rect -4276 -3813 -4260 -3779
rect -4216 -3813 -4200 -3779
rect -4098 -3813 -4082 -3779
rect -4038 -3813 -4022 -3779
rect -3920 -3813 -3904 -3779
rect -3860 -3813 -3844 -3779
rect -3742 -3813 -3726 -3779
rect -3682 -3813 -3666 -3779
rect -3564 -3813 -3548 -3779
rect -3504 -3813 -3488 -3779
rect -1454 -3784 -1420 -3768
rect -6302 -3872 -6268 -3856
rect -6302 -4144 -6268 -4128
rect -6124 -3872 -6090 -3856
rect -6124 -4144 -6090 -4128
rect -5946 -3872 -5912 -3856
rect -5946 -4144 -5912 -4128
rect -5768 -3872 -5734 -3856
rect -5768 -4144 -5734 -4128
rect -5590 -3872 -5556 -3856
rect -5590 -4144 -5556 -4128
rect -5412 -3872 -5378 -3856
rect -5412 -4144 -5378 -4128
rect -5234 -3872 -5200 -3856
rect -5234 -4144 -5200 -4128
rect -5056 -3872 -5022 -3856
rect -5056 -4144 -5022 -4128
rect -4878 -3872 -4844 -3856
rect -4878 -4144 -4844 -4128
rect -4700 -3872 -4666 -3856
rect -4700 -4144 -4666 -4128
rect -4522 -3872 -4488 -3856
rect -4522 -4144 -4488 -4128
rect -4344 -3872 -4310 -3856
rect -4344 -4144 -4310 -4128
rect -4166 -3872 -4132 -3856
rect -4166 -4144 -4132 -4128
rect -3988 -3872 -3954 -3856
rect -3988 -4144 -3954 -4128
rect -3810 -3872 -3776 -3856
rect -3810 -4144 -3776 -4128
rect -3632 -3872 -3598 -3856
rect -3632 -4144 -3598 -4128
rect -3454 -3872 -3420 -3856
rect -1454 -4056 -1420 -4040
rect -1276 -3784 -1242 -3768
rect -1276 -4056 -1242 -4040
rect -1098 -3784 -1064 -3768
rect -1098 -4056 -1064 -4040
rect -920 -3784 -886 -3768
rect -920 -4056 -886 -4040
rect -742 -3784 -708 -3768
rect -742 -4056 -708 -4040
rect -564 -3784 -530 -3768
rect -564 -4056 -530 -4040
rect -386 -3784 -352 -3768
rect -386 -4056 -352 -4040
rect -208 -3784 -174 -3768
rect -208 -4056 -174 -4040
rect -30 -3784 4 -3768
rect -30 -4056 4 -4040
rect 148 -3784 182 -3768
rect 148 -4056 182 -4040
rect 326 -3784 360 -3768
rect 326 -4056 360 -4040
rect 504 -3784 538 -3768
rect 504 -4056 538 -4040
rect 682 -3784 716 -3768
rect 682 -4056 716 -4040
rect 860 -3784 894 -3768
rect 860 -4056 894 -4040
rect 1038 -3784 1072 -3768
rect 1038 -4056 1072 -4040
rect 1216 -3784 1250 -3768
rect 1216 -4056 1250 -4040
rect 1394 -3784 1428 -3768
rect 1394 -4056 1428 -4040
rect 1572 -3784 1606 -3768
rect 1572 -4056 1606 -4040
rect 1750 -3784 1784 -3768
rect 1750 -4056 1784 -4040
rect 1928 -3784 1962 -3768
rect 1928 -4056 1962 -4040
rect 2106 -3784 2140 -3768
rect 2106 -4056 2140 -4040
rect 2284 -3784 2318 -3768
rect 2284 -4056 2318 -4040
rect 2462 -3784 2496 -3768
rect 2462 -4056 2496 -4040
rect 2640 -3784 2674 -3768
rect 2640 -4056 2674 -4040
rect -3454 -4144 -3420 -4128
rect -1386 -4133 -1370 -4099
rect -1326 -4133 -1310 -4099
rect -1208 -4133 -1192 -4099
rect -1148 -4133 -1132 -4099
rect -1030 -4133 -1014 -4099
rect -970 -4133 -954 -4099
rect -852 -4133 -836 -4099
rect -792 -4133 -776 -4099
rect -674 -4133 -658 -4099
rect -614 -4133 -598 -4099
rect -496 -4133 -480 -4099
rect -436 -4133 -420 -4099
rect -318 -4133 -302 -4099
rect -258 -4133 -242 -4099
rect -140 -4133 -124 -4099
rect -80 -4133 -64 -4099
rect 38 -4133 54 -4099
rect 98 -4133 114 -4099
rect 216 -4133 232 -4099
rect 276 -4133 292 -4099
rect 394 -4133 410 -4099
rect 454 -4133 470 -4099
rect 572 -4133 588 -4099
rect 632 -4133 648 -4099
rect 750 -4133 766 -4099
rect 810 -4133 826 -4099
rect 928 -4133 944 -4099
rect 988 -4133 1004 -4099
rect 1106 -4133 1122 -4099
rect 1166 -4133 1182 -4099
rect 1284 -4133 1300 -4099
rect 1344 -4133 1360 -4099
rect 1462 -4133 1478 -4099
rect 1522 -4133 1538 -4099
rect 1640 -4133 1656 -4099
rect 1700 -4133 1716 -4099
rect 1818 -4133 1834 -4099
rect 1878 -4133 1894 -4099
rect 1996 -4133 2012 -4099
rect 2056 -4133 2072 -4099
rect 2174 -4133 2190 -4099
rect 2234 -4133 2250 -4099
rect 2352 -4133 2368 -4099
rect 2412 -4133 2428 -4099
rect 2530 -4133 2546 -4099
rect 2590 -4133 2606 -4099
rect -6234 -4221 -6218 -4187
rect -6174 -4221 -6158 -4187
rect -6056 -4221 -6040 -4187
rect -5996 -4221 -5980 -4187
rect -5878 -4221 -5862 -4187
rect -5818 -4221 -5802 -4187
rect -5700 -4221 -5684 -4187
rect -5640 -4221 -5624 -4187
rect -5522 -4221 -5506 -4187
rect -5462 -4221 -5446 -4187
rect -5344 -4221 -5328 -4187
rect -5284 -4221 -5268 -4187
rect -5166 -4221 -5150 -4187
rect -5106 -4221 -5090 -4187
rect -4988 -4221 -4972 -4187
rect -4928 -4221 -4912 -4187
rect -4810 -4221 -4794 -4187
rect -4750 -4221 -4734 -4187
rect -4632 -4221 -4616 -4187
rect -4572 -4221 -4556 -4187
rect -4454 -4221 -4438 -4187
rect -4394 -4221 -4378 -4187
rect -4276 -4221 -4260 -4187
rect -4216 -4221 -4200 -4187
rect -4098 -4221 -4082 -4187
rect -4038 -4221 -4022 -4187
rect -3920 -4221 -3904 -4187
rect -3860 -4221 -3844 -4187
rect -3742 -4221 -3726 -4187
rect -3682 -4221 -3666 -4187
rect -3564 -4221 -3548 -4187
rect -3504 -4221 -3488 -4187
rect -1386 -4625 -1370 -4591
rect -1326 -4625 -1310 -4591
rect -1208 -4625 -1192 -4591
rect -1148 -4625 -1132 -4591
rect -1030 -4625 -1014 -4591
rect -970 -4625 -954 -4591
rect -852 -4625 -836 -4591
rect -792 -4625 -776 -4591
rect -674 -4625 -658 -4591
rect -614 -4625 -598 -4591
rect -496 -4625 -480 -4591
rect -436 -4625 -420 -4591
rect -318 -4625 -302 -4591
rect -258 -4625 -242 -4591
rect -140 -4625 -124 -4591
rect -80 -4625 -64 -4591
rect 38 -4625 54 -4591
rect 98 -4625 114 -4591
rect 216 -4625 232 -4591
rect 276 -4625 292 -4591
rect 394 -4625 410 -4591
rect 454 -4625 470 -4591
rect 572 -4625 588 -4591
rect 632 -4625 648 -4591
rect 750 -4625 766 -4591
rect 810 -4625 826 -4591
rect 928 -4625 944 -4591
rect 988 -4625 1004 -4591
rect 1106 -4625 1122 -4591
rect 1166 -4625 1182 -4591
rect 1284 -4625 1300 -4591
rect 1344 -4625 1360 -4591
rect 1462 -4625 1478 -4591
rect 1522 -4625 1538 -4591
rect 1640 -4625 1656 -4591
rect 1700 -4625 1716 -4591
rect 1818 -4625 1834 -4591
rect 1878 -4625 1894 -4591
rect 1996 -4625 2012 -4591
rect 2056 -4625 2072 -4591
rect 2174 -4625 2190 -4591
rect 2234 -4625 2250 -4591
rect 2352 -4625 2368 -4591
rect 2412 -4625 2428 -4591
rect 2530 -4625 2546 -4591
rect 2590 -4625 2606 -4591
rect -6234 -4683 -6218 -4649
rect -6174 -4683 -6158 -4649
rect -6056 -4683 -6040 -4649
rect -5996 -4683 -5980 -4649
rect -5878 -4683 -5862 -4649
rect -5818 -4683 -5802 -4649
rect -5700 -4683 -5684 -4649
rect -5640 -4683 -5624 -4649
rect -5522 -4683 -5506 -4649
rect -5462 -4683 -5446 -4649
rect -5344 -4683 -5328 -4649
rect -5284 -4683 -5268 -4649
rect -5166 -4683 -5150 -4649
rect -5106 -4683 -5090 -4649
rect -4988 -4683 -4972 -4649
rect -4928 -4683 -4912 -4649
rect -4810 -4683 -4794 -4649
rect -4750 -4683 -4734 -4649
rect -4632 -4683 -4616 -4649
rect -4572 -4683 -4556 -4649
rect -4454 -4683 -4438 -4649
rect -4394 -4683 -4378 -4649
rect -4276 -4683 -4260 -4649
rect -4216 -4683 -4200 -4649
rect -4098 -4683 -4082 -4649
rect -4038 -4683 -4022 -4649
rect -3920 -4683 -3904 -4649
rect -3860 -4683 -3844 -4649
rect -3742 -4683 -3726 -4649
rect -3682 -4683 -3666 -4649
rect -3564 -4683 -3548 -4649
rect -3504 -4683 -3488 -4649
rect -1454 -4684 -1420 -4668
rect -6302 -4742 -6268 -4726
rect -6302 -5014 -6268 -4998
rect -6124 -4742 -6090 -4726
rect -6124 -5014 -6090 -4998
rect -5946 -4742 -5912 -4726
rect -5946 -5014 -5912 -4998
rect -5768 -4742 -5734 -4726
rect -5768 -5014 -5734 -4998
rect -5590 -4742 -5556 -4726
rect -5590 -5014 -5556 -4998
rect -5412 -4742 -5378 -4726
rect -5412 -5014 -5378 -4998
rect -5234 -4742 -5200 -4726
rect -5234 -5014 -5200 -4998
rect -5056 -4742 -5022 -4726
rect -5056 -5014 -5022 -4998
rect -4878 -4742 -4844 -4726
rect -4878 -5014 -4844 -4998
rect -4700 -4742 -4666 -4726
rect -4700 -5014 -4666 -4998
rect -4522 -4742 -4488 -4726
rect -4522 -5014 -4488 -4998
rect -4344 -4742 -4310 -4726
rect -4344 -5014 -4310 -4998
rect -4166 -4742 -4132 -4726
rect -4166 -5014 -4132 -4998
rect -3988 -4742 -3954 -4726
rect -3988 -5014 -3954 -4998
rect -3810 -4742 -3776 -4726
rect -3810 -5014 -3776 -4998
rect -3632 -4742 -3598 -4726
rect -3632 -5014 -3598 -4998
rect -3454 -4742 -3420 -4726
rect -1454 -4956 -1420 -4940
rect -1276 -4684 -1242 -4668
rect -1276 -4956 -1242 -4940
rect -1098 -4684 -1064 -4668
rect -1098 -4956 -1064 -4940
rect -920 -4684 -886 -4668
rect -920 -4956 -886 -4940
rect -742 -4684 -708 -4668
rect -742 -4956 -708 -4940
rect -564 -4684 -530 -4668
rect -564 -4956 -530 -4940
rect -386 -4684 -352 -4668
rect -386 -4956 -352 -4940
rect -208 -4684 -174 -4668
rect -208 -4956 -174 -4940
rect -30 -4684 4 -4668
rect -30 -4956 4 -4940
rect 148 -4684 182 -4668
rect 148 -4956 182 -4940
rect 326 -4684 360 -4668
rect 326 -4956 360 -4940
rect 504 -4684 538 -4668
rect 504 -4956 538 -4940
rect 682 -4684 716 -4668
rect 682 -4956 716 -4940
rect 860 -4684 894 -4668
rect 860 -4956 894 -4940
rect 1038 -4684 1072 -4668
rect 1038 -4956 1072 -4940
rect 1216 -4684 1250 -4668
rect 1216 -4956 1250 -4940
rect 1394 -4684 1428 -4668
rect 1394 -4956 1428 -4940
rect 1572 -4684 1606 -4668
rect 1572 -4956 1606 -4940
rect 1750 -4684 1784 -4668
rect 1750 -4956 1784 -4940
rect 1928 -4684 1962 -4668
rect 1928 -4956 1962 -4940
rect 2106 -4684 2140 -4668
rect 2106 -4956 2140 -4940
rect 2284 -4684 2318 -4668
rect 2284 -4956 2318 -4940
rect 2462 -4684 2496 -4668
rect 2462 -4956 2496 -4940
rect 2640 -4684 2674 -4668
rect 2640 -4956 2674 -4940
rect -3454 -5014 -3420 -4998
rect -1386 -5033 -1370 -4999
rect -1326 -5033 -1310 -4999
rect -1208 -5033 -1192 -4999
rect -1148 -5033 -1132 -4999
rect -1030 -5033 -1014 -4999
rect -970 -5033 -954 -4999
rect -852 -5033 -836 -4999
rect -792 -5033 -776 -4999
rect -674 -5033 -658 -4999
rect -614 -5033 -598 -4999
rect -496 -5033 -480 -4999
rect -436 -5033 -420 -4999
rect -318 -5033 -302 -4999
rect -258 -5033 -242 -4999
rect -140 -5033 -124 -4999
rect -80 -5033 -64 -4999
rect 38 -5033 54 -4999
rect 98 -5033 114 -4999
rect 216 -5033 232 -4999
rect 276 -5033 292 -4999
rect 394 -5033 410 -4999
rect 454 -5033 470 -4999
rect 572 -5033 588 -4999
rect 632 -5033 648 -4999
rect 750 -5033 766 -4999
rect 810 -5033 826 -4999
rect 928 -5033 944 -4999
rect 988 -5033 1004 -4999
rect 1106 -5033 1122 -4999
rect 1166 -5033 1182 -4999
rect 1284 -5033 1300 -4999
rect 1344 -5033 1360 -4999
rect 1462 -5033 1478 -4999
rect 1522 -5033 1538 -4999
rect 1640 -5033 1656 -4999
rect 1700 -5033 1716 -4999
rect 1818 -5033 1834 -4999
rect 1878 -5033 1894 -4999
rect 1996 -5033 2012 -4999
rect 2056 -5033 2072 -4999
rect 2174 -5033 2190 -4999
rect 2234 -5033 2250 -4999
rect 2352 -5033 2368 -4999
rect 2412 -5033 2428 -4999
rect 2530 -5033 2546 -4999
rect 2590 -5033 2606 -4999
rect -6234 -5091 -6218 -5057
rect -6174 -5091 -6158 -5057
rect -6056 -5091 -6040 -5057
rect -5996 -5091 -5980 -5057
rect -5878 -5091 -5862 -5057
rect -5818 -5091 -5802 -5057
rect -5700 -5091 -5684 -5057
rect -5640 -5091 -5624 -5057
rect -5522 -5091 -5506 -5057
rect -5462 -5091 -5446 -5057
rect -5344 -5091 -5328 -5057
rect -5284 -5091 -5268 -5057
rect -5166 -5091 -5150 -5057
rect -5106 -5091 -5090 -5057
rect -4988 -5091 -4972 -5057
rect -4928 -5091 -4912 -5057
rect -4810 -5091 -4794 -5057
rect -4750 -5091 -4734 -5057
rect -4632 -5091 -4616 -5057
rect -4572 -5091 -4556 -5057
rect -4454 -5091 -4438 -5057
rect -4394 -5091 -4378 -5057
rect -4276 -5091 -4260 -5057
rect -4216 -5091 -4200 -5057
rect -4098 -5091 -4082 -5057
rect -4038 -5091 -4022 -5057
rect -3920 -5091 -3904 -5057
rect -3860 -5091 -3844 -5057
rect -3742 -5091 -3726 -5057
rect -3682 -5091 -3666 -5057
rect -3564 -5091 -3548 -5057
rect -3504 -5091 -3488 -5057
rect -6234 -5553 -6218 -5519
rect -6174 -5553 -6158 -5519
rect -6056 -5553 -6040 -5519
rect -5996 -5553 -5980 -5519
rect -5878 -5553 -5862 -5519
rect -5818 -5553 -5802 -5519
rect -5700 -5553 -5684 -5519
rect -5640 -5553 -5624 -5519
rect -5522 -5553 -5506 -5519
rect -5462 -5553 -5446 -5519
rect -5344 -5553 -5328 -5519
rect -5284 -5553 -5268 -5519
rect -5166 -5553 -5150 -5519
rect -5106 -5553 -5090 -5519
rect -4988 -5553 -4972 -5519
rect -4928 -5553 -4912 -5519
rect -4810 -5553 -4794 -5519
rect -4750 -5553 -4734 -5519
rect -4632 -5553 -4616 -5519
rect -4572 -5553 -4556 -5519
rect -4454 -5553 -4438 -5519
rect -4394 -5553 -4378 -5519
rect -4276 -5553 -4260 -5519
rect -4216 -5553 -4200 -5519
rect -4098 -5553 -4082 -5519
rect -4038 -5553 -4022 -5519
rect -3920 -5553 -3904 -5519
rect -3860 -5553 -3844 -5519
rect -3742 -5553 -3726 -5519
rect -3682 -5553 -3666 -5519
rect -3564 -5553 -3548 -5519
rect -3504 -5553 -3488 -5519
rect -1386 -5525 -1370 -5491
rect -1326 -5525 -1310 -5491
rect -1208 -5525 -1192 -5491
rect -1148 -5525 -1132 -5491
rect -1030 -5525 -1014 -5491
rect -970 -5525 -954 -5491
rect -852 -5525 -836 -5491
rect -792 -5525 -776 -5491
rect -674 -5525 -658 -5491
rect -614 -5525 -598 -5491
rect -496 -5525 -480 -5491
rect -436 -5525 -420 -5491
rect -318 -5525 -302 -5491
rect -258 -5525 -242 -5491
rect -140 -5525 -124 -5491
rect -80 -5525 -64 -5491
rect 38 -5525 54 -5491
rect 98 -5525 114 -5491
rect 216 -5525 232 -5491
rect 276 -5525 292 -5491
rect 394 -5525 410 -5491
rect 454 -5525 470 -5491
rect 572 -5525 588 -5491
rect 632 -5525 648 -5491
rect 750 -5525 766 -5491
rect 810 -5525 826 -5491
rect 928 -5525 944 -5491
rect 988 -5525 1004 -5491
rect 1106 -5525 1122 -5491
rect 1166 -5525 1182 -5491
rect 1284 -5525 1300 -5491
rect 1344 -5525 1360 -5491
rect 1462 -5525 1478 -5491
rect 1522 -5525 1538 -5491
rect 1640 -5525 1656 -5491
rect 1700 -5525 1716 -5491
rect 1818 -5525 1834 -5491
rect 1878 -5525 1894 -5491
rect 1996 -5525 2012 -5491
rect 2056 -5525 2072 -5491
rect 2174 -5525 2190 -5491
rect 2234 -5525 2250 -5491
rect 2352 -5525 2368 -5491
rect 2412 -5525 2428 -5491
rect 2530 -5525 2546 -5491
rect 2590 -5525 2606 -5491
rect -1454 -5584 -1420 -5568
rect -6302 -5612 -6268 -5596
rect -6302 -5884 -6268 -5868
rect -6124 -5612 -6090 -5596
rect -6124 -5884 -6090 -5868
rect -5946 -5612 -5912 -5596
rect -5946 -5884 -5912 -5868
rect -5768 -5612 -5734 -5596
rect -5768 -5884 -5734 -5868
rect -5590 -5612 -5556 -5596
rect -5590 -5884 -5556 -5868
rect -5412 -5612 -5378 -5596
rect -5412 -5884 -5378 -5868
rect -5234 -5612 -5200 -5596
rect -5234 -5884 -5200 -5868
rect -5056 -5612 -5022 -5596
rect -5056 -5884 -5022 -5868
rect -4878 -5612 -4844 -5596
rect -4878 -5884 -4844 -5868
rect -4700 -5612 -4666 -5596
rect -4700 -5884 -4666 -5868
rect -4522 -5612 -4488 -5596
rect -4522 -5884 -4488 -5868
rect -4344 -5612 -4310 -5596
rect -4344 -5884 -4310 -5868
rect -4166 -5612 -4132 -5596
rect -4166 -5884 -4132 -5868
rect -3988 -5612 -3954 -5596
rect -3988 -5884 -3954 -5868
rect -3810 -5612 -3776 -5596
rect -3810 -5884 -3776 -5868
rect -3632 -5612 -3598 -5596
rect -3632 -5884 -3598 -5868
rect -3454 -5612 -3420 -5596
rect -3058 -5662 -2832 -5638
rect -3058 -5840 -3034 -5662
rect -2856 -5840 -2832 -5662
rect -3058 -5864 -2832 -5840
rect -1454 -5856 -1420 -5840
rect -1276 -5584 -1242 -5568
rect -1276 -5856 -1242 -5840
rect -1098 -5584 -1064 -5568
rect -1098 -5856 -1064 -5840
rect -920 -5584 -886 -5568
rect -920 -5856 -886 -5840
rect -742 -5584 -708 -5568
rect -742 -5856 -708 -5840
rect -564 -5584 -530 -5568
rect -564 -5856 -530 -5840
rect -386 -5584 -352 -5568
rect -386 -5856 -352 -5840
rect -208 -5584 -174 -5568
rect -208 -5856 -174 -5840
rect -30 -5584 4 -5568
rect -30 -5856 4 -5840
rect 148 -5584 182 -5568
rect 148 -5856 182 -5840
rect 326 -5584 360 -5568
rect 326 -5856 360 -5840
rect 504 -5584 538 -5568
rect 504 -5856 538 -5840
rect 682 -5584 716 -5568
rect 682 -5856 716 -5840
rect 860 -5584 894 -5568
rect 860 -5856 894 -5840
rect 1038 -5584 1072 -5568
rect 1038 -5856 1072 -5840
rect 1216 -5584 1250 -5568
rect 1216 -5856 1250 -5840
rect 1394 -5584 1428 -5568
rect 1394 -5856 1428 -5840
rect 1572 -5584 1606 -5568
rect 1572 -5856 1606 -5840
rect 1750 -5584 1784 -5568
rect 1750 -5856 1784 -5840
rect 1928 -5584 1962 -5568
rect 1928 -5856 1962 -5840
rect 2106 -5584 2140 -5568
rect 2106 -5856 2140 -5840
rect 2284 -5584 2318 -5568
rect 2284 -5856 2318 -5840
rect 2462 -5584 2496 -5568
rect 2462 -5856 2496 -5840
rect 2640 -5584 2674 -5568
rect 2640 -5856 2674 -5840
rect -3454 -5884 -3420 -5868
rect -6234 -5961 -6218 -5927
rect -6174 -5961 -6158 -5927
rect -6056 -5961 -6040 -5927
rect -5996 -5961 -5980 -5927
rect -5878 -5961 -5862 -5927
rect -5818 -5961 -5802 -5927
rect -5700 -5961 -5684 -5927
rect -5640 -5961 -5624 -5927
rect -5522 -5961 -5506 -5927
rect -5462 -5961 -5446 -5927
rect -5344 -5961 -5328 -5927
rect -5284 -5961 -5268 -5927
rect -5166 -5961 -5150 -5927
rect -5106 -5961 -5090 -5927
rect -4988 -5961 -4972 -5927
rect -4928 -5961 -4912 -5927
rect -4810 -5961 -4794 -5927
rect -4750 -5961 -4734 -5927
rect -4632 -5961 -4616 -5927
rect -4572 -5961 -4556 -5927
rect -4454 -5961 -4438 -5927
rect -4394 -5961 -4378 -5927
rect -4276 -5961 -4260 -5927
rect -4216 -5961 -4200 -5927
rect -4098 -5961 -4082 -5927
rect -4038 -5961 -4022 -5927
rect -3920 -5961 -3904 -5927
rect -3860 -5961 -3844 -5927
rect -3742 -5961 -3726 -5927
rect -3682 -5961 -3666 -5927
rect -3564 -5961 -3548 -5927
rect -3504 -5961 -3488 -5927
rect -1386 -5933 -1370 -5899
rect -1326 -5933 -1310 -5899
rect -1208 -5933 -1192 -5899
rect -1148 -5933 -1132 -5899
rect -1030 -5933 -1014 -5899
rect -970 -5933 -954 -5899
rect -852 -5933 -836 -5899
rect -792 -5933 -776 -5899
rect -674 -5933 -658 -5899
rect -614 -5933 -598 -5899
rect -496 -5933 -480 -5899
rect -436 -5933 -420 -5899
rect -318 -5933 -302 -5899
rect -258 -5933 -242 -5899
rect -140 -5933 -124 -5899
rect -80 -5933 -64 -5899
rect 38 -5933 54 -5899
rect 98 -5933 114 -5899
rect 216 -5933 232 -5899
rect 276 -5933 292 -5899
rect 394 -5933 410 -5899
rect 454 -5933 470 -5899
rect 572 -5933 588 -5899
rect 632 -5933 648 -5899
rect 750 -5933 766 -5899
rect 810 -5933 826 -5899
rect 928 -5933 944 -5899
rect 988 -5933 1004 -5899
rect 1106 -5933 1122 -5899
rect 1166 -5933 1182 -5899
rect 1284 -5933 1300 -5899
rect 1344 -5933 1360 -5899
rect 1462 -5933 1478 -5899
rect 1522 -5933 1538 -5899
rect 1640 -5933 1656 -5899
rect 1700 -5933 1716 -5899
rect 1818 -5933 1834 -5899
rect 1878 -5933 1894 -5899
rect 1996 -5933 2012 -5899
rect 2056 -5933 2072 -5899
rect 2174 -5933 2190 -5899
rect 2234 -5933 2250 -5899
rect 2352 -5933 2368 -5899
rect 2412 -5933 2428 -5899
rect 2530 -5933 2546 -5899
rect 2590 -5933 2606 -5899
rect -7605 -7140 -7512 -6976
rect 7040 -1477 7136 -1443
rect 8166 -1477 8262 -1443
rect 7040 -1537 7074 -1477
rect 8228 -1539 8262 -1477
rect 7154 -1567 7188 -1551
rect 7154 -1663 7188 -1647
rect 7250 -1567 7284 -1551
rect 7250 -1663 7284 -1647
rect 7346 -1567 7380 -1551
rect 7346 -1663 7380 -1647
rect 7442 -1567 7476 -1551
rect 7442 -1663 7476 -1647
rect 7538 -1567 7572 -1551
rect 7538 -1663 7572 -1647
rect 7634 -1567 7668 -1551
rect 7634 -1663 7668 -1647
rect 7730 -1567 7764 -1551
rect 7730 -1663 7764 -1647
rect 7826 -1567 7860 -1551
rect 7826 -1663 7860 -1647
rect 7922 -1567 7956 -1551
rect 7922 -1663 7956 -1647
rect 8018 -1567 8052 -1551
rect 8018 -1663 8052 -1647
rect 8114 -1567 8148 -1551
rect 8114 -1663 8148 -1647
rect 7138 -1735 7154 -1701
rect 7188 -1735 7204 -1701
rect 7330 -1735 7346 -1701
rect 7380 -1735 7396 -1701
rect 7522 -1735 7538 -1701
rect 7572 -1735 7588 -1701
rect 7714 -1735 7730 -1701
rect 7764 -1735 7780 -1701
rect 7906 -1735 7922 -1701
rect 7956 -1735 7972 -1701
rect 8098 -1735 8114 -1701
rect 8148 -1735 8164 -1701
rect 7040 -1799 7074 -1737
rect 8228 -1799 8262 -1737
rect 7040 -1833 7136 -1799
rect 8166 -1833 8262 -1799
rect 16040 -1477 16136 -1443
rect 17166 -1477 17262 -1443
rect 16040 -1537 16074 -1477
rect 17228 -1539 17262 -1477
rect 16154 -1567 16188 -1551
rect 16154 -1663 16188 -1647
rect 16250 -1567 16284 -1551
rect 16250 -1663 16284 -1647
rect 16346 -1567 16380 -1551
rect 16346 -1663 16380 -1647
rect 16442 -1567 16476 -1551
rect 16442 -1663 16476 -1647
rect 16538 -1567 16572 -1551
rect 16538 -1663 16572 -1647
rect 16634 -1567 16668 -1551
rect 16634 -1663 16668 -1647
rect 16730 -1567 16764 -1551
rect 16730 -1663 16764 -1647
rect 16826 -1567 16860 -1551
rect 16826 -1663 16860 -1647
rect 16922 -1567 16956 -1551
rect 16922 -1663 16956 -1647
rect 17018 -1567 17052 -1551
rect 17018 -1663 17052 -1647
rect 17114 -1567 17148 -1551
rect 17114 -1663 17148 -1647
rect 16138 -1735 16154 -1701
rect 16188 -1735 16204 -1701
rect 16330 -1735 16346 -1701
rect 16380 -1735 16396 -1701
rect 16522 -1735 16538 -1701
rect 16572 -1735 16588 -1701
rect 16714 -1735 16730 -1701
rect 16764 -1735 16780 -1701
rect 16906 -1735 16922 -1701
rect 16956 -1735 16972 -1701
rect 17098 -1735 17114 -1701
rect 17148 -1735 17164 -1701
rect 16040 -1799 16074 -1737
rect 17228 -1799 17262 -1737
rect 16040 -1833 16136 -1799
rect 17166 -1833 17262 -1799
rect 7040 -2625 7136 -2591
rect 8166 -2625 8262 -2591
rect 7040 -2687 7074 -2625
rect 8228 -2687 8262 -2625
rect 7138 -2727 7154 -2693
rect 7188 -2727 7204 -2693
rect 7330 -2727 7346 -2693
rect 7380 -2727 7396 -2693
rect 7522 -2727 7538 -2693
rect 7572 -2727 7588 -2693
rect 7714 -2727 7730 -2693
rect 7764 -2727 7780 -2693
rect 7906 -2727 7922 -2693
rect 7956 -2727 7972 -2693
rect 8098 -2727 8114 -2693
rect 8148 -2727 8164 -2693
rect 7154 -2787 7188 -2771
rect 7154 -3051 7188 -3035
rect 7250 -2787 7284 -2771
rect 7250 -3051 7284 -3035
rect 7346 -2787 7380 -2771
rect 7346 -3051 7380 -3035
rect 7442 -2787 7476 -2771
rect 7442 -3051 7476 -3035
rect 7538 -2787 7572 -2771
rect 7538 -3051 7572 -3035
rect 7634 -2787 7668 -2771
rect 7634 -3051 7668 -3035
rect 7730 -2787 7764 -2771
rect 7730 -3051 7764 -3035
rect 7826 -2787 7860 -2771
rect 7826 -3051 7860 -3035
rect 7922 -2787 7956 -2771
rect 7922 -3051 7956 -3035
rect 8018 -2787 8052 -2771
rect 8018 -3051 8052 -3035
rect 8114 -2787 8148 -2771
rect 8114 -3051 8148 -3035
rect 7040 -3135 7074 -3073
rect 8228 -3135 8262 -3073
rect 7040 -3169 7136 -3135
rect 8166 -3169 8262 -3135
rect 16040 -2625 16136 -2591
rect 17166 -2625 17262 -2591
rect 16040 -2687 16074 -2625
rect 17228 -2687 17262 -2625
rect 16138 -2727 16154 -2693
rect 16188 -2727 16204 -2693
rect 16330 -2727 16346 -2693
rect 16380 -2727 16396 -2693
rect 16522 -2727 16538 -2693
rect 16572 -2727 16588 -2693
rect 16714 -2727 16730 -2693
rect 16764 -2727 16780 -2693
rect 16906 -2727 16922 -2693
rect 16956 -2727 16972 -2693
rect 17098 -2727 17114 -2693
rect 17148 -2727 17164 -2693
rect 16154 -2787 16188 -2771
rect 16154 -3051 16188 -3035
rect 16250 -2787 16284 -2771
rect 16250 -3051 16284 -3035
rect 16346 -2787 16380 -2771
rect 16346 -3051 16380 -3035
rect 16442 -2787 16476 -2771
rect 16442 -3051 16476 -3035
rect 16538 -2787 16572 -2771
rect 16538 -3051 16572 -3035
rect 16634 -2787 16668 -2771
rect 16634 -3051 16668 -3035
rect 16730 -2787 16764 -2771
rect 16730 -3051 16764 -3035
rect 16826 -2787 16860 -2771
rect 16826 -3051 16860 -3035
rect 16922 -2787 16956 -2771
rect 16922 -3051 16956 -3035
rect 17018 -2787 17052 -2771
rect 17018 -3051 17052 -3035
rect 17114 -2787 17148 -2771
rect 17114 -3051 17148 -3035
rect 16040 -3135 16074 -3073
rect 17228 -3135 17262 -3073
rect 16040 -3169 16136 -3135
rect 17166 -3169 17262 -3135
rect 7040 -3277 7136 -3243
rect 8166 -3277 8262 -3243
rect 7040 -3337 7074 -3277
rect 8228 -3339 8262 -3277
rect 7154 -3367 7188 -3351
rect 7154 -3463 7188 -3447
rect 7250 -3367 7284 -3351
rect 7250 -3463 7284 -3447
rect 7346 -3367 7380 -3351
rect 7346 -3463 7380 -3447
rect 7442 -3367 7476 -3351
rect 7442 -3463 7476 -3447
rect 7538 -3367 7572 -3351
rect 7538 -3463 7572 -3447
rect 7634 -3367 7668 -3351
rect 7634 -3463 7668 -3447
rect 7730 -3367 7764 -3351
rect 7730 -3463 7764 -3447
rect 7826 -3367 7860 -3351
rect 7826 -3463 7860 -3447
rect 7922 -3367 7956 -3351
rect 7922 -3463 7956 -3447
rect 8018 -3367 8052 -3351
rect 8018 -3463 8052 -3447
rect 8114 -3367 8148 -3351
rect 8114 -3463 8148 -3447
rect 7138 -3535 7154 -3501
rect 7188 -3535 7204 -3501
rect 7330 -3535 7346 -3501
rect 7380 -3535 7396 -3501
rect 7522 -3535 7538 -3501
rect 7572 -3535 7588 -3501
rect 7714 -3535 7730 -3501
rect 7764 -3535 7780 -3501
rect 7906 -3535 7922 -3501
rect 7956 -3535 7972 -3501
rect 8098 -3535 8114 -3501
rect 8148 -3535 8164 -3501
rect 7040 -3599 7074 -3537
rect 8228 -3599 8262 -3537
rect 7040 -3633 7136 -3599
rect 8166 -3633 8262 -3599
rect 16040 -3277 16136 -3243
rect 17166 -3277 17262 -3243
rect 16040 -3337 16074 -3277
rect 17228 -3339 17262 -3277
rect 16154 -3367 16188 -3351
rect 16154 -3463 16188 -3447
rect 16250 -3367 16284 -3351
rect 16250 -3463 16284 -3447
rect 16346 -3367 16380 -3351
rect 16346 -3463 16380 -3447
rect 16442 -3367 16476 -3351
rect 16442 -3463 16476 -3447
rect 16538 -3367 16572 -3351
rect 16538 -3463 16572 -3447
rect 16634 -3367 16668 -3351
rect 16634 -3463 16668 -3447
rect 16730 -3367 16764 -3351
rect 16730 -3463 16764 -3447
rect 16826 -3367 16860 -3351
rect 16826 -3463 16860 -3447
rect 16922 -3367 16956 -3351
rect 16922 -3463 16956 -3447
rect 17018 -3367 17052 -3351
rect 17018 -3463 17052 -3447
rect 17114 -3367 17148 -3351
rect 17114 -3463 17148 -3447
rect 16138 -3535 16154 -3501
rect 16188 -3535 16204 -3501
rect 16330 -3535 16346 -3501
rect 16380 -3535 16396 -3501
rect 16522 -3535 16538 -3501
rect 16572 -3535 16588 -3501
rect 16714 -3535 16730 -3501
rect 16764 -3535 16780 -3501
rect 16906 -3535 16922 -3501
rect 16956 -3535 16972 -3501
rect 17098 -3535 17114 -3501
rect 17148 -3535 17164 -3501
rect 16040 -3599 16074 -3537
rect 17228 -3599 17262 -3537
rect 16040 -3633 16136 -3599
rect 17166 -3633 17262 -3599
rect 7040 -4425 7136 -4391
rect 8166 -4425 8262 -4391
rect 7040 -4487 7074 -4425
rect 8228 -4487 8262 -4425
rect 7138 -4527 7154 -4493
rect 7188 -4527 7204 -4493
rect 7330 -4527 7346 -4493
rect 7380 -4527 7396 -4493
rect 7522 -4527 7538 -4493
rect 7572 -4527 7588 -4493
rect 7714 -4527 7730 -4493
rect 7764 -4527 7780 -4493
rect 7906 -4527 7922 -4493
rect 7956 -4527 7972 -4493
rect 8098 -4527 8114 -4493
rect 8148 -4527 8164 -4493
rect 7154 -4587 7188 -4571
rect 7154 -4851 7188 -4835
rect 7250 -4587 7284 -4571
rect 7250 -4851 7284 -4835
rect 7346 -4587 7380 -4571
rect 7346 -4851 7380 -4835
rect 7442 -4587 7476 -4571
rect 7442 -4851 7476 -4835
rect 7538 -4587 7572 -4571
rect 7538 -4851 7572 -4835
rect 7634 -4587 7668 -4571
rect 7634 -4851 7668 -4835
rect 7730 -4587 7764 -4571
rect 7730 -4851 7764 -4835
rect 7826 -4587 7860 -4571
rect 7826 -4851 7860 -4835
rect 7922 -4587 7956 -4571
rect 7922 -4851 7956 -4835
rect 8018 -4587 8052 -4571
rect 8018 -4851 8052 -4835
rect 8114 -4587 8148 -4571
rect 8114 -4851 8148 -4835
rect 7040 -4935 7074 -4873
rect 8228 -4935 8262 -4873
rect 7040 -4969 7136 -4935
rect 8166 -4969 8262 -4935
rect 16040 -4425 16136 -4391
rect 17166 -4425 17262 -4391
rect 16040 -4487 16074 -4425
rect 17228 -4487 17262 -4425
rect 16138 -4527 16154 -4493
rect 16188 -4527 16204 -4493
rect 16330 -4527 16346 -4493
rect 16380 -4527 16396 -4493
rect 16522 -4527 16538 -4493
rect 16572 -4527 16588 -4493
rect 16714 -4527 16730 -4493
rect 16764 -4527 16780 -4493
rect 16906 -4527 16922 -4493
rect 16956 -4527 16972 -4493
rect 17098 -4527 17114 -4493
rect 17148 -4527 17164 -4493
rect 16154 -4587 16188 -4571
rect 16154 -4851 16188 -4835
rect 16250 -4587 16284 -4571
rect 16250 -4851 16284 -4835
rect 16346 -4587 16380 -4571
rect 16346 -4851 16380 -4835
rect 16442 -4587 16476 -4571
rect 16442 -4851 16476 -4835
rect 16538 -4587 16572 -4571
rect 16538 -4851 16572 -4835
rect 16634 -4587 16668 -4571
rect 16634 -4851 16668 -4835
rect 16730 -4587 16764 -4571
rect 16730 -4851 16764 -4835
rect 16826 -4587 16860 -4571
rect 16826 -4851 16860 -4835
rect 16922 -4587 16956 -4571
rect 16922 -4851 16956 -4835
rect 17018 -4587 17052 -4571
rect 17018 -4851 17052 -4835
rect 17114 -4587 17148 -4571
rect 17114 -4851 17148 -4835
rect 16040 -4935 16074 -4873
rect 17228 -4935 17262 -4873
rect 16040 -4969 16136 -4935
rect 17166 -4969 17262 -4935
rect 7040 -5077 7136 -5043
rect 8166 -5077 8262 -5043
rect 7040 -5137 7074 -5077
rect 8228 -5139 8262 -5077
rect 7154 -5167 7188 -5151
rect 7154 -5263 7188 -5247
rect 7250 -5167 7284 -5151
rect 7250 -5263 7284 -5247
rect 7346 -5167 7380 -5151
rect 7346 -5263 7380 -5247
rect 7442 -5167 7476 -5151
rect 7442 -5263 7476 -5247
rect 7538 -5167 7572 -5151
rect 7538 -5263 7572 -5247
rect 7634 -5167 7668 -5151
rect 7634 -5263 7668 -5247
rect 7730 -5167 7764 -5151
rect 7730 -5263 7764 -5247
rect 7826 -5167 7860 -5151
rect 7826 -5263 7860 -5247
rect 7922 -5167 7956 -5151
rect 7922 -5263 7956 -5247
rect 8018 -5167 8052 -5151
rect 8018 -5263 8052 -5247
rect 8114 -5167 8148 -5151
rect 8114 -5263 8148 -5247
rect 7138 -5335 7154 -5301
rect 7188 -5335 7204 -5301
rect 7330 -5335 7346 -5301
rect 7380 -5335 7396 -5301
rect 7522 -5335 7538 -5301
rect 7572 -5335 7588 -5301
rect 7714 -5335 7730 -5301
rect 7764 -5335 7780 -5301
rect 7906 -5335 7922 -5301
rect 7956 -5335 7972 -5301
rect 8098 -5335 8114 -5301
rect 8148 -5335 8164 -5301
rect 7040 -5399 7074 -5337
rect 8228 -5399 8262 -5337
rect 7040 -5433 7136 -5399
rect 8166 -5433 8262 -5399
rect 16040 -5077 16136 -5043
rect 17166 -5077 17262 -5043
rect 16040 -5137 16074 -5077
rect 17228 -5139 17262 -5077
rect 16154 -5167 16188 -5151
rect 16154 -5263 16188 -5247
rect 16250 -5167 16284 -5151
rect 16250 -5263 16284 -5247
rect 16346 -5167 16380 -5151
rect 16346 -5263 16380 -5247
rect 16442 -5167 16476 -5151
rect 16442 -5263 16476 -5247
rect 16538 -5167 16572 -5151
rect 16538 -5263 16572 -5247
rect 16634 -5167 16668 -5151
rect 16634 -5263 16668 -5247
rect 16730 -5167 16764 -5151
rect 16730 -5263 16764 -5247
rect 16826 -5167 16860 -5151
rect 16826 -5263 16860 -5247
rect 16922 -5167 16956 -5151
rect 16922 -5263 16956 -5247
rect 17018 -5167 17052 -5151
rect 17018 -5263 17052 -5247
rect 17114 -5167 17148 -5151
rect 17114 -5263 17148 -5247
rect 16138 -5335 16154 -5301
rect 16188 -5335 16204 -5301
rect 16330 -5335 16346 -5301
rect 16380 -5335 16396 -5301
rect 16522 -5335 16538 -5301
rect 16572 -5335 16588 -5301
rect 16714 -5335 16730 -5301
rect 16764 -5335 16780 -5301
rect 16906 -5335 16922 -5301
rect 16956 -5335 16972 -5301
rect 17098 -5335 17114 -5301
rect 17148 -5335 17164 -5301
rect 16040 -5399 16074 -5337
rect 17228 -5399 17262 -5337
rect 16040 -5433 16136 -5399
rect 17166 -5433 17262 -5399
rect 7040 -6225 7136 -6191
rect 8166 -6225 8262 -6191
rect 7040 -6287 7074 -6225
rect 8228 -6287 8262 -6225
rect 7138 -6327 7154 -6293
rect 7188 -6327 7204 -6293
rect 7330 -6327 7346 -6293
rect 7380 -6327 7396 -6293
rect 7522 -6327 7538 -6293
rect 7572 -6327 7588 -6293
rect 7714 -6327 7730 -6293
rect 7764 -6327 7780 -6293
rect 7906 -6327 7922 -6293
rect 7956 -6327 7972 -6293
rect 8098 -6327 8114 -6293
rect 8148 -6327 8164 -6293
rect 7154 -6387 7188 -6371
rect 7154 -6651 7188 -6635
rect 7250 -6387 7284 -6371
rect 7250 -6651 7284 -6635
rect 7346 -6387 7380 -6371
rect 7346 -6651 7380 -6635
rect 7442 -6387 7476 -6371
rect 7442 -6651 7476 -6635
rect 7538 -6387 7572 -6371
rect 7538 -6651 7572 -6635
rect 7634 -6387 7668 -6371
rect 7634 -6651 7668 -6635
rect 7730 -6387 7764 -6371
rect 7730 -6651 7764 -6635
rect 7826 -6387 7860 -6371
rect 7826 -6651 7860 -6635
rect 7922 -6387 7956 -6371
rect 7922 -6651 7956 -6635
rect 8018 -6387 8052 -6371
rect 8018 -6651 8052 -6635
rect 8114 -6387 8148 -6371
rect 8114 -6651 8148 -6635
rect 7040 -6735 7074 -6673
rect 8228 -6735 8262 -6673
rect 7040 -6769 7136 -6735
rect 8166 -6769 8262 -6735
rect 16040 -6225 16136 -6191
rect 17166 -6225 17262 -6191
rect 16040 -6287 16074 -6225
rect 17228 -6287 17262 -6225
rect 16138 -6327 16154 -6293
rect 16188 -6327 16204 -6293
rect 16330 -6327 16346 -6293
rect 16380 -6327 16396 -6293
rect 16522 -6327 16538 -6293
rect 16572 -6327 16588 -6293
rect 16714 -6327 16730 -6293
rect 16764 -6327 16780 -6293
rect 16906 -6327 16922 -6293
rect 16956 -6327 16972 -6293
rect 17098 -6327 17114 -6293
rect 17148 -6327 17164 -6293
rect 16154 -6387 16188 -6371
rect 16154 -6651 16188 -6635
rect 16250 -6387 16284 -6371
rect 16250 -6651 16284 -6635
rect 16346 -6387 16380 -6371
rect 16346 -6651 16380 -6635
rect 16442 -6387 16476 -6371
rect 16442 -6651 16476 -6635
rect 16538 -6387 16572 -6371
rect 16538 -6651 16572 -6635
rect 16634 -6387 16668 -6371
rect 16634 -6651 16668 -6635
rect 16730 -6387 16764 -6371
rect 16730 -6651 16764 -6635
rect 16826 -6387 16860 -6371
rect 16826 -6651 16860 -6635
rect 16922 -6387 16956 -6371
rect 16922 -6651 16956 -6635
rect 17018 -6387 17052 -6371
rect 17018 -6651 17052 -6635
rect 17114 -6387 17148 -6371
rect 17114 -6651 17148 -6635
rect 16040 -6735 16074 -6673
rect 17228 -6735 17262 -6673
rect 16040 -6769 16136 -6735
rect 17166 -6769 17262 -6735
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
rect 7040 -6877 7136 -6843
rect 8166 -6877 8262 -6843
rect 7040 -6937 7074 -6877
rect 8228 -6939 8262 -6877
rect 7154 -6967 7188 -6951
rect 7154 -7063 7188 -7047
rect 7250 -6967 7284 -6951
rect 7250 -7063 7284 -7047
rect 7346 -6967 7380 -6951
rect 7346 -7063 7380 -7047
rect 7442 -6967 7476 -6951
rect 7442 -7063 7476 -7047
rect 7538 -6967 7572 -6951
rect 7538 -7063 7572 -7047
rect 7634 -6967 7668 -6951
rect 7634 -7063 7668 -7047
rect 7730 -6967 7764 -6951
rect 7730 -7063 7764 -7047
rect 7826 -6967 7860 -6951
rect 7826 -7063 7860 -7047
rect 7922 -6967 7956 -6951
rect 7922 -7063 7956 -7047
rect 8018 -6967 8052 -6951
rect 8018 -7063 8052 -7047
rect 8114 -6967 8148 -6951
rect 8114 -7063 8148 -7047
rect 7138 -7135 7154 -7101
rect 7188 -7135 7204 -7101
rect 7330 -7135 7346 -7101
rect 7380 -7135 7396 -7101
rect 7522 -7135 7538 -7101
rect 7572 -7135 7588 -7101
rect 7714 -7135 7730 -7101
rect 7764 -7135 7780 -7101
rect 7906 -7135 7922 -7101
rect 7956 -7135 7972 -7101
rect 8098 -7135 8114 -7101
rect 8148 -7135 8164 -7101
rect 7040 -7199 7074 -7137
rect 8228 -7199 8262 -7137
rect 7040 -7233 7136 -7199
rect 8166 -7233 8262 -7199
rect 16040 -6877 16136 -6843
rect 17166 -6877 17262 -6843
rect 16040 -6937 16074 -6877
rect 17228 -6939 17262 -6877
rect 16154 -6967 16188 -6951
rect 16154 -7063 16188 -7047
rect 16250 -6967 16284 -6951
rect 16250 -7063 16284 -7047
rect 16346 -6967 16380 -6951
rect 16346 -7063 16380 -7047
rect 16442 -6967 16476 -6951
rect 16442 -7063 16476 -7047
rect 16538 -6967 16572 -6951
rect 16538 -7063 16572 -7047
rect 16634 -6967 16668 -6951
rect 16634 -7063 16668 -7047
rect 16730 -6967 16764 -6951
rect 16730 -7063 16764 -7047
rect 16826 -6967 16860 -6951
rect 16826 -7063 16860 -7047
rect 16922 -6967 16956 -6951
rect 16922 -7063 16956 -7047
rect 17018 -6967 17052 -6951
rect 17018 -7063 17052 -7047
rect 17114 -6967 17148 -6951
rect 17114 -7063 17148 -7047
rect 16138 -7135 16154 -7101
rect 16188 -7135 16204 -7101
rect 16330 -7135 16346 -7101
rect 16380 -7135 16396 -7101
rect 16522 -7135 16538 -7101
rect 16572 -7135 16588 -7101
rect 16714 -7135 16730 -7101
rect 16764 -7135 16780 -7101
rect 16906 -7135 16922 -7101
rect 16956 -7135 16972 -7101
rect 17098 -7135 17114 -7101
rect 17148 -7135 17164 -7101
rect 16040 -7199 16074 -7137
rect 17228 -7199 17262 -7137
rect 16040 -7233 16136 -7199
rect 17166 -7233 17262 -7199
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect 13619 -7731 13719 -7621
rect -5560 -7824 -5544 -7790
rect -5500 -7824 -5484 -7790
rect -5382 -7824 -5366 -7790
rect -5322 -7824 -5306 -7790
rect -5204 -7824 -5188 -7790
rect -5144 -7824 -5128 -7790
rect -5026 -7824 -5010 -7790
rect -4966 -7824 -4950 -7790
rect -4848 -7824 -4832 -7790
rect -4788 -7824 -4772 -7790
rect -4670 -7824 -4654 -7790
rect -4610 -7824 -4594 -7790
rect -4492 -7824 -4476 -7790
rect -4432 -7824 -4416 -7790
rect -4314 -7824 -4298 -7790
rect -4254 -7824 -4238 -7790
rect -4136 -7824 -4120 -7790
rect -4076 -7824 -4060 -7790
rect -5628 -7874 -5594 -7858
rect -5628 -8146 -5594 -8130
rect -5450 -7874 -5416 -7858
rect -5450 -8146 -5416 -8130
rect -5272 -7874 -5238 -7858
rect -5272 -8146 -5238 -8130
rect -5094 -7874 -5060 -7858
rect -5094 -8146 -5060 -8130
rect -4916 -7874 -4882 -7858
rect -4916 -8146 -4882 -8130
rect -4738 -7874 -4704 -7858
rect -4738 -8146 -4704 -8130
rect -4560 -7874 -4526 -7858
rect -4560 -8146 -4526 -8130
rect -4382 -7874 -4348 -7858
rect -4382 -8146 -4348 -8130
rect -4204 -7874 -4170 -7858
rect -4204 -8146 -4170 -8130
rect -4026 -7874 -3992 -7858
rect -2105 -8082 -2089 -8048
rect -2045 -8082 -2029 -8048
rect -1927 -8082 -1911 -8048
rect -1867 -8082 -1851 -8048
rect -1749 -8082 -1733 -8048
rect -1689 -8082 -1673 -8048
rect -1571 -8082 -1555 -8048
rect -1511 -8082 -1495 -8048
rect -1393 -8082 -1377 -8048
rect -1333 -8082 -1317 -8048
rect -1215 -8082 -1199 -8048
rect -1155 -8082 -1139 -8048
rect -1037 -8082 -1021 -8048
rect -977 -8082 -961 -8048
rect -859 -8082 -843 -8048
rect -799 -8082 -783 -8048
rect -681 -8082 -665 -8048
rect -621 -8082 -605 -8048
rect -503 -8082 -487 -8048
rect -443 -8082 -427 -8048
rect -325 -8082 -309 -8048
rect -265 -8082 -249 -8048
rect -147 -8082 -131 -8048
rect -87 -8082 -71 -8048
rect 31 -8082 47 -8048
rect 91 -8082 107 -8048
rect 209 -8082 225 -8048
rect 269 -8082 285 -8048
rect 387 -8082 403 -8048
rect 447 -8082 463 -8048
rect 565 -8082 581 -8048
rect 625 -8082 641 -8048
rect 743 -8082 759 -8048
rect 803 -8082 819 -8048
rect 921 -8082 937 -8048
rect 981 -8082 997 -8048
rect 1099 -8082 1115 -8048
rect 1159 -8082 1175 -8048
rect 1277 -8082 1293 -8048
rect 1337 -8082 1353 -8048
rect 1455 -8082 1471 -8048
rect 1515 -8082 1531 -8048
rect 1633 -8082 1649 -8048
rect 1693 -8082 1709 -8048
rect 1811 -8082 1827 -8048
rect 1871 -8082 1887 -8048
rect 1989 -8082 2005 -8048
rect 2049 -8082 2065 -8048
rect 2167 -8082 2183 -8048
rect 2227 -8082 2243 -8048
rect 2345 -8082 2361 -8048
rect 2405 -8082 2421 -8048
rect 2523 -8082 2539 -8048
rect 2583 -8082 2599 -8048
rect 2701 -8082 2717 -8048
rect 2761 -8082 2777 -8048
rect 2879 -8082 2895 -8048
rect 2939 -8082 2955 -8048
rect 3057 -8082 3073 -8048
rect 3117 -8082 3133 -8048
rect 3235 -8082 3251 -8048
rect 3295 -8082 3311 -8048
rect 3413 -8082 3429 -8048
rect 3473 -8082 3489 -8048
rect 3591 -8082 3607 -8048
rect 3651 -8082 3667 -8048
rect 3769 -8082 3785 -8048
rect 3829 -8082 3845 -8048
rect 3947 -8082 3963 -8048
rect 4007 -8082 4023 -8048
rect -4026 -8146 -3992 -8130
rect -2173 -8132 -2139 -8116
rect -5560 -8214 -5544 -8180
rect -5500 -8214 -5484 -8180
rect -5382 -8214 -5366 -8180
rect -5322 -8214 -5306 -8180
rect -5204 -8214 -5188 -8180
rect -5144 -8214 -5128 -8180
rect -5026 -8214 -5010 -8180
rect -4966 -8214 -4950 -8180
rect -4848 -8214 -4832 -8180
rect -4788 -8214 -4772 -8180
rect -4670 -8214 -4654 -8180
rect -4610 -8214 -4594 -8180
rect -4492 -8214 -4476 -8180
rect -4432 -8214 -4416 -8180
rect -4314 -8214 -4298 -8180
rect -4254 -8214 -4238 -8180
rect -4136 -8214 -4120 -8180
rect -4076 -8214 -4060 -8180
rect -5560 -8374 -5544 -8340
rect -5500 -8374 -5484 -8340
rect -5382 -8374 -5366 -8340
rect -5322 -8374 -5306 -8340
rect -5204 -8374 -5188 -8340
rect -5144 -8374 -5128 -8340
rect -5026 -8374 -5010 -8340
rect -4966 -8374 -4950 -8340
rect -4848 -8374 -4832 -8340
rect -4788 -8374 -4772 -8340
rect -4670 -8374 -4654 -8340
rect -4610 -8374 -4594 -8340
rect -4492 -8374 -4476 -8340
rect -4432 -8374 -4416 -8340
rect -4314 -8374 -4298 -8340
rect -4254 -8374 -4238 -8340
rect -4136 -8374 -4120 -8340
rect -4076 -8374 -4060 -8340
rect -2173 -8404 -2139 -8388
rect -1995 -8132 -1961 -8116
rect -1995 -8404 -1961 -8388
rect -1817 -8132 -1783 -8116
rect -1817 -8404 -1783 -8388
rect -1639 -8132 -1605 -8116
rect -1639 -8404 -1605 -8388
rect -1461 -8132 -1427 -8116
rect -1461 -8404 -1427 -8388
rect -1283 -8132 -1249 -8116
rect -1283 -8404 -1249 -8388
rect -1105 -8132 -1071 -8116
rect -1105 -8404 -1071 -8388
rect -927 -8132 -893 -8116
rect -927 -8404 -893 -8388
rect -749 -8132 -715 -8116
rect -749 -8404 -715 -8388
rect -571 -8132 -537 -8116
rect -571 -8404 -537 -8388
rect -393 -8132 -359 -8116
rect -393 -8404 -359 -8388
rect -215 -8132 -181 -8116
rect -215 -8404 -181 -8388
rect -37 -8132 -3 -8116
rect -37 -8404 -3 -8388
rect 141 -8132 175 -8116
rect 141 -8404 175 -8388
rect 319 -8132 353 -8116
rect 319 -8404 353 -8388
rect 497 -8132 531 -8116
rect 497 -8404 531 -8388
rect 675 -8132 709 -8116
rect 675 -8404 709 -8388
rect 853 -8132 887 -8116
rect 853 -8404 887 -8388
rect 1031 -8132 1065 -8116
rect 1031 -8404 1065 -8388
rect 1209 -8132 1243 -8116
rect 1209 -8404 1243 -8388
rect 1387 -8132 1421 -8116
rect 1387 -8404 1421 -8388
rect 1565 -8132 1599 -8116
rect 1565 -8404 1599 -8388
rect 1743 -8132 1777 -8116
rect 1743 -8404 1777 -8388
rect 1921 -8132 1955 -8116
rect 1921 -8404 1955 -8388
rect 2099 -8132 2133 -8116
rect 2099 -8404 2133 -8388
rect 2277 -8132 2311 -8116
rect 2277 -8404 2311 -8388
rect 2455 -8132 2489 -8116
rect 2455 -8404 2489 -8388
rect 2633 -8132 2667 -8116
rect 2633 -8404 2667 -8388
rect 2811 -8132 2845 -8116
rect 2811 -8404 2845 -8388
rect 2989 -8132 3023 -8116
rect 2989 -8404 3023 -8388
rect 3167 -8132 3201 -8116
rect 3167 -8404 3201 -8388
rect 3345 -8132 3379 -8116
rect 3345 -8404 3379 -8388
rect 3523 -8132 3557 -8116
rect 3523 -8404 3557 -8388
rect 3701 -8132 3735 -8116
rect 3701 -8404 3735 -8388
rect 3879 -8132 3913 -8116
rect 3879 -8404 3913 -8388
rect 4057 -8132 4091 -8116
rect 4057 -8404 4091 -8388
rect -5628 -8424 -5594 -8408
rect -5628 -8696 -5594 -8680
rect -5450 -8424 -5416 -8408
rect -5450 -8696 -5416 -8680
rect -5272 -8424 -5238 -8408
rect -5272 -8696 -5238 -8680
rect -5094 -8424 -5060 -8408
rect -5094 -8696 -5060 -8680
rect -4916 -8424 -4882 -8408
rect -4916 -8696 -4882 -8680
rect -4738 -8424 -4704 -8408
rect -4738 -8696 -4704 -8680
rect -4560 -8424 -4526 -8408
rect -4560 -8696 -4526 -8680
rect -4382 -8424 -4348 -8408
rect -4382 -8696 -4348 -8680
rect -4204 -8424 -4170 -8408
rect -4204 -8696 -4170 -8680
rect -4026 -8424 -3992 -8408
rect -2105 -8472 -2089 -8438
rect -2045 -8472 -2029 -8438
rect -1927 -8472 -1911 -8438
rect -1867 -8472 -1851 -8438
rect -1749 -8472 -1733 -8438
rect -1689 -8472 -1673 -8438
rect -1571 -8472 -1555 -8438
rect -1511 -8472 -1495 -8438
rect -1393 -8472 -1377 -8438
rect -1333 -8472 -1317 -8438
rect -1215 -8472 -1199 -8438
rect -1155 -8472 -1139 -8438
rect -1037 -8472 -1021 -8438
rect -977 -8472 -961 -8438
rect -859 -8472 -843 -8438
rect -799 -8472 -783 -8438
rect -681 -8472 -665 -8438
rect -621 -8472 -605 -8438
rect -503 -8472 -487 -8438
rect -443 -8472 -427 -8438
rect -325 -8472 -309 -8438
rect -265 -8472 -249 -8438
rect -147 -8472 -131 -8438
rect -87 -8472 -71 -8438
rect 31 -8472 47 -8438
rect 91 -8472 107 -8438
rect 209 -8472 225 -8438
rect 269 -8472 285 -8438
rect 387 -8472 403 -8438
rect 447 -8472 463 -8438
rect 565 -8472 581 -8438
rect 625 -8472 641 -8438
rect 743 -8472 759 -8438
rect 803 -8472 819 -8438
rect 921 -8472 937 -8438
rect 981 -8472 997 -8438
rect 1099 -8472 1115 -8438
rect 1159 -8472 1175 -8438
rect 1277 -8472 1293 -8438
rect 1337 -8472 1353 -8438
rect 1455 -8472 1471 -8438
rect 1515 -8472 1531 -8438
rect 1633 -8472 1649 -8438
rect 1693 -8472 1709 -8438
rect 1811 -8472 1827 -8438
rect 1871 -8472 1887 -8438
rect 1989 -8472 2005 -8438
rect 2049 -8472 2065 -8438
rect 2167 -8472 2183 -8438
rect 2227 -8472 2243 -8438
rect 2345 -8472 2361 -8438
rect 2405 -8472 2421 -8438
rect 2523 -8472 2539 -8438
rect 2583 -8472 2599 -8438
rect 2701 -8472 2717 -8438
rect 2761 -8472 2777 -8438
rect 2879 -8472 2895 -8438
rect 2939 -8472 2955 -8438
rect 3057 -8472 3073 -8438
rect 3117 -8472 3133 -8438
rect 3235 -8472 3251 -8438
rect 3295 -8472 3311 -8438
rect 3413 -8472 3429 -8438
rect 3473 -8472 3489 -8438
rect 3591 -8472 3607 -8438
rect 3651 -8472 3667 -8438
rect 3769 -8472 3785 -8438
rect 3829 -8472 3845 -8438
rect 3947 -8472 3963 -8438
rect 4007 -8472 4023 -8438
rect -4026 -8696 -3992 -8680
rect -5560 -8764 -5544 -8730
rect -5500 -8764 -5484 -8730
rect -5382 -8764 -5366 -8730
rect -5322 -8764 -5306 -8730
rect -5204 -8764 -5188 -8730
rect -5144 -8764 -5128 -8730
rect -5026 -8764 -5010 -8730
rect -4966 -8764 -4950 -8730
rect -4848 -8764 -4832 -8730
rect -4788 -8764 -4772 -8730
rect -4670 -8764 -4654 -8730
rect -4610 -8764 -4594 -8730
rect -4492 -8764 -4476 -8730
rect -4432 -8764 -4416 -8730
rect -4314 -8764 -4298 -8730
rect -4254 -8764 -4238 -8730
rect -4136 -8764 -4120 -8730
rect -4076 -8764 -4060 -8730
rect 6580 -8844 6596 -8810
rect 6640 -8844 6656 -8810
rect 6758 -8844 6774 -8810
rect 6818 -8844 6834 -8810
rect 6936 -8844 6952 -8810
rect 6996 -8844 7012 -8810
rect 7114 -8844 7130 -8810
rect 7174 -8844 7190 -8810
rect 7292 -8844 7308 -8810
rect 7352 -8844 7368 -8810
rect 7470 -8844 7486 -8810
rect 7530 -8844 7546 -8810
rect 7648 -8844 7664 -8810
rect 7708 -8844 7724 -8810
rect 7826 -8844 7842 -8810
rect 7886 -8844 7902 -8810
rect 8004 -8844 8020 -8810
rect 8064 -8844 8080 -8810
rect 8182 -8844 8198 -8810
rect 8242 -8844 8258 -8810
rect 8360 -8844 8376 -8810
rect 8420 -8844 8436 -8810
rect 8538 -8844 8554 -8810
rect 8598 -8844 8614 -8810
rect 8716 -8844 8732 -8810
rect 8776 -8844 8792 -8810
rect 8894 -8844 8910 -8810
rect 8954 -8844 8970 -8810
rect 9072 -8844 9088 -8810
rect 9132 -8844 9148 -8810
rect 9250 -8844 9266 -8810
rect 9310 -8844 9326 -8810
rect 10840 -8874 10856 -8840
rect 10900 -8874 10916 -8840
rect 11132 -8874 11148 -8840
rect 11192 -8874 11208 -8840
rect 11424 -8874 11440 -8840
rect 11484 -8874 11500 -8840
rect 11716 -8874 11732 -8840
rect 11776 -8874 11792 -8840
rect 12008 -8874 12024 -8840
rect 12068 -8874 12084 -8840
rect 12300 -8874 12316 -8840
rect 12360 -8874 12376 -8840
rect 12592 -8874 12608 -8840
rect 12652 -8874 12668 -8840
rect -5560 -8924 -5544 -8890
rect -5500 -8924 -5484 -8890
rect -5382 -8924 -5366 -8890
rect -5322 -8924 -5306 -8890
rect -5204 -8924 -5188 -8890
rect -5144 -8924 -5128 -8890
rect -5026 -8924 -5010 -8890
rect -4966 -8924 -4950 -8890
rect -4848 -8924 -4832 -8890
rect -4788 -8924 -4772 -8890
rect -4670 -8924 -4654 -8890
rect -4610 -8924 -4594 -8890
rect -4492 -8924 -4476 -8890
rect -4432 -8924 -4416 -8890
rect -4314 -8924 -4298 -8890
rect -4254 -8924 -4238 -8890
rect -4136 -8924 -4120 -8890
rect -4076 -8924 -4060 -8890
rect 6512 -8894 6546 -8878
rect -5628 -8974 -5594 -8958
rect -5628 -9246 -5594 -9230
rect -5450 -8974 -5416 -8958
rect -5450 -9246 -5416 -9230
rect -5272 -8974 -5238 -8958
rect -5272 -9246 -5238 -9230
rect -5094 -8974 -5060 -8958
rect -5094 -9246 -5060 -9230
rect -4916 -8974 -4882 -8958
rect -4916 -9246 -4882 -9230
rect -4738 -8974 -4704 -8958
rect -4738 -9246 -4704 -9230
rect -4560 -8974 -4526 -8958
rect -4560 -9246 -4526 -9230
rect -4382 -8974 -4348 -8958
rect -4382 -9246 -4348 -9230
rect -4204 -8974 -4170 -8958
rect -4204 -9246 -4170 -9230
rect -4026 -8974 -3992 -8958
rect -2105 -9082 -2089 -9048
rect -2045 -9082 -2029 -9048
rect -1927 -9082 -1911 -9048
rect -1867 -9082 -1851 -9048
rect -1749 -9082 -1733 -9048
rect -1689 -9082 -1673 -9048
rect -1571 -9082 -1555 -9048
rect -1511 -9082 -1495 -9048
rect -1393 -9082 -1377 -9048
rect -1333 -9082 -1317 -9048
rect -1215 -9082 -1199 -9048
rect -1155 -9082 -1139 -9048
rect -1037 -9082 -1021 -9048
rect -977 -9082 -961 -9048
rect -859 -9082 -843 -9048
rect -799 -9082 -783 -9048
rect -681 -9082 -665 -9048
rect -621 -9082 -605 -9048
rect -503 -9082 -487 -9048
rect -443 -9082 -427 -9048
rect -325 -9082 -309 -9048
rect -265 -9082 -249 -9048
rect -147 -9082 -131 -9048
rect -87 -9082 -71 -9048
rect 31 -9082 47 -9048
rect 91 -9082 107 -9048
rect 209 -9082 225 -9048
rect 269 -9082 285 -9048
rect 387 -9082 403 -9048
rect 447 -9082 463 -9048
rect 565 -9082 581 -9048
rect 625 -9082 641 -9048
rect 743 -9082 759 -9048
rect 803 -9082 819 -9048
rect 921 -9082 937 -9048
rect 981 -9082 997 -9048
rect 1099 -9082 1115 -9048
rect 1159 -9082 1175 -9048
rect 1277 -9082 1293 -9048
rect 1337 -9082 1353 -9048
rect 1455 -9082 1471 -9048
rect 1515 -9082 1531 -9048
rect 1633 -9082 1649 -9048
rect 1693 -9082 1709 -9048
rect 1811 -9082 1827 -9048
rect 1871 -9082 1887 -9048
rect 1989 -9082 2005 -9048
rect 2049 -9082 2065 -9048
rect 2167 -9082 2183 -9048
rect 2227 -9082 2243 -9048
rect 2345 -9082 2361 -9048
rect 2405 -9082 2421 -9048
rect 2523 -9082 2539 -9048
rect 2583 -9082 2599 -9048
rect 2701 -9082 2717 -9048
rect 2761 -9082 2777 -9048
rect 2879 -9082 2895 -9048
rect 2939 -9082 2955 -9048
rect 3057 -9082 3073 -9048
rect 3117 -9082 3133 -9048
rect 3235 -9082 3251 -9048
rect 3295 -9082 3311 -9048
rect 3413 -9082 3429 -9048
rect 3473 -9082 3489 -9048
rect 3591 -9082 3607 -9048
rect 3651 -9082 3667 -9048
rect 3769 -9082 3785 -9048
rect 3829 -9082 3845 -9048
rect 3947 -9082 3963 -9048
rect 4007 -9082 4023 -9048
rect -4026 -9246 -3992 -9230
rect -2173 -9132 -2139 -9116
rect -3009 -9276 -2783 -9252
rect -5560 -9314 -5544 -9280
rect -5500 -9314 -5484 -9280
rect -5382 -9314 -5366 -9280
rect -5322 -9314 -5306 -9280
rect -5204 -9314 -5188 -9280
rect -5144 -9314 -5128 -9280
rect -5026 -9314 -5010 -9280
rect -4966 -9314 -4950 -9280
rect -4848 -9314 -4832 -9280
rect -4788 -9314 -4772 -9280
rect -4670 -9314 -4654 -9280
rect -4610 -9314 -4594 -9280
rect -4492 -9314 -4476 -9280
rect -4432 -9314 -4416 -9280
rect -4314 -9314 -4298 -9280
rect -4254 -9314 -4238 -9280
rect -4136 -9314 -4120 -9280
rect -4076 -9314 -4060 -9280
rect -5560 -9474 -5544 -9440
rect -5500 -9474 -5484 -9440
rect -5382 -9474 -5366 -9440
rect -5322 -9474 -5306 -9440
rect -5204 -9474 -5188 -9440
rect -5144 -9474 -5128 -9440
rect -5026 -9474 -5010 -9440
rect -4966 -9474 -4950 -9440
rect -4848 -9474 -4832 -9440
rect -4788 -9474 -4772 -9440
rect -4670 -9474 -4654 -9440
rect -4610 -9474 -4594 -9440
rect -4492 -9474 -4476 -9440
rect -4432 -9474 -4416 -9440
rect -4314 -9474 -4298 -9440
rect -4254 -9474 -4238 -9440
rect -4136 -9474 -4120 -9440
rect -4076 -9474 -4060 -9440
rect -3009 -9454 -2985 -9276
rect -2807 -9454 -2783 -9276
rect -2173 -9404 -2139 -9388
rect -1995 -9132 -1961 -9116
rect -1995 -9404 -1961 -9388
rect -1817 -9132 -1783 -9116
rect -1817 -9404 -1783 -9388
rect -1639 -9132 -1605 -9116
rect -1639 -9404 -1605 -9388
rect -1461 -9132 -1427 -9116
rect -1461 -9404 -1427 -9388
rect -1283 -9132 -1249 -9116
rect -1283 -9404 -1249 -9388
rect -1105 -9132 -1071 -9116
rect -1105 -9404 -1071 -9388
rect -927 -9132 -893 -9116
rect -927 -9404 -893 -9388
rect -749 -9132 -715 -9116
rect -749 -9404 -715 -9388
rect -571 -9132 -537 -9116
rect -571 -9404 -537 -9388
rect -393 -9132 -359 -9116
rect -393 -9404 -359 -9388
rect -215 -9132 -181 -9116
rect -215 -9404 -181 -9388
rect -37 -9132 -3 -9116
rect -37 -9404 -3 -9388
rect 141 -9132 175 -9116
rect 141 -9404 175 -9388
rect 319 -9132 353 -9116
rect 319 -9404 353 -9388
rect 497 -9132 531 -9116
rect 497 -9404 531 -9388
rect 675 -9132 709 -9116
rect 675 -9404 709 -9388
rect 853 -9132 887 -9116
rect 853 -9404 887 -9388
rect 1031 -9132 1065 -9116
rect 1031 -9404 1065 -9388
rect 1209 -9132 1243 -9116
rect 1209 -9404 1243 -9388
rect 1387 -9132 1421 -9116
rect 1387 -9404 1421 -9388
rect 1565 -9132 1599 -9116
rect 1565 -9404 1599 -9388
rect 1743 -9132 1777 -9116
rect 1743 -9404 1777 -9388
rect 1921 -9132 1955 -9116
rect 1921 -9404 1955 -9388
rect 2099 -9132 2133 -9116
rect 2099 -9404 2133 -9388
rect 2277 -9132 2311 -9116
rect 2277 -9404 2311 -9388
rect 2455 -9132 2489 -9116
rect 2455 -9404 2489 -9388
rect 2633 -9132 2667 -9116
rect 2633 -9404 2667 -9388
rect 2811 -9132 2845 -9116
rect 2811 -9404 2845 -9388
rect 2989 -9132 3023 -9116
rect 2989 -9404 3023 -9388
rect 3167 -9132 3201 -9116
rect 3167 -9404 3201 -9388
rect 3345 -9132 3379 -9116
rect 3345 -9404 3379 -9388
rect 3523 -9132 3557 -9116
rect 3523 -9404 3557 -9388
rect 3701 -9132 3735 -9116
rect 3701 -9404 3735 -9388
rect 3879 -9132 3913 -9116
rect 3879 -9404 3913 -9388
rect 4057 -9132 4091 -9116
rect 6512 -9166 6546 -9150
rect 6690 -8894 6724 -8878
rect 6690 -9166 6724 -9150
rect 6868 -8894 6902 -8878
rect 6868 -9166 6902 -9150
rect 7046 -8894 7080 -8878
rect 7046 -9166 7080 -9150
rect 7224 -8894 7258 -8878
rect 7224 -9166 7258 -9150
rect 7402 -8894 7436 -8878
rect 7402 -9166 7436 -9150
rect 7580 -8894 7614 -8878
rect 7580 -9166 7614 -9150
rect 7758 -8894 7792 -8878
rect 7758 -9166 7792 -9150
rect 7936 -8894 7970 -8878
rect 7936 -9166 7970 -9150
rect 8114 -8894 8148 -8878
rect 8114 -9166 8148 -9150
rect 8292 -8894 8326 -8878
rect 8292 -9166 8326 -9150
rect 8470 -8894 8504 -8878
rect 8470 -9166 8504 -9150
rect 8648 -8894 8682 -8878
rect 8648 -9166 8682 -9150
rect 8826 -8894 8860 -8878
rect 8826 -9166 8860 -9150
rect 9004 -8894 9038 -8878
rect 9004 -9166 9038 -9150
rect 9182 -8894 9216 -8878
rect 9182 -9166 9216 -9150
rect 9360 -8894 9394 -8878
rect 9360 -9166 9394 -9150
rect 10772 -8924 10806 -8908
rect 9958 -9191 10184 -9167
rect 6580 -9234 6596 -9200
rect 6640 -9234 6656 -9200
rect 6758 -9234 6774 -9200
rect 6818 -9234 6834 -9200
rect 6936 -9234 6952 -9200
rect 6996 -9234 7012 -9200
rect 7114 -9234 7130 -9200
rect 7174 -9234 7190 -9200
rect 7292 -9234 7308 -9200
rect 7352 -9234 7368 -9200
rect 7470 -9234 7486 -9200
rect 7530 -9234 7546 -9200
rect 7648 -9234 7664 -9200
rect 7708 -9234 7724 -9200
rect 7826 -9234 7842 -9200
rect 7886 -9234 7902 -9200
rect 8004 -9234 8020 -9200
rect 8064 -9234 8080 -9200
rect 8182 -9234 8198 -9200
rect 8242 -9234 8258 -9200
rect 8360 -9234 8376 -9200
rect 8420 -9234 8436 -9200
rect 8538 -9234 8554 -9200
rect 8598 -9234 8614 -9200
rect 8716 -9234 8732 -9200
rect 8776 -9234 8792 -9200
rect 8894 -9234 8910 -9200
rect 8954 -9234 8970 -9200
rect 9072 -9234 9088 -9200
rect 9132 -9234 9148 -9200
rect 9250 -9234 9266 -9200
rect 9310 -9234 9326 -9200
rect 4057 -9404 4091 -9388
rect 9958 -9369 9982 -9191
rect 10160 -9369 10184 -9191
rect 10772 -9196 10806 -9180
rect 10950 -8924 10984 -8908
rect 10950 -9196 10984 -9180
rect 11064 -8924 11098 -8908
rect 11064 -9196 11098 -9180
rect 11242 -8924 11276 -8908
rect 11242 -9196 11276 -9180
rect 11356 -8924 11390 -8908
rect 11356 -9196 11390 -9180
rect 11534 -8924 11568 -8908
rect 11534 -9196 11568 -9180
rect 11648 -8924 11682 -8908
rect 11648 -9196 11682 -9180
rect 11826 -8924 11860 -8908
rect 11826 -9196 11860 -9180
rect 11940 -8924 11974 -8908
rect 11940 -9196 11974 -9180
rect 12118 -8924 12152 -8908
rect 12118 -9196 12152 -9180
rect 12232 -8924 12266 -8908
rect 12232 -9196 12266 -9180
rect 12410 -8924 12444 -8908
rect 12410 -9196 12444 -9180
rect 12524 -8924 12558 -8908
rect 12524 -9196 12558 -9180
rect 12702 -8924 12736 -8908
rect 12702 -9196 12736 -9180
rect 10840 -9264 10856 -9230
rect 10900 -9264 10916 -9230
rect 11132 -9264 11148 -9230
rect 11192 -9264 11208 -9230
rect 11424 -9264 11440 -9230
rect 11484 -9264 11500 -9230
rect 11716 -9264 11732 -9230
rect 11776 -9264 11792 -9230
rect 12008 -9264 12024 -9230
rect 12068 -9264 12084 -9230
rect 12300 -9264 12316 -9230
rect 12360 -9264 12376 -9230
rect 12592 -9264 12608 -9230
rect 12652 -9264 12668 -9230
rect 9958 -9393 10184 -9369
rect -3009 -9478 -2783 -9454
rect -2105 -9472 -2089 -9438
rect -2045 -9472 -2029 -9438
rect -1927 -9472 -1911 -9438
rect -1867 -9472 -1851 -9438
rect -1749 -9472 -1733 -9438
rect -1689 -9472 -1673 -9438
rect -1571 -9472 -1555 -9438
rect -1511 -9472 -1495 -9438
rect -1393 -9472 -1377 -9438
rect -1333 -9472 -1317 -9438
rect -1215 -9472 -1199 -9438
rect -1155 -9472 -1139 -9438
rect -1037 -9472 -1021 -9438
rect -977 -9472 -961 -9438
rect -859 -9472 -843 -9438
rect -799 -9472 -783 -9438
rect -681 -9472 -665 -9438
rect -621 -9472 -605 -9438
rect -503 -9472 -487 -9438
rect -443 -9472 -427 -9438
rect -325 -9472 -309 -9438
rect -265 -9472 -249 -9438
rect -147 -9472 -131 -9438
rect -87 -9472 -71 -9438
rect 31 -9472 47 -9438
rect 91 -9472 107 -9438
rect 209 -9472 225 -9438
rect 269 -9472 285 -9438
rect 387 -9472 403 -9438
rect 447 -9472 463 -9438
rect 565 -9472 581 -9438
rect 625 -9472 641 -9438
rect 743 -9472 759 -9438
rect 803 -9472 819 -9438
rect 921 -9472 937 -9438
rect 981 -9472 997 -9438
rect 1099 -9472 1115 -9438
rect 1159 -9472 1175 -9438
rect 1277 -9472 1293 -9438
rect 1337 -9472 1353 -9438
rect 1455 -9472 1471 -9438
rect 1515 -9472 1531 -9438
rect 1633 -9472 1649 -9438
rect 1693 -9472 1709 -9438
rect 1811 -9472 1827 -9438
rect 1871 -9472 1887 -9438
rect 1989 -9472 2005 -9438
rect 2049 -9472 2065 -9438
rect 2167 -9472 2183 -9438
rect 2227 -9472 2243 -9438
rect 2345 -9472 2361 -9438
rect 2405 -9472 2421 -9438
rect 2523 -9472 2539 -9438
rect 2583 -9472 2599 -9438
rect 2701 -9472 2717 -9438
rect 2761 -9472 2777 -9438
rect 2879 -9472 2895 -9438
rect 2939 -9472 2955 -9438
rect 3057 -9472 3073 -9438
rect 3117 -9472 3133 -9438
rect 3235 -9472 3251 -9438
rect 3295 -9472 3311 -9438
rect 3413 -9472 3429 -9438
rect 3473 -9472 3489 -9438
rect 3591 -9472 3607 -9438
rect 3651 -9472 3667 -9438
rect 3769 -9472 3785 -9438
rect 3829 -9472 3845 -9438
rect 3947 -9472 3963 -9438
rect 4007 -9472 4023 -9438
rect -5628 -9524 -5594 -9508
rect -5628 -9796 -5594 -9780
rect -5450 -9524 -5416 -9508
rect -5450 -9796 -5416 -9780
rect -5272 -9524 -5238 -9508
rect -5272 -9796 -5238 -9780
rect -5094 -9524 -5060 -9508
rect -5094 -9796 -5060 -9780
rect -4916 -9524 -4882 -9508
rect -4916 -9796 -4882 -9780
rect -4738 -9524 -4704 -9508
rect -4738 -9796 -4704 -9780
rect -4560 -9524 -4526 -9508
rect -4560 -9796 -4526 -9780
rect -4382 -9524 -4348 -9508
rect -4382 -9796 -4348 -9780
rect -4204 -9524 -4170 -9508
rect -4204 -9796 -4170 -9780
rect -4026 -9524 -3992 -9508
rect 10840 -9644 10856 -9610
rect 10900 -9644 10916 -9610
rect 11132 -9644 11148 -9610
rect 11192 -9644 11208 -9610
rect 11424 -9644 11440 -9610
rect 11484 -9644 11500 -9610
rect 11716 -9644 11732 -9610
rect 11776 -9644 11792 -9610
rect 12008 -9644 12024 -9610
rect 12068 -9644 12084 -9610
rect 12300 -9644 12316 -9610
rect 12360 -9644 12376 -9610
rect 12592 -9644 12608 -9610
rect 12652 -9644 12668 -9610
rect 10772 -9694 10806 -9678
rect 6580 -9744 6596 -9710
rect 6640 -9744 6656 -9710
rect 6758 -9744 6774 -9710
rect 6818 -9744 6834 -9710
rect 6936 -9744 6952 -9710
rect 6996 -9744 7012 -9710
rect 7114 -9744 7130 -9710
rect 7174 -9744 7190 -9710
rect 7292 -9744 7308 -9710
rect 7352 -9744 7368 -9710
rect 7470 -9744 7486 -9710
rect 7530 -9744 7546 -9710
rect 7648 -9744 7664 -9710
rect 7708 -9744 7724 -9710
rect 7826 -9744 7842 -9710
rect 7886 -9744 7902 -9710
rect 8004 -9744 8020 -9710
rect 8064 -9744 8080 -9710
rect 8182 -9744 8198 -9710
rect 8242 -9744 8258 -9710
rect 8360 -9744 8376 -9710
rect 8420 -9744 8436 -9710
rect 8538 -9744 8554 -9710
rect 8598 -9744 8614 -9710
rect 8716 -9744 8732 -9710
rect 8776 -9744 8792 -9710
rect 8894 -9744 8910 -9710
rect 8954 -9744 8970 -9710
rect 9072 -9744 9088 -9710
rect 9132 -9744 9148 -9710
rect 9250 -9744 9266 -9710
rect 9310 -9744 9326 -9710
rect -4026 -9796 -3992 -9780
rect 6512 -9794 6546 -9778
rect -5560 -9864 -5544 -9830
rect -5500 -9864 -5484 -9830
rect -5382 -9864 -5366 -9830
rect -5322 -9864 -5306 -9830
rect -5204 -9864 -5188 -9830
rect -5144 -9864 -5128 -9830
rect -5026 -9864 -5010 -9830
rect -4966 -9864 -4950 -9830
rect -4848 -9864 -4832 -9830
rect -4788 -9864 -4772 -9830
rect -4670 -9864 -4654 -9830
rect -4610 -9864 -4594 -9830
rect -4492 -9864 -4476 -9830
rect -4432 -9864 -4416 -9830
rect -4314 -9864 -4298 -9830
rect -4254 -9864 -4238 -9830
rect -4136 -9864 -4120 -9830
rect -4076 -9864 -4060 -9830
rect -5560 -10024 -5544 -9990
rect -5500 -10024 -5484 -9990
rect -5382 -10024 -5366 -9990
rect -5322 -10024 -5306 -9990
rect -5204 -10024 -5188 -9990
rect -5144 -10024 -5128 -9990
rect -5026 -10024 -5010 -9990
rect -4966 -10024 -4950 -9990
rect -4848 -10024 -4832 -9990
rect -4788 -10024 -4772 -9990
rect -4670 -10024 -4654 -9990
rect -4610 -10024 -4594 -9990
rect -4492 -10024 -4476 -9990
rect -4432 -10024 -4416 -9990
rect -4314 -10024 -4298 -9990
rect -4254 -10024 -4238 -9990
rect -4136 -10024 -4120 -9990
rect -4076 -10024 -4060 -9990
rect -5628 -10074 -5594 -10058
rect -5628 -10346 -5594 -10330
rect -5450 -10074 -5416 -10058
rect -5450 -10346 -5416 -10330
rect -5272 -10074 -5238 -10058
rect -5272 -10346 -5238 -10330
rect -5094 -10074 -5060 -10058
rect -5094 -10346 -5060 -10330
rect -4916 -10074 -4882 -10058
rect -4916 -10346 -4882 -10330
rect -4738 -10074 -4704 -10058
rect -4738 -10346 -4704 -10330
rect -4560 -10074 -4526 -10058
rect -4560 -10346 -4526 -10330
rect -4382 -10074 -4348 -10058
rect -4382 -10346 -4348 -10330
rect -4204 -10074 -4170 -10058
rect -4204 -10346 -4170 -10330
rect -4026 -10074 -3992 -10058
rect -2105 -10082 -2089 -10048
rect -2045 -10082 -2029 -10048
rect -1927 -10082 -1911 -10048
rect -1867 -10082 -1851 -10048
rect -1749 -10082 -1733 -10048
rect -1689 -10082 -1673 -10048
rect -1571 -10082 -1555 -10048
rect -1511 -10082 -1495 -10048
rect -1393 -10082 -1377 -10048
rect -1333 -10082 -1317 -10048
rect -1215 -10082 -1199 -10048
rect -1155 -10082 -1139 -10048
rect -1037 -10082 -1021 -10048
rect -977 -10082 -961 -10048
rect -859 -10082 -843 -10048
rect -799 -10082 -783 -10048
rect -681 -10082 -665 -10048
rect -621 -10082 -605 -10048
rect -503 -10082 -487 -10048
rect -443 -10082 -427 -10048
rect -325 -10082 -309 -10048
rect -265 -10082 -249 -10048
rect -147 -10082 -131 -10048
rect -87 -10082 -71 -10048
rect 31 -10082 47 -10048
rect 91 -10082 107 -10048
rect 209 -10082 225 -10048
rect 269 -10082 285 -10048
rect 387 -10082 403 -10048
rect 447 -10082 463 -10048
rect 565 -10082 581 -10048
rect 625 -10082 641 -10048
rect 743 -10082 759 -10048
rect 803 -10082 819 -10048
rect 921 -10082 937 -10048
rect 981 -10082 997 -10048
rect 1099 -10082 1115 -10048
rect 1159 -10082 1175 -10048
rect 1277 -10082 1293 -10048
rect 1337 -10082 1353 -10048
rect 1455 -10082 1471 -10048
rect 1515 -10082 1531 -10048
rect 1633 -10082 1649 -10048
rect 1693 -10082 1709 -10048
rect 1811 -10082 1827 -10048
rect 1871 -10082 1887 -10048
rect 1989 -10082 2005 -10048
rect 2049 -10082 2065 -10048
rect 2167 -10082 2183 -10048
rect 2227 -10082 2243 -10048
rect 2345 -10082 2361 -10048
rect 2405 -10082 2421 -10048
rect 2523 -10082 2539 -10048
rect 2583 -10082 2599 -10048
rect 2701 -10082 2717 -10048
rect 2761 -10082 2777 -10048
rect 2879 -10082 2895 -10048
rect 2939 -10082 2955 -10048
rect 3057 -10082 3073 -10048
rect 3117 -10082 3133 -10048
rect 3235 -10082 3251 -10048
rect 3295 -10082 3311 -10048
rect 3413 -10082 3429 -10048
rect 3473 -10082 3489 -10048
rect 3591 -10082 3607 -10048
rect 3651 -10082 3667 -10048
rect 3769 -10082 3785 -10048
rect 3829 -10082 3845 -10048
rect 3947 -10082 3963 -10048
rect 4007 -10082 4023 -10048
rect 6512 -10066 6546 -10050
rect 6690 -9794 6724 -9778
rect 6690 -10066 6724 -10050
rect 6868 -9794 6902 -9778
rect 6868 -10066 6902 -10050
rect 7046 -9794 7080 -9778
rect 7046 -10066 7080 -10050
rect 7224 -9794 7258 -9778
rect 7224 -10066 7258 -10050
rect 7402 -9794 7436 -9778
rect 7402 -10066 7436 -10050
rect 7580 -9794 7614 -9778
rect 7580 -10066 7614 -10050
rect 7758 -9794 7792 -9778
rect 7758 -10066 7792 -10050
rect 7936 -9794 7970 -9778
rect 7936 -10066 7970 -10050
rect 8114 -9794 8148 -9778
rect 8114 -10066 8148 -10050
rect 8292 -9794 8326 -9778
rect 8292 -10066 8326 -10050
rect 8470 -9794 8504 -9778
rect 8470 -10066 8504 -10050
rect 8648 -9794 8682 -9778
rect 8648 -10066 8682 -10050
rect 8826 -9794 8860 -9778
rect 8826 -10066 8860 -10050
rect 9004 -9794 9038 -9778
rect 9004 -10066 9038 -10050
rect 9182 -9794 9216 -9778
rect 9182 -10066 9216 -10050
rect 9360 -9794 9394 -9778
rect 10772 -9966 10806 -9950
rect 10950 -9694 10984 -9678
rect 10950 -9966 10984 -9950
rect 11064 -9694 11098 -9678
rect 11064 -9966 11098 -9950
rect 11242 -9694 11276 -9678
rect 11242 -9966 11276 -9950
rect 11356 -9694 11390 -9678
rect 11356 -9966 11390 -9950
rect 11534 -9694 11568 -9678
rect 11534 -9966 11568 -9950
rect 11648 -9694 11682 -9678
rect 11648 -9966 11682 -9950
rect 11826 -9694 11860 -9678
rect 11826 -9966 11860 -9950
rect 11940 -9694 11974 -9678
rect 11940 -9966 11974 -9950
rect 12118 -9694 12152 -9678
rect 12118 -9966 12152 -9950
rect 12232 -9694 12266 -9678
rect 12232 -9966 12266 -9950
rect 12410 -9694 12444 -9678
rect 12410 -9966 12444 -9950
rect 12524 -9694 12558 -9678
rect 12524 -9966 12558 -9950
rect 12702 -9694 12736 -9678
rect 12702 -9966 12736 -9950
rect 10840 -10034 10856 -10000
rect 10900 -10034 10916 -10000
rect 11132 -10034 11148 -10000
rect 11192 -10034 11208 -10000
rect 11424 -10034 11440 -10000
rect 11484 -10034 11500 -10000
rect 11716 -10034 11732 -10000
rect 11776 -10034 11792 -10000
rect 12008 -10034 12024 -10000
rect 12068 -10034 12084 -10000
rect 12300 -10034 12316 -10000
rect 12360 -10034 12376 -10000
rect 12592 -10034 12608 -10000
rect 12652 -10034 12668 -10000
rect 9360 -10066 9394 -10050
rect -4026 -10346 -3992 -10330
rect -2173 -10132 -2139 -10116
rect -5560 -10414 -5544 -10380
rect -5500 -10414 -5484 -10380
rect -5382 -10414 -5366 -10380
rect -5322 -10414 -5306 -10380
rect -5204 -10414 -5188 -10380
rect -5144 -10414 -5128 -10380
rect -5026 -10414 -5010 -10380
rect -4966 -10414 -4950 -10380
rect -4848 -10414 -4832 -10380
rect -4788 -10414 -4772 -10380
rect -4670 -10414 -4654 -10380
rect -4610 -10414 -4594 -10380
rect -4492 -10414 -4476 -10380
rect -4432 -10414 -4416 -10380
rect -4314 -10414 -4298 -10380
rect -4254 -10414 -4238 -10380
rect -4136 -10414 -4120 -10380
rect -4076 -10414 -4060 -10380
rect -2173 -10404 -2139 -10388
rect -1995 -10132 -1961 -10116
rect -1995 -10404 -1961 -10388
rect -1817 -10132 -1783 -10116
rect -1817 -10404 -1783 -10388
rect -1639 -10132 -1605 -10116
rect -1639 -10404 -1605 -10388
rect -1461 -10132 -1427 -10116
rect -1461 -10404 -1427 -10388
rect -1283 -10132 -1249 -10116
rect -1283 -10404 -1249 -10388
rect -1105 -10132 -1071 -10116
rect -1105 -10404 -1071 -10388
rect -927 -10132 -893 -10116
rect -927 -10404 -893 -10388
rect -749 -10132 -715 -10116
rect -749 -10404 -715 -10388
rect -571 -10132 -537 -10116
rect -571 -10404 -537 -10388
rect -393 -10132 -359 -10116
rect -393 -10404 -359 -10388
rect -215 -10132 -181 -10116
rect -215 -10404 -181 -10388
rect -37 -10132 -3 -10116
rect -37 -10404 -3 -10388
rect 141 -10132 175 -10116
rect 141 -10404 175 -10388
rect 319 -10132 353 -10116
rect 319 -10404 353 -10388
rect 497 -10132 531 -10116
rect 497 -10404 531 -10388
rect 675 -10132 709 -10116
rect 675 -10404 709 -10388
rect 853 -10132 887 -10116
rect 853 -10404 887 -10388
rect 1031 -10132 1065 -10116
rect 1031 -10404 1065 -10388
rect 1209 -10132 1243 -10116
rect 1209 -10404 1243 -10388
rect 1387 -10132 1421 -10116
rect 1387 -10404 1421 -10388
rect 1565 -10132 1599 -10116
rect 1565 -10404 1599 -10388
rect 1743 -10132 1777 -10116
rect 1743 -10404 1777 -10388
rect 1921 -10132 1955 -10116
rect 1921 -10404 1955 -10388
rect 2099 -10132 2133 -10116
rect 2099 -10404 2133 -10388
rect 2277 -10132 2311 -10116
rect 2277 -10404 2311 -10388
rect 2455 -10132 2489 -10116
rect 2455 -10404 2489 -10388
rect 2633 -10132 2667 -10116
rect 2633 -10404 2667 -10388
rect 2811 -10132 2845 -10116
rect 2811 -10404 2845 -10388
rect 2989 -10132 3023 -10116
rect 2989 -10404 3023 -10388
rect 3167 -10132 3201 -10116
rect 3167 -10404 3201 -10388
rect 3345 -10132 3379 -10116
rect 3345 -10404 3379 -10388
rect 3523 -10132 3557 -10116
rect 3523 -10404 3557 -10388
rect 3701 -10132 3735 -10116
rect 3701 -10404 3735 -10388
rect 3879 -10132 3913 -10116
rect 3879 -10404 3913 -10388
rect 4057 -10132 4091 -10116
rect 6580 -10134 6596 -10100
rect 6640 -10134 6656 -10100
rect 6758 -10134 6774 -10100
rect 6818 -10134 6834 -10100
rect 6936 -10134 6952 -10100
rect 6996 -10134 7012 -10100
rect 7114 -10134 7130 -10100
rect 7174 -10134 7190 -10100
rect 7292 -10134 7308 -10100
rect 7352 -10134 7368 -10100
rect 7470 -10134 7486 -10100
rect 7530 -10134 7546 -10100
rect 7648 -10134 7664 -10100
rect 7708 -10134 7724 -10100
rect 7826 -10134 7842 -10100
rect 7886 -10134 7902 -10100
rect 8004 -10134 8020 -10100
rect 8064 -10134 8080 -10100
rect 8182 -10134 8198 -10100
rect 8242 -10134 8258 -10100
rect 8360 -10134 8376 -10100
rect 8420 -10134 8436 -10100
rect 8538 -10134 8554 -10100
rect 8598 -10134 8614 -10100
rect 8716 -10134 8732 -10100
rect 8776 -10134 8792 -10100
rect 8894 -10134 8910 -10100
rect 8954 -10134 8970 -10100
rect 9072 -10134 9088 -10100
rect 9132 -10134 9148 -10100
rect 9250 -10134 9266 -10100
rect 9310 -10134 9326 -10100
rect 4057 -10404 4091 -10388
rect 10840 -10414 10856 -10380
rect 10900 -10414 10916 -10380
rect 11132 -10414 11148 -10380
rect 11192 -10414 11208 -10380
rect 11424 -10414 11440 -10380
rect 11484 -10414 11500 -10380
rect 11716 -10414 11732 -10380
rect 11776 -10414 11792 -10380
rect 12008 -10414 12024 -10380
rect 12068 -10414 12084 -10380
rect 12300 -10414 12316 -10380
rect 12360 -10414 12376 -10380
rect 12592 -10414 12608 -10380
rect 12652 -10414 12668 -10380
rect -2105 -10472 -2089 -10438
rect -2045 -10472 -2029 -10438
rect -1927 -10472 -1911 -10438
rect -1867 -10472 -1851 -10438
rect -1749 -10472 -1733 -10438
rect -1689 -10472 -1673 -10438
rect -1571 -10472 -1555 -10438
rect -1511 -10472 -1495 -10438
rect -1393 -10472 -1377 -10438
rect -1333 -10472 -1317 -10438
rect -1215 -10472 -1199 -10438
rect -1155 -10472 -1139 -10438
rect -1037 -10472 -1021 -10438
rect -977 -10472 -961 -10438
rect -859 -10472 -843 -10438
rect -799 -10472 -783 -10438
rect -681 -10472 -665 -10438
rect -621 -10472 -605 -10438
rect -503 -10472 -487 -10438
rect -443 -10472 -427 -10438
rect -325 -10472 -309 -10438
rect -265 -10472 -249 -10438
rect -147 -10472 -131 -10438
rect -87 -10472 -71 -10438
rect 31 -10472 47 -10438
rect 91 -10472 107 -10438
rect 209 -10472 225 -10438
rect 269 -10472 285 -10438
rect 387 -10472 403 -10438
rect 447 -10472 463 -10438
rect 565 -10472 581 -10438
rect 625 -10472 641 -10438
rect 743 -10472 759 -10438
rect 803 -10472 819 -10438
rect 921 -10472 937 -10438
rect 981 -10472 997 -10438
rect 1099 -10472 1115 -10438
rect 1159 -10472 1175 -10438
rect 1277 -10472 1293 -10438
rect 1337 -10472 1353 -10438
rect 1455 -10472 1471 -10438
rect 1515 -10472 1531 -10438
rect 1633 -10472 1649 -10438
rect 1693 -10472 1709 -10438
rect 1811 -10472 1827 -10438
rect 1871 -10472 1887 -10438
rect 1989 -10472 2005 -10438
rect 2049 -10472 2065 -10438
rect 2167 -10472 2183 -10438
rect 2227 -10472 2243 -10438
rect 2345 -10472 2361 -10438
rect 2405 -10472 2421 -10438
rect 2523 -10472 2539 -10438
rect 2583 -10472 2599 -10438
rect 2701 -10472 2717 -10438
rect 2761 -10472 2777 -10438
rect 2879 -10472 2895 -10438
rect 2939 -10472 2955 -10438
rect 3057 -10472 3073 -10438
rect 3117 -10472 3133 -10438
rect 3235 -10472 3251 -10438
rect 3295 -10472 3311 -10438
rect 3413 -10472 3429 -10438
rect 3473 -10472 3489 -10438
rect 3591 -10472 3607 -10438
rect 3651 -10472 3667 -10438
rect 3769 -10472 3785 -10438
rect 3829 -10472 3845 -10438
rect 3947 -10472 3963 -10438
rect 4007 -10472 4023 -10438
rect 10772 -10464 10806 -10448
rect -5560 -10574 -5544 -10540
rect -5500 -10574 -5484 -10540
rect -5382 -10574 -5366 -10540
rect -5322 -10574 -5306 -10540
rect -5204 -10574 -5188 -10540
rect -5144 -10574 -5128 -10540
rect -5026 -10574 -5010 -10540
rect -4966 -10574 -4950 -10540
rect -4848 -10574 -4832 -10540
rect -4788 -10574 -4772 -10540
rect -4670 -10574 -4654 -10540
rect -4610 -10574 -4594 -10540
rect -4492 -10574 -4476 -10540
rect -4432 -10574 -4416 -10540
rect -4314 -10574 -4298 -10540
rect -4254 -10574 -4238 -10540
rect -4136 -10574 -4120 -10540
rect -4076 -10574 -4060 -10540
rect -5628 -10624 -5594 -10608
rect -5628 -10896 -5594 -10880
rect -5450 -10624 -5416 -10608
rect -5450 -10896 -5416 -10880
rect -5272 -10624 -5238 -10608
rect -5272 -10896 -5238 -10880
rect -5094 -10624 -5060 -10608
rect -5094 -10896 -5060 -10880
rect -4916 -10624 -4882 -10608
rect -4916 -10896 -4882 -10880
rect -4738 -10624 -4704 -10608
rect -4738 -10896 -4704 -10880
rect -4560 -10624 -4526 -10608
rect -4560 -10896 -4526 -10880
rect -4382 -10624 -4348 -10608
rect -4382 -10896 -4348 -10880
rect -4204 -10624 -4170 -10608
rect -4204 -10896 -4170 -10880
rect -4026 -10624 -3992 -10608
rect 6580 -10644 6596 -10610
rect 6640 -10644 6656 -10610
rect 6758 -10644 6774 -10610
rect 6818 -10644 6834 -10610
rect 6936 -10644 6952 -10610
rect 6996 -10644 7012 -10610
rect 7114 -10644 7130 -10610
rect 7174 -10644 7190 -10610
rect 7292 -10644 7308 -10610
rect 7352 -10644 7368 -10610
rect 7470 -10644 7486 -10610
rect 7530 -10644 7546 -10610
rect 7648 -10644 7664 -10610
rect 7708 -10644 7724 -10610
rect 7826 -10644 7842 -10610
rect 7886 -10644 7902 -10610
rect 8004 -10644 8020 -10610
rect 8064 -10644 8080 -10610
rect 8182 -10644 8198 -10610
rect 8242 -10644 8258 -10610
rect 8360 -10644 8376 -10610
rect 8420 -10644 8436 -10610
rect 8538 -10644 8554 -10610
rect 8598 -10644 8614 -10610
rect 8716 -10644 8732 -10610
rect 8776 -10644 8792 -10610
rect 8894 -10644 8910 -10610
rect 8954 -10644 8970 -10610
rect 9072 -10644 9088 -10610
rect 9132 -10644 9148 -10610
rect 9250 -10644 9266 -10610
rect 9310 -10644 9326 -10610
rect -4026 -10896 -3992 -10880
rect 6512 -10694 6546 -10678
rect -5560 -10964 -5544 -10930
rect -5500 -10964 -5484 -10930
rect -5382 -10964 -5366 -10930
rect -5322 -10964 -5306 -10930
rect -5204 -10964 -5188 -10930
rect -5144 -10964 -5128 -10930
rect -5026 -10964 -5010 -10930
rect -4966 -10964 -4950 -10930
rect -4848 -10964 -4832 -10930
rect -4788 -10964 -4772 -10930
rect -4670 -10964 -4654 -10930
rect -4610 -10964 -4594 -10930
rect -4492 -10964 -4476 -10930
rect -4432 -10964 -4416 -10930
rect -4314 -10964 -4298 -10930
rect -4254 -10964 -4238 -10930
rect -4136 -10964 -4120 -10930
rect -4076 -10964 -4060 -10930
rect 6512 -10966 6546 -10950
rect 6690 -10694 6724 -10678
rect 6690 -10966 6724 -10950
rect 6868 -10694 6902 -10678
rect 6868 -10966 6902 -10950
rect 7046 -10694 7080 -10678
rect 7046 -10966 7080 -10950
rect 7224 -10694 7258 -10678
rect 7224 -10966 7258 -10950
rect 7402 -10694 7436 -10678
rect 7402 -10966 7436 -10950
rect 7580 -10694 7614 -10678
rect 7580 -10966 7614 -10950
rect 7758 -10694 7792 -10678
rect 7758 -10966 7792 -10950
rect 7936 -10694 7970 -10678
rect 7936 -10966 7970 -10950
rect 8114 -10694 8148 -10678
rect 8114 -10966 8148 -10950
rect 8292 -10694 8326 -10678
rect 8292 -10966 8326 -10950
rect 8470 -10694 8504 -10678
rect 8470 -10966 8504 -10950
rect 8648 -10694 8682 -10678
rect 8648 -10966 8682 -10950
rect 8826 -10694 8860 -10678
rect 8826 -10966 8860 -10950
rect 9004 -10694 9038 -10678
rect 9004 -10966 9038 -10950
rect 9182 -10694 9216 -10678
rect 9182 -10966 9216 -10950
rect 9360 -10694 9394 -10678
rect 10772 -10736 10806 -10720
rect 10950 -10464 10984 -10448
rect 10950 -10736 10984 -10720
rect 11064 -10464 11098 -10448
rect 11064 -10736 11098 -10720
rect 11242 -10464 11276 -10448
rect 11242 -10736 11276 -10720
rect 11356 -10464 11390 -10448
rect 11356 -10736 11390 -10720
rect 11534 -10464 11568 -10448
rect 11534 -10736 11568 -10720
rect 11648 -10464 11682 -10448
rect 11648 -10736 11682 -10720
rect 11826 -10464 11860 -10448
rect 11826 -10736 11860 -10720
rect 11940 -10464 11974 -10448
rect 11940 -10736 11974 -10720
rect 12118 -10464 12152 -10448
rect 12118 -10736 12152 -10720
rect 12232 -10464 12266 -10448
rect 12232 -10736 12266 -10720
rect 12410 -10464 12444 -10448
rect 12410 -10736 12444 -10720
rect 12524 -10464 12558 -10448
rect 12524 -10736 12558 -10720
rect 12702 -10464 12736 -10448
rect 12702 -10736 12736 -10720
rect 10840 -10804 10856 -10770
rect 10900 -10804 10916 -10770
rect 11132 -10804 11148 -10770
rect 11192 -10804 11208 -10770
rect 11424 -10804 11440 -10770
rect 11484 -10804 11500 -10770
rect 11716 -10804 11732 -10770
rect 11776 -10804 11792 -10770
rect 12008 -10804 12024 -10770
rect 12068 -10804 12084 -10770
rect 12300 -10804 12316 -10770
rect 12360 -10804 12376 -10770
rect 12592 -10804 12608 -10770
rect 12652 -10804 12668 -10770
rect 9360 -10966 9394 -10950
rect 6580 -11034 6596 -11000
rect 6640 -11034 6656 -11000
rect 6758 -11034 6774 -11000
rect 6818 -11034 6834 -11000
rect 6936 -11034 6952 -11000
rect 6996 -11034 7012 -11000
rect 7114 -11034 7130 -11000
rect 7174 -11034 7190 -11000
rect 7292 -11034 7308 -11000
rect 7352 -11034 7368 -11000
rect 7470 -11034 7486 -11000
rect 7530 -11034 7546 -11000
rect 7648 -11034 7664 -11000
rect 7708 -11034 7724 -11000
rect 7826 -11034 7842 -11000
rect 7886 -11034 7902 -11000
rect 8004 -11034 8020 -11000
rect 8064 -11034 8080 -11000
rect 8182 -11034 8198 -11000
rect 8242 -11034 8258 -11000
rect 8360 -11034 8376 -11000
rect 8420 -11034 8436 -11000
rect 8538 -11034 8554 -11000
rect 8598 -11034 8614 -11000
rect 8716 -11034 8732 -11000
rect 8776 -11034 8792 -11000
rect 8894 -11034 8910 -11000
rect 8954 -11034 8970 -11000
rect 9072 -11034 9088 -11000
rect 9132 -11034 9148 -11000
rect 9250 -11034 9266 -11000
rect 9310 -11034 9326 -11000
rect -2105 -11082 -2089 -11048
rect -2045 -11082 -2029 -11048
rect -1927 -11082 -1911 -11048
rect -1867 -11082 -1851 -11048
rect -1749 -11082 -1733 -11048
rect -1689 -11082 -1673 -11048
rect -1571 -11082 -1555 -11048
rect -1511 -11082 -1495 -11048
rect -1393 -11082 -1377 -11048
rect -1333 -11082 -1317 -11048
rect -1215 -11082 -1199 -11048
rect -1155 -11082 -1139 -11048
rect -1037 -11082 -1021 -11048
rect -977 -11082 -961 -11048
rect -859 -11082 -843 -11048
rect -799 -11082 -783 -11048
rect -681 -11082 -665 -11048
rect -621 -11082 -605 -11048
rect -503 -11082 -487 -11048
rect -443 -11082 -427 -11048
rect -325 -11082 -309 -11048
rect -265 -11082 -249 -11048
rect -147 -11082 -131 -11048
rect -87 -11082 -71 -11048
rect 31 -11082 47 -11048
rect 91 -11082 107 -11048
rect 209 -11082 225 -11048
rect 269 -11082 285 -11048
rect 387 -11082 403 -11048
rect 447 -11082 463 -11048
rect 565 -11082 581 -11048
rect 625 -11082 641 -11048
rect 743 -11082 759 -11048
rect 803 -11082 819 -11048
rect 921 -11082 937 -11048
rect 981 -11082 997 -11048
rect 1099 -11082 1115 -11048
rect 1159 -11082 1175 -11048
rect 1277 -11082 1293 -11048
rect 1337 -11082 1353 -11048
rect 1455 -11082 1471 -11048
rect 1515 -11082 1531 -11048
rect 1633 -11082 1649 -11048
rect 1693 -11082 1709 -11048
rect 1811 -11082 1827 -11048
rect 1871 -11082 1887 -11048
rect 1989 -11082 2005 -11048
rect 2049 -11082 2065 -11048
rect 2167 -11082 2183 -11048
rect 2227 -11082 2243 -11048
rect 2345 -11082 2361 -11048
rect 2405 -11082 2421 -11048
rect 2523 -11082 2539 -11048
rect 2583 -11082 2599 -11048
rect 2701 -11082 2717 -11048
rect 2761 -11082 2777 -11048
rect 2879 -11082 2895 -11048
rect 2939 -11082 2955 -11048
rect 3057 -11082 3073 -11048
rect 3117 -11082 3133 -11048
rect 3235 -11082 3251 -11048
rect 3295 -11082 3311 -11048
rect 3413 -11082 3429 -11048
rect 3473 -11082 3489 -11048
rect 3591 -11082 3607 -11048
rect 3651 -11082 3667 -11048
rect 3769 -11082 3785 -11048
rect 3829 -11082 3845 -11048
rect 3947 -11082 3963 -11048
rect 4007 -11082 4023 -11048
rect -5560 -11124 -5544 -11090
rect -5500 -11124 -5484 -11090
rect -5382 -11124 -5366 -11090
rect -5322 -11124 -5306 -11090
rect -5204 -11124 -5188 -11090
rect -5144 -11124 -5128 -11090
rect -5026 -11124 -5010 -11090
rect -4966 -11124 -4950 -11090
rect -4848 -11124 -4832 -11090
rect -4788 -11124 -4772 -11090
rect -4670 -11124 -4654 -11090
rect -4610 -11124 -4594 -11090
rect -4492 -11124 -4476 -11090
rect -4432 -11124 -4416 -11090
rect -4314 -11124 -4298 -11090
rect -4254 -11124 -4238 -11090
rect -4136 -11124 -4120 -11090
rect -4076 -11124 -4060 -11090
rect -2173 -11132 -2139 -11116
rect -5628 -11174 -5594 -11158
rect -5628 -11446 -5594 -11430
rect -5450 -11174 -5416 -11158
rect -5450 -11446 -5416 -11430
rect -5272 -11174 -5238 -11158
rect -5272 -11446 -5238 -11430
rect -5094 -11174 -5060 -11158
rect -5094 -11446 -5060 -11430
rect -4916 -11174 -4882 -11158
rect -4916 -11446 -4882 -11430
rect -4738 -11174 -4704 -11158
rect -4738 -11446 -4704 -11430
rect -4560 -11174 -4526 -11158
rect -4560 -11446 -4526 -11430
rect -4382 -11174 -4348 -11158
rect -4382 -11446 -4348 -11430
rect -4204 -11174 -4170 -11158
rect -4204 -11446 -4170 -11430
rect -4026 -11174 -3992 -11158
rect -4026 -11446 -3992 -11430
rect -3009 -11276 -2783 -11252
rect -3009 -11454 -2985 -11276
rect -2807 -11454 -2783 -11276
rect -2173 -11404 -2139 -11388
rect -1995 -11132 -1961 -11116
rect -1995 -11404 -1961 -11388
rect -1817 -11132 -1783 -11116
rect -1817 -11404 -1783 -11388
rect -1639 -11132 -1605 -11116
rect -1639 -11404 -1605 -11388
rect -1461 -11132 -1427 -11116
rect -1461 -11404 -1427 -11388
rect -1283 -11132 -1249 -11116
rect -1283 -11404 -1249 -11388
rect -1105 -11132 -1071 -11116
rect -1105 -11404 -1071 -11388
rect -927 -11132 -893 -11116
rect -927 -11404 -893 -11388
rect -749 -11132 -715 -11116
rect -749 -11404 -715 -11388
rect -571 -11132 -537 -11116
rect -571 -11404 -537 -11388
rect -393 -11132 -359 -11116
rect -393 -11404 -359 -11388
rect -215 -11132 -181 -11116
rect -215 -11404 -181 -11388
rect -37 -11132 -3 -11116
rect -37 -11404 -3 -11388
rect 141 -11132 175 -11116
rect 141 -11404 175 -11388
rect 319 -11132 353 -11116
rect 319 -11404 353 -11388
rect 497 -11132 531 -11116
rect 497 -11404 531 -11388
rect 675 -11132 709 -11116
rect 675 -11404 709 -11388
rect 853 -11132 887 -11116
rect 853 -11404 887 -11388
rect 1031 -11132 1065 -11116
rect 1031 -11404 1065 -11388
rect 1209 -11132 1243 -11116
rect 1209 -11404 1243 -11388
rect 1387 -11132 1421 -11116
rect 1387 -11404 1421 -11388
rect 1565 -11132 1599 -11116
rect 1565 -11404 1599 -11388
rect 1743 -11132 1777 -11116
rect 1743 -11404 1777 -11388
rect 1921 -11132 1955 -11116
rect 1921 -11404 1955 -11388
rect 2099 -11132 2133 -11116
rect 2099 -11404 2133 -11388
rect 2277 -11132 2311 -11116
rect 2277 -11404 2311 -11388
rect 2455 -11132 2489 -11116
rect 2455 -11404 2489 -11388
rect 2633 -11132 2667 -11116
rect 2633 -11404 2667 -11388
rect 2811 -11132 2845 -11116
rect 2811 -11404 2845 -11388
rect 2989 -11132 3023 -11116
rect 2989 -11404 3023 -11388
rect 3167 -11132 3201 -11116
rect 3167 -11404 3201 -11388
rect 3345 -11132 3379 -11116
rect 3345 -11404 3379 -11388
rect 3523 -11132 3557 -11116
rect 3523 -11404 3557 -11388
rect 3701 -11132 3735 -11116
rect 3701 -11404 3735 -11388
rect 3879 -11132 3913 -11116
rect 3879 -11404 3913 -11388
rect 4057 -11132 4091 -11116
rect 5662 -11151 5888 -11127
rect 5662 -11329 5686 -11151
rect 5864 -11329 5888 -11151
rect 5662 -11353 5888 -11329
rect 9958 -11191 10184 -11167
rect 10840 -11184 10856 -11150
rect 10900 -11184 10916 -11150
rect 11132 -11184 11148 -11150
rect 11192 -11184 11208 -11150
rect 11424 -11184 11440 -11150
rect 11484 -11184 11500 -11150
rect 11716 -11184 11732 -11150
rect 11776 -11184 11792 -11150
rect 12008 -11184 12024 -11150
rect 12068 -11184 12084 -11150
rect 12300 -11184 12316 -11150
rect 12360 -11184 12376 -11150
rect 12592 -11184 12608 -11150
rect 12652 -11184 12668 -11150
rect 4057 -11404 4091 -11388
rect 9958 -11369 9982 -11191
rect 10160 -11369 10184 -11191
rect 9958 -11393 10184 -11369
rect 10772 -11234 10806 -11218
rect -3009 -11478 -2783 -11454
rect -2105 -11472 -2089 -11438
rect -2045 -11472 -2029 -11438
rect -1927 -11472 -1911 -11438
rect -1867 -11472 -1851 -11438
rect -1749 -11472 -1733 -11438
rect -1689 -11472 -1673 -11438
rect -1571 -11472 -1555 -11438
rect -1511 -11472 -1495 -11438
rect -1393 -11472 -1377 -11438
rect -1333 -11472 -1317 -11438
rect -1215 -11472 -1199 -11438
rect -1155 -11472 -1139 -11438
rect -1037 -11472 -1021 -11438
rect -977 -11472 -961 -11438
rect -859 -11472 -843 -11438
rect -799 -11472 -783 -11438
rect -681 -11472 -665 -11438
rect -621 -11472 -605 -11438
rect -503 -11472 -487 -11438
rect -443 -11472 -427 -11438
rect -325 -11472 -309 -11438
rect -265 -11472 -249 -11438
rect -147 -11472 -131 -11438
rect -87 -11472 -71 -11438
rect 31 -11472 47 -11438
rect 91 -11472 107 -11438
rect 209 -11472 225 -11438
rect 269 -11472 285 -11438
rect 387 -11472 403 -11438
rect 447 -11472 463 -11438
rect 565 -11472 581 -11438
rect 625 -11472 641 -11438
rect 743 -11472 759 -11438
rect 803 -11472 819 -11438
rect 921 -11472 937 -11438
rect 981 -11472 997 -11438
rect 1099 -11472 1115 -11438
rect 1159 -11472 1175 -11438
rect 1277 -11472 1293 -11438
rect 1337 -11472 1353 -11438
rect 1455 -11472 1471 -11438
rect 1515 -11472 1531 -11438
rect 1633 -11472 1649 -11438
rect 1693 -11472 1709 -11438
rect 1811 -11472 1827 -11438
rect 1871 -11472 1887 -11438
rect 1989 -11472 2005 -11438
rect 2049 -11472 2065 -11438
rect 2167 -11472 2183 -11438
rect 2227 -11472 2243 -11438
rect 2345 -11472 2361 -11438
rect 2405 -11472 2421 -11438
rect 2523 -11472 2539 -11438
rect 2583 -11472 2599 -11438
rect 2701 -11472 2717 -11438
rect 2761 -11472 2777 -11438
rect 2879 -11472 2895 -11438
rect 2939 -11472 2955 -11438
rect 3057 -11472 3073 -11438
rect 3117 -11472 3133 -11438
rect 3235 -11472 3251 -11438
rect 3295 -11472 3311 -11438
rect 3413 -11472 3429 -11438
rect 3473 -11472 3489 -11438
rect 3591 -11472 3607 -11438
rect 3651 -11472 3667 -11438
rect 3769 -11472 3785 -11438
rect 3829 -11472 3845 -11438
rect 3947 -11472 3963 -11438
rect 4007 -11472 4023 -11438
rect -5560 -11514 -5544 -11480
rect -5500 -11514 -5484 -11480
rect -5382 -11514 -5366 -11480
rect -5322 -11514 -5306 -11480
rect -5204 -11514 -5188 -11480
rect -5144 -11514 -5128 -11480
rect -5026 -11514 -5010 -11480
rect -4966 -11514 -4950 -11480
rect -4848 -11514 -4832 -11480
rect -4788 -11514 -4772 -11480
rect -4670 -11514 -4654 -11480
rect -4610 -11514 -4594 -11480
rect -4492 -11514 -4476 -11480
rect -4432 -11514 -4416 -11480
rect -4314 -11514 -4298 -11480
rect -4254 -11514 -4238 -11480
rect -4136 -11514 -4120 -11480
rect -4076 -11514 -4060 -11480
rect 10772 -11506 10806 -11490
rect 10950 -11234 10984 -11218
rect 10950 -11506 10984 -11490
rect 11064 -11234 11098 -11218
rect 11064 -11506 11098 -11490
rect 11242 -11234 11276 -11218
rect 11242 -11506 11276 -11490
rect 11356 -11234 11390 -11218
rect 11356 -11506 11390 -11490
rect 11534 -11234 11568 -11218
rect 11534 -11506 11568 -11490
rect 11648 -11234 11682 -11218
rect 11648 -11506 11682 -11490
rect 11826 -11234 11860 -11218
rect 11826 -11506 11860 -11490
rect 11940 -11234 11974 -11218
rect 11940 -11506 11974 -11490
rect 12118 -11234 12152 -11218
rect 12118 -11506 12152 -11490
rect 12232 -11234 12266 -11218
rect 12232 -11506 12266 -11490
rect 12410 -11234 12444 -11218
rect 12410 -11506 12444 -11490
rect 12524 -11234 12558 -11218
rect 12524 -11506 12558 -11490
rect 12702 -11234 12736 -11218
rect 12702 -11506 12736 -11490
rect 6580 -11544 6596 -11510
rect 6640 -11544 6656 -11510
rect 6758 -11544 6774 -11510
rect 6818 -11544 6834 -11510
rect 6936 -11544 6952 -11510
rect 6996 -11544 7012 -11510
rect 7114 -11544 7130 -11510
rect 7174 -11544 7190 -11510
rect 7292 -11544 7308 -11510
rect 7352 -11544 7368 -11510
rect 7470 -11544 7486 -11510
rect 7530 -11544 7546 -11510
rect 7648 -11544 7664 -11510
rect 7708 -11544 7724 -11510
rect 7826 -11544 7842 -11510
rect 7886 -11544 7902 -11510
rect 8004 -11544 8020 -11510
rect 8064 -11544 8080 -11510
rect 8182 -11544 8198 -11510
rect 8242 -11544 8258 -11510
rect 8360 -11544 8376 -11510
rect 8420 -11544 8436 -11510
rect 8538 -11544 8554 -11510
rect 8598 -11544 8614 -11510
rect 8716 -11544 8732 -11510
rect 8776 -11544 8792 -11510
rect 8894 -11544 8910 -11510
rect 8954 -11544 8970 -11510
rect 9072 -11544 9088 -11510
rect 9132 -11544 9148 -11510
rect 9250 -11544 9266 -11510
rect 9310 -11544 9326 -11510
rect 10840 -11574 10856 -11540
rect 10900 -11574 10916 -11540
rect 11132 -11574 11148 -11540
rect 11192 -11574 11208 -11540
rect 11424 -11574 11440 -11540
rect 11484 -11574 11500 -11540
rect 11716 -11574 11732 -11540
rect 11776 -11574 11792 -11540
rect 12008 -11574 12024 -11540
rect 12068 -11574 12084 -11540
rect 12300 -11574 12316 -11540
rect 12360 -11574 12376 -11540
rect 12592 -11574 12608 -11540
rect 12652 -11574 12668 -11540
rect 6512 -11594 6546 -11578
rect -5560 -11674 -5544 -11640
rect -5500 -11674 -5484 -11640
rect -5382 -11674 -5366 -11640
rect -5322 -11674 -5306 -11640
rect -5204 -11674 -5188 -11640
rect -5144 -11674 -5128 -11640
rect -5026 -11674 -5010 -11640
rect -4966 -11674 -4950 -11640
rect -4848 -11674 -4832 -11640
rect -4788 -11674 -4772 -11640
rect -4670 -11674 -4654 -11640
rect -4610 -11674 -4594 -11640
rect -4492 -11674 -4476 -11640
rect -4432 -11674 -4416 -11640
rect -4314 -11674 -4298 -11640
rect -4254 -11674 -4238 -11640
rect -4136 -11674 -4120 -11640
rect -4076 -11674 -4060 -11640
rect -5628 -11724 -5594 -11708
rect -5628 -11996 -5594 -11980
rect -5450 -11724 -5416 -11708
rect -5450 -11996 -5416 -11980
rect -5272 -11724 -5238 -11708
rect -5272 -11996 -5238 -11980
rect -5094 -11724 -5060 -11708
rect -5094 -11996 -5060 -11980
rect -4916 -11724 -4882 -11708
rect -4916 -11996 -4882 -11980
rect -4738 -11724 -4704 -11708
rect -4738 -11996 -4704 -11980
rect -4560 -11724 -4526 -11708
rect -4560 -11996 -4526 -11980
rect -4382 -11724 -4348 -11708
rect -4382 -11996 -4348 -11980
rect -4204 -11724 -4170 -11708
rect -4204 -11996 -4170 -11980
rect -4026 -11724 -3992 -11708
rect 6512 -11866 6546 -11850
rect 6690 -11594 6724 -11578
rect 6690 -11866 6724 -11850
rect 6868 -11594 6902 -11578
rect 6868 -11866 6902 -11850
rect 7046 -11594 7080 -11578
rect 7046 -11866 7080 -11850
rect 7224 -11594 7258 -11578
rect 7224 -11866 7258 -11850
rect 7402 -11594 7436 -11578
rect 7402 -11866 7436 -11850
rect 7580 -11594 7614 -11578
rect 7580 -11866 7614 -11850
rect 7758 -11594 7792 -11578
rect 7758 -11866 7792 -11850
rect 7936 -11594 7970 -11578
rect 7936 -11866 7970 -11850
rect 8114 -11594 8148 -11578
rect 8114 -11866 8148 -11850
rect 8292 -11594 8326 -11578
rect 8292 -11866 8326 -11850
rect 8470 -11594 8504 -11578
rect 8470 -11866 8504 -11850
rect 8648 -11594 8682 -11578
rect 8648 -11866 8682 -11850
rect 8826 -11594 8860 -11578
rect 8826 -11866 8860 -11850
rect 9004 -11594 9038 -11578
rect 9004 -11866 9038 -11850
rect 9182 -11594 9216 -11578
rect 9182 -11866 9216 -11850
rect 9360 -11594 9394 -11578
rect 9360 -11866 9394 -11850
rect 6580 -11934 6596 -11900
rect 6640 -11934 6656 -11900
rect 6758 -11934 6774 -11900
rect 6818 -11934 6834 -11900
rect 6936 -11934 6952 -11900
rect 6996 -11934 7012 -11900
rect 7114 -11934 7130 -11900
rect 7174 -11934 7190 -11900
rect 7292 -11934 7308 -11900
rect 7352 -11934 7368 -11900
rect 7470 -11934 7486 -11900
rect 7530 -11934 7546 -11900
rect 7648 -11934 7664 -11900
rect 7708 -11934 7724 -11900
rect 7826 -11934 7842 -11900
rect 7886 -11934 7902 -11900
rect 8004 -11934 8020 -11900
rect 8064 -11934 8080 -11900
rect 8182 -11934 8198 -11900
rect 8242 -11934 8258 -11900
rect 8360 -11934 8376 -11900
rect 8420 -11934 8436 -11900
rect 8538 -11934 8554 -11900
rect 8598 -11934 8614 -11900
rect 8716 -11934 8732 -11900
rect 8776 -11934 8792 -11900
rect 8894 -11934 8910 -11900
rect 8954 -11934 8970 -11900
rect 9072 -11934 9088 -11900
rect 9132 -11934 9148 -11900
rect 9250 -11934 9266 -11900
rect 9310 -11934 9326 -11900
rect -4026 -11996 -3992 -11980
rect -5560 -12064 -5544 -12030
rect -5500 -12064 -5484 -12030
rect -5382 -12064 -5366 -12030
rect -5322 -12064 -5306 -12030
rect -5204 -12064 -5188 -12030
rect -5144 -12064 -5128 -12030
rect -5026 -12064 -5010 -12030
rect -4966 -12064 -4950 -12030
rect -4848 -12064 -4832 -12030
rect -4788 -12064 -4772 -12030
rect -4670 -12064 -4654 -12030
rect -4610 -12064 -4594 -12030
rect -4492 -12064 -4476 -12030
rect -4432 -12064 -4416 -12030
rect -4314 -12064 -4298 -12030
rect -4254 -12064 -4238 -12030
rect -4136 -12064 -4120 -12030
rect -4076 -12064 -4060 -12030
rect -2105 -12082 -2089 -12048
rect -2045 -12082 -2029 -12048
rect -1927 -12082 -1911 -12048
rect -1867 -12082 -1851 -12048
rect -1749 -12082 -1733 -12048
rect -1689 -12082 -1673 -12048
rect -1571 -12082 -1555 -12048
rect -1511 -12082 -1495 -12048
rect -1393 -12082 -1377 -12048
rect -1333 -12082 -1317 -12048
rect -1215 -12082 -1199 -12048
rect -1155 -12082 -1139 -12048
rect -1037 -12082 -1021 -12048
rect -977 -12082 -961 -12048
rect -859 -12082 -843 -12048
rect -799 -12082 -783 -12048
rect -681 -12082 -665 -12048
rect -621 -12082 -605 -12048
rect -503 -12082 -487 -12048
rect -443 -12082 -427 -12048
rect -325 -12082 -309 -12048
rect -265 -12082 -249 -12048
rect -147 -12082 -131 -12048
rect -87 -12082 -71 -12048
rect 31 -12082 47 -12048
rect 91 -12082 107 -12048
rect 209 -12082 225 -12048
rect 269 -12082 285 -12048
rect 387 -12082 403 -12048
rect 447 -12082 463 -12048
rect 565 -12082 581 -12048
rect 625 -12082 641 -12048
rect 743 -12082 759 -12048
rect 803 -12082 819 -12048
rect 921 -12082 937 -12048
rect 981 -12082 997 -12048
rect 1099 -12082 1115 -12048
rect 1159 -12082 1175 -12048
rect 1277 -12082 1293 -12048
rect 1337 -12082 1353 -12048
rect 1455 -12082 1471 -12048
rect 1515 -12082 1531 -12048
rect 1633 -12082 1649 -12048
rect 1693 -12082 1709 -12048
rect 1811 -12082 1827 -12048
rect 1871 -12082 1887 -12048
rect 1989 -12082 2005 -12048
rect 2049 -12082 2065 -12048
rect 2167 -12082 2183 -12048
rect 2227 -12082 2243 -12048
rect 2345 -12082 2361 -12048
rect 2405 -12082 2421 -12048
rect 2523 -12082 2539 -12048
rect 2583 -12082 2599 -12048
rect 2701 -12082 2717 -12048
rect 2761 -12082 2777 -12048
rect 2879 -12082 2895 -12048
rect 2939 -12082 2955 -12048
rect 3057 -12082 3073 -12048
rect 3117 -12082 3133 -12048
rect 3235 -12082 3251 -12048
rect 3295 -12082 3311 -12048
rect 3413 -12082 3429 -12048
rect 3473 -12082 3489 -12048
rect 3591 -12082 3607 -12048
rect 3651 -12082 3667 -12048
rect 3769 -12082 3785 -12048
rect 3829 -12082 3845 -12048
rect 3947 -12082 3963 -12048
rect 4007 -12082 4023 -12048
rect -2173 -12132 -2139 -12116
rect -2173 -12404 -2139 -12388
rect -1995 -12132 -1961 -12116
rect -1995 -12404 -1961 -12388
rect -1817 -12132 -1783 -12116
rect -1817 -12404 -1783 -12388
rect -1639 -12132 -1605 -12116
rect -1639 -12404 -1605 -12388
rect -1461 -12132 -1427 -12116
rect -1461 -12404 -1427 -12388
rect -1283 -12132 -1249 -12116
rect -1283 -12404 -1249 -12388
rect -1105 -12132 -1071 -12116
rect -1105 -12404 -1071 -12388
rect -927 -12132 -893 -12116
rect -927 -12404 -893 -12388
rect -749 -12132 -715 -12116
rect -749 -12404 -715 -12388
rect -571 -12132 -537 -12116
rect -571 -12404 -537 -12388
rect -393 -12132 -359 -12116
rect -393 -12404 -359 -12388
rect -215 -12132 -181 -12116
rect -215 -12404 -181 -12388
rect -37 -12132 -3 -12116
rect -37 -12404 -3 -12388
rect 141 -12132 175 -12116
rect 141 -12404 175 -12388
rect 319 -12132 353 -12116
rect 319 -12404 353 -12388
rect 497 -12132 531 -12116
rect 497 -12404 531 -12388
rect 675 -12132 709 -12116
rect 675 -12404 709 -12388
rect 853 -12132 887 -12116
rect 853 -12404 887 -12388
rect 1031 -12132 1065 -12116
rect 1031 -12404 1065 -12388
rect 1209 -12132 1243 -12116
rect 1209 -12404 1243 -12388
rect 1387 -12132 1421 -12116
rect 1387 -12404 1421 -12388
rect 1565 -12132 1599 -12116
rect 1565 -12404 1599 -12388
rect 1743 -12132 1777 -12116
rect 1743 -12404 1777 -12388
rect 1921 -12132 1955 -12116
rect 1921 -12404 1955 -12388
rect 2099 -12132 2133 -12116
rect 2099 -12404 2133 -12388
rect 2277 -12132 2311 -12116
rect 2277 -12404 2311 -12388
rect 2455 -12132 2489 -12116
rect 2455 -12404 2489 -12388
rect 2633 -12132 2667 -12116
rect 2633 -12404 2667 -12388
rect 2811 -12132 2845 -12116
rect 2811 -12404 2845 -12388
rect 2989 -12132 3023 -12116
rect 2989 -12404 3023 -12388
rect 3167 -12132 3201 -12116
rect 3167 -12404 3201 -12388
rect 3345 -12132 3379 -12116
rect 3345 -12404 3379 -12388
rect 3523 -12132 3557 -12116
rect 3523 -12404 3557 -12388
rect 3701 -12132 3735 -12116
rect 3701 -12404 3735 -12388
rect 3879 -12132 3913 -12116
rect 3879 -12404 3913 -12388
rect 4057 -12132 4091 -12116
rect 4057 -12404 4091 -12388
rect -2105 -12472 -2089 -12438
rect -2045 -12472 -2029 -12438
rect -1927 -12472 -1911 -12438
rect -1867 -12472 -1851 -12438
rect -1749 -12472 -1733 -12438
rect -1689 -12472 -1673 -12438
rect -1571 -12472 -1555 -12438
rect -1511 -12472 -1495 -12438
rect -1393 -12472 -1377 -12438
rect -1333 -12472 -1317 -12438
rect -1215 -12472 -1199 -12438
rect -1155 -12472 -1139 -12438
rect -1037 -12472 -1021 -12438
rect -977 -12472 -961 -12438
rect -859 -12472 -843 -12438
rect -799 -12472 -783 -12438
rect -681 -12472 -665 -12438
rect -621 -12472 -605 -12438
rect -503 -12472 -487 -12438
rect -443 -12472 -427 -12438
rect -325 -12472 -309 -12438
rect -265 -12472 -249 -12438
rect -147 -12472 -131 -12438
rect -87 -12472 -71 -12438
rect 31 -12472 47 -12438
rect 91 -12472 107 -12438
rect 209 -12472 225 -12438
rect 269 -12472 285 -12438
rect 387 -12472 403 -12438
rect 447 -12472 463 -12438
rect 565 -12472 581 -12438
rect 625 -12472 641 -12438
rect 743 -12472 759 -12438
rect 803 -12472 819 -12438
rect 921 -12472 937 -12438
rect 981 -12472 997 -12438
rect 1099 -12472 1115 -12438
rect 1159 -12472 1175 -12438
rect 1277 -12472 1293 -12438
rect 1337 -12472 1353 -12438
rect 1455 -12472 1471 -12438
rect 1515 -12472 1531 -12438
rect 1633 -12472 1649 -12438
rect 1693 -12472 1709 -12438
rect 1811 -12472 1827 -12438
rect 1871 -12472 1887 -12438
rect 1989 -12472 2005 -12438
rect 2049 -12472 2065 -12438
rect 2167 -12472 2183 -12438
rect 2227 -12472 2243 -12438
rect 2345 -12472 2361 -12438
rect 2405 -12472 2421 -12438
rect 2523 -12472 2539 -12438
rect 2583 -12472 2599 -12438
rect 2701 -12472 2717 -12438
rect 2761 -12472 2777 -12438
rect 2879 -12472 2895 -12438
rect 2939 -12472 2955 -12438
rect 3057 -12472 3073 -12438
rect 3117 -12472 3133 -12438
rect 3235 -12472 3251 -12438
rect 3295 -12472 3311 -12438
rect 3413 -12472 3429 -12438
rect 3473 -12472 3489 -12438
rect 3591 -12472 3607 -12438
rect 3651 -12472 3667 -12438
rect 3769 -12472 3785 -12438
rect 3829 -12472 3845 -12438
rect 3947 -12472 3963 -12438
rect 4007 -12472 4023 -12438
rect 8413 -12554 8639 -12530
rect -5883 -12662 -5867 -12628
rect -5833 -12662 -5817 -12628
rect -5633 -12662 -5617 -12628
rect -5583 -12662 -5567 -12628
rect -5383 -12662 -5367 -12628
rect -5333 -12662 -5317 -12628
rect -5133 -12662 -5117 -12628
rect -5083 -12662 -5067 -12628
rect -4883 -12662 -4867 -12628
rect -4833 -12662 -4817 -12628
rect -4633 -12662 -4617 -12628
rect -4583 -12662 -4567 -12628
rect -4383 -12662 -4367 -12628
rect -4333 -12662 -4317 -12628
rect -4133 -12662 -4117 -12628
rect -4083 -12662 -4067 -12628
rect -5917 -12712 -5883 -12696
rect -5917 -12944 -5883 -12928
rect -5817 -12712 -5783 -12696
rect -5817 -12944 -5783 -12928
rect -5667 -12712 -5633 -12696
rect -5667 -12944 -5633 -12928
rect -5567 -12712 -5533 -12696
rect -5567 -12944 -5533 -12928
rect -5417 -12712 -5383 -12696
rect -5417 -12944 -5383 -12928
rect -5317 -12712 -5283 -12696
rect -5317 -12944 -5283 -12928
rect -5167 -12712 -5133 -12696
rect -5167 -12944 -5133 -12928
rect -5067 -12712 -5033 -12696
rect -5067 -12944 -5033 -12928
rect -4917 -12712 -4883 -12696
rect -4917 -12944 -4883 -12928
rect -4817 -12712 -4783 -12696
rect -4817 -12944 -4783 -12928
rect -4667 -12712 -4633 -12696
rect -4667 -12944 -4633 -12928
rect -4567 -12712 -4533 -12696
rect -4567 -12944 -4533 -12928
rect -4417 -12712 -4383 -12696
rect -4417 -12944 -4383 -12928
rect -4317 -12712 -4283 -12696
rect -4317 -12944 -4283 -12928
rect -4167 -12712 -4133 -12696
rect -4167 -12944 -4133 -12928
rect -4067 -12712 -4033 -12696
rect 8413 -12732 8437 -12554
rect 8615 -12732 8639 -12554
rect 8413 -12756 8639 -12732
rect 11413 -12554 11639 -12530
rect 11413 -12732 11437 -12554
rect 11615 -12732 11639 -12554
rect 11413 -12756 11639 -12732
rect -4067 -12944 -4033 -12928
rect -5883 -13012 -5867 -12978
rect -5833 -13012 -5817 -12978
rect -5633 -13012 -5617 -12978
rect -5583 -13012 -5567 -12978
rect -5383 -13012 -5367 -12978
rect -5333 -13012 -5317 -12978
rect -5133 -13012 -5117 -12978
rect -5083 -13012 -5067 -12978
rect -4883 -13012 -4867 -12978
rect -4833 -13012 -4817 -12978
rect -4633 -13012 -4617 -12978
rect -4583 -13012 -4567 -12978
rect -4383 -13012 -4367 -12978
rect -4333 -13012 -4317 -12978
rect -4133 -13012 -4117 -12978
rect -4083 -13012 -4067 -12978
rect -2105 -13082 -2089 -13048
rect -2045 -13082 -2029 -13048
rect -1927 -13082 -1911 -13048
rect -1867 -13082 -1851 -13048
rect -1749 -13082 -1733 -13048
rect -1689 -13082 -1673 -13048
rect -1571 -13082 -1555 -13048
rect -1511 -13082 -1495 -13048
rect -1393 -13082 -1377 -13048
rect -1333 -13082 -1317 -13048
rect -1215 -13082 -1199 -13048
rect -1155 -13082 -1139 -13048
rect -1037 -13082 -1021 -13048
rect -977 -13082 -961 -13048
rect -859 -13082 -843 -13048
rect -799 -13082 -783 -13048
rect -681 -13082 -665 -13048
rect -621 -13082 -605 -13048
rect -503 -13082 -487 -13048
rect -443 -13082 -427 -13048
rect -325 -13082 -309 -13048
rect -265 -13082 -249 -13048
rect -147 -13082 -131 -13048
rect -87 -13082 -71 -13048
rect 31 -13082 47 -13048
rect 91 -13082 107 -13048
rect 209 -13082 225 -13048
rect 269 -13082 285 -13048
rect 387 -13082 403 -13048
rect 447 -13082 463 -13048
rect 565 -13082 581 -13048
rect 625 -13082 641 -13048
rect 743 -13082 759 -13048
rect 803 -13082 819 -13048
rect 921 -13082 937 -13048
rect 981 -13082 997 -13048
rect 1099 -13082 1115 -13048
rect 1159 -13082 1175 -13048
rect 1277 -13082 1293 -13048
rect 1337 -13082 1353 -13048
rect 1455 -13082 1471 -13048
rect 1515 -13082 1531 -13048
rect 1633 -13082 1649 -13048
rect 1693 -13082 1709 -13048
rect 1811 -13082 1827 -13048
rect 1871 -13082 1887 -13048
rect 1989 -13082 2005 -13048
rect 2049 -13082 2065 -13048
rect 2167 -13082 2183 -13048
rect 2227 -13082 2243 -13048
rect 2345 -13082 2361 -13048
rect 2405 -13082 2421 -13048
rect 2523 -13082 2539 -13048
rect 2583 -13082 2599 -13048
rect 2701 -13082 2717 -13048
rect 2761 -13082 2777 -13048
rect 2879 -13082 2895 -13048
rect 2939 -13082 2955 -13048
rect 3057 -13082 3073 -13048
rect 3117 -13082 3133 -13048
rect 3235 -13082 3251 -13048
rect 3295 -13082 3311 -13048
rect 3413 -13082 3429 -13048
rect 3473 -13082 3489 -13048
rect 3591 -13082 3607 -13048
rect 3651 -13082 3667 -13048
rect 3769 -13082 3785 -13048
rect 3829 -13082 3845 -13048
rect 3947 -13082 3963 -13048
rect 4007 -13082 4023 -13048
rect -2173 -13132 -2139 -13116
rect -3009 -13276 -2783 -13252
rect -5883 -13342 -5867 -13308
rect -5833 -13342 -5817 -13308
rect -5633 -13342 -5617 -13308
rect -5583 -13342 -5567 -13308
rect -5383 -13342 -5367 -13308
rect -5333 -13342 -5317 -13308
rect -5133 -13342 -5117 -13308
rect -5083 -13342 -5067 -13308
rect -4883 -13342 -4867 -13308
rect -4833 -13342 -4817 -13308
rect -4633 -13342 -4617 -13308
rect -4583 -13342 -4567 -13308
rect -4383 -13342 -4367 -13308
rect -4333 -13342 -4317 -13308
rect -4133 -13342 -4117 -13308
rect -4083 -13342 -4067 -13308
rect -5917 -13392 -5883 -13376
rect -5917 -13624 -5883 -13608
rect -5817 -13392 -5783 -13376
rect -5817 -13624 -5783 -13608
rect -5667 -13392 -5633 -13376
rect -5667 -13624 -5633 -13608
rect -5567 -13392 -5533 -13376
rect -5567 -13624 -5533 -13608
rect -5417 -13392 -5383 -13376
rect -5417 -13624 -5383 -13608
rect -5317 -13392 -5283 -13376
rect -5317 -13624 -5283 -13608
rect -5167 -13392 -5133 -13376
rect -5167 -13624 -5133 -13608
rect -5067 -13392 -5033 -13376
rect -5067 -13624 -5033 -13608
rect -4917 -13392 -4883 -13376
rect -4917 -13624 -4883 -13608
rect -4817 -13392 -4783 -13376
rect -4817 -13624 -4783 -13608
rect -4667 -13392 -4633 -13376
rect -4667 -13624 -4633 -13608
rect -4567 -13392 -4533 -13376
rect -4567 -13624 -4533 -13608
rect -4417 -13392 -4383 -13376
rect -4417 -13624 -4383 -13608
rect -4317 -13392 -4283 -13376
rect -4317 -13624 -4283 -13608
rect -4167 -13392 -4133 -13376
rect -4167 -13624 -4133 -13608
rect -4067 -13392 -4033 -13376
rect -3009 -13454 -2985 -13276
rect -2807 -13454 -2783 -13276
rect -2173 -13404 -2139 -13388
rect -1995 -13132 -1961 -13116
rect -1995 -13404 -1961 -13388
rect -1817 -13132 -1783 -13116
rect -1817 -13404 -1783 -13388
rect -1639 -13132 -1605 -13116
rect -1639 -13404 -1605 -13388
rect -1461 -13132 -1427 -13116
rect -1461 -13404 -1427 -13388
rect -1283 -13132 -1249 -13116
rect -1283 -13404 -1249 -13388
rect -1105 -13132 -1071 -13116
rect -1105 -13404 -1071 -13388
rect -927 -13132 -893 -13116
rect -927 -13404 -893 -13388
rect -749 -13132 -715 -13116
rect -749 -13404 -715 -13388
rect -571 -13132 -537 -13116
rect -571 -13404 -537 -13388
rect -393 -13132 -359 -13116
rect -393 -13404 -359 -13388
rect -215 -13132 -181 -13116
rect -215 -13404 -181 -13388
rect -37 -13132 -3 -13116
rect -37 -13404 -3 -13388
rect 141 -13132 175 -13116
rect 141 -13404 175 -13388
rect 319 -13132 353 -13116
rect 319 -13404 353 -13388
rect 497 -13132 531 -13116
rect 497 -13404 531 -13388
rect 675 -13132 709 -13116
rect 675 -13404 709 -13388
rect 853 -13132 887 -13116
rect 853 -13404 887 -13388
rect 1031 -13132 1065 -13116
rect 1031 -13404 1065 -13388
rect 1209 -13132 1243 -13116
rect 1209 -13404 1243 -13388
rect 1387 -13132 1421 -13116
rect 1387 -13404 1421 -13388
rect 1565 -13132 1599 -13116
rect 1565 -13404 1599 -13388
rect 1743 -13132 1777 -13116
rect 1743 -13404 1777 -13388
rect 1921 -13132 1955 -13116
rect 1921 -13404 1955 -13388
rect 2099 -13132 2133 -13116
rect 2099 -13404 2133 -13388
rect 2277 -13132 2311 -13116
rect 2277 -13404 2311 -13388
rect 2455 -13132 2489 -13116
rect 2455 -13404 2489 -13388
rect 2633 -13132 2667 -13116
rect 2633 -13404 2667 -13388
rect 2811 -13132 2845 -13116
rect 2811 -13404 2845 -13388
rect 2989 -13132 3023 -13116
rect 2989 -13404 3023 -13388
rect 3167 -13132 3201 -13116
rect 3167 -13404 3201 -13388
rect 3345 -13132 3379 -13116
rect 3345 -13404 3379 -13388
rect 3523 -13132 3557 -13116
rect 3523 -13404 3557 -13388
rect 3701 -13132 3735 -13116
rect 3701 -13404 3735 -13388
rect 3879 -13132 3913 -13116
rect 3879 -13404 3913 -13388
rect 4057 -13132 4091 -13116
rect 4057 -13404 4091 -13388
rect -3009 -13478 -2783 -13454
rect -2105 -13472 -2089 -13438
rect -2045 -13472 -2029 -13438
rect -1927 -13472 -1911 -13438
rect -1867 -13472 -1851 -13438
rect -1749 -13472 -1733 -13438
rect -1689 -13472 -1673 -13438
rect -1571 -13472 -1555 -13438
rect -1511 -13472 -1495 -13438
rect -1393 -13472 -1377 -13438
rect -1333 -13472 -1317 -13438
rect -1215 -13472 -1199 -13438
rect -1155 -13472 -1139 -13438
rect -1037 -13472 -1021 -13438
rect -977 -13472 -961 -13438
rect -859 -13472 -843 -13438
rect -799 -13472 -783 -13438
rect -681 -13472 -665 -13438
rect -621 -13472 -605 -13438
rect -503 -13472 -487 -13438
rect -443 -13472 -427 -13438
rect -325 -13472 -309 -13438
rect -265 -13472 -249 -13438
rect -147 -13472 -131 -13438
rect -87 -13472 -71 -13438
rect 31 -13472 47 -13438
rect 91 -13472 107 -13438
rect 209 -13472 225 -13438
rect 269 -13472 285 -13438
rect 387 -13472 403 -13438
rect 447 -13472 463 -13438
rect 565 -13472 581 -13438
rect 625 -13472 641 -13438
rect 743 -13472 759 -13438
rect 803 -13472 819 -13438
rect 921 -13472 937 -13438
rect 981 -13472 997 -13438
rect 1099 -13472 1115 -13438
rect 1159 -13472 1175 -13438
rect 1277 -13472 1293 -13438
rect 1337 -13472 1353 -13438
rect 1455 -13472 1471 -13438
rect 1515 -13472 1531 -13438
rect 1633 -13472 1649 -13438
rect 1693 -13472 1709 -13438
rect 1811 -13472 1827 -13438
rect 1871 -13472 1887 -13438
rect 1989 -13472 2005 -13438
rect 2049 -13472 2065 -13438
rect 2167 -13472 2183 -13438
rect 2227 -13472 2243 -13438
rect 2345 -13472 2361 -13438
rect 2405 -13472 2421 -13438
rect 2523 -13472 2539 -13438
rect 2583 -13472 2599 -13438
rect 2701 -13472 2717 -13438
rect 2761 -13472 2777 -13438
rect 2879 -13472 2895 -13438
rect 2939 -13472 2955 -13438
rect 3057 -13472 3073 -13438
rect 3117 -13472 3133 -13438
rect 3235 -13472 3251 -13438
rect 3295 -13472 3311 -13438
rect 3413 -13472 3429 -13438
rect 3473 -13472 3489 -13438
rect 3591 -13472 3607 -13438
rect 3651 -13472 3667 -13438
rect 3769 -13472 3785 -13438
rect 3829 -13472 3845 -13438
rect 3947 -13472 3963 -13438
rect 4007 -13472 4023 -13438
rect -4067 -13624 -4033 -13608
rect -5883 -13692 -5867 -13658
rect -5833 -13692 -5817 -13658
rect -5633 -13692 -5617 -13658
rect -5583 -13692 -5567 -13658
rect -5383 -13692 -5367 -13658
rect -5333 -13692 -5317 -13658
rect -5133 -13692 -5117 -13658
rect -5083 -13692 -5067 -13658
rect -4883 -13692 -4867 -13658
rect -4833 -13692 -4817 -13658
rect -4633 -13692 -4617 -13658
rect -4583 -13692 -4567 -13658
rect -4383 -13692 -4367 -13658
rect -4333 -13692 -4317 -13658
rect -4133 -13692 -4117 -13658
rect -4083 -13692 -4067 -13658
rect -2105 -14082 -2089 -14048
rect -2045 -14082 -2029 -14048
rect -1927 -14082 -1911 -14048
rect -1867 -14082 -1851 -14048
rect -1749 -14082 -1733 -14048
rect -1689 -14082 -1673 -14048
rect -1571 -14082 -1555 -14048
rect -1511 -14082 -1495 -14048
rect -1393 -14082 -1377 -14048
rect -1333 -14082 -1317 -14048
rect -1215 -14082 -1199 -14048
rect -1155 -14082 -1139 -14048
rect -1037 -14082 -1021 -14048
rect -977 -14082 -961 -14048
rect -859 -14082 -843 -14048
rect -799 -14082 -783 -14048
rect -681 -14082 -665 -14048
rect -621 -14082 -605 -14048
rect -503 -14082 -487 -14048
rect -443 -14082 -427 -14048
rect -325 -14082 -309 -14048
rect -265 -14082 -249 -14048
rect -147 -14082 -131 -14048
rect -87 -14082 -71 -14048
rect 31 -14082 47 -14048
rect 91 -14082 107 -14048
rect 209 -14082 225 -14048
rect 269 -14082 285 -14048
rect 387 -14082 403 -14048
rect 447 -14082 463 -14048
rect 565 -14082 581 -14048
rect 625 -14082 641 -14048
rect 743 -14082 759 -14048
rect 803 -14082 819 -14048
rect 921 -14082 937 -14048
rect 981 -14082 997 -14048
rect 1099 -14082 1115 -14048
rect 1159 -14082 1175 -14048
rect 1277 -14082 1293 -14048
rect 1337 -14082 1353 -14048
rect 1455 -14082 1471 -14048
rect 1515 -14082 1531 -14048
rect 1633 -14082 1649 -14048
rect 1693 -14082 1709 -14048
rect 1811 -14082 1827 -14048
rect 1871 -14082 1887 -14048
rect 1989 -14082 2005 -14048
rect 2049 -14082 2065 -14048
rect 2167 -14082 2183 -14048
rect 2227 -14082 2243 -14048
rect 2345 -14082 2361 -14048
rect 2405 -14082 2421 -14048
rect 2523 -14082 2539 -14048
rect 2583 -14082 2599 -14048
rect 2701 -14082 2717 -14048
rect 2761 -14082 2777 -14048
rect 2879 -14082 2895 -14048
rect 2939 -14082 2955 -14048
rect 3057 -14082 3073 -14048
rect 3117 -14082 3133 -14048
rect 3235 -14082 3251 -14048
rect 3295 -14082 3311 -14048
rect 3413 -14082 3429 -14048
rect 3473 -14082 3489 -14048
rect 3591 -14082 3607 -14048
rect 3651 -14082 3667 -14048
rect 3769 -14082 3785 -14048
rect 3829 -14082 3845 -14048
rect 3947 -14082 3963 -14048
rect 4007 -14082 4023 -14048
rect 5645 -14082 5661 -14048
rect 5705 -14082 5721 -14048
rect 5823 -14082 5839 -14048
rect 5883 -14082 5899 -14048
rect 6001 -14082 6017 -14048
rect 6061 -14082 6077 -14048
rect 6179 -14082 6195 -14048
rect 6239 -14082 6255 -14048
rect 6357 -14082 6373 -14048
rect 6417 -14082 6433 -14048
rect 6535 -14082 6551 -14048
rect 6595 -14082 6611 -14048
rect 6713 -14082 6729 -14048
rect 6773 -14082 6789 -14048
rect 6891 -14082 6907 -14048
rect 6951 -14082 6967 -14048
rect 7069 -14082 7085 -14048
rect 7129 -14082 7145 -14048
rect 7247 -14082 7263 -14048
rect 7307 -14082 7323 -14048
rect 7425 -14082 7441 -14048
rect 7485 -14082 7501 -14048
rect 7603 -14082 7619 -14048
rect 7663 -14082 7679 -14048
rect 7781 -14082 7797 -14048
rect 7841 -14082 7857 -14048
rect 7959 -14082 7975 -14048
rect 8019 -14082 8035 -14048
rect 8137 -14082 8153 -14048
rect 8197 -14082 8213 -14048
rect 8315 -14082 8331 -14048
rect 8375 -14082 8391 -14048
rect 8493 -14082 8509 -14048
rect 8553 -14082 8569 -14048
rect 8671 -14082 8687 -14048
rect 8731 -14082 8747 -14048
rect 8849 -14082 8865 -14048
rect 8909 -14082 8925 -14048
rect 9027 -14082 9043 -14048
rect 9087 -14082 9103 -14048
rect 9205 -14082 9221 -14048
rect 9265 -14082 9281 -14048
rect 9383 -14082 9399 -14048
rect 9443 -14082 9459 -14048
rect 9561 -14082 9577 -14048
rect 9621 -14082 9637 -14048
rect 9739 -14082 9755 -14048
rect 9799 -14082 9815 -14048
rect 9917 -14082 9933 -14048
rect 9977 -14082 9993 -14048
rect 10095 -14082 10111 -14048
rect 10155 -14082 10171 -14048
rect 10273 -14082 10289 -14048
rect 10333 -14082 10349 -14048
rect 10451 -14082 10467 -14048
rect 10511 -14082 10527 -14048
rect 10629 -14082 10645 -14048
rect 10689 -14082 10705 -14048
rect 10807 -14082 10823 -14048
rect 10867 -14082 10883 -14048
rect 10985 -14082 11001 -14048
rect 11045 -14082 11061 -14048
rect 11163 -14082 11179 -14048
rect 11223 -14082 11239 -14048
rect 11341 -14082 11357 -14048
rect 11401 -14082 11417 -14048
rect 11519 -14082 11535 -14048
rect 11579 -14082 11595 -14048
rect 11697 -14082 11713 -14048
rect 11757 -14082 11773 -14048
rect 11875 -14082 11891 -14048
rect 11935 -14082 11951 -14048
rect 12053 -14082 12069 -14048
rect 12113 -14082 12129 -14048
rect 12231 -14082 12247 -14048
rect 12291 -14082 12307 -14048
rect 12409 -14082 12425 -14048
rect 12469 -14082 12485 -14048
rect 12587 -14082 12603 -14048
rect 12647 -14082 12663 -14048
rect -2173 -14132 -2139 -14116
rect -5960 -14344 -5944 -14310
rect -5900 -14344 -5884 -14310
rect -5782 -14344 -5766 -14310
rect -5722 -14344 -5706 -14310
rect -5604 -14344 -5588 -14310
rect -5544 -14344 -5528 -14310
rect -5426 -14344 -5410 -14310
rect -5366 -14344 -5350 -14310
rect -5248 -14344 -5232 -14310
rect -5188 -14344 -5172 -14310
rect -5070 -14344 -5054 -14310
rect -5010 -14344 -4994 -14310
rect -4892 -14344 -4876 -14310
rect -4832 -14344 -4816 -14310
rect -4714 -14344 -4698 -14310
rect -4654 -14344 -4638 -14310
rect -4536 -14344 -4520 -14310
rect -4476 -14344 -4460 -14310
rect -4358 -14344 -4342 -14310
rect -4298 -14344 -4282 -14310
rect -4180 -14344 -4164 -14310
rect -4120 -14344 -4104 -14310
rect -6028 -14394 -5994 -14378
rect -6028 -14666 -5994 -14650
rect -5850 -14394 -5816 -14378
rect -5850 -14666 -5816 -14650
rect -5672 -14394 -5638 -14378
rect -5672 -14666 -5638 -14650
rect -5494 -14394 -5460 -14378
rect -5494 -14666 -5460 -14650
rect -5316 -14394 -5282 -14378
rect -5316 -14666 -5282 -14650
rect -5138 -14394 -5104 -14378
rect -5138 -14666 -5104 -14650
rect -4960 -14394 -4926 -14378
rect -4960 -14666 -4926 -14650
rect -4782 -14394 -4748 -14378
rect -4782 -14666 -4748 -14650
rect -4604 -14394 -4570 -14378
rect -4604 -14666 -4570 -14650
rect -4426 -14394 -4392 -14378
rect -4426 -14666 -4392 -14650
rect -4248 -14394 -4214 -14378
rect -4248 -14666 -4214 -14650
rect -4070 -14394 -4036 -14378
rect -2173 -14404 -2139 -14388
rect -1995 -14132 -1961 -14116
rect -1995 -14404 -1961 -14388
rect -1817 -14132 -1783 -14116
rect -1817 -14404 -1783 -14388
rect -1639 -14132 -1605 -14116
rect -1639 -14404 -1605 -14388
rect -1461 -14132 -1427 -14116
rect -1461 -14404 -1427 -14388
rect -1283 -14132 -1249 -14116
rect -1283 -14404 -1249 -14388
rect -1105 -14132 -1071 -14116
rect -1105 -14404 -1071 -14388
rect -927 -14132 -893 -14116
rect -927 -14404 -893 -14388
rect -749 -14132 -715 -14116
rect -749 -14404 -715 -14388
rect -571 -14132 -537 -14116
rect -571 -14404 -537 -14388
rect -393 -14132 -359 -14116
rect -393 -14404 -359 -14388
rect -215 -14132 -181 -14116
rect -215 -14404 -181 -14388
rect -37 -14132 -3 -14116
rect -37 -14404 -3 -14388
rect 141 -14132 175 -14116
rect 141 -14404 175 -14388
rect 319 -14132 353 -14116
rect 319 -14404 353 -14388
rect 497 -14132 531 -14116
rect 497 -14404 531 -14388
rect 675 -14132 709 -14116
rect 675 -14404 709 -14388
rect 853 -14132 887 -14116
rect 853 -14404 887 -14388
rect 1031 -14132 1065 -14116
rect 1031 -14404 1065 -14388
rect 1209 -14132 1243 -14116
rect 1209 -14404 1243 -14388
rect 1387 -14132 1421 -14116
rect 1387 -14404 1421 -14388
rect 1565 -14132 1599 -14116
rect 1565 -14404 1599 -14388
rect 1743 -14132 1777 -14116
rect 1743 -14404 1777 -14388
rect 1921 -14132 1955 -14116
rect 1921 -14404 1955 -14388
rect 2099 -14132 2133 -14116
rect 2099 -14404 2133 -14388
rect 2277 -14132 2311 -14116
rect 2277 -14404 2311 -14388
rect 2455 -14132 2489 -14116
rect 2455 -14404 2489 -14388
rect 2633 -14132 2667 -14116
rect 2633 -14404 2667 -14388
rect 2811 -14132 2845 -14116
rect 2811 -14404 2845 -14388
rect 2989 -14132 3023 -14116
rect 2989 -14404 3023 -14388
rect 3167 -14132 3201 -14116
rect 3167 -14404 3201 -14388
rect 3345 -14132 3379 -14116
rect 3345 -14404 3379 -14388
rect 3523 -14132 3557 -14116
rect 3523 -14404 3557 -14388
rect 3701 -14132 3735 -14116
rect 3701 -14404 3735 -14388
rect 3879 -14132 3913 -14116
rect 3879 -14404 3913 -14388
rect 4057 -14132 4091 -14116
rect 4057 -14404 4091 -14388
rect 5577 -14132 5611 -14116
rect 5577 -14404 5611 -14388
rect 5755 -14132 5789 -14116
rect 5755 -14404 5789 -14388
rect 5933 -14132 5967 -14116
rect 5933 -14404 5967 -14388
rect 6111 -14132 6145 -14116
rect 6111 -14404 6145 -14388
rect 6289 -14132 6323 -14116
rect 6289 -14404 6323 -14388
rect 6467 -14132 6501 -14116
rect 6467 -14404 6501 -14388
rect 6645 -14132 6679 -14116
rect 6645 -14404 6679 -14388
rect 6823 -14132 6857 -14116
rect 6823 -14404 6857 -14388
rect 7001 -14132 7035 -14116
rect 7001 -14404 7035 -14388
rect 7179 -14132 7213 -14116
rect 7179 -14404 7213 -14388
rect 7357 -14132 7391 -14116
rect 7357 -14404 7391 -14388
rect 7535 -14132 7569 -14116
rect 7535 -14404 7569 -14388
rect 7713 -14132 7747 -14116
rect 7713 -14404 7747 -14388
rect 7891 -14132 7925 -14116
rect 7891 -14404 7925 -14388
rect 8069 -14132 8103 -14116
rect 8069 -14404 8103 -14388
rect 8247 -14132 8281 -14116
rect 8247 -14404 8281 -14388
rect 8425 -14132 8459 -14116
rect 8425 -14404 8459 -14388
rect 8603 -14132 8637 -14116
rect 8603 -14404 8637 -14388
rect 8781 -14132 8815 -14116
rect 8781 -14404 8815 -14388
rect 8959 -14132 8993 -14116
rect 8959 -14404 8993 -14388
rect 9137 -14132 9171 -14116
rect 9137 -14404 9171 -14388
rect 9315 -14132 9349 -14116
rect 9315 -14404 9349 -14388
rect 9493 -14132 9527 -14116
rect 9493 -14404 9527 -14388
rect 9671 -14132 9705 -14116
rect 9671 -14404 9705 -14388
rect 9849 -14132 9883 -14116
rect 9849 -14404 9883 -14388
rect 10027 -14132 10061 -14116
rect 10027 -14404 10061 -14388
rect 10205 -14132 10239 -14116
rect 10205 -14404 10239 -14388
rect 10383 -14132 10417 -14116
rect 10383 -14404 10417 -14388
rect 10561 -14132 10595 -14116
rect 10561 -14404 10595 -14388
rect 10739 -14132 10773 -14116
rect 10739 -14404 10773 -14388
rect 10917 -14132 10951 -14116
rect 10917 -14404 10951 -14388
rect 11095 -14132 11129 -14116
rect 11095 -14404 11129 -14388
rect 11273 -14132 11307 -14116
rect 11273 -14404 11307 -14388
rect 11451 -14132 11485 -14116
rect 11451 -14404 11485 -14388
rect 11629 -14132 11663 -14116
rect 11629 -14404 11663 -14388
rect 11807 -14132 11841 -14116
rect 11807 -14404 11841 -14388
rect 11985 -14132 12019 -14116
rect 11985 -14404 12019 -14388
rect 12163 -14132 12197 -14116
rect 12163 -14404 12197 -14388
rect 12341 -14132 12375 -14116
rect 12341 -14404 12375 -14388
rect 12519 -14132 12553 -14116
rect 12519 -14404 12553 -14388
rect 12697 -14132 12731 -14116
rect 12697 -14404 12731 -14388
rect -2105 -14472 -2089 -14438
rect -2045 -14472 -2029 -14438
rect -1927 -14472 -1911 -14438
rect -1867 -14472 -1851 -14438
rect -1749 -14472 -1733 -14438
rect -1689 -14472 -1673 -14438
rect -1571 -14472 -1555 -14438
rect -1511 -14472 -1495 -14438
rect -1393 -14472 -1377 -14438
rect -1333 -14472 -1317 -14438
rect -1215 -14472 -1199 -14438
rect -1155 -14472 -1139 -14438
rect -1037 -14472 -1021 -14438
rect -977 -14472 -961 -14438
rect -859 -14472 -843 -14438
rect -799 -14472 -783 -14438
rect -681 -14472 -665 -14438
rect -621 -14472 -605 -14438
rect -503 -14472 -487 -14438
rect -443 -14472 -427 -14438
rect -325 -14472 -309 -14438
rect -265 -14472 -249 -14438
rect -147 -14472 -131 -14438
rect -87 -14472 -71 -14438
rect 31 -14472 47 -14438
rect 91 -14472 107 -14438
rect 209 -14472 225 -14438
rect 269 -14472 285 -14438
rect 387 -14472 403 -14438
rect 447 -14472 463 -14438
rect 565 -14472 581 -14438
rect 625 -14472 641 -14438
rect 743 -14472 759 -14438
rect 803 -14472 819 -14438
rect 921 -14472 937 -14438
rect 981 -14472 997 -14438
rect 1099 -14472 1115 -14438
rect 1159 -14472 1175 -14438
rect 1277 -14472 1293 -14438
rect 1337 -14472 1353 -14438
rect 1455 -14472 1471 -14438
rect 1515 -14472 1531 -14438
rect 1633 -14472 1649 -14438
rect 1693 -14472 1709 -14438
rect 1811 -14472 1827 -14438
rect 1871 -14472 1887 -14438
rect 1989 -14472 2005 -14438
rect 2049 -14472 2065 -14438
rect 2167 -14472 2183 -14438
rect 2227 -14472 2243 -14438
rect 2345 -14472 2361 -14438
rect 2405 -14472 2421 -14438
rect 2523 -14472 2539 -14438
rect 2583 -14472 2599 -14438
rect 2701 -14472 2717 -14438
rect 2761 -14472 2777 -14438
rect 2879 -14472 2895 -14438
rect 2939 -14472 2955 -14438
rect 3057 -14472 3073 -14438
rect 3117 -14472 3133 -14438
rect 3235 -14472 3251 -14438
rect 3295 -14472 3311 -14438
rect 3413 -14472 3429 -14438
rect 3473 -14472 3489 -14438
rect 3591 -14472 3607 -14438
rect 3651 -14472 3667 -14438
rect 3769 -14472 3785 -14438
rect 3829 -14472 3845 -14438
rect 3947 -14472 3963 -14438
rect 4007 -14472 4023 -14438
rect 5645 -14472 5661 -14438
rect 5705 -14472 5721 -14438
rect 5823 -14472 5839 -14438
rect 5883 -14472 5899 -14438
rect 6001 -14472 6017 -14438
rect 6061 -14472 6077 -14438
rect 6179 -14472 6195 -14438
rect 6239 -14472 6255 -14438
rect 6357 -14472 6373 -14438
rect 6417 -14472 6433 -14438
rect 6535 -14472 6551 -14438
rect 6595 -14472 6611 -14438
rect 6713 -14472 6729 -14438
rect 6773 -14472 6789 -14438
rect 6891 -14472 6907 -14438
rect 6951 -14472 6967 -14438
rect 7069 -14472 7085 -14438
rect 7129 -14472 7145 -14438
rect 7247 -14472 7263 -14438
rect 7307 -14472 7323 -14438
rect 7425 -14472 7441 -14438
rect 7485 -14472 7501 -14438
rect 7603 -14472 7619 -14438
rect 7663 -14472 7679 -14438
rect 7781 -14472 7797 -14438
rect 7841 -14472 7857 -14438
rect 7959 -14472 7975 -14438
rect 8019 -14472 8035 -14438
rect 8137 -14472 8153 -14438
rect 8197 -14472 8213 -14438
rect 8315 -14472 8331 -14438
rect 8375 -14472 8391 -14438
rect 8493 -14472 8509 -14438
rect 8553 -14472 8569 -14438
rect 8671 -14472 8687 -14438
rect 8731 -14472 8747 -14438
rect 8849 -14472 8865 -14438
rect 8909 -14472 8925 -14438
rect 9027 -14472 9043 -14438
rect 9087 -14472 9103 -14438
rect 9205 -14472 9221 -14438
rect 9265 -14472 9281 -14438
rect 9383 -14472 9399 -14438
rect 9443 -14472 9459 -14438
rect 9561 -14472 9577 -14438
rect 9621 -14472 9637 -14438
rect 9739 -14472 9755 -14438
rect 9799 -14472 9815 -14438
rect 9917 -14472 9933 -14438
rect 9977 -14472 9993 -14438
rect 10095 -14472 10111 -14438
rect 10155 -14472 10171 -14438
rect 10273 -14472 10289 -14438
rect 10333 -14472 10349 -14438
rect 10451 -14472 10467 -14438
rect 10511 -14472 10527 -14438
rect 10629 -14472 10645 -14438
rect 10689 -14472 10705 -14438
rect 10807 -14472 10823 -14438
rect 10867 -14472 10883 -14438
rect 10985 -14472 11001 -14438
rect 11045 -14472 11061 -14438
rect 11163 -14472 11179 -14438
rect 11223 -14472 11239 -14438
rect 11341 -14472 11357 -14438
rect 11401 -14472 11417 -14438
rect 11519 -14472 11535 -14438
rect 11579 -14472 11595 -14438
rect 11697 -14472 11713 -14438
rect 11757 -14472 11773 -14438
rect 11875 -14472 11891 -14438
rect 11935 -14472 11951 -14438
rect 12053 -14472 12069 -14438
rect 12113 -14472 12129 -14438
rect 12231 -14472 12247 -14438
rect 12291 -14472 12307 -14438
rect 12409 -14472 12425 -14438
rect 12469 -14472 12485 -14438
rect 12587 -14472 12603 -14438
rect 12647 -14472 12663 -14438
rect -4070 -14666 -4036 -14650
rect -5960 -14734 -5944 -14700
rect -5900 -14734 -5884 -14700
rect -5782 -14734 -5766 -14700
rect -5722 -14734 -5706 -14700
rect -5604 -14734 -5588 -14700
rect -5544 -14734 -5528 -14700
rect -5426 -14734 -5410 -14700
rect -5366 -14734 -5350 -14700
rect -5248 -14734 -5232 -14700
rect -5188 -14734 -5172 -14700
rect -5070 -14734 -5054 -14700
rect -5010 -14734 -4994 -14700
rect -4892 -14734 -4876 -14700
rect -4832 -14734 -4816 -14700
rect -4714 -14734 -4698 -14700
rect -4654 -14734 -4638 -14700
rect -4536 -14734 -4520 -14700
rect -4476 -14734 -4460 -14700
rect -4358 -14734 -4342 -14700
rect -4298 -14734 -4282 -14700
rect -4180 -14734 -4164 -14700
rect -4120 -14734 -4104 -14700
rect 4519 -14869 4745 -14845
rect -5960 -15044 -5944 -15010
rect -5900 -15044 -5884 -15010
rect -5782 -15044 -5766 -15010
rect -5722 -15044 -5706 -15010
rect -5604 -15044 -5588 -15010
rect -5544 -15044 -5528 -15010
rect -5426 -15044 -5410 -15010
rect -5366 -15044 -5350 -15010
rect -5248 -15044 -5232 -15010
rect -5188 -15044 -5172 -15010
rect -5070 -15044 -5054 -15010
rect -5010 -15044 -4994 -15010
rect -4892 -15044 -4876 -15010
rect -4832 -15044 -4816 -15010
rect -4714 -15044 -4698 -15010
rect -4654 -15044 -4638 -15010
rect -4536 -15044 -4520 -15010
rect -4476 -15044 -4460 -15010
rect -4358 -15044 -4342 -15010
rect -4298 -15044 -4282 -15010
rect -4180 -15044 -4164 -15010
rect -4120 -15044 -4104 -15010
rect 4519 -15047 4543 -14869
rect 4721 -15047 4745 -14869
rect -6028 -15094 -5994 -15078
rect -6028 -15366 -5994 -15350
rect -5850 -15094 -5816 -15078
rect -5850 -15366 -5816 -15350
rect -5672 -15094 -5638 -15078
rect -5672 -15366 -5638 -15350
rect -5494 -15094 -5460 -15078
rect -5494 -15366 -5460 -15350
rect -5316 -15094 -5282 -15078
rect -5316 -15366 -5282 -15350
rect -5138 -15094 -5104 -15078
rect -5138 -15366 -5104 -15350
rect -4960 -15094 -4926 -15078
rect -4960 -15366 -4926 -15350
rect -4782 -15094 -4748 -15078
rect -4782 -15366 -4748 -15350
rect -4604 -15094 -4570 -15078
rect -4604 -15366 -4570 -15350
rect -4426 -15094 -4392 -15078
rect -4426 -15366 -4392 -15350
rect -4248 -15094 -4214 -15078
rect -4248 -15366 -4214 -15350
rect -4070 -15094 -4036 -15078
rect -2105 -15082 -2089 -15048
rect -2045 -15082 -2029 -15048
rect -1927 -15082 -1911 -15048
rect -1867 -15082 -1851 -15048
rect -1749 -15082 -1733 -15048
rect -1689 -15082 -1673 -15048
rect -1571 -15082 -1555 -15048
rect -1511 -15082 -1495 -15048
rect -1393 -15082 -1377 -15048
rect -1333 -15082 -1317 -15048
rect -1215 -15082 -1199 -15048
rect -1155 -15082 -1139 -15048
rect -1037 -15082 -1021 -15048
rect -977 -15082 -961 -15048
rect -859 -15082 -843 -15048
rect -799 -15082 -783 -15048
rect -681 -15082 -665 -15048
rect -621 -15082 -605 -15048
rect -503 -15082 -487 -15048
rect -443 -15082 -427 -15048
rect -325 -15082 -309 -15048
rect -265 -15082 -249 -15048
rect -147 -15082 -131 -15048
rect -87 -15082 -71 -15048
rect 31 -15082 47 -15048
rect 91 -15082 107 -15048
rect 209 -15082 225 -15048
rect 269 -15082 285 -15048
rect 387 -15082 403 -15048
rect 447 -15082 463 -15048
rect 565 -15082 581 -15048
rect 625 -15082 641 -15048
rect 743 -15082 759 -15048
rect 803 -15082 819 -15048
rect 921 -15082 937 -15048
rect 981 -15082 997 -15048
rect 1099 -15082 1115 -15048
rect 1159 -15082 1175 -15048
rect 1277 -15082 1293 -15048
rect 1337 -15082 1353 -15048
rect 1455 -15082 1471 -15048
rect 1515 -15082 1531 -15048
rect 1633 -15082 1649 -15048
rect 1693 -15082 1709 -15048
rect 1811 -15082 1827 -15048
rect 1871 -15082 1887 -15048
rect 1989 -15082 2005 -15048
rect 2049 -15082 2065 -15048
rect 2167 -15082 2183 -15048
rect 2227 -15082 2243 -15048
rect 2345 -15082 2361 -15048
rect 2405 -15082 2421 -15048
rect 2523 -15082 2539 -15048
rect 2583 -15082 2599 -15048
rect 2701 -15082 2717 -15048
rect 2761 -15082 2777 -15048
rect 2879 -15082 2895 -15048
rect 2939 -15082 2955 -15048
rect 3057 -15082 3073 -15048
rect 3117 -15082 3133 -15048
rect 3235 -15082 3251 -15048
rect 3295 -15082 3311 -15048
rect 3413 -15082 3429 -15048
rect 3473 -15082 3489 -15048
rect 3591 -15082 3607 -15048
rect 3651 -15082 3667 -15048
rect 3769 -15082 3785 -15048
rect 3829 -15082 3845 -15048
rect 3947 -15082 3963 -15048
rect 4007 -15082 4023 -15048
rect 4519 -15071 4745 -15047
rect 5645 -15082 5661 -15048
rect 5705 -15082 5721 -15048
rect 5823 -15082 5839 -15048
rect 5883 -15082 5899 -15048
rect 6001 -15082 6017 -15048
rect 6061 -15082 6077 -15048
rect 6179 -15082 6195 -15048
rect 6239 -15082 6255 -15048
rect 6357 -15082 6373 -15048
rect 6417 -15082 6433 -15048
rect 6535 -15082 6551 -15048
rect 6595 -15082 6611 -15048
rect 6713 -15082 6729 -15048
rect 6773 -15082 6789 -15048
rect 6891 -15082 6907 -15048
rect 6951 -15082 6967 -15048
rect 7069 -15082 7085 -15048
rect 7129 -15082 7145 -15048
rect 7247 -15082 7263 -15048
rect 7307 -15082 7323 -15048
rect 7425 -15082 7441 -15048
rect 7485 -15082 7501 -15048
rect 7603 -15082 7619 -15048
rect 7663 -15082 7679 -15048
rect 7781 -15082 7797 -15048
rect 7841 -15082 7857 -15048
rect 7959 -15082 7975 -15048
rect 8019 -15082 8035 -15048
rect 8137 -15082 8153 -15048
rect 8197 -15082 8213 -15048
rect 8315 -15082 8331 -15048
rect 8375 -15082 8391 -15048
rect 8493 -15082 8509 -15048
rect 8553 -15082 8569 -15048
rect 8671 -15082 8687 -15048
rect 8731 -15082 8747 -15048
rect 8849 -15082 8865 -15048
rect 8909 -15082 8925 -15048
rect 9027 -15082 9043 -15048
rect 9087 -15082 9103 -15048
rect 9205 -15082 9221 -15048
rect 9265 -15082 9281 -15048
rect 9383 -15082 9399 -15048
rect 9443 -15082 9459 -15048
rect 9561 -15082 9577 -15048
rect 9621 -15082 9637 -15048
rect 9739 -15082 9755 -15048
rect 9799 -15082 9815 -15048
rect 9917 -15082 9933 -15048
rect 9977 -15082 9993 -15048
rect 10095 -15082 10111 -15048
rect 10155 -15082 10171 -15048
rect 10273 -15082 10289 -15048
rect 10333 -15082 10349 -15048
rect 10451 -15082 10467 -15048
rect 10511 -15082 10527 -15048
rect 10629 -15082 10645 -15048
rect 10689 -15082 10705 -15048
rect 10807 -15082 10823 -15048
rect 10867 -15082 10883 -15048
rect 10985 -15082 11001 -15048
rect 11045 -15082 11061 -15048
rect 11163 -15082 11179 -15048
rect 11223 -15082 11239 -15048
rect 11341 -15082 11357 -15048
rect 11401 -15082 11417 -15048
rect 11519 -15082 11535 -15048
rect 11579 -15082 11595 -15048
rect 11697 -15082 11713 -15048
rect 11757 -15082 11773 -15048
rect 11875 -15082 11891 -15048
rect 11935 -15082 11951 -15048
rect 12053 -15082 12069 -15048
rect 12113 -15082 12129 -15048
rect 12231 -15082 12247 -15048
rect 12291 -15082 12307 -15048
rect 12409 -15082 12425 -15048
rect 12469 -15082 12485 -15048
rect 12587 -15082 12603 -15048
rect 12647 -15082 12663 -15048
rect -2173 -15132 -2139 -15116
rect -4070 -15366 -4036 -15350
rect -3009 -15276 -2783 -15252
rect -5960 -15434 -5944 -15400
rect -5900 -15434 -5884 -15400
rect -5782 -15434 -5766 -15400
rect -5722 -15434 -5706 -15400
rect -5604 -15434 -5588 -15400
rect -5544 -15434 -5528 -15400
rect -5426 -15434 -5410 -15400
rect -5366 -15434 -5350 -15400
rect -5248 -15434 -5232 -15400
rect -5188 -15434 -5172 -15400
rect -5070 -15434 -5054 -15400
rect -5010 -15434 -4994 -15400
rect -4892 -15434 -4876 -15400
rect -4832 -15434 -4816 -15400
rect -4714 -15434 -4698 -15400
rect -4654 -15434 -4638 -15400
rect -4536 -15434 -4520 -15400
rect -4476 -15434 -4460 -15400
rect -4358 -15434 -4342 -15400
rect -4298 -15434 -4282 -15400
rect -4180 -15434 -4164 -15400
rect -4120 -15434 -4104 -15400
rect -3009 -15454 -2985 -15276
rect -2807 -15454 -2783 -15276
rect -2173 -15404 -2139 -15388
rect -1995 -15132 -1961 -15116
rect -1995 -15404 -1961 -15388
rect -1817 -15132 -1783 -15116
rect -1817 -15404 -1783 -15388
rect -1639 -15132 -1605 -15116
rect -1639 -15404 -1605 -15388
rect -1461 -15132 -1427 -15116
rect -1461 -15404 -1427 -15388
rect -1283 -15132 -1249 -15116
rect -1283 -15404 -1249 -15388
rect -1105 -15132 -1071 -15116
rect -1105 -15404 -1071 -15388
rect -927 -15132 -893 -15116
rect -927 -15404 -893 -15388
rect -749 -15132 -715 -15116
rect -749 -15404 -715 -15388
rect -571 -15132 -537 -15116
rect -571 -15404 -537 -15388
rect -393 -15132 -359 -15116
rect -393 -15404 -359 -15388
rect -215 -15132 -181 -15116
rect -215 -15404 -181 -15388
rect -37 -15132 -3 -15116
rect -37 -15404 -3 -15388
rect 141 -15132 175 -15116
rect 141 -15404 175 -15388
rect 319 -15132 353 -15116
rect 319 -15404 353 -15388
rect 497 -15132 531 -15116
rect 497 -15404 531 -15388
rect 675 -15132 709 -15116
rect 675 -15404 709 -15388
rect 853 -15132 887 -15116
rect 853 -15404 887 -15388
rect 1031 -15132 1065 -15116
rect 1031 -15404 1065 -15388
rect 1209 -15132 1243 -15116
rect 1209 -15404 1243 -15388
rect 1387 -15132 1421 -15116
rect 1387 -15404 1421 -15388
rect 1565 -15132 1599 -15116
rect 1565 -15404 1599 -15388
rect 1743 -15132 1777 -15116
rect 1743 -15404 1777 -15388
rect 1921 -15132 1955 -15116
rect 1921 -15404 1955 -15388
rect 2099 -15132 2133 -15116
rect 2099 -15404 2133 -15388
rect 2277 -15132 2311 -15116
rect 2277 -15404 2311 -15388
rect 2455 -15132 2489 -15116
rect 2455 -15404 2489 -15388
rect 2633 -15132 2667 -15116
rect 2633 -15404 2667 -15388
rect 2811 -15132 2845 -15116
rect 2811 -15404 2845 -15388
rect 2989 -15132 3023 -15116
rect 2989 -15404 3023 -15388
rect 3167 -15132 3201 -15116
rect 3167 -15404 3201 -15388
rect 3345 -15132 3379 -15116
rect 3345 -15404 3379 -15388
rect 3523 -15132 3557 -15116
rect 3523 -15404 3557 -15388
rect 3701 -15132 3735 -15116
rect 3701 -15404 3735 -15388
rect 3879 -15132 3913 -15116
rect 3879 -15404 3913 -15388
rect 4057 -15132 4091 -15116
rect 4057 -15404 4091 -15388
rect 5577 -15132 5611 -15116
rect 5577 -15404 5611 -15388
rect 5755 -15132 5789 -15116
rect 5755 -15404 5789 -15388
rect 5933 -15132 5967 -15116
rect 5933 -15404 5967 -15388
rect 6111 -15132 6145 -15116
rect 6111 -15404 6145 -15388
rect 6289 -15132 6323 -15116
rect 6289 -15404 6323 -15388
rect 6467 -15132 6501 -15116
rect 6467 -15404 6501 -15388
rect 6645 -15132 6679 -15116
rect 6645 -15404 6679 -15388
rect 6823 -15132 6857 -15116
rect 6823 -15404 6857 -15388
rect 7001 -15132 7035 -15116
rect 7001 -15404 7035 -15388
rect 7179 -15132 7213 -15116
rect 7179 -15404 7213 -15388
rect 7357 -15132 7391 -15116
rect 7357 -15404 7391 -15388
rect 7535 -15132 7569 -15116
rect 7535 -15404 7569 -15388
rect 7713 -15132 7747 -15116
rect 7713 -15404 7747 -15388
rect 7891 -15132 7925 -15116
rect 7891 -15404 7925 -15388
rect 8069 -15132 8103 -15116
rect 8069 -15404 8103 -15388
rect 8247 -15132 8281 -15116
rect 8247 -15404 8281 -15388
rect 8425 -15132 8459 -15116
rect 8425 -15404 8459 -15388
rect 8603 -15132 8637 -15116
rect 8603 -15404 8637 -15388
rect 8781 -15132 8815 -15116
rect 8781 -15404 8815 -15388
rect 8959 -15132 8993 -15116
rect 8959 -15404 8993 -15388
rect 9137 -15132 9171 -15116
rect 9137 -15404 9171 -15388
rect 9315 -15132 9349 -15116
rect 9315 -15404 9349 -15388
rect 9493 -15132 9527 -15116
rect 9493 -15404 9527 -15388
rect 9671 -15132 9705 -15116
rect 9671 -15404 9705 -15388
rect 9849 -15132 9883 -15116
rect 9849 -15404 9883 -15388
rect 10027 -15132 10061 -15116
rect 10027 -15404 10061 -15388
rect 10205 -15132 10239 -15116
rect 10205 -15404 10239 -15388
rect 10383 -15132 10417 -15116
rect 10383 -15404 10417 -15388
rect 10561 -15132 10595 -15116
rect 10561 -15404 10595 -15388
rect 10739 -15132 10773 -15116
rect 10739 -15404 10773 -15388
rect 10917 -15132 10951 -15116
rect 10917 -15404 10951 -15388
rect 11095 -15132 11129 -15116
rect 11095 -15404 11129 -15388
rect 11273 -15132 11307 -15116
rect 11273 -15404 11307 -15388
rect 11451 -15132 11485 -15116
rect 11451 -15404 11485 -15388
rect 11629 -15132 11663 -15116
rect 11629 -15404 11663 -15388
rect 11807 -15132 11841 -15116
rect 11807 -15404 11841 -15388
rect 11985 -15132 12019 -15116
rect 11985 -15404 12019 -15388
rect 12163 -15132 12197 -15116
rect 12163 -15404 12197 -15388
rect 12341 -15132 12375 -15116
rect 12341 -15404 12375 -15388
rect 12519 -15132 12553 -15116
rect 12519 -15404 12553 -15388
rect 12697 -15132 12731 -15116
rect 12697 -15404 12731 -15388
rect -3009 -15478 -2783 -15454
rect -2105 -15472 -2089 -15438
rect -2045 -15472 -2029 -15438
rect -1927 -15472 -1911 -15438
rect -1867 -15472 -1851 -15438
rect -1749 -15472 -1733 -15438
rect -1689 -15472 -1673 -15438
rect -1571 -15472 -1555 -15438
rect -1511 -15472 -1495 -15438
rect -1393 -15472 -1377 -15438
rect -1333 -15472 -1317 -15438
rect -1215 -15472 -1199 -15438
rect -1155 -15472 -1139 -15438
rect -1037 -15472 -1021 -15438
rect -977 -15472 -961 -15438
rect -859 -15472 -843 -15438
rect -799 -15472 -783 -15438
rect -681 -15472 -665 -15438
rect -621 -15472 -605 -15438
rect -503 -15472 -487 -15438
rect -443 -15472 -427 -15438
rect -325 -15472 -309 -15438
rect -265 -15472 -249 -15438
rect -147 -15472 -131 -15438
rect -87 -15472 -71 -15438
rect 31 -15472 47 -15438
rect 91 -15472 107 -15438
rect 209 -15472 225 -15438
rect 269 -15472 285 -15438
rect 387 -15472 403 -15438
rect 447 -15472 463 -15438
rect 565 -15472 581 -15438
rect 625 -15472 641 -15438
rect 743 -15472 759 -15438
rect 803 -15472 819 -15438
rect 921 -15472 937 -15438
rect 981 -15472 997 -15438
rect 1099 -15472 1115 -15438
rect 1159 -15472 1175 -15438
rect 1277 -15472 1293 -15438
rect 1337 -15472 1353 -15438
rect 1455 -15472 1471 -15438
rect 1515 -15472 1531 -15438
rect 1633 -15472 1649 -15438
rect 1693 -15472 1709 -15438
rect 1811 -15472 1827 -15438
rect 1871 -15472 1887 -15438
rect 1989 -15472 2005 -15438
rect 2049 -15472 2065 -15438
rect 2167 -15472 2183 -15438
rect 2227 -15472 2243 -15438
rect 2345 -15472 2361 -15438
rect 2405 -15472 2421 -15438
rect 2523 -15472 2539 -15438
rect 2583 -15472 2599 -15438
rect 2701 -15472 2717 -15438
rect 2761 -15472 2777 -15438
rect 2879 -15472 2895 -15438
rect 2939 -15472 2955 -15438
rect 3057 -15472 3073 -15438
rect 3117 -15472 3133 -15438
rect 3235 -15472 3251 -15438
rect 3295 -15472 3311 -15438
rect 3413 -15472 3429 -15438
rect 3473 -15472 3489 -15438
rect 3591 -15472 3607 -15438
rect 3651 -15472 3667 -15438
rect 3769 -15472 3785 -15438
rect 3829 -15472 3845 -15438
rect 3947 -15472 3963 -15438
rect 4007 -15472 4023 -15438
rect 5645 -15472 5661 -15438
rect 5705 -15472 5721 -15438
rect 5823 -15472 5839 -15438
rect 5883 -15472 5899 -15438
rect 6001 -15472 6017 -15438
rect 6061 -15472 6077 -15438
rect 6179 -15472 6195 -15438
rect 6239 -15472 6255 -15438
rect 6357 -15472 6373 -15438
rect 6417 -15472 6433 -15438
rect 6535 -15472 6551 -15438
rect 6595 -15472 6611 -15438
rect 6713 -15472 6729 -15438
rect 6773 -15472 6789 -15438
rect 6891 -15472 6907 -15438
rect 6951 -15472 6967 -15438
rect 7069 -15472 7085 -15438
rect 7129 -15472 7145 -15438
rect 7247 -15472 7263 -15438
rect 7307 -15472 7323 -15438
rect 7425 -15472 7441 -15438
rect 7485 -15472 7501 -15438
rect 7603 -15472 7619 -15438
rect 7663 -15472 7679 -15438
rect 7781 -15472 7797 -15438
rect 7841 -15472 7857 -15438
rect 7959 -15472 7975 -15438
rect 8019 -15472 8035 -15438
rect 8137 -15472 8153 -15438
rect 8197 -15472 8213 -15438
rect 8315 -15472 8331 -15438
rect 8375 -15472 8391 -15438
rect 8493 -15472 8509 -15438
rect 8553 -15472 8569 -15438
rect 8671 -15472 8687 -15438
rect 8731 -15472 8747 -15438
rect 8849 -15472 8865 -15438
rect 8909 -15472 8925 -15438
rect 9027 -15472 9043 -15438
rect 9087 -15472 9103 -15438
rect 9205 -15472 9221 -15438
rect 9265 -15472 9281 -15438
rect 9383 -15472 9399 -15438
rect 9443 -15472 9459 -15438
rect 9561 -15472 9577 -15438
rect 9621 -15472 9637 -15438
rect 9739 -15472 9755 -15438
rect 9799 -15472 9815 -15438
rect 9917 -15472 9933 -15438
rect 9977 -15472 9993 -15438
rect 10095 -15472 10111 -15438
rect 10155 -15472 10171 -15438
rect 10273 -15472 10289 -15438
rect 10333 -15472 10349 -15438
rect 10451 -15472 10467 -15438
rect 10511 -15472 10527 -15438
rect 10629 -15472 10645 -15438
rect 10689 -15472 10705 -15438
rect 10807 -15472 10823 -15438
rect 10867 -15472 10883 -15438
rect 10985 -15472 11001 -15438
rect 11045 -15472 11061 -15438
rect 11163 -15472 11179 -15438
rect 11223 -15472 11239 -15438
rect 11341 -15472 11357 -15438
rect 11401 -15472 11417 -15438
rect 11519 -15472 11535 -15438
rect 11579 -15472 11595 -15438
rect 11697 -15472 11713 -15438
rect 11757 -15472 11773 -15438
rect 11875 -15472 11891 -15438
rect 11935 -15472 11951 -15438
rect 12053 -15472 12069 -15438
rect 12113 -15472 12129 -15438
rect 12231 -15472 12247 -15438
rect 12291 -15472 12307 -15438
rect 12409 -15472 12425 -15438
rect 12469 -15472 12485 -15438
rect 12587 -15472 12603 -15438
rect 12647 -15472 12663 -15438
rect -5960 -15744 -5944 -15710
rect -5900 -15744 -5884 -15710
rect -5782 -15744 -5766 -15710
rect -5722 -15744 -5706 -15710
rect -5604 -15744 -5588 -15710
rect -5544 -15744 -5528 -15710
rect -5426 -15744 -5410 -15710
rect -5366 -15744 -5350 -15710
rect -5248 -15744 -5232 -15710
rect -5188 -15744 -5172 -15710
rect -5070 -15744 -5054 -15710
rect -5010 -15744 -4994 -15710
rect -4892 -15744 -4876 -15710
rect -4832 -15744 -4816 -15710
rect -4714 -15744 -4698 -15710
rect -4654 -15744 -4638 -15710
rect -4536 -15744 -4520 -15710
rect -4476 -15744 -4460 -15710
rect -4358 -15744 -4342 -15710
rect -4298 -15744 -4282 -15710
rect -4180 -15744 -4164 -15710
rect -4120 -15744 -4104 -15710
rect -6028 -15794 -5994 -15778
rect -6028 -16066 -5994 -16050
rect -5850 -15794 -5816 -15778
rect -5850 -16066 -5816 -16050
rect -5672 -15794 -5638 -15778
rect -5672 -16066 -5638 -16050
rect -5494 -15794 -5460 -15778
rect -5494 -16066 -5460 -16050
rect -5316 -15794 -5282 -15778
rect -5316 -16066 -5282 -16050
rect -5138 -15794 -5104 -15778
rect -5138 -16066 -5104 -16050
rect -4960 -15794 -4926 -15778
rect -4960 -16066 -4926 -16050
rect -4782 -15794 -4748 -15778
rect -4782 -16066 -4748 -16050
rect -4604 -15794 -4570 -15778
rect -4604 -16066 -4570 -16050
rect -4426 -15794 -4392 -15778
rect -4426 -16066 -4392 -16050
rect -4248 -15794 -4214 -15778
rect -4248 -16066 -4214 -16050
rect -4070 -15794 -4036 -15778
rect -4070 -16066 -4036 -16050
rect -2105 -16082 -2089 -16048
rect -2045 -16082 -2029 -16048
rect -1927 -16082 -1911 -16048
rect -1867 -16082 -1851 -16048
rect -1749 -16082 -1733 -16048
rect -1689 -16082 -1673 -16048
rect -1571 -16082 -1555 -16048
rect -1511 -16082 -1495 -16048
rect -1393 -16082 -1377 -16048
rect -1333 -16082 -1317 -16048
rect -1215 -16082 -1199 -16048
rect -1155 -16082 -1139 -16048
rect -1037 -16082 -1021 -16048
rect -977 -16082 -961 -16048
rect -859 -16082 -843 -16048
rect -799 -16082 -783 -16048
rect -681 -16082 -665 -16048
rect -621 -16082 -605 -16048
rect -503 -16082 -487 -16048
rect -443 -16082 -427 -16048
rect -325 -16082 -309 -16048
rect -265 -16082 -249 -16048
rect -147 -16082 -131 -16048
rect -87 -16082 -71 -16048
rect 31 -16082 47 -16048
rect 91 -16082 107 -16048
rect 209 -16082 225 -16048
rect 269 -16082 285 -16048
rect 387 -16082 403 -16048
rect 447 -16082 463 -16048
rect 565 -16082 581 -16048
rect 625 -16082 641 -16048
rect 743 -16082 759 -16048
rect 803 -16082 819 -16048
rect 921 -16082 937 -16048
rect 981 -16082 997 -16048
rect 1099 -16082 1115 -16048
rect 1159 -16082 1175 -16048
rect 1277 -16082 1293 -16048
rect 1337 -16082 1353 -16048
rect 1455 -16082 1471 -16048
rect 1515 -16082 1531 -16048
rect 1633 -16082 1649 -16048
rect 1693 -16082 1709 -16048
rect 1811 -16082 1827 -16048
rect 1871 -16082 1887 -16048
rect 1989 -16082 2005 -16048
rect 2049 -16082 2065 -16048
rect 2167 -16082 2183 -16048
rect 2227 -16082 2243 -16048
rect 2345 -16082 2361 -16048
rect 2405 -16082 2421 -16048
rect 2523 -16082 2539 -16048
rect 2583 -16082 2599 -16048
rect 2701 -16082 2717 -16048
rect 2761 -16082 2777 -16048
rect 2879 -16082 2895 -16048
rect 2939 -16082 2955 -16048
rect 3057 -16082 3073 -16048
rect 3117 -16082 3133 -16048
rect 3235 -16082 3251 -16048
rect 3295 -16082 3311 -16048
rect 3413 -16082 3429 -16048
rect 3473 -16082 3489 -16048
rect 3591 -16082 3607 -16048
rect 3651 -16082 3667 -16048
rect 3769 -16082 3785 -16048
rect 3829 -16082 3845 -16048
rect 3947 -16082 3963 -16048
rect 4007 -16082 4023 -16048
rect 5645 -16082 5661 -16048
rect 5705 -16082 5721 -16048
rect 5823 -16082 5839 -16048
rect 5883 -16082 5899 -16048
rect 6001 -16082 6017 -16048
rect 6061 -16082 6077 -16048
rect 6179 -16082 6195 -16048
rect 6239 -16082 6255 -16048
rect 6357 -16082 6373 -16048
rect 6417 -16082 6433 -16048
rect 6535 -16082 6551 -16048
rect 6595 -16082 6611 -16048
rect 6713 -16082 6729 -16048
rect 6773 -16082 6789 -16048
rect 6891 -16082 6907 -16048
rect 6951 -16082 6967 -16048
rect 7069 -16082 7085 -16048
rect 7129 -16082 7145 -16048
rect 7247 -16082 7263 -16048
rect 7307 -16082 7323 -16048
rect 7425 -16082 7441 -16048
rect 7485 -16082 7501 -16048
rect 7603 -16082 7619 -16048
rect 7663 -16082 7679 -16048
rect 7781 -16082 7797 -16048
rect 7841 -16082 7857 -16048
rect 7959 -16082 7975 -16048
rect 8019 -16082 8035 -16048
rect 8137 -16082 8153 -16048
rect 8197 -16082 8213 -16048
rect 8315 -16082 8331 -16048
rect 8375 -16082 8391 -16048
rect 8493 -16082 8509 -16048
rect 8553 -16082 8569 -16048
rect 8671 -16082 8687 -16048
rect 8731 -16082 8747 -16048
rect 8849 -16082 8865 -16048
rect 8909 -16082 8925 -16048
rect 9027 -16082 9043 -16048
rect 9087 -16082 9103 -16048
rect 9205 -16082 9221 -16048
rect 9265 -16082 9281 -16048
rect 9383 -16082 9399 -16048
rect 9443 -16082 9459 -16048
rect 9561 -16082 9577 -16048
rect 9621 -16082 9637 -16048
rect 9739 -16082 9755 -16048
rect 9799 -16082 9815 -16048
rect 9917 -16082 9933 -16048
rect 9977 -16082 9993 -16048
rect 10095 -16082 10111 -16048
rect 10155 -16082 10171 -16048
rect 10273 -16082 10289 -16048
rect 10333 -16082 10349 -16048
rect 10451 -16082 10467 -16048
rect 10511 -16082 10527 -16048
rect 10629 -16082 10645 -16048
rect 10689 -16082 10705 -16048
rect 10807 -16082 10823 -16048
rect 10867 -16082 10883 -16048
rect 10985 -16082 11001 -16048
rect 11045 -16082 11061 -16048
rect 11163 -16082 11179 -16048
rect 11223 -16082 11239 -16048
rect 11341 -16082 11357 -16048
rect 11401 -16082 11417 -16048
rect 11519 -16082 11535 -16048
rect 11579 -16082 11595 -16048
rect 11697 -16082 11713 -16048
rect 11757 -16082 11773 -16048
rect 11875 -16082 11891 -16048
rect 11935 -16082 11951 -16048
rect 12053 -16082 12069 -16048
rect 12113 -16082 12129 -16048
rect 12231 -16082 12247 -16048
rect 12291 -16082 12307 -16048
rect 12409 -16082 12425 -16048
rect 12469 -16082 12485 -16048
rect 12587 -16082 12603 -16048
rect 12647 -16082 12663 -16048
rect -5960 -16134 -5944 -16100
rect -5900 -16134 -5884 -16100
rect -5782 -16134 -5766 -16100
rect -5722 -16134 -5706 -16100
rect -5604 -16134 -5588 -16100
rect -5544 -16134 -5528 -16100
rect -5426 -16134 -5410 -16100
rect -5366 -16134 -5350 -16100
rect -5248 -16134 -5232 -16100
rect -5188 -16134 -5172 -16100
rect -5070 -16134 -5054 -16100
rect -5010 -16134 -4994 -16100
rect -4892 -16134 -4876 -16100
rect -4832 -16134 -4816 -16100
rect -4714 -16134 -4698 -16100
rect -4654 -16134 -4638 -16100
rect -4536 -16134 -4520 -16100
rect -4476 -16134 -4460 -16100
rect -4358 -16134 -4342 -16100
rect -4298 -16134 -4282 -16100
rect -4180 -16134 -4164 -16100
rect -4120 -16134 -4104 -16100
rect -2173 -16132 -2139 -16116
rect -2173 -16404 -2139 -16388
rect -1995 -16132 -1961 -16116
rect -1995 -16404 -1961 -16388
rect -1817 -16132 -1783 -16116
rect -1817 -16404 -1783 -16388
rect -1639 -16132 -1605 -16116
rect -1639 -16404 -1605 -16388
rect -1461 -16132 -1427 -16116
rect -1461 -16404 -1427 -16388
rect -1283 -16132 -1249 -16116
rect -1283 -16404 -1249 -16388
rect -1105 -16132 -1071 -16116
rect -1105 -16404 -1071 -16388
rect -927 -16132 -893 -16116
rect -927 -16404 -893 -16388
rect -749 -16132 -715 -16116
rect -749 -16404 -715 -16388
rect -571 -16132 -537 -16116
rect -571 -16404 -537 -16388
rect -393 -16132 -359 -16116
rect -393 -16404 -359 -16388
rect -215 -16132 -181 -16116
rect -215 -16404 -181 -16388
rect -37 -16132 -3 -16116
rect -37 -16404 -3 -16388
rect 141 -16132 175 -16116
rect 141 -16404 175 -16388
rect 319 -16132 353 -16116
rect 319 -16404 353 -16388
rect 497 -16132 531 -16116
rect 497 -16404 531 -16388
rect 675 -16132 709 -16116
rect 675 -16404 709 -16388
rect 853 -16132 887 -16116
rect 853 -16404 887 -16388
rect 1031 -16132 1065 -16116
rect 1031 -16404 1065 -16388
rect 1209 -16132 1243 -16116
rect 1209 -16404 1243 -16388
rect 1387 -16132 1421 -16116
rect 1387 -16404 1421 -16388
rect 1565 -16132 1599 -16116
rect 1565 -16404 1599 -16388
rect 1743 -16132 1777 -16116
rect 1743 -16404 1777 -16388
rect 1921 -16132 1955 -16116
rect 1921 -16404 1955 -16388
rect 2099 -16132 2133 -16116
rect 2099 -16404 2133 -16388
rect 2277 -16132 2311 -16116
rect 2277 -16404 2311 -16388
rect 2455 -16132 2489 -16116
rect 2455 -16404 2489 -16388
rect 2633 -16132 2667 -16116
rect 2633 -16404 2667 -16388
rect 2811 -16132 2845 -16116
rect 2811 -16404 2845 -16388
rect 2989 -16132 3023 -16116
rect 2989 -16404 3023 -16388
rect 3167 -16132 3201 -16116
rect 3167 -16404 3201 -16388
rect 3345 -16132 3379 -16116
rect 3345 -16404 3379 -16388
rect 3523 -16132 3557 -16116
rect 3523 -16404 3557 -16388
rect 3701 -16132 3735 -16116
rect 3701 -16404 3735 -16388
rect 3879 -16132 3913 -16116
rect 3879 -16404 3913 -16388
rect 4057 -16132 4091 -16116
rect 4057 -16404 4091 -16388
rect 5577 -16132 5611 -16116
rect 5577 -16404 5611 -16388
rect 5755 -16132 5789 -16116
rect 5755 -16404 5789 -16388
rect 5933 -16132 5967 -16116
rect 5933 -16404 5967 -16388
rect 6111 -16132 6145 -16116
rect 6111 -16404 6145 -16388
rect 6289 -16132 6323 -16116
rect 6289 -16404 6323 -16388
rect 6467 -16132 6501 -16116
rect 6467 -16404 6501 -16388
rect 6645 -16132 6679 -16116
rect 6645 -16404 6679 -16388
rect 6823 -16132 6857 -16116
rect 6823 -16404 6857 -16388
rect 7001 -16132 7035 -16116
rect 7001 -16404 7035 -16388
rect 7179 -16132 7213 -16116
rect 7179 -16404 7213 -16388
rect 7357 -16132 7391 -16116
rect 7357 -16404 7391 -16388
rect 7535 -16132 7569 -16116
rect 7535 -16404 7569 -16388
rect 7713 -16132 7747 -16116
rect 7713 -16404 7747 -16388
rect 7891 -16132 7925 -16116
rect 7891 -16404 7925 -16388
rect 8069 -16132 8103 -16116
rect 8069 -16404 8103 -16388
rect 8247 -16132 8281 -16116
rect 8247 -16404 8281 -16388
rect 8425 -16132 8459 -16116
rect 8425 -16404 8459 -16388
rect 8603 -16132 8637 -16116
rect 8603 -16404 8637 -16388
rect 8781 -16132 8815 -16116
rect 8781 -16404 8815 -16388
rect 8959 -16132 8993 -16116
rect 8959 -16404 8993 -16388
rect 9137 -16132 9171 -16116
rect 9137 -16404 9171 -16388
rect 9315 -16132 9349 -16116
rect 9315 -16404 9349 -16388
rect 9493 -16132 9527 -16116
rect 9493 -16404 9527 -16388
rect 9671 -16132 9705 -16116
rect 9671 -16404 9705 -16388
rect 9849 -16132 9883 -16116
rect 9849 -16404 9883 -16388
rect 10027 -16132 10061 -16116
rect 10027 -16404 10061 -16388
rect 10205 -16132 10239 -16116
rect 10205 -16404 10239 -16388
rect 10383 -16132 10417 -16116
rect 10383 -16404 10417 -16388
rect 10561 -16132 10595 -16116
rect 10561 -16404 10595 -16388
rect 10739 -16132 10773 -16116
rect 10739 -16404 10773 -16388
rect 10917 -16132 10951 -16116
rect 10917 -16404 10951 -16388
rect 11095 -16132 11129 -16116
rect 11095 -16404 11129 -16388
rect 11273 -16132 11307 -16116
rect 11273 -16404 11307 -16388
rect 11451 -16132 11485 -16116
rect 11451 -16404 11485 -16388
rect 11629 -16132 11663 -16116
rect 11629 -16404 11663 -16388
rect 11807 -16132 11841 -16116
rect 11807 -16404 11841 -16388
rect 11985 -16132 12019 -16116
rect 11985 -16404 12019 -16388
rect 12163 -16132 12197 -16116
rect 12163 -16404 12197 -16388
rect 12341 -16132 12375 -16116
rect 12341 -16404 12375 -16388
rect 12519 -16132 12553 -16116
rect 12519 -16404 12553 -16388
rect 12697 -16132 12731 -16116
rect 12697 -16404 12731 -16388
rect -5960 -16444 -5944 -16410
rect -5900 -16444 -5884 -16410
rect -5782 -16444 -5766 -16410
rect -5722 -16444 -5706 -16410
rect -5604 -16444 -5588 -16410
rect -5544 -16444 -5528 -16410
rect -5426 -16444 -5410 -16410
rect -5366 -16444 -5350 -16410
rect -5248 -16444 -5232 -16410
rect -5188 -16444 -5172 -16410
rect -5070 -16444 -5054 -16410
rect -5010 -16444 -4994 -16410
rect -4892 -16444 -4876 -16410
rect -4832 -16444 -4816 -16410
rect -4714 -16444 -4698 -16410
rect -4654 -16444 -4638 -16410
rect -4536 -16444 -4520 -16410
rect -4476 -16444 -4460 -16410
rect -4358 -16444 -4342 -16410
rect -4298 -16444 -4282 -16410
rect -4180 -16444 -4164 -16410
rect -4120 -16444 -4104 -16410
rect -2105 -16472 -2089 -16438
rect -2045 -16472 -2029 -16438
rect -1927 -16472 -1911 -16438
rect -1867 -16472 -1851 -16438
rect -1749 -16472 -1733 -16438
rect -1689 -16472 -1673 -16438
rect -1571 -16472 -1555 -16438
rect -1511 -16472 -1495 -16438
rect -1393 -16472 -1377 -16438
rect -1333 -16472 -1317 -16438
rect -1215 -16472 -1199 -16438
rect -1155 -16472 -1139 -16438
rect -1037 -16472 -1021 -16438
rect -977 -16472 -961 -16438
rect -859 -16472 -843 -16438
rect -799 -16472 -783 -16438
rect -681 -16472 -665 -16438
rect -621 -16472 -605 -16438
rect -503 -16472 -487 -16438
rect -443 -16472 -427 -16438
rect -325 -16472 -309 -16438
rect -265 -16472 -249 -16438
rect -147 -16472 -131 -16438
rect -87 -16472 -71 -16438
rect 31 -16472 47 -16438
rect 91 -16472 107 -16438
rect 209 -16472 225 -16438
rect 269 -16472 285 -16438
rect 387 -16472 403 -16438
rect 447 -16472 463 -16438
rect 565 -16472 581 -16438
rect 625 -16472 641 -16438
rect 743 -16472 759 -16438
rect 803 -16472 819 -16438
rect 921 -16472 937 -16438
rect 981 -16472 997 -16438
rect 1099 -16472 1115 -16438
rect 1159 -16472 1175 -16438
rect 1277 -16472 1293 -16438
rect 1337 -16472 1353 -16438
rect 1455 -16472 1471 -16438
rect 1515 -16472 1531 -16438
rect 1633 -16472 1649 -16438
rect 1693 -16472 1709 -16438
rect 1811 -16472 1827 -16438
rect 1871 -16472 1887 -16438
rect 1989 -16472 2005 -16438
rect 2049 -16472 2065 -16438
rect 2167 -16472 2183 -16438
rect 2227 -16472 2243 -16438
rect 2345 -16472 2361 -16438
rect 2405 -16472 2421 -16438
rect 2523 -16472 2539 -16438
rect 2583 -16472 2599 -16438
rect 2701 -16472 2717 -16438
rect 2761 -16472 2777 -16438
rect 2879 -16472 2895 -16438
rect 2939 -16472 2955 -16438
rect 3057 -16472 3073 -16438
rect 3117 -16472 3133 -16438
rect 3235 -16472 3251 -16438
rect 3295 -16472 3311 -16438
rect 3413 -16472 3429 -16438
rect 3473 -16472 3489 -16438
rect 3591 -16472 3607 -16438
rect 3651 -16472 3667 -16438
rect 3769 -16472 3785 -16438
rect 3829 -16472 3845 -16438
rect 3947 -16472 3963 -16438
rect 4007 -16472 4023 -16438
rect 5645 -16472 5661 -16438
rect 5705 -16472 5721 -16438
rect 5823 -16472 5839 -16438
rect 5883 -16472 5899 -16438
rect 6001 -16472 6017 -16438
rect 6061 -16472 6077 -16438
rect 6179 -16472 6195 -16438
rect 6239 -16472 6255 -16438
rect 6357 -16472 6373 -16438
rect 6417 -16472 6433 -16438
rect 6535 -16472 6551 -16438
rect 6595 -16472 6611 -16438
rect 6713 -16472 6729 -16438
rect 6773 -16472 6789 -16438
rect 6891 -16472 6907 -16438
rect 6951 -16472 6967 -16438
rect 7069 -16472 7085 -16438
rect 7129 -16472 7145 -16438
rect 7247 -16472 7263 -16438
rect 7307 -16472 7323 -16438
rect 7425 -16472 7441 -16438
rect 7485 -16472 7501 -16438
rect 7603 -16472 7619 -16438
rect 7663 -16472 7679 -16438
rect 7781 -16472 7797 -16438
rect 7841 -16472 7857 -16438
rect 7959 -16472 7975 -16438
rect 8019 -16472 8035 -16438
rect 8137 -16472 8153 -16438
rect 8197 -16472 8213 -16438
rect 8315 -16472 8331 -16438
rect 8375 -16472 8391 -16438
rect 8493 -16472 8509 -16438
rect 8553 -16472 8569 -16438
rect 8671 -16472 8687 -16438
rect 8731 -16472 8747 -16438
rect 8849 -16472 8865 -16438
rect 8909 -16472 8925 -16438
rect 9027 -16472 9043 -16438
rect 9087 -16472 9103 -16438
rect 9205 -16472 9221 -16438
rect 9265 -16472 9281 -16438
rect 9383 -16472 9399 -16438
rect 9443 -16472 9459 -16438
rect 9561 -16472 9577 -16438
rect 9621 -16472 9637 -16438
rect 9739 -16472 9755 -16438
rect 9799 -16472 9815 -16438
rect 9917 -16472 9933 -16438
rect 9977 -16472 9993 -16438
rect 10095 -16472 10111 -16438
rect 10155 -16472 10171 -16438
rect 10273 -16472 10289 -16438
rect 10333 -16472 10349 -16438
rect 10451 -16472 10467 -16438
rect 10511 -16472 10527 -16438
rect 10629 -16472 10645 -16438
rect 10689 -16472 10705 -16438
rect 10807 -16472 10823 -16438
rect 10867 -16472 10883 -16438
rect 10985 -16472 11001 -16438
rect 11045 -16472 11061 -16438
rect 11163 -16472 11179 -16438
rect 11223 -16472 11239 -16438
rect 11341 -16472 11357 -16438
rect 11401 -16472 11417 -16438
rect 11519 -16472 11535 -16438
rect 11579 -16472 11595 -16438
rect 11697 -16472 11713 -16438
rect 11757 -16472 11773 -16438
rect 11875 -16472 11891 -16438
rect 11935 -16472 11951 -16438
rect 12053 -16472 12069 -16438
rect 12113 -16472 12129 -16438
rect 12231 -16472 12247 -16438
rect 12291 -16472 12307 -16438
rect 12409 -16472 12425 -16438
rect 12469 -16472 12485 -16438
rect 12587 -16472 12603 -16438
rect 12647 -16472 12663 -16438
rect -6028 -16494 -5994 -16478
rect -6028 -16766 -5994 -16750
rect -5850 -16494 -5816 -16478
rect -5850 -16766 -5816 -16750
rect -5672 -16494 -5638 -16478
rect -5672 -16766 -5638 -16750
rect -5494 -16494 -5460 -16478
rect -5494 -16766 -5460 -16750
rect -5316 -16494 -5282 -16478
rect -5316 -16766 -5282 -16750
rect -5138 -16494 -5104 -16478
rect -5138 -16766 -5104 -16750
rect -4960 -16494 -4926 -16478
rect -4960 -16766 -4926 -16750
rect -4782 -16494 -4748 -16478
rect -4782 -16766 -4748 -16750
rect -4604 -16494 -4570 -16478
rect -4604 -16766 -4570 -16750
rect -4426 -16494 -4392 -16478
rect -4426 -16766 -4392 -16750
rect -4248 -16494 -4214 -16478
rect -4248 -16766 -4214 -16750
rect -4070 -16494 -4036 -16478
rect -4070 -16766 -4036 -16750
rect -5960 -16834 -5944 -16800
rect -5900 -16834 -5884 -16800
rect -5782 -16834 -5766 -16800
rect -5722 -16834 -5706 -16800
rect -5604 -16834 -5588 -16800
rect -5544 -16834 -5528 -16800
rect -5426 -16834 -5410 -16800
rect -5366 -16834 -5350 -16800
rect -5248 -16834 -5232 -16800
rect -5188 -16834 -5172 -16800
rect -5070 -16834 -5054 -16800
rect -5010 -16834 -4994 -16800
rect -4892 -16834 -4876 -16800
rect -4832 -16834 -4816 -16800
rect -4714 -16834 -4698 -16800
rect -4654 -16834 -4638 -16800
rect -4536 -16834 -4520 -16800
rect -4476 -16834 -4460 -16800
rect -4358 -16834 -4342 -16800
rect -4298 -16834 -4282 -16800
rect -4180 -16834 -4164 -16800
rect -4120 -16834 -4104 -16800
rect -7605 -17459 -7505 -17268
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< viali >>
rect 7040 2327 7074 2713
rect 7154 2673 7188 2707
rect 7346 2673 7380 2707
rect 7538 2673 7572 2707
rect 7730 2673 7764 2707
rect 7922 2673 7956 2707
rect 8114 2673 8148 2707
rect 7154 2365 7188 2613
rect 7250 2365 7284 2613
rect 7346 2365 7380 2613
rect 7442 2365 7476 2613
rect 7538 2365 7572 2613
rect 7634 2365 7668 2613
rect 7730 2365 7764 2613
rect 7826 2365 7860 2613
rect 7922 2365 7956 2613
rect 8018 2365 8052 2613
rect 8114 2365 8148 2613
rect 16040 2327 16074 2713
rect 16154 2673 16188 2707
rect 16346 2673 16380 2707
rect 16538 2673 16572 2707
rect 16730 2673 16764 2707
rect 16922 2673 16956 2707
rect 17114 2673 17148 2707
rect 16154 2365 16188 2613
rect 16250 2365 16284 2613
rect 16346 2365 16380 2613
rect 16442 2365 16476 2613
rect 16538 2365 16572 2613
rect 16634 2365 16668 2613
rect 16730 2365 16764 2613
rect 16826 2365 16860 2613
rect 16922 2365 16956 2613
rect 17018 2365 17052 2613
rect 17114 2365 17148 2613
rect 7040 2061 7074 2063
rect 7040 1863 7074 2061
rect 7154 1953 7188 2033
rect 7250 1953 7284 2033
rect 7346 1953 7380 2033
rect 7442 1953 7476 2033
rect 7538 1953 7572 2033
rect 7634 1953 7668 2033
rect 7730 1953 7764 2033
rect 7826 1953 7860 2033
rect 7922 1953 7956 2033
rect 8018 1953 8052 2033
rect 8114 1953 8148 2033
rect 7154 1865 7188 1899
rect 7346 1865 7380 1899
rect 7538 1865 7572 1899
rect 7730 1865 7764 1899
rect 7922 1865 7956 1899
rect 8114 1865 8148 1899
rect 16040 2061 16074 2063
rect 16040 1863 16074 2061
rect 16154 1953 16188 2033
rect 16250 1953 16284 2033
rect 16346 1953 16380 2033
rect 16442 1953 16476 2033
rect 16538 1953 16572 2033
rect 16634 1953 16668 2033
rect 16730 1953 16764 2033
rect 16826 1953 16860 2033
rect 16922 1953 16956 2033
rect 17018 1953 17052 2033
rect 17114 1953 17148 2033
rect 16154 1865 16188 1899
rect 16346 1865 16380 1899
rect 16538 1865 16572 1899
rect 16730 1865 16764 1899
rect 16922 1865 16956 1899
rect 17114 1865 17148 1899
rect 7040 527 7074 913
rect 7154 873 7188 907
rect 7346 873 7380 907
rect 7538 873 7572 907
rect 7730 873 7764 907
rect 7922 873 7956 907
rect 8114 873 8148 907
rect 7154 565 7188 813
rect 7250 565 7284 813
rect 7346 565 7380 813
rect 7442 565 7476 813
rect 7538 565 7572 813
rect 7634 565 7668 813
rect 7730 565 7764 813
rect 7826 565 7860 813
rect 7922 565 7956 813
rect 8018 565 8052 813
rect 8114 565 8148 813
rect 16040 527 16074 913
rect 16154 873 16188 907
rect 16346 873 16380 907
rect 16538 873 16572 907
rect 16730 873 16764 907
rect 16922 873 16956 907
rect 17114 873 17148 907
rect 16154 565 16188 813
rect 16250 565 16284 813
rect 16346 565 16380 813
rect 16442 565 16476 813
rect 16538 565 16572 813
rect 16634 565 16668 813
rect 16730 565 16764 813
rect 16826 565 16860 813
rect 16922 565 16956 813
rect 17018 565 17052 813
rect 17114 565 17148 813
rect 7040 261 7074 263
rect 7040 63 7074 261
rect 7154 153 7188 233
rect 7250 153 7284 233
rect 7346 153 7380 233
rect 7442 153 7476 233
rect 7538 153 7572 233
rect 7634 153 7668 233
rect 7730 153 7764 233
rect 7826 153 7860 233
rect 7922 153 7956 233
rect 8018 153 8052 233
rect 8114 153 8148 233
rect 7154 65 7188 99
rect 7346 65 7380 99
rect 7538 65 7572 99
rect 7730 65 7764 99
rect 7922 65 7956 99
rect 8114 65 8148 99
rect 16040 261 16074 263
rect 16040 63 16074 261
rect 16154 153 16188 233
rect 16250 153 16284 233
rect 16346 153 16380 233
rect 16442 153 16476 233
rect 16538 153 16572 233
rect 16634 153 16668 233
rect 16730 153 16764 233
rect 16826 153 16860 233
rect 16922 153 16956 233
rect 17018 153 17052 233
rect 17114 153 17148 233
rect 16154 65 16188 99
rect 16346 65 16380 99
rect 16538 65 16572 99
rect 16730 65 16764 99
rect 16922 65 16956 99
rect 17114 65 17148 99
rect -7379 -1353 3329 -1260
rect 7040 -1273 7074 -887
rect 7154 -927 7188 -893
rect 7346 -927 7380 -893
rect 7538 -927 7572 -893
rect 7730 -927 7764 -893
rect 7922 -927 7956 -893
rect 8114 -927 8148 -893
rect 7154 -1235 7188 -987
rect 7250 -1235 7284 -987
rect 7346 -1235 7380 -987
rect 7442 -1235 7476 -987
rect 7538 -1235 7572 -987
rect 7634 -1235 7668 -987
rect 7730 -1235 7764 -987
rect 7826 -1235 7860 -987
rect 7922 -1235 7956 -987
rect 8018 -1235 8052 -987
rect 8114 -1235 8148 -987
rect 16040 -1273 16074 -887
rect 16154 -927 16188 -893
rect 16346 -927 16380 -893
rect 16538 -927 16572 -893
rect 16730 -927 16764 -893
rect 16922 -927 16956 -893
rect 17114 -927 17148 -893
rect 16154 -1235 16188 -987
rect 16250 -1235 16284 -987
rect 16346 -1235 16380 -987
rect 16442 -1235 16476 -987
rect 16538 -1235 16572 -987
rect 16634 -1235 16668 -987
rect 16730 -1235 16764 -987
rect 16826 -1235 16860 -987
rect 16922 -1235 16956 -987
rect 17018 -1235 17052 -987
rect 17114 -1235 17148 -987
rect -6218 -2073 -6174 -2039
rect -6040 -2073 -5996 -2039
rect -5862 -2073 -5818 -2039
rect -5684 -2073 -5640 -2039
rect -5506 -2073 -5462 -2039
rect -5328 -2073 -5284 -2039
rect -5150 -2073 -5106 -2039
rect -4972 -2073 -4928 -2039
rect -4794 -2073 -4750 -2039
rect -4616 -2073 -4572 -2039
rect -4438 -2073 -4394 -2039
rect -4260 -2073 -4216 -2039
rect -4082 -2073 -4038 -2039
rect -3904 -2073 -3860 -2039
rect -3726 -2073 -3682 -2039
rect -3548 -2073 -3504 -2039
rect -6302 -2388 -6268 -2132
rect -6124 -2388 -6090 -2132
rect -5946 -2388 -5912 -2132
rect -5768 -2388 -5734 -2132
rect -5590 -2388 -5556 -2132
rect -5412 -2388 -5378 -2132
rect -5234 -2388 -5200 -2132
rect -5056 -2388 -5022 -2132
rect -4878 -2388 -4844 -2132
rect -4700 -2388 -4666 -2132
rect -4522 -2388 -4488 -2132
rect -4344 -2388 -4310 -2132
rect -4166 -2388 -4132 -2132
rect -3988 -2388 -3954 -2132
rect -3810 -2388 -3776 -2132
rect -3632 -2388 -3598 -2132
rect -3454 -2388 -3420 -2132
rect -6218 -2481 -6174 -2447
rect -6040 -2481 -5996 -2447
rect -5862 -2481 -5818 -2447
rect -5684 -2481 -5640 -2447
rect -5506 -2481 -5462 -2447
rect -5328 -2481 -5284 -2447
rect -5150 -2481 -5106 -2447
rect -4972 -2481 -4928 -2447
rect -4794 -2481 -4750 -2447
rect -4616 -2481 -4572 -2447
rect -4438 -2481 -4394 -2447
rect -4260 -2481 -4216 -2447
rect -4082 -2481 -4038 -2447
rect -3904 -2481 -3860 -2447
rect -3726 -2481 -3682 -2447
rect -3548 -2481 -3504 -2447
rect -1370 -2825 -1326 -2791
rect -1192 -2825 -1148 -2791
rect -1014 -2825 -970 -2791
rect -836 -2825 -792 -2791
rect -658 -2825 -614 -2791
rect -480 -2825 -436 -2791
rect -302 -2825 -258 -2791
rect -124 -2825 -80 -2791
rect 54 -2825 98 -2791
rect 232 -2825 276 -2791
rect 410 -2825 454 -2791
rect 588 -2825 632 -2791
rect 766 -2825 810 -2791
rect 944 -2825 988 -2791
rect 1122 -2825 1166 -2791
rect 1300 -2825 1344 -2791
rect 1478 -2825 1522 -2791
rect 1656 -2825 1700 -2791
rect 1834 -2825 1878 -2791
rect 2012 -2825 2056 -2791
rect 2190 -2825 2234 -2791
rect 2368 -2825 2412 -2791
rect 2546 -2825 2590 -2791
rect -6218 -2943 -6174 -2909
rect -6040 -2943 -5996 -2909
rect -5862 -2943 -5818 -2909
rect -5684 -2943 -5640 -2909
rect -5506 -2943 -5462 -2909
rect -5328 -2943 -5284 -2909
rect -5150 -2943 -5106 -2909
rect -4972 -2943 -4928 -2909
rect -4794 -2943 -4750 -2909
rect -4616 -2943 -4572 -2909
rect -4438 -2943 -4394 -2909
rect -4260 -2943 -4216 -2909
rect -4082 -2943 -4038 -2909
rect -3904 -2943 -3860 -2909
rect -3726 -2943 -3682 -2909
rect -3548 -2943 -3504 -2909
rect -6302 -3258 -6268 -3002
rect -6124 -3258 -6090 -3002
rect -5946 -3258 -5912 -3002
rect -5768 -3258 -5734 -3002
rect -5590 -3258 -5556 -3002
rect -5412 -3258 -5378 -3002
rect -5234 -3258 -5200 -3002
rect -5056 -3258 -5022 -3002
rect -4878 -3258 -4844 -3002
rect -4700 -3258 -4666 -3002
rect -4522 -3258 -4488 -3002
rect -4344 -3258 -4310 -3002
rect -4166 -3258 -4132 -3002
rect -3988 -3258 -3954 -3002
rect -3810 -3258 -3776 -3002
rect -3632 -3258 -3598 -3002
rect -3454 -3258 -3420 -3002
rect -2186 -3221 -2008 -3043
rect -1454 -3140 -1420 -2884
rect -1276 -3140 -1242 -2884
rect -1098 -3140 -1064 -2884
rect -920 -3140 -886 -2884
rect -742 -3140 -708 -2884
rect -564 -3140 -530 -2884
rect -386 -3140 -352 -2884
rect -208 -3140 -174 -2884
rect -30 -3140 4 -2884
rect 148 -3140 182 -2884
rect 326 -3140 360 -2884
rect 504 -3140 538 -2884
rect 682 -3140 716 -2884
rect 860 -3140 894 -2884
rect 1038 -3140 1072 -2884
rect 1216 -3140 1250 -2884
rect 1394 -3140 1428 -2884
rect 1572 -3140 1606 -2884
rect 1750 -3140 1784 -2884
rect 1928 -3140 1962 -2884
rect 2106 -3140 2140 -2884
rect 2284 -3140 2318 -2884
rect 2462 -3140 2496 -2884
rect 2640 -3140 2674 -2884
rect -1370 -3233 -1326 -3199
rect -1192 -3233 -1148 -3199
rect -1014 -3233 -970 -3199
rect -836 -3233 -792 -3199
rect -658 -3233 -614 -3199
rect -480 -3233 -436 -3199
rect -302 -3233 -258 -3199
rect -124 -3233 -80 -3199
rect 54 -3233 98 -3199
rect 232 -3233 276 -3199
rect 410 -3233 454 -3199
rect 588 -3233 632 -3199
rect 766 -3233 810 -3199
rect 944 -3233 988 -3199
rect 1122 -3233 1166 -3199
rect 1300 -3233 1344 -3199
rect 1478 -3233 1522 -3199
rect 1656 -3233 1700 -3199
rect 1834 -3233 1878 -3199
rect 2012 -3233 2056 -3199
rect 2190 -3233 2234 -3199
rect 2368 -3233 2412 -3199
rect 2546 -3233 2590 -3199
rect -6218 -3351 -6174 -3317
rect -6040 -3351 -5996 -3317
rect -5862 -3351 -5818 -3317
rect -5684 -3351 -5640 -3317
rect -5506 -3351 -5462 -3317
rect -5328 -3351 -5284 -3317
rect -5150 -3351 -5106 -3317
rect -4972 -3351 -4928 -3317
rect -4794 -3351 -4750 -3317
rect -4616 -3351 -4572 -3317
rect -4438 -3351 -4394 -3317
rect -4260 -3351 -4216 -3317
rect -4082 -3351 -4038 -3317
rect -3904 -3351 -3860 -3317
rect -3726 -3351 -3682 -3317
rect -3548 -3351 -3504 -3317
rect -1370 -3725 -1326 -3691
rect -1192 -3725 -1148 -3691
rect -1014 -3725 -970 -3691
rect -836 -3725 -792 -3691
rect -658 -3725 -614 -3691
rect -480 -3725 -436 -3691
rect -302 -3725 -258 -3691
rect -124 -3725 -80 -3691
rect 54 -3725 98 -3691
rect 232 -3725 276 -3691
rect 410 -3725 454 -3691
rect 588 -3725 632 -3691
rect 766 -3725 810 -3691
rect 944 -3725 988 -3691
rect 1122 -3725 1166 -3691
rect 1300 -3725 1344 -3691
rect 1478 -3725 1522 -3691
rect 1656 -3725 1700 -3691
rect 1834 -3725 1878 -3691
rect 2012 -3725 2056 -3691
rect 2190 -3725 2234 -3691
rect 2368 -3725 2412 -3691
rect 2546 -3725 2590 -3691
rect -6218 -3813 -6174 -3779
rect -6040 -3813 -5996 -3779
rect -5862 -3813 -5818 -3779
rect -5684 -3813 -5640 -3779
rect -5506 -3813 -5462 -3779
rect -5328 -3813 -5284 -3779
rect -5150 -3813 -5106 -3779
rect -4972 -3813 -4928 -3779
rect -4794 -3813 -4750 -3779
rect -4616 -3813 -4572 -3779
rect -4438 -3813 -4394 -3779
rect -4260 -3813 -4216 -3779
rect -4082 -3813 -4038 -3779
rect -3904 -3813 -3860 -3779
rect -3726 -3813 -3682 -3779
rect -3548 -3813 -3504 -3779
rect -6302 -4128 -6268 -3872
rect -6124 -4128 -6090 -3872
rect -5946 -4128 -5912 -3872
rect -5768 -4128 -5734 -3872
rect -5590 -4128 -5556 -3872
rect -5412 -4128 -5378 -3872
rect -5234 -4128 -5200 -3872
rect -5056 -4128 -5022 -3872
rect -4878 -4128 -4844 -3872
rect -4700 -4128 -4666 -3872
rect -4522 -4128 -4488 -3872
rect -4344 -4128 -4310 -3872
rect -4166 -4128 -4132 -3872
rect -3988 -4128 -3954 -3872
rect -3810 -4128 -3776 -3872
rect -3632 -4128 -3598 -3872
rect -3454 -4128 -3420 -3872
rect -1454 -4040 -1420 -3784
rect -1276 -4040 -1242 -3784
rect -1098 -4040 -1064 -3784
rect -920 -4040 -886 -3784
rect -742 -4040 -708 -3784
rect -564 -4040 -530 -3784
rect -386 -4040 -352 -3784
rect -208 -4040 -174 -3784
rect -30 -4040 4 -3784
rect 148 -4040 182 -3784
rect 326 -4040 360 -3784
rect 504 -4040 538 -3784
rect 682 -4040 716 -3784
rect 860 -4040 894 -3784
rect 1038 -4040 1072 -3784
rect 1216 -4040 1250 -3784
rect 1394 -4040 1428 -3784
rect 1572 -4040 1606 -3784
rect 1750 -4040 1784 -3784
rect 1928 -4040 1962 -3784
rect 2106 -4040 2140 -3784
rect 2284 -4040 2318 -3784
rect 2462 -4040 2496 -3784
rect 2640 -4040 2674 -3784
rect -1370 -4133 -1326 -4099
rect -1192 -4133 -1148 -4099
rect -1014 -4133 -970 -4099
rect -836 -4133 -792 -4099
rect -658 -4133 -614 -4099
rect -480 -4133 -436 -4099
rect -302 -4133 -258 -4099
rect -124 -4133 -80 -4099
rect 54 -4133 98 -4099
rect 232 -4133 276 -4099
rect 410 -4133 454 -4099
rect 588 -4133 632 -4099
rect 766 -4133 810 -4099
rect 944 -4133 988 -4099
rect 1122 -4133 1166 -4099
rect 1300 -4133 1344 -4099
rect 1478 -4133 1522 -4099
rect 1656 -4133 1700 -4099
rect 1834 -4133 1878 -4099
rect 2012 -4133 2056 -4099
rect 2190 -4133 2234 -4099
rect 2368 -4133 2412 -4099
rect 2546 -4133 2590 -4099
rect -6218 -4221 -6174 -4187
rect -6040 -4221 -5996 -4187
rect -5862 -4221 -5818 -4187
rect -5684 -4221 -5640 -4187
rect -5506 -4221 -5462 -4187
rect -5328 -4221 -5284 -4187
rect -5150 -4221 -5106 -4187
rect -4972 -4221 -4928 -4187
rect -4794 -4221 -4750 -4187
rect -4616 -4221 -4572 -4187
rect -4438 -4221 -4394 -4187
rect -4260 -4221 -4216 -4187
rect -4082 -4221 -4038 -4187
rect -3904 -4221 -3860 -4187
rect -3726 -4221 -3682 -4187
rect -3548 -4221 -3504 -4187
rect -1370 -4625 -1326 -4591
rect -1192 -4625 -1148 -4591
rect -1014 -4625 -970 -4591
rect -836 -4625 -792 -4591
rect -658 -4625 -614 -4591
rect -480 -4625 -436 -4591
rect -302 -4625 -258 -4591
rect -124 -4625 -80 -4591
rect 54 -4625 98 -4591
rect 232 -4625 276 -4591
rect 410 -4625 454 -4591
rect 588 -4625 632 -4591
rect 766 -4625 810 -4591
rect 944 -4625 988 -4591
rect 1122 -4625 1166 -4591
rect 1300 -4625 1344 -4591
rect 1478 -4625 1522 -4591
rect 1656 -4625 1700 -4591
rect 1834 -4625 1878 -4591
rect 2012 -4625 2056 -4591
rect 2190 -4625 2234 -4591
rect 2368 -4625 2412 -4591
rect 2546 -4625 2590 -4591
rect -6218 -4683 -6174 -4649
rect -6040 -4683 -5996 -4649
rect -5862 -4683 -5818 -4649
rect -5684 -4683 -5640 -4649
rect -5506 -4683 -5462 -4649
rect -5328 -4683 -5284 -4649
rect -5150 -4683 -5106 -4649
rect -4972 -4683 -4928 -4649
rect -4794 -4683 -4750 -4649
rect -4616 -4683 -4572 -4649
rect -4438 -4683 -4394 -4649
rect -4260 -4683 -4216 -4649
rect -4082 -4683 -4038 -4649
rect -3904 -4683 -3860 -4649
rect -3726 -4683 -3682 -4649
rect -3548 -4683 -3504 -4649
rect -6302 -4998 -6268 -4742
rect -6124 -4998 -6090 -4742
rect -5946 -4998 -5912 -4742
rect -5768 -4998 -5734 -4742
rect -5590 -4998 -5556 -4742
rect -5412 -4998 -5378 -4742
rect -5234 -4998 -5200 -4742
rect -5056 -4998 -5022 -4742
rect -4878 -4998 -4844 -4742
rect -4700 -4998 -4666 -4742
rect -4522 -4998 -4488 -4742
rect -4344 -4998 -4310 -4742
rect -4166 -4998 -4132 -4742
rect -3988 -4998 -3954 -4742
rect -3810 -4998 -3776 -4742
rect -3632 -4998 -3598 -4742
rect -3454 -4998 -3420 -4742
rect -1454 -4940 -1420 -4684
rect -1276 -4940 -1242 -4684
rect -1098 -4940 -1064 -4684
rect -920 -4940 -886 -4684
rect -742 -4940 -708 -4684
rect -564 -4940 -530 -4684
rect -386 -4940 -352 -4684
rect -208 -4940 -174 -4684
rect -30 -4940 4 -4684
rect 148 -4940 182 -4684
rect 326 -4940 360 -4684
rect 504 -4940 538 -4684
rect 682 -4940 716 -4684
rect 860 -4940 894 -4684
rect 1038 -4940 1072 -4684
rect 1216 -4940 1250 -4684
rect 1394 -4940 1428 -4684
rect 1572 -4940 1606 -4684
rect 1750 -4940 1784 -4684
rect 1928 -4940 1962 -4684
rect 2106 -4940 2140 -4684
rect 2284 -4940 2318 -4684
rect 2462 -4940 2496 -4684
rect 2640 -4940 2674 -4684
rect -1370 -5033 -1326 -4999
rect -1192 -5033 -1148 -4999
rect -1014 -5033 -970 -4999
rect -836 -5033 -792 -4999
rect -658 -5033 -614 -4999
rect -480 -5033 -436 -4999
rect -302 -5033 -258 -4999
rect -124 -5033 -80 -4999
rect 54 -5033 98 -4999
rect 232 -5033 276 -4999
rect 410 -5033 454 -4999
rect 588 -5033 632 -4999
rect 766 -5033 810 -4999
rect 944 -5033 988 -4999
rect 1122 -5033 1166 -4999
rect 1300 -5033 1344 -4999
rect 1478 -5033 1522 -4999
rect 1656 -5033 1700 -4999
rect 1834 -5033 1878 -4999
rect 2012 -5033 2056 -4999
rect 2190 -5033 2234 -4999
rect 2368 -5033 2412 -4999
rect 2546 -5033 2590 -4999
rect -6218 -5091 -6174 -5057
rect -6040 -5091 -5996 -5057
rect -5862 -5091 -5818 -5057
rect -5684 -5091 -5640 -5057
rect -5506 -5091 -5462 -5057
rect -5328 -5091 -5284 -5057
rect -5150 -5091 -5106 -5057
rect -4972 -5091 -4928 -5057
rect -4794 -5091 -4750 -5057
rect -4616 -5091 -4572 -5057
rect -4438 -5091 -4394 -5057
rect -4260 -5091 -4216 -5057
rect -4082 -5091 -4038 -5057
rect -3904 -5091 -3860 -5057
rect -3726 -5091 -3682 -5057
rect -3548 -5091 -3504 -5057
rect -6218 -5553 -6174 -5519
rect -6040 -5553 -5996 -5519
rect -5862 -5553 -5818 -5519
rect -5684 -5553 -5640 -5519
rect -5506 -5553 -5462 -5519
rect -5328 -5553 -5284 -5519
rect -5150 -5553 -5106 -5519
rect -4972 -5553 -4928 -5519
rect -4794 -5553 -4750 -5519
rect -4616 -5553 -4572 -5519
rect -4438 -5553 -4394 -5519
rect -4260 -5553 -4216 -5519
rect -4082 -5553 -4038 -5519
rect -3904 -5553 -3860 -5519
rect -3726 -5553 -3682 -5519
rect -3548 -5553 -3504 -5519
rect -1370 -5525 -1326 -5491
rect -1192 -5525 -1148 -5491
rect -1014 -5525 -970 -5491
rect -836 -5525 -792 -5491
rect -658 -5525 -614 -5491
rect -480 -5525 -436 -5491
rect -302 -5525 -258 -5491
rect -124 -5525 -80 -5491
rect 54 -5525 98 -5491
rect 232 -5525 276 -5491
rect 410 -5525 454 -5491
rect 588 -5525 632 -5491
rect 766 -5525 810 -5491
rect 944 -5525 988 -5491
rect 1122 -5525 1166 -5491
rect 1300 -5525 1344 -5491
rect 1478 -5525 1522 -5491
rect 1656 -5525 1700 -5491
rect 1834 -5525 1878 -5491
rect 2012 -5525 2056 -5491
rect 2190 -5525 2234 -5491
rect 2368 -5525 2412 -5491
rect 2546 -5525 2590 -5491
rect -6302 -5868 -6268 -5612
rect -6124 -5868 -6090 -5612
rect -5946 -5868 -5912 -5612
rect -5768 -5868 -5734 -5612
rect -5590 -5868 -5556 -5612
rect -5412 -5868 -5378 -5612
rect -5234 -5868 -5200 -5612
rect -5056 -5868 -5022 -5612
rect -4878 -5868 -4844 -5612
rect -4700 -5868 -4666 -5612
rect -4522 -5868 -4488 -5612
rect -4344 -5868 -4310 -5612
rect -4166 -5868 -4132 -5612
rect -3988 -5868 -3954 -5612
rect -3810 -5868 -3776 -5612
rect -3632 -5868 -3598 -5612
rect -3454 -5868 -3420 -5612
rect -3034 -5840 -2856 -5662
rect -1454 -5840 -1420 -5584
rect -1276 -5840 -1242 -5584
rect -1098 -5840 -1064 -5584
rect -920 -5840 -886 -5584
rect -742 -5840 -708 -5584
rect -564 -5840 -530 -5584
rect -386 -5840 -352 -5584
rect -208 -5840 -174 -5584
rect -30 -5840 4 -5584
rect 148 -5840 182 -5584
rect 326 -5840 360 -5584
rect 504 -5840 538 -5584
rect 682 -5840 716 -5584
rect 860 -5840 894 -5584
rect 1038 -5840 1072 -5584
rect 1216 -5840 1250 -5584
rect 1394 -5840 1428 -5584
rect 1572 -5840 1606 -5584
rect 1750 -5840 1784 -5584
rect 1928 -5840 1962 -5584
rect 2106 -5840 2140 -5584
rect 2284 -5840 2318 -5584
rect 2462 -5840 2496 -5584
rect 2640 -5840 2674 -5584
rect -6218 -5961 -6174 -5927
rect -6040 -5961 -5996 -5927
rect -5862 -5961 -5818 -5927
rect -5684 -5961 -5640 -5927
rect -5506 -5961 -5462 -5927
rect -5328 -5961 -5284 -5927
rect -5150 -5961 -5106 -5927
rect -4972 -5961 -4928 -5927
rect -4794 -5961 -4750 -5927
rect -4616 -5961 -4572 -5927
rect -4438 -5961 -4394 -5927
rect -4260 -5961 -4216 -5927
rect -4082 -5961 -4038 -5927
rect -3904 -5961 -3860 -5927
rect -3726 -5961 -3682 -5927
rect -3548 -5961 -3504 -5927
rect -1370 -5933 -1326 -5899
rect -1192 -5933 -1148 -5899
rect -1014 -5933 -970 -5899
rect -836 -5933 -792 -5899
rect -658 -5933 -614 -5899
rect -480 -5933 -436 -5899
rect -302 -5933 -258 -5899
rect -124 -5933 -80 -5899
rect 54 -5933 98 -5899
rect 232 -5933 276 -5899
rect 410 -5933 454 -5899
rect 588 -5933 632 -5899
rect 766 -5933 810 -5899
rect 944 -5933 988 -5899
rect 1122 -5933 1166 -5899
rect 1300 -5933 1344 -5899
rect 1478 -5933 1522 -5899
rect 1656 -5933 1700 -5899
rect 1834 -5933 1878 -5899
rect 2012 -5933 2056 -5899
rect 2190 -5933 2234 -5899
rect 2368 -5933 2412 -5899
rect 2546 -5933 2590 -5899
rect 7040 -1539 7074 -1537
rect 7040 -1737 7074 -1539
rect 7154 -1647 7188 -1567
rect 7250 -1647 7284 -1567
rect 7346 -1647 7380 -1567
rect 7442 -1647 7476 -1567
rect 7538 -1647 7572 -1567
rect 7634 -1647 7668 -1567
rect 7730 -1647 7764 -1567
rect 7826 -1647 7860 -1567
rect 7922 -1647 7956 -1567
rect 8018 -1647 8052 -1567
rect 8114 -1647 8148 -1567
rect 7154 -1735 7188 -1701
rect 7346 -1735 7380 -1701
rect 7538 -1735 7572 -1701
rect 7730 -1735 7764 -1701
rect 7922 -1735 7956 -1701
rect 8114 -1735 8148 -1701
rect 16040 -1539 16074 -1537
rect 16040 -1737 16074 -1539
rect 16154 -1647 16188 -1567
rect 16250 -1647 16284 -1567
rect 16346 -1647 16380 -1567
rect 16442 -1647 16476 -1567
rect 16538 -1647 16572 -1567
rect 16634 -1647 16668 -1567
rect 16730 -1647 16764 -1567
rect 16826 -1647 16860 -1567
rect 16922 -1647 16956 -1567
rect 17018 -1647 17052 -1567
rect 17114 -1647 17148 -1567
rect 16154 -1735 16188 -1701
rect 16346 -1735 16380 -1701
rect 16538 -1735 16572 -1701
rect 16730 -1735 16764 -1701
rect 16922 -1735 16956 -1701
rect 17114 -1735 17148 -1701
rect 7040 -3073 7074 -2687
rect 7154 -2727 7188 -2693
rect 7346 -2727 7380 -2693
rect 7538 -2727 7572 -2693
rect 7730 -2727 7764 -2693
rect 7922 -2727 7956 -2693
rect 8114 -2727 8148 -2693
rect 7154 -3035 7188 -2787
rect 7250 -3035 7284 -2787
rect 7346 -3035 7380 -2787
rect 7442 -3035 7476 -2787
rect 7538 -3035 7572 -2787
rect 7634 -3035 7668 -2787
rect 7730 -3035 7764 -2787
rect 7826 -3035 7860 -2787
rect 7922 -3035 7956 -2787
rect 8018 -3035 8052 -2787
rect 8114 -3035 8148 -2787
rect 16040 -3073 16074 -2687
rect 16154 -2727 16188 -2693
rect 16346 -2727 16380 -2693
rect 16538 -2727 16572 -2693
rect 16730 -2727 16764 -2693
rect 16922 -2727 16956 -2693
rect 17114 -2727 17148 -2693
rect 16154 -3035 16188 -2787
rect 16250 -3035 16284 -2787
rect 16346 -3035 16380 -2787
rect 16442 -3035 16476 -2787
rect 16538 -3035 16572 -2787
rect 16634 -3035 16668 -2787
rect 16730 -3035 16764 -2787
rect 16826 -3035 16860 -2787
rect 16922 -3035 16956 -2787
rect 17018 -3035 17052 -2787
rect 17114 -3035 17148 -2787
rect 7040 -3339 7074 -3337
rect 7040 -3537 7074 -3339
rect 7154 -3447 7188 -3367
rect 7250 -3447 7284 -3367
rect 7346 -3447 7380 -3367
rect 7442 -3447 7476 -3367
rect 7538 -3447 7572 -3367
rect 7634 -3447 7668 -3367
rect 7730 -3447 7764 -3367
rect 7826 -3447 7860 -3367
rect 7922 -3447 7956 -3367
rect 8018 -3447 8052 -3367
rect 8114 -3447 8148 -3367
rect 7154 -3535 7188 -3501
rect 7346 -3535 7380 -3501
rect 7538 -3535 7572 -3501
rect 7730 -3535 7764 -3501
rect 7922 -3535 7956 -3501
rect 8114 -3535 8148 -3501
rect 16040 -3339 16074 -3337
rect 16040 -3537 16074 -3339
rect 16154 -3447 16188 -3367
rect 16250 -3447 16284 -3367
rect 16346 -3447 16380 -3367
rect 16442 -3447 16476 -3367
rect 16538 -3447 16572 -3367
rect 16634 -3447 16668 -3367
rect 16730 -3447 16764 -3367
rect 16826 -3447 16860 -3367
rect 16922 -3447 16956 -3367
rect 17018 -3447 17052 -3367
rect 17114 -3447 17148 -3367
rect 16154 -3535 16188 -3501
rect 16346 -3535 16380 -3501
rect 16538 -3535 16572 -3501
rect 16730 -3535 16764 -3501
rect 16922 -3535 16956 -3501
rect 17114 -3535 17148 -3501
rect 7040 -4873 7074 -4487
rect 7154 -4527 7188 -4493
rect 7346 -4527 7380 -4493
rect 7538 -4527 7572 -4493
rect 7730 -4527 7764 -4493
rect 7922 -4527 7956 -4493
rect 8114 -4527 8148 -4493
rect 7154 -4835 7188 -4587
rect 7250 -4835 7284 -4587
rect 7346 -4835 7380 -4587
rect 7442 -4835 7476 -4587
rect 7538 -4835 7572 -4587
rect 7634 -4835 7668 -4587
rect 7730 -4835 7764 -4587
rect 7826 -4835 7860 -4587
rect 7922 -4835 7956 -4587
rect 8018 -4835 8052 -4587
rect 8114 -4835 8148 -4587
rect 16040 -4873 16074 -4487
rect 16154 -4527 16188 -4493
rect 16346 -4527 16380 -4493
rect 16538 -4527 16572 -4493
rect 16730 -4527 16764 -4493
rect 16922 -4527 16956 -4493
rect 17114 -4527 17148 -4493
rect 16154 -4835 16188 -4587
rect 16250 -4835 16284 -4587
rect 16346 -4835 16380 -4587
rect 16442 -4835 16476 -4587
rect 16538 -4835 16572 -4587
rect 16634 -4835 16668 -4587
rect 16730 -4835 16764 -4587
rect 16826 -4835 16860 -4587
rect 16922 -4835 16956 -4587
rect 17018 -4835 17052 -4587
rect 17114 -4835 17148 -4587
rect 7040 -5139 7074 -5137
rect 7040 -5337 7074 -5139
rect 7154 -5247 7188 -5167
rect 7250 -5247 7284 -5167
rect 7346 -5247 7380 -5167
rect 7442 -5247 7476 -5167
rect 7538 -5247 7572 -5167
rect 7634 -5247 7668 -5167
rect 7730 -5247 7764 -5167
rect 7826 -5247 7860 -5167
rect 7922 -5247 7956 -5167
rect 8018 -5247 8052 -5167
rect 8114 -5247 8148 -5167
rect 7154 -5335 7188 -5301
rect 7346 -5335 7380 -5301
rect 7538 -5335 7572 -5301
rect 7730 -5335 7764 -5301
rect 7922 -5335 7956 -5301
rect 8114 -5335 8148 -5301
rect 16040 -5139 16074 -5137
rect 16040 -5337 16074 -5139
rect 16154 -5247 16188 -5167
rect 16250 -5247 16284 -5167
rect 16346 -5247 16380 -5167
rect 16442 -5247 16476 -5167
rect 16538 -5247 16572 -5167
rect 16634 -5247 16668 -5167
rect 16730 -5247 16764 -5167
rect 16826 -5247 16860 -5167
rect 16922 -5247 16956 -5167
rect 17018 -5247 17052 -5167
rect 17114 -5247 17148 -5167
rect 16154 -5335 16188 -5301
rect 16346 -5335 16380 -5301
rect 16538 -5335 16572 -5301
rect 16730 -5335 16764 -5301
rect 16922 -5335 16956 -5301
rect 17114 -5335 17148 -5301
rect 7040 -6673 7074 -6287
rect 7154 -6327 7188 -6293
rect 7346 -6327 7380 -6293
rect 7538 -6327 7572 -6293
rect 7730 -6327 7764 -6293
rect 7922 -6327 7956 -6293
rect 8114 -6327 8148 -6293
rect 7154 -6635 7188 -6387
rect 7250 -6635 7284 -6387
rect 7346 -6635 7380 -6387
rect 7442 -6635 7476 -6387
rect 7538 -6635 7572 -6387
rect 7634 -6635 7668 -6387
rect 7730 -6635 7764 -6387
rect 7826 -6635 7860 -6387
rect 7922 -6635 7956 -6387
rect 8018 -6635 8052 -6387
rect 8114 -6635 8148 -6387
rect 16040 -6673 16074 -6287
rect 16154 -6327 16188 -6293
rect 16346 -6327 16380 -6293
rect 16538 -6327 16572 -6293
rect 16730 -6327 16764 -6293
rect 16922 -6327 16956 -6293
rect 17114 -6327 17148 -6293
rect 16154 -6635 16188 -6387
rect 16250 -6635 16284 -6387
rect 16346 -6635 16380 -6387
rect 16442 -6635 16476 -6387
rect 16538 -6635 16572 -6387
rect 16634 -6635 16668 -6387
rect 16730 -6635 16764 -6387
rect 16826 -6635 16860 -6387
rect 16922 -6635 16956 -6387
rect 17018 -6635 17052 -6387
rect 17114 -6635 17148 -6387
rect 7040 -6939 7074 -6937
rect 7040 -7137 7074 -6939
rect 7154 -7047 7188 -6967
rect 7250 -7047 7284 -6967
rect 7346 -7047 7380 -6967
rect 7442 -7047 7476 -6967
rect 7538 -7047 7572 -6967
rect 7634 -7047 7668 -6967
rect 7730 -7047 7764 -6967
rect 7826 -7047 7860 -6967
rect 7922 -7047 7956 -6967
rect 8018 -7047 8052 -6967
rect 8114 -7047 8148 -6967
rect 7154 -7135 7188 -7101
rect 7346 -7135 7380 -7101
rect 7538 -7135 7572 -7101
rect 7730 -7135 7764 -7101
rect 7922 -7135 7956 -7101
rect 8114 -7135 8148 -7101
rect 16040 -6939 16074 -6937
rect 16040 -7137 16074 -6939
rect 16154 -7047 16188 -6967
rect 16250 -7047 16284 -6967
rect 16346 -7047 16380 -6967
rect 16442 -7047 16476 -6967
rect 16538 -7047 16572 -6967
rect 16634 -7047 16668 -6967
rect 16730 -7047 16764 -6967
rect 16826 -7047 16860 -6967
rect 16922 -7047 16956 -6967
rect 17018 -7047 17052 -6967
rect 17114 -7047 17148 -6967
rect 16154 -7135 16188 -7101
rect 16346 -7135 16380 -7101
rect 16538 -7135 16572 -7101
rect 16730 -7135 16764 -7101
rect 16922 -7135 16956 -7101
rect 17114 -7135 17148 -7101
rect -5544 -7824 -5500 -7790
rect -5366 -7824 -5322 -7790
rect -5188 -7824 -5144 -7790
rect -5010 -7824 -4966 -7790
rect -4832 -7824 -4788 -7790
rect -4654 -7824 -4610 -7790
rect -4476 -7824 -4432 -7790
rect -4298 -7824 -4254 -7790
rect -4120 -7824 -4076 -7790
rect -5628 -8130 -5594 -7874
rect -5450 -8130 -5416 -7874
rect -5272 -8130 -5238 -7874
rect -5094 -8130 -5060 -7874
rect -4916 -8130 -4882 -7874
rect -4738 -8130 -4704 -7874
rect -4560 -8130 -4526 -7874
rect -4382 -8130 -4348 -7874
rect -4204 -8130 -4170 -7874
rect -4026 -8130 -3992 -7874
rect -2089 -8082 -2045 -8048
rect -1911 -8082 -1867 -8048
rect -1733 -8082 -1689 -8048
rect -1555 -8082 -1511 -8048
rect -1377 -8082 -1333 -8048
rect -1199 -8082 -1155 -8048
rect -1021 -8082 -977 -8048
rect -843 -8082 -799 -8048
rect -665 -8082 -621 -8048
rect -487 -8082 -443 -8048
rect -309 -8082 -265 -8048
rect -131 -8082 -87 -8048
rect 47 -8082 91 -8048
rect 225 -8082 269 -8048
rect 403 -8082 447 -8048
rect 581 -8082 625 -8048
rect 759 -8082 803 -8048
rect 937 -8082 981 -8048
rect 1115 -8082 1159 -8048
rect 1293 -8082 1337 -8048
rect 1471 -8082 1515 -8048
rect 1649 -8082 1693 -8048
rect 1827 -8082 1871 -8048
rect 2005 -8082 2049 -8048
rect 2183 -8082 2227 -8048
rect 2361 -8082 2405 -8048
rect 2539 -8082 2583 -8048
rect 2717 -8082 2761 -8048
rect 2895 -8082 2939 -8048
rect 3073 -8082 3117 -8048
rect 3251 -8082 3295 -8048
rect 3429 -8082 3473 -8048
rect 3607 -8082 3651 -8048
rect 3785 -8082 3829 -8048
rect 3963 -8082 4007 -8048
rect -5544 -8214 -5500 -8180
rect -5366 -8214 -5322 -8180
rect -5188 -8214 -5144 -8180
rect -5010 -8214 -4966 -8180
rect -4832 -8214 -4788 -8180
rect -4654 -8214 -4610 -8180
rect -4476 -8214 -4432 -8180
rect -4298 -8214 -4254 -8180
rect -4120 -8214 -4076 -8180
rect -5544 -8374 -5500 -8340
rect -5366 -8374 -5322 -8340
rect -5188 -8374 -5144 -8340
rect -5010 -8374 -4966 -8340
rect -4832 -8374 -4788 -8340
rect -4654 -8374 -4610 -8340
rect -4476 -8374 -4432 -8340
rect -4298 -8374 -4254 -8340
rect -4120 -8374 -4076 -8340
rect -2173 -8388 -2139 -8132
rect -1995 -8388 -1961 -8132
rect -1817 -8388 -1783 -8132
rect -1639 -8388 -1605 -8132
rect -1461 -8388 -1427 -8132
rect -1283 -8388 -1249 -8132
rect -1105 -8388 -1071 -8132
rect -927 -8388 -893 -8132
rect -749 -8388 -715 -8132
rect -571 -8388 -537 -8132
rect -393 -8388 -359 -8132
rect -215 -8388 -181 -8132
rect -37 -8388 -3 -8132
rect 141 -8388 175 -8132
rect 319 -8388 353 -8132
rect 497 -8388 531 -8132
rect 675 -8388 709 -8132
rect 853 -8388 887 -8132
rect 1031 -8388 1065 -8132
rect 1209 -8388 1243 -8132
rect 1387 -8388 1421 -8132
rect 1565 -8388 1599 -8132
rect 1743 -8388 1777 -8132
rect 1921 -8388 1955 -8132
rect 2099 -8388 2133 -8132
rect 2277 -8388 2311 -8132
rect 2455 -8388 2489 -8132
rect 2633 -8388 2667 -8132
rect 2811 -8388 2845 -8132
rect 2989 -8388 3023 -8132
rect 3167 -8388 3201 -8132
rect 3345 -8388 3379 -8132
rect 3523 -8388 3557 -8132
rect 3701 -8388 3735 -8132
rect 3879 -8388 3913 -8132
rect 4057 -8388 4091 -8132
rect -5628 -8680 -5594 -8424
rect -5450 -8680 -5416 -8424
rect -5272 -8680 -5238 -8424
rect -5094 -8680 -5060 -8424
rect -4916 -8680 -4882 -8424
rect -4738 -8680 -4704 -8424
rect -4560 -8680 -4526 -8424
rect -4382 -8680 -4348 -8424
rect -4204 -8680 -4170 -8424
rect -4026 -8680 -3992 -8424
rect -2089 -8472 -2045 -8438
rect -1911 -8472 -1867 -8438
rect -1733 -8472 -1689 -8438
rect -1555 -8472 -1511 -8438
rect -1377 -8472 -1333 -8438
rect -1199 -8472 -1155 -8438
rect -1021 -8472 -977 -8438
rect -843 -8472 -799 -8438
rect -665 -8472 -621 -8438
rect -487 -8472 -443 -8438
rect -309 -8472 -265 -8438
rect -131 -8472 -87 -8438
rect 47 -8472 91 -8438
rect 225 -8472 269 -8438
rect 403 -8472 447 -8438
rect 581 -8472 625 -8438
rect 759 -8472 803 -8438
rect 937 -8472 981 -8438
rect 1115 -8472 1159 -8438
rect 1293 -8472 1337 -8438
rect 1471 -8472 1515 -8438
rect 1649 -8472 1693 -8438
rect 1827 -8472 1871 -8438
rect 2005 -8472 2049 -8438
rect 2183 -8472 2227 -8438
rect 2361 -8472 2405 -8438
rect 2539 -8472 2583 -8438
rect 2717 -8472 2761 -8438
rect 2895 -8472 2939 -8438
rect 3073 -8472 3117 -8438
rect 3251 -8472 3295 -8438
rect 3429 -8472 3473 -8438
rect 3607 -8472 3651 -8438
rect 3785 -8472 3829 -8438
rect 3963 -8472 4007 -8438
rect -5544 -8764 -5500 -8730
rect -5366 -8764 -5322 -8730
rect -5188 -8764 -5144 -8730
rect -5010 -8764 -4966 -8730
rect -4832 -8764 -4788 -8730
rect -4654 -8764 -4610 -8730
rect -4476 -8764 -4432 -8730
rect -4298 -8764 -4254 -8730
rect -4120 -8764 -4076 -8730
rect 6596 -8844 6640 -8810
rect 6774 -8844 6818 -8810
rect 6952 -8844 6996 -8810
rect 7130 -8844 7174 -8810
rect 7308 -8844 7352 -8810
rect 7486 -8844 7530 -8810
rect 7664 -8844 7708 -8810
rect 7842 -8844 7886 -8810
rect 8020 -8844 8064 -8810
rect 8198 -8844 8242 -8810
rect 8376 -8844 8420 -8810
rect 8554 -8844 8598 -8810
rect 8732 -8844 8776 -8810
rect 8910 -8844 8954 -8810
rect 9088 -8844 9132 -8810
rect 9266 -8844 9310 -8810
rect 10856 -8874 10900 -8840
rect 11148 -8874 11192 -8840
rect 11440 -8874 11484 -8840
rect 11732 -8874 11776 -8840
rect 12024 -8874 12068 -8840
rect 12316 -8874 12360 -8840
rect 12608 -8874 12652 -8840
rect -5544 -8924 -5500 -8890
rect -5366 -8924 -5322 -8890
rect -5188 -8924 -5144 -8890
rect -5010 -8924 -4966 -8890
rect -4832 -8924 -4788 -8890
rect -4654 -8924 -4610 -8890
rect -4476 -8924 -4432 -8890
rect -4298 -8924 -4254 -8890
rect -4120 -8924 -4076 -8890
rect -5628 -9230 -5594 -8974
rect -5450 -9230 -5416 -8974
rect -5272 -9230 -5238 -8974
rect -5094 -9230 -5060 -8974
rect -4916 -9230 -4882 -8974
rect -4738 -9230 -4704 -8974
rect -4560 -9230 -4526 -8974
rect -4382 -9230 -4348 -8974
rect -4204 -9230 -4170 -8974
rect -4026 -9230 -3992 -8974
rect -2089 -9082 -2045 -9048
rect -1911 -9082 -1867 -9048
rect -1733 -9082 -1689 -9048
rect -1555 -9082 -1511 -9048
rect -1377 -9082 -1333 -9048
rect -1199 -9082 -1155 -9048
rect -1021 -9082 -977 -9048
rect -843 -9082 -799 -9048
rect -665 -9082 -621 -9048
rect -487 -9082 -443 -9048
rect -309 -9082 -265 -9048
rect -131 -9082 -87 -9048
rect 47 -9082 91 -9048
rect 225 -9082 269 -9048
rect 403 -9082 447 -9048
rect 581 -9082 625 -9048
rect 759 -9082 803 -9048
rect 937 -9082 981 -9048
rect 1115 -9082 1159 -9048
rect 1293 -9082 1337 -9048
rect 1471 -9082 1515 -9048
rect 1649 -9082 1693 -9048
rect 1827 -9082 1871 -9048
rect 2005 -9082 2049 -9048
rect 2183 -9082 2227 -9048
rect 2361 -9082 2405 -9048
rect 2539 -9082 2583 -9048
rect 2717 -9082 2761 -9048
rect 2895 -9082 2939 -9048
rect 3073 -9082 3117 -9048
rect 3251 -9082 3295 -9048
rect 3429 -9082 3473 -9048
rect 3607 -9082 3651 -9048
rect 3785 -9082 3829 -9048
rect 3963 -9082 4007 -9048
rect -5544 -9314 -5500 -9280
rect -5366 -9314 -5322 -9280
rect -5188 -9314 -5144 -9280
rect -5010 -9314 -4966 -9280
rect -4832 -9314 -4788 -9280
rect -4654 -9314 -4610 -9280
rect -4476 -9314 -4432 -9280
rect -4298 -9314 -4254 -9280
rect -4120 -9314 -4076 -9280
rect -5544 -9474 -5500 -9440
rect -5366 -9474 -5322 -9440
rect -5188 -9474 -5144 -9440
rect -5010 -9474 -4966 -9440
rect -4832 -9474 -4788 -9440
rect -4654 -9474 -4610 -9440
rect -4476 -9474 -4432 -9440
rect -4298 -9474 -4254 -9440
rect -4120 -9474 -4076 -9440
rect -2985 -9454 -2807 -9276
rect -2173 -9388 -2139 -9132
rect -1995 -9388 -1961 -9132
rect -1817 -9388 -1783 -9132
rect -1639 -9388 -1605 -9132
rect -1461 -9388 -1427 -9132
rect -1283 -9388 -1249 -9132
rect -1105 -9388 -1071 -9132
rect -927 -9388 -893 -9132
rect -749 -9388 -715 -9132
rect -571 -9388 -537 -9132
rect -393 -9388 -359 -9132
rect -215 -9388 -181 -9132
rect -37 -9388 -3 -9132
rect 141 -9388 175 -9132
rect 319 -9388 353 -9132
rect 497 -9388 531 -9132
rect 675 -9388 709 -9132
rect 853 -9388 887 -9132
rect 1031 -9388 1065 -9132
rect 1209 -9388 1243 -9132
rect 1387 -9388 1421 -9132
rect 1565 -9388 1599 -9132
rect 1743 -9388 1777 -9132
rect 1921 -9388 1955 -9132
rect 2099 -9388 2133 -9132
rect 2277 -9388 2311 -9132
rect 2455 -9388 2489 -9132
rect 2633 -9388 2667 -9132
rect 2811 -9388 2845 -9132
rect 2989 -9388 3023 -9132
rect 3167 -9388 3201 -9132
rect 3345 -9388 3379 -9132
rect 3523 -9388 3557 -9132
rect 3701 -9388 3735 -9132
rect 3879 -9388 3913 -9132
rect 4057 -9388 4091 -9132
rect 6512 -9150 6546 -8894
rect 6690 -9150 6724 -8894
rect 6868 -9150 6902 -8894
rect 7046 -9150 7080 -8894
rect 7224 -9150 7258 -8894
rect 7402 -9150 7436 -8894
rect 7580 -9150 7614 -8894
rect 7758 -9150 7792 -8894
rect 7936 -9150 7970 -8894
rect 8114 -9150 8148 -8894
rect 8292 -9150 8326 -8894
rect 8470 -9150 8504 -8894
rect 8648 -9150 8682 -8894
rect 8826 -9150 8860 -8894
rect 9004 -9150 9038 -8894
rect 9182 -9150 9216 -8894
rect 9360 -9150 9394 -8894
rect 6596 -9234 6640 -9200
rect 6774 -9234 6818 -9200
rect 6952 -9234 6996 -9200
rect 7130 -9234 7174 -9200
rect 7308 -9234 7352 -9200
rect 7486 -9234 7530 -9200
rect 7664 -9234 7708 -9200
rect 7842 -9234 7886 -9200
rect 8020 -9234 8064 -9200
rect 8198 -9234 8242 -9200
rect 8376 -9234 8420 -9200
rect 8554 -9234 8598 -9200
rect 8732 -9234 8776 -9200
rect 8910 -9234 8954 -9200
rect 9088 -9234 9132 -9200
rect 9266 -9234 9310 -9200
rect 9982 -9369 10160 -9191
rect 10772 -9180 10806 -8924
rect 10950 -9180 10984 -8924
rect 11064 -9180 11098 -8924
rect 11242 -9180 11276 -8924
rect 11356 -9180 11390 -8924
rect 11534 -9180 11568 -8924
rect 11648 -9180 11682 -8924
rect 11826 -9180 11860 -8924
rect 11940 -9180 11974 -8924
rect 12118 -9180 12152 -8924
rect 12232 -9180 12266 -8924
rect 12410 -9180 12444 -8924
rect 12524 -9180 12558 -8924
rect 12702 -9180 12736 -8924
rect 10856 -9264 10900 -9230
rect 11148 -9264 11192 -9230
rect 11440 -9264 11484 -9230
rect 11732 -9264 11776 -9230
rect 12024 -9264 12068 -9230
rect 12316 -9264 12360 -9230
rect 12608 -9264 12652 -9230
rect -2089 -9472 -2045 -9438
rect -1911 -9472 -1867 -9438
rect -1733 -9472 -1689 -9438
rect -1555 -9472 -1511 -9438
rect -1377 -9472 -1333 -9438
rect -1199 -9472 -1155 -9438
rect -1021 -9472 -977 -9438
rect -843 -9472 -799 -9438
rect -665 -9472 -621 -9438
rect -487 -9472 -443 -9438
rect -309 -9472 -265 -9438
rect -131 -9472 -87 -9438
rect 47 -9472 91 -9438
rect 225 -9472 269 -9438
rect 403 -9472 447 -9438
rect 581 -9472 625 -9438
rect 759 -9472 803 -9438
rect 937 -9472 981 -9438
rect 1115 -9472 1159 -9438
rect 1293 -9472 1337 -9438
rect 1471 -9472 1515 -9438
rect 1649 -9472 1693 -9438
rect 1827 -9472 1871 -9438
rect 2005 -9472 2049 -9438
rect 2183 -9472 2227 -9438
rect 2361 -9472 2405 -9438
rect 2539 -9472 2583 -9438
rect 2717 -9472 2761 -9438
rect 2895 -9472 2939 -9438
rect 3073 -9472 3117 -9438
rect 3251 -9472 3295 -9438
rect 3429 -9472 3473 -9438
rect 3607 -9472 3651 -9438
rect 3785 -9472 3829 -9438
rect 3963 -9472 4007 -9438
rect -5628 -9780 -5594 -9524
rect -5450 -9780 -5416 -9524
rect -5272 -9780 -5238 -9524
rect -5094 -9780 -5060 -9524
rect -4916 -9780 -4882 -9524
rect -4738 -9780 -4704 -9524
rect -4560 -9780 -4526 -9524
rect -4382 -9780 -4348 -9524
rect -4204 -9780 -4170 -9524
rect -4026 -9780 -3992 -9524
rect 10856 -9644 10900 -9610
rect 11148 -9644 11192 -9610
rect 11440 -9644 11484 -9610
rect 11732 -9644 11776 -9610
rect 12024 -9644 12068 -9610
rect 12316 -9644 12360 -9610
rect 12608 -9644 12652 -9610
rect 6596 -9744 6640 -9710
rect 6774 -9744 6818 -9710
rect 6952 -9744 6996 -9710
rect 7130 -9744 7174 -9710
rect 7308 -9744 7352 -9710
rect 7486 -9744 7530 -9710
rect 7664 -9744 7708 -9710
rect 7842 -9744 7886 -9710
rect 8020 -9744 8064 -9710
rect 8198 -9744 8242 -9710
rect 8376 -9744 8420 -9710
rect 8554 -9744 8598 -9710
rect 8732 -9744 8776 -9710
rect 8910 -9744 8954 -9710
rect 9088 -9744 9132 -9710
rect 9266 -9744 9310 -9710
rect -5544 -9864 -5500 -9830
rect -5366 -9864 -5322 -9830
rect -5188 -9864 -5144 -9830
rect -5010 -9864 -4966 -9830
rect -4832 -9864 -4788 -9830
rect -4654 -9864 -4610 -9830
rect -4476 -9864 -4432 -9830
rect -4298 -9864 -4254 -9830
rect -4120 -9864 -4076 -9830
rect -5544 -10024 -5500 -9990
rect -5366 -10024 -5322 -9990
rect -5188 -10024 -5144 -9990
rect -5010 -10024 -4966 -9990
rect -4832 -10024 -4788 -9990
rect -4654 -10024 -4610 -9990
rect -4476 -10024 -4432 -9990
rect -4298 -10024 -4254 -9990
rect -4120 -10024 -4076 -9990
rect -5628 -10330 -5594 -10074
rect -5450 -10330 -5416 -10074
rect -5272 -10330 -5238 -10074
rect -5094 -10330 -5060 -10074
rect -4916 -10330 -4882 -10074
rect -4738 -10330 -4704 -10074
rect -4560 -10330 -4526 -10074
rect -4382 -10330 -4348 -10074
rect -4204 -10330 -4170 -10074
rect -4026 -10330 -3992 -10074
rect -2089 -10082 -2045 -10048
rect -1911 -10082 -1867 -10048
rect -1733 -10082 -1689 -10048
rect -1555 -10082 -1511 -10048
rect -1377 -10082 -1333 -10048
rect -1199 -10082 -1155 -10048
rect -1021 -10082 -977 -10048
rect -843 -10082 -799 -10048
rect -665 -10082 -621 -10048
rect -487 -10082 -443 -10048
rect -309 -10082 -265 -10048
rect -131 -10082 -87 -10048
rect 47 -10082 91 -10048
rect 225 -10082 269 -10048
rect 403 -10082 447 -10048
rect 581 -10082 625 -10048
rect 759 -10082 803 -10048
rect 937 -10082 981 -10048
rect 1115 -10082 1159 -10048
rect 1293 -10082 1337 -10048
rect 1471 -10082 1515 -10048
rect 1649 -10082 1693 -10048
rect 1827 -10082 1871 -10048
rect 2005 -10082 2049 -10048
rect 2183 -10082 2227 -10048
rect 2361 -10082 2405 -10048
rect 2539 -10082 2583 -10048
rect 2717 -10082 2761 -10048
rect 2895 -10082 2939 -10048
rect 3073 -10082 3117 -10048
rect 3251 -10082 3295 -10048
rect 3429 -10082 3473 -10048
rect 3607 -10082 3651 -10048
rect 3785 -10082 3829 -10048
rect 3963 -10082 4007 -10048
rect 6512 -10050 6546 -9794
rect 6690 -10050 6724 -9794
rect 6868 -10050 6902 -9794
rect 7046 -10050 7080 -9794
rect 7224 -10050 7258 -9794
rect 7402 -10050 7436 -9794
rect 7580 -10050 7614 -9794
rect 7758 -10050 7792 -9794
rect 7936 -10050 7970 -9794
rect 8114 -10050 8148 -9794
rect 8292 -10050 8326 -9794
rect 8470 -10050 8504 -9794
rect 8648 -10050 8682 -9794
rect 8826 -10050 8860 -9794
rect 9004 -10050 9038 -9794
rect 9182 -10050 9216 -9794
rect 9360 -10050 9394 -9794
rect 10772 -9950 10806 -9694
rect 10950 -9950 10984 -9694
rect 11064 -9950 11098 -9694
rect 11242 -9950 11276 -9694
rect 11356 -9950 11390 -9694
rect 11534 -9950 11568 -9694
rect 11648 -9950 11682 -9694
rect 11826 -9950 11860 -9694
rect 11940 -9950 11974 -9694
rect 12118 -9950 12152 -9694
rect 12232 -9950 12266 -9694
rect 12410 -9950 12444 -9694
rect 12524 -9950 12558 -9694
rect 12702 -9950 12736 -9694
rect 10856 -10034 10900 -10000
rect 11148 -10034 11192 -10000
rect 11440 -10034 11484 -10000
rect 11732 -10034 11776 -10000
rect 12024 -10034 12068 -10000
rect 12316 -10034 12360 -10000
rect 12608 -10034 12652 -10000
rect -5544 -10414 -5500 -10380
rect -5366 -10414 -5322 -10380
rect -5188 -10414 -5144 -10380
rect -5010 -10414 -4966 -10380
rect -4832 -10414 -4788 -10380
rect -4654 -10414 -4610 -10380
rect -4476 -10414 -4432 -10380
rect -4298 -10414 -4254 -10380
rect -4120 -10414 -4076 -10380
rect -2173 -10388 -2139 -10132
rect -1995 -10388 -1961 -10132
rect -1817 -10388 -1783 -10132
rect -1639 -10388 -1605 -10132
rect -1461 -10388 -1427 -10132
rect -1283 -10388 -1249 -10132
rect -1105 -10388 -1071 -10132
rect -927 -10388 -893 -10132
rect -749 -10388 -715 -10132
rect -571 -10388 -537 -10132
rect -393 -10388 -359 -10132
rect -215 -10388 -181 -10132
rect -37 -10388 -3 -10132
rect 141 -10388 175 -10132
rect 319 -10388 353 -10132
rect 497 -10388 531 -10132
rect 675 -10388 709 -10132
rect 853 -10388 887 -10132
rect 1031 -10388 1065 -10132
rect 1209 -10388 1243 -10132
rect 1387 -10388 1421 -10132
rect 1565 -10388 1599 -10132
rect 1743 -10388 1777 -10132
rect 1921 -10388 1955 -10132
rect 2099 -10388 2133 -10132
rect 2277 -10388 2311 -10132
rect 2455 -10388 2489 -10132
rect 2633 -10388 2667 -10132
rect 2811 -10388 2845 -10132
rect 2989 -10388 3023 -10132
rect 3167 -10388 3201 -10132
rect 3345 -10388 3379 -10132
rect 3523 -10388 3557 -10132
rect 3701 -10388 3735 -10132
rect 3879 -10388 3913 -10132
rect 4057 -10388 4091 -10132
rect 6596 -10134 6640 -10100
rect 6774 -10134 6818 -10100
rect 6952 -10134 6996 -10100
rect 7130 -10134 7174 -10100
rect 7308 -10134 7352 -10100
rect 7486 -10134 7530 -10100
rect 7664 -10134 7708 -10100
rect 7842 -10134 7886 -10100
rect 8020 -10134 8064 -10100
rect 8198 -10134 8242 -10100
rect 8376 -10134 8420 -10100
rect 8554 -10134 8598 -10100
rect 8732 -10134 8776 -10100
rect 8910 -10134 8954 -10100
rect 9088 -10134 9132 -10100
rect 9266 -10134 9310 -10100
rect 10856 -10414 10900 -10380
rect 11148 -10414 11192 -10380
rect 11440 -10414 11484 -10380
rect 11732 -10414 11776 -10380
rect 12024 -10414 12068 -10380
rect 12316 -10414 12360 -10380
rect 12608 -10414 12652 -10380
rect -2089 -10472 -2045 -10438
rect -1911 -10472 -1867 -10438
rect -1733 -10472 -1689 -10438
rect -1555 -10472 -1511 -10438
rect -1377 -10472 -1333 -10438
rect -1199 -10472 -1155 -10438
rect -1021 -10472 -977 -10438
rect -843 -10472 -799 -10438
rect -665 -10472 -621 -10438
rect -487 -10472 -443 -10438
rect -309 -10472 -265 -10438
rect -131 -10472 -87 -10438
rect 47 -10472 91 -10438
rect 225 -10472 269 -10438
rect 403 -10472 447 -10438
rect 581 -10472 625 -10438
rect 759 -10472 803 -10438
rect 937 -10472 981 -10438
rect 1115 -10472 1159 -10438
rect 1293 -10472 1337 -10438
rect 1471 -10472 1515 -10438
rect 1649 -10472 1693 -10438
rect 1827 -10472 1871 -10438
rect 2005 -10472 2049 -10438
rect 2183 -10472 2227 -10438
rect 2361 -10472 2405 -10438
rect 2539 -10472 2583 -10438
rect 2717 -10472 2761 -10438
rect 2895 -10472 2939 -10438
rect 3073 -10472 3117 -10438
rect 3251 -10472 3295 -10438
rect 3429 -10472 3473 -10438
rect 3607 -10472 3651 -10438
rect 3785 -10472 3829 -10438
rect 3963 -10472 4007 -10438
rect -5544 -10574 -5500 -10540
rect -5366 -10574 -5322 -10540
rect -5188 -10574 -5144 -10540
rect -5010 -10574 -4966 -10540
rect -4832 -10574 -4788 -10540
rect -4654 -10574 -4610 -10540
rect -4476 -10574 -4432 -10540
rect -4298 -10574 -4254 -10540
rect -4120 -10574 -4076 -10540
rect -5628 -10880 -5594 -10624
rect -5450 -10880 -5416 -10624
rect -5272 -10880 -5238 -10624
rect -5094 -10880 -5060 -10624
rect -4916 -10880 -4882 -10624
rect -4738 -10880 -4704 -10624
rect -4560 -10880 -4526 -10624
rect -4382 -10880 -4348 -10624
rect -4204 -10880 -4170 -10624
rect -4026 -10880 -3992 -10624
rect 6596 -10644 6640 -10610
rect 6774 -10644 6818 -10610
rect 6952 -10644 6996 -10610
rect 7130 -10644 7174 -10610
rect 7308 -10644 7352 -10610
rect 7486 -10644 7530 -10610
rect 7664 -10644 7708 -10610
rect 7842 -10644 7886 -10610
rect 8020 -10644 8064 -10610
rect 8198 -10644 8242 -10610
rect 8376 -10644 8420 -10610
rect 8554 -10644 8598 -10610
rect 8732 -10644 8776 -10610
rect 8910 -10644 8954 -10610
rect 9088 -10644 9132 -10610
rect 9266 -10644 9310 -10610
rect -5544 -10964 -5500 -10930
rect -5366 -10964 -5322 -10930
rect -5188 -10964 -5144 -10930
rect -5010 -10964 -4966 -10930
rect -4832 -10964 -4788 -10930
rect -4654 -10964 -4610 -10930
rect -4476 -10964 -4432 -10930
rect -4298 -10964 -4254 -10930
rect -4120 -10964 -4076 -10930
rect 6512 -10950 6546 -10694
rect 6690 -10950 6724 -10694
rect 6868 -10950 6902 -10694
rect 7046 -10950 7080 -10694
rect 7224 -10950 7258 -10694
rect 7402 -10950 7436 -10694
rect 7580 -10950 7614 -10694
rect 7758 -10950 7792 -10694
rect 7936 -10950 7970 -10694
rect 8114 -10950 8148 -10694
rect 8292 -10950 8326 -10694
rect 8470 -10950 8504 -10694
rect 8648 -10950 8682 -10694
rect 8826 -10950 8860 -10694
rect 9004 -10950 9038 -10694
rect 9182 -10950 9216 -10694
rect 9360 -10950 9394 -10694
rect 10772 -10720 10806 -10464
rect 10950 -10720 10984 -10464
rect 11064 -10720 11098 -10464
rect 11242 -10720 11276 -10464
rect 11356 -10720 11390 -10464
rect 11534 -10720 11568 -10464
rect 11648 -10720 11682 -10464
rect 11826 -10720 11860 -10464
rect 11940 -10720 11974 -10464
rect 12118 -10720 12152 -10464
rect 12232 -10720 12266 -10464
rect 12410 -10720 12444 -10464
rect 12524 -10720 12558 -10464
rect 12702 -10720 12736 -10464
rect 10856 -10804 10900 -10770
rect 11148 -10804 11192 -10770
rect 11440 -10804 11484 -10770
rect 11732 -10804 11776 -10770
rect 12024 -10804 12068 -10770
rect 12316 -10804 12360 -10770
rect 12608 -10804 12652 -10770
rect 6596 -11034 6640 -11000
rect 6774 -11034 6818 -11000
rect 6952 -11034 6996 -11000
rect 7130 -11034 7174 -11000
rect 7308 -11034 7352 -11000
rect 7486 -11034 7530 -11000
rect 7664 -11034 7708 -11000
rect 7842 -11034 7886 -11000
rect 8020 -11034 8064 -11000
rect 8198 -11034 8242 -11000
rect 8376 -11034 8420 -11000
rect 8554 -11034 8598 -11000
rect 8732 -11034 8776 -11000
rect 8910 -11034 8954 -11000
rect 9088 -11034 9132 -11000
rect 9266 -11034 9310 -11000
rect -2089 -11082 -2045 -11048
rect -1911 -11082 -1867 -11048
rect -1733 -11082 -1689 -11048
rect -1555 -11082 -1511 -11048
rect -1377 -11082 -1333 -11048
rect -1199 -11082 -1155 -11048
rect -1021 -11082 -977 -11048
rect -843 -11082 -799 -11048
rect -665 -11082 -621 -11048
rect -487 -11082 -443 -11048
rect -309 -11082 -265 -11048
rect -131 -11082 -87 -11048
rect 47 -11082 91 -11048
rect 225 -11082 269 -11048
rect 403 -11082 447 -11048
rect 581 -11082 625 -11048
rect 759 -11082 803 -11048
rect 937 -11082 981 -11048
rect 1115 -11082 1159 -11048
rect 1293 -11082 1337 -11048
rect 1471 -11082 1515 -11048
rect 1649 -11082 1693 -11048
rect 1827 -11082 1871 -11048
rect 2005 -11082 2049 -11048
rect 2183 -11082 2227 -11048
rect 2361 -11082 2405 -11048
rect 2539 -11082 2583 -11048
rect 2717 -11082 2761 -11048
rect 2895 -11082 2939 -11048
rect 3073 -11082 3117 -11048
rect 3251 -11082 3295 -11048
rect 3429 -11082 3473 -11048
rect 3607 -11082 3651 -11048
rect 3785 -11082 3829 -11048
rect 3963 -11082 4007 -11048
rect -5544 -11124 -5500 -11090
rect -5366 -11124 -5322 -11090
rect -5188 -11124 -5144 -11090
rect -5010 -11124 -4966 -11090
rect -4832 -11124 -4788 -11090
rect -4654 -11124 -4610 -11090
rect -4476 -11124 -4432 -11090
rect -4298 -11124 -4254 -11090
rect -4120 -11124 -4076 -11090
rect -5628 -11430 -5594 -11174
rect -5450 -11430 -5416 -11174
rect -5272 -11430 -5238 -11174
rect -5094 -11430 -5060 -11174
rect -4916 -11430 -4882 -11174
rect -4738 -11430 -4704 -11174
rect -4560 -11430 -4526 -11174
rect -4382 -11430 -4348 -11174
rect -4204 -11430 -4170 -11174
rect -4026 -11430 -3992 -11174
rect -2985 -11454 -2807 -11276
rect -2173 -11388 -2139 -11132
rect -1995 -11388 -1961 -11132
rect -1817 -11388 -1783 -11132
rect -1639 -11388 -1605 -11132
rect -1461 -11388 -1427 -11132
rect -1283 -11388 -1249 -11132
rect -1105 -11388 -1071 -11132
rect -927 -11388 -893 -11132
rect -749 -11388 -715 -11132
rect -571 -11388 -537 -11132
rect -393 -11388 -359 -11132
rect -215 -11388 -181 -11132
rect -37 -11388 -3 -11132
rect 141 -11388 175 -11132
rect 319 -11388 353 -11132
rect 497 -11388 531 -11132
rect 675 -11388 709 -11132
rect 853 -11388 887 -11132
rect 1031 -11388 1065 -11132
rect 1209 -11388 1243 -11132
rect 1387 -11388 1421 -11132
rect 1565 -11388 1599 -11132
rect 1743 -11388 1777 -11132
rect 1921 -11388 1955 -11132
rect 2099 -11388 2133 -11132
rect 2277 -11388 2311 -11132
rect 2455 -11388 2489 -11132
rect 2633 -11388 2667 -11132
rect 2811 -11388 2845 -11132
rect 2989 -11388 3023 -11132
rect 3167 -11388 3201 -11132
rect 3345 -11388 3379 -11132
rect 3523 -11388 3557 -11132
rect 3701 -11388 3735 -11132
rect 3879 -11388 3913 -11132
rect 4057 -11388 4091 -11132
rect 5686 -11329 5864 -11151
rect 10856 -11184 10900 -11150
rect 11148 -11184 11192 -11150
rect 11440 -11184 11484 -11150
rect 11732 -11184 11776 -11150
rect 12024 -11184 12068 -11150
rect 12316 -11184 12360 -11150
rect 12608 -11184 12652 -11150
rect 9982 -11369 10160 -11191
rect -2089 -11472 -2045 -11438
rect -1911 -11472 -1867 -11438
rect -1733 -11472 -1689 -11438
rect -1555 -11472 -1511 -11438
rect -1377 -11472 -1333 -11438
rect -1199 -11472 -1155 -11438
rect -1021 -11472 -977 -11438
rect -843 -11472 -799 -11438
rect -665 -11472 -621 -11438
rect -487 -11472 -443 -11438
rect -309 -11472 -265 -11438
rect -131 -11472 -87 -11438
rect 47 -11472 91 -11438
rect 225 -11472 269 -11438
rect 403 -11472 447 -11438
rect 581 -11472 625 -11438
rect 759 -11472 803 -11438
rect 937 -11472 981 -11438
rect 1115 -11472 1159 -11438
rect 1293 -11472 1337 -11438
rect 1471 -11472 1515 -11438
rect 1649 -11472 1693 -11438
rect 1827 -11472 1871 -11438
rect 2005 -11472 2049 -11438
rect 2183 -11472 2227 -11438
rect 2361 -11472 2405 -11438
rect 2539 -11472 2583 -11438
rect 2717 -11472 2761 -11438
rect 2895 -11472 2939 -11438
rect 3073 -11472 3117 -11438
rect 3251 -11472 3295 -11438
rect 3429 -11472 3473 -11438
rect 3607 -11472 3651 -11438
rect 3785 -11472 3829 -11438
rect 3963 -11472 4007 -11438
rect -5544 -11514 -5500 -11480
rect -5366 -11514 -5322 -11480
rect -5188 -11514 -5144 -11480
rect -5010 -11514 -4966 -11480
rect -4832 -11514 -4788 -11480
rect -4654 -11514 -4610 -11480
rect -4476 -11514 -4432 -11480
rect -4298 -11514 -4254 -11480
rect -4120 -11514 -4076 -11480
rect 10772 -11490 10806 -11234
rect 10950 -11490 10984 -11234
rect 11064 -11490 11098 -11234
rect 11242 -11490 11276 -11234
rect 11356 -11490 11390 -11234
rect 11534 -11490 11568 -11234
rect 11648 -11490 11682 -11234
rect 11826 -11490 11860 -11234
rect 11940 -11490 11974 -11234
rect 12118 -11490 12152 -11234
rect 12232 -11490 12266 -11234
rect 12410 -11490 12444 -11234
rect 12524 -11490 12558 -11234
rect 12702 -11490 12736 -11234
rect 6596 -11544 6640 -11510
rect 6774 -11544 6818 -11510
rect 6952 -11544 6996 -11510
rect 7130 -11544 7174 -11510
rect 7308 -11544 7352 -11510
rect 7486 -11544 7530 -11510
rect 7664 -11544 7708 -11510
rect 7842 -11544 7886 -11510
rect 8020 -11544 8064 -11510
rect 8198 -11544 8242 -11510
rect 8376 -11544 8420 -11510
rect 8554 -11544 8598 -11510
rect 8732 -11544 8776 -11510
rect 8910 -11544 8954 -11510
rect 9088 -11544 9132 -11510
rect 9266 -11544 9310 -11510
rect 10856 -11574 10900 -11540
rect 11148 -11574 11192 -11540
rect 11440 -11574 11484 -11540
rect 11732 -11574 11776 -11540
rect 12024 -11574 12068 -11540
rect 12316 -11574 12360 -11540
rect 12608 -11574 12652 -11540
rect -5544 -11674 -5500 -11640
rect -5366 -11674 -5322 -11640
rect -5188 -11674 -5144 -11640
rect -5010 -11674 -4966 -11640
rect -4832 -11674 -4788 -11640
rect -4654 -11674 -4610 -11640
rect -4476 -11674 -4432 -11640
rect -4298 -11674 -4254 -11640
rect -4120 -11674 -4076 -11640
rect -5628 -11980 -5594 -11724
rect -5450 -11980 -5416 -11724
rect -5272 -11980 -5238 -11724
rect -5094 -11980 -5060 -11724
rect -4916 -11980 -4882 -11724
rect -4738 -11980 -4704 -11724
rect -4560 -11980 -4526 -11724
rect -4382 -11980 -4348 -11724
rect -4204 -11980 -4170 -11724
rect -4026 -11980 -3992 -11724
rect 6512 -11850 6546 -11594
rect 6690 -11850 6724 -11594
rect 6868 -11850 6902 -11594
rect 7046 -11850 7080 -11594
rect 7224 -11850 7258 -11594
rect 7402 -11850 7436 -11594
rect 7580 -11850 7614 -11594
rect 7758 -11850 7792 -11594
rect 7936 -11850 7970 -11594
rect 8114 -11850 8148 -11594
rect 8292 -11850 8326 -11594
rect 8470 -11850 8504 -11594
rect 8648 -11850 8682 -11594
rect 8826 -11850 8860 -11594
rect 9004 -11850 9038 -11594
rect 9182 -11850 9216 -11594
rect 9360 -11850 9394 -11594
rect 6596 -11934 6640 -11900
rect 6774 -11934 6818 -11900
rect 6952 -11934 6996 -11900
rect 7130 -11934 7174 -11900
rect 7308 -11934 7352 -11900
rect 7486 -11934 7530 -11900
rect 7664 -11934 7708 -11900
rect 7842 -11934 7886 -11900
rect 8020 -11934 8064 -11900
rect 8198 -11934 8242 -11900
rect 8376 -11934 8420 -11900
rect 8554 -11934 8598 -11900
rect 8732 -11934 8776 -11900
rect 8910 -11934 8954 -11900
rect 9088 -11934 9132 -11900
rect 9266 -11934 9310 -11900
rect -5544 -12064 -5500 -12030
rect -5366 -12064 -5322 -12030
rect -5188 -12064 -5144 -12030
rect -5010 -12064 -4966 -12030
rect -4832 -12064 -4788 -12030
rect -4654 -12064 -4610 -12030
rect -4476 -12064 -4432 -12030
rect -4298 -12064 -4254 -12030
rect -4120 -12064 -4076 -12030
rect -2089 -12082 -2045 -12048
rect -1911 -12082 -1867 -12048
rect -1733 -12082 -1689 -12048
rect -1555 -12082 -1511 -12048
rect -1377 -12082 -1333 -12048
rect -1199 -12082 -1155 -12048
rect -1021 -12082 -977 -12048
rect -843 -12082 -799 -12048
rect -665 -12082 -621 -12048
rect -487 -12082 -443 -12048
rect -309 -12082 -265 -12048
rect -131 -12082 -87 -12048
rect 47 -12082 91 -12048
rect 225 -12082 269 -12048
rect 403 -12082 447 -12048
rect 581 -12082 625 -12048
rect 759 -12082 803 -12048
rect 937 -12082 981 -12048
rect 1115 -12082 1159 -12048
rect 1293 -12082 1337 -12048
rect 1471 -12082 1515 -12048
rect 1649 -12082 1693 -12048
rect 1827 -12082 1871 -12048
rect 2005 -12082 2049 -12048
rect 2183 -12082 2227 -12048
rect 2361 -12082 2405 -12048
rect 2539 -12082 2583 -12048
rect 2717 -12082 2761 -12048
rect 2895 -12082 2939 -12048
rect 3073 -12082 3117 -12048
rect 3251 -12082 3295 -12048
rect 3429 -12082 3473 -12048
rect 3607 -12082 3651 -12048
rect 3785 -12082 3829 -12048
rect 3963 -12082 4007 -12048
rect -2173 -12388 -2139 -12132
rect -1995 -12388 -1961 -12132
rect -1817 -12388 -1783 -12132
rect -1639 -12388 -1605 -12132
rect -1461 -12388 -1427 -12132
rect -1283 -12388 -1249 -12132
rect -1105 -12388 -1071 -12132
rect -927 -12388 -893 -12132
rect -749 -12388 -715 -12132
rect -571 -12388 -537 -12132
rect -393 -12388 -359 -12132
rect -215 -12388 -181 -12132
rect -37 -12388 -3 -12132
rect 141 -12388 175 -12132
rect 319 -12388 353 -12132
rect 497 -12388 531 -12132
rect 675 -12388 709 -12132
rect 853 -12388 887 -12132
rect 1031 -12388 1065 -12132
rect 1209 -12388 1243 -12132
rect 1387 -12388 1421 -12132
rect 1565 -12388 1599 -12132
rect 1743 -12388 1777 -12132
rect 1921 -12388 1955 -12132
rect 2099 -12388 2133 -12132
rect 2277 -12388 2311 -12132
rect 2455 -12388 2489 -12132
rect 2633 -12388 2667 -12132
rect 2811 -12388 2845 -12132
rect 2989 -12388 3023 -12132
rect 3167 -12388 3201 -12132
rect 3345 -12388 3379 -12132
rect 3523 -12388 3557 -12132
rect 3701 -12388 3735 -12132
rect 3879 -12388 3913 -12132
rect 4057 -12388 4091 -12132
rect -2089 -12472 -2045 -12438
rect -1911 -12472 -1867 -12438
rect -1733 -12472 -1689 -12438
rect -1555 -12472 -1511 -12438
rect -1377 -12472 -1333 -12438
rect -1199 -12472 -1155 -12438
rect -1021 -12472 -977 -12438
rect -843 -12472 -799 -12438
rect -665 -12472 -621 -12438
rect -487 -12472 -443 -12438
rect -309 -12472 -265 -12438
rect -131 -12472 -87 -12438
rect 47 -12472 91 -12438
rect 225 -12472 269 -12438
rect 403 -12472 447 -12438
rect 581 -12472 625 -12438
rect 759 -12472 803 -12438
rect 937 -12472 981 -12438
rect 1115 -12472 1159 -12438
rect 1293 -12472 1337 -12438
rect 1471 -12472 1515 -12438
rect 1649 -12472 1693 -12438
rect 1827 -12472 1871 -12438
rect 2005 -12472 2049 -12438
rect 2183 -12472 2227 -12438
rect 2361 -12472 2405 -12438
rect 2539 -12472 2583 -12438
rect 2717 -12472 2761 -12438
rect 2895 -12472 2939 -12438
rect 3073 -12472 3117 -12438
rect 3251 -12472 3295 -12438
rect 3429 -12472 3473 -12438
rect 3607 -12472 3651 -12438
rect 3785 -12472 3829 -12438
rect 3963 -12472 4007 -12438
rect -5867 -12662 -5833 -12628
rect -5617 -12662 -5583 -12628
rect -5367 -12662 -5333 -12628
rect -5117 -12662 -5083 -12628
rect -4867 -12662 -4833 -12628
rect -4617 -12662 -4583 -12628
rect -4367 -12662 -4333 -12628
rect -4117 -12662 -4083 -12628
rect -5917 -12928 -5883 -12712
rect -5817 -12928 -5783 -12712
rect -5667 -12928 -5633 -12712
rect -5567 -12928 -5533 -12712
rect -5417 -12928 -5383 -12712
rect -5317 -12928 -5283 -12712
rect -5167 -12928 -5133 -12712
rect -5067 -12928 -5033 -12712
rect -4917 -12928 -4883 -12712
rect -4817 -12928 -4783 -12712
rect -4667 -12928 -4633 -12712
rect -4567 -12928 -4533 -12712
rect -4417 -12928 -4383 -12712
rect -4317 -12928 -4283 -12712
rect -4167 -12928 -4133 -12712
rect -4067 -12928 -4033 -12712
rect 8437 -12732 8615 -12554
rect 11437 -12732 11615 -12554
rect -5867 -13012 -5833 -12978
rect -5617 -13012 -5583 -12978
rect -5367 -13012 -5333 -12978
rect -5117 -13012 -5083 -12978
rect -4867 -13012 -4833 -12978
rect -4617 -13012 -4583 -12978
rect -4367 -13012 -4333 -12978
rect -4117 -13012 -4083 -12978
rect -2089 -13082 -2045 -13048
rect -1911 -13082 -1867 -13048
rect -1733 -13082 -1689 -13048
rect -1555 -13082 -1511 -13048
rect -1377 -13082 -1333 -13048
rect -1199 -13082 -1155 -13048
rect -1021 -13082 -977 -13048
rect -843 -13082 -799 -13048
rect -665 -13082 -621 -13048
rect -487 -13082 -443 -13048
rect -309 -13082 -265 -13048
rect -131 -13082 -87 -13048
rect 47 -13082 91 -13048
rect 225 -13082 269 -13048
rect 403 -13082 447 -13048
rect 581 -13082 625 -13048
rect 759 -13082 803 -13048
rect 937 -13082 981 -13048
rect 1115 -13082 1159 -13048
rect 1293 -13082 1337 -13048
rect 1471 -13082 1515 -13048
rect 1649 -13082 1693 -13048
rect 1827 -13082 1871 -13048
rect 2005 -13082 2049 -13048
rect 2183 -13082 2227 -13048
rect 2361 -13082 2405 -13048
rect 2539 -13082 2583 -13048
rect 2717 -13082 2761 -13048
rect 2895 -13082 2939 -13048
rect 3073 -13082 3117 -13048
rect 3251 -13082 3295 -13048
rect 3429 -13082 3473 -13048
rect 3607 -13082 3651 -13048
rect 3785 -13082 3829 -13048
rect 3963 -13082 4007 -13048
rect -5867 -13342 -5833 -13308
rect -5617 -13342 -5583 -13308
rect -5367 -13342 -5333 -13308
rect -5117 -13342 -5083 -13308
rect -4867 -13342 -4833 -13308
rect -4617 -13342 -4583 -13308
rect -4367 -13342 -4333 -13308
rect -4117 -13342 -4083 -13308
rect -5917 -13608 -5883 -13392
rect -5817 -13608 -5783 -13392
rect -5667 -13608 -5633 -13392
rect -5567 -13608 -5533 -13392
rect -5417 -13608 -5383 -13392
rect -5317 -13608 -5283 -13392
rect -5167 -13608 -5133 -13392
rect -5067 -13608 -5033 -13392
rect -4917 -13608 -4883 -13392
rect -4817 -13608 -4783 -13392
rect -4667 -13608 -4633 -13392
rect -4567 -13608 -4533 -13392
rect -4417 -13608 -4383 -13392
rect -4317 -13608 -4283 -13392
rect -4167 -13608 -4133 -13392
rect -4067 -13608 -4033 -13392
rect -2985 -13454 -2807 -13276
rect -2173 -13388 -2139 -13132
rect -1995 -13388 -1961 -13132
rect -1817 -13388 -1783 -13132
rect -1639 -13388 -1605 -13132
rect -1461 -13388 -1427 -13132
rect -1283 -13388 -1249 -13132
rect -1105 -13388 -1071 -13132
rect -927 -13388 -893 -13132
rect -749 -13388 -715 -13132
rect -571 -13388 -537 -13132
rect -393 -13388 -359 -13132
rect -215 -13388 -181 -13132
rect -37 -13388 -3 -13132
rect 141 -13388 175 -13132
rect 319 -13388 353 -13132
rect 497 -13388 531 -13132
rect 675 -13388 709 -13132
rect 853 -13388 887 -13132
rect 1031 -13388 1065 -13132
rect 1209 -13388 1243 -13132
rect 1387 -13388 1421 -13132
rect 1565 -13388 1599 -13132
rect 1743 -13388 1777 -13132
rect 1921 -13388 1955 -13132
rect 2099 -13388 2133 -13132
rect 2277 -13388 2311 -13132
rect 2455 -13388 2489 -13132
rect 2633 -13388 2667 -13132
rect 2811 -13388 2845 -13132
rect 2989 -13388 3023 -13132
rect 3167 -13388 3201 -13132
rect 3345 -13388 3379 -13132
rect 3523 -13388 3557 -13132
rect 3701 -13388 3735 -13132
rect 3879 -13388 3913 -13132
rect 4057 -13388 4091 -13132
rect -2089 -13472 -2045 -13438
rect -1911 -13472 -1867 -13438
rect -1733 -13472 -1689 -13438
rect -1555 -13472 -1511 -13438
rect -1377 -13472 -1333 -13438
rect -1199 -13472 -1155 -13438
rect -1021 -13472 -977 -13438
rect -843 -13472 -799 -13438
rect -665 -13472 -621 -13438
rect -487 -13472 -443 -13438
rect -309 -13472 -265 -13438
rect -131 -13472 -87 -13438
rect 47 -13472 91 -13438
rect 225 -13472 269 -13438
rect 403 -13472 447 -13438
rect 581 -13472 625 -13438
rect 759 -13472 803 -13438
rect 937 -13472 981 -13438
rect 1115 -13472 1159 -13438
rect 1293 -13472 1337 -13438
rect 1471 -13472 1515 -13438
rect 1649 -13472 1693 -13438
rect 1827 -13472 1871 -13438
rect 2005 -13472 2049 -13438
rect 2183 -13472 2227 -13438
rect 2361 -13472 2405 -13438
rect 2539 -13472 2583 -13438
rect 2717 -13472 2761 -13438
rect 2895 -13472 2939 -13438
rect 3073 -13472 3117 -13438
rect 3251 -13472 3295 -13438
rect 3429 -13472 3473 -13438
rect 3607 -13472 3651 -13438
rect 3785 -13472 3829 -13438
rect 3963 -13472 4007 -13438
rect -5867 -13692 -5833 -13658
rect -5617 -13692 -5583 -13658
rect -5367 -13692 -5333 -13658
rect -5117 -13692 -5083 -13658
rect -4867 -13692 -4833 -13658
rect -4617 -13692 -4583 -13658
rect -4367 -13692 -4333 -13658
rect -4117 -13692 -4083 -13658
rect -2089 -14082 -2045 -14048
rect -1911 -14082 -1867 -14048
rect -1733 -14082 -1689 -14048
rect -1555 -14082 -1511 -14048
rect -1377 -14082 -1333 -14048
rect -1199 -14082 -1155 -14048
rect -1021 -14082 -977 -14048
rect -843 -14082 -799 -14048
rect -665 -14082 -621 -14048
rect -487 -14082 -443 -14048
rect -309 -14082 -265 -14048
rect -131 -14082 -87 -14048
rect 47 -14082 91 -14048
rect 225 -14082 269 -14048
rect 403 -14082 447 -14048
rect 581 -14082 625 -14048
rect 759 -14082 803 -14048
rect 937 -14082 981 -14048
rect 1115 -14082 1159 -14048
rect 1293 -14082 1337 -14048
rect 1471 -14082 1515 -14048
rect 1649 -14082 1693 -14048
rect 1827 -14082 1871 -14048
rect 2005 -14082 2049 -14048
rect 2183 -14082 2227 -14048
rect 2361 -14082 2405 -14048
rect 2539 -14082 2583 -14048
rect 2717 -14082 2761 -14048
rect 2895 -14082 2939 -14048
rect 3073 -14082 3117 -14048
rect 3251 -14082 3295 -14048
rect 3429 -14082 3473 -14048
rect 3607 -14082 3651 -14048
rect 3785 -14082 3829 -14048
rect 3963 -14082 4007 -14048
rect 5661 -14082 5705 -14048
rect 5839 -14082 5883 -14048
rect 6017 -14082 6061 -14048
rect 6195 -14082 6239 -14048
rect 6373 -14082 6417 -14048
rect 6551 -14082 6595 -14048
rect 6729 -14082 6773 -14048
rect 6907 -14082 6951 -14048
rect 7085 -14082 7129 -14048
rect 7263 -14082 7307 -14048
rect 7441 -14082 7485 -14048
rect 7619 -14082 7663 -14048
rect 7797 -14082 7841 -14048
rect 7975 -14082 8019 -14048
rect 8153 -14082 8197 -14048
rect 8331 -14082 8375 -14048
rect 8509 -14082 8553 -14048
rect 8687 -14082 8731 -14048
rect 8865 -14082 8909 -14048
rect 9043 -14082 9087 -14048
rect 9221 -14082 9265 -14048
rect 9399 -14082 9443 -14048
rect 9577 -14082 9621 -14048
rect 9755 -14082 9799 -14048
rect 9933 -14082 9977 -14048
rect 10111 -14082 10155 -14048
rect 10289 -14082 10333 -14048
rect 10467 -14082 10511 -14048
rect 10645 -14082 10689 -14048
rect 10823 -14082 10867 -14048
rect 11001 -14082 11045 -14048
rect 11179 -14082 11223 -14048
rect 11357 -14082 11401 -14048
rect 11535 -14082 11579 -14048
rect 11713 -14082 11757 -14048
rect 11891 -14082 11935 -14048
rect 12069 -14082 12113 -14048
rect 12247 -14082 12291 -14048
rect 12425 -14082 12469 -14048
rect 12603 -14082 12647 -14048
rect -5944 -14344 -5900 -14310
rect -5766 -14344 -5722 -14310
rect -5588 -14344 -5544 -14310
rect -5410 -14344 -5366 -14310
rect -5232 -14344 -5188 -14310
rect -5054 -14344 -5010 -14310
rect -4876 -14344 -4832 -14310
rect -4698 -14344 -4654 -14310
rect -4520 -14344 -4476 -14310
rect -4342 -14344 -4298 -14310
rect -4164 -14344 -4120 -14310
rect -6028 -14650 -5994 -14394
rect -5850 -14650 -5816 -14394
rect -5672 -14650 -5638 -14394
rect -5494 -14650 -5460 -14394
rect -5316 -14650 -5282 -14394
rect -5138 -14650 -5104 -14394
rect -4960 -14650 -4926 -14394
rect -4782 -14650 -4748 -14394
rect -4604 -14650 -4570 -14394
rect -4426 -14650 -4392 -14394
rect -4248 -14650 -4214 -14394
rect -4070 -14650 -4036 -14394
rect -2173 -14388 -2139 -14132
rect -1995 -14388 -1961 -14132
rect -1817 -14388 -1783 -14132
rect -1639 -14388 -1605 -14132
rect -1461 -14388 -1427 -14132
rect -1283 -14388 -1249 -14132
rect -1105 -14388 -1071 -14132
rect -927 -14388 -893 -14132
rect -749 -14388 -715 -14132
rect -571 -14388 -537 -14132
rect -393 -14388 -359 -14132
rect -215 -14388 -181 -14132
rect -37 -14388 -3 -14132
rect 141 -14388 175 -14132
rect 319 -14388 353 -14132
rect 497 -14388 531 -14132
rect 675 -14388 709 -14132
rect 853 -14388 887 -14132
rect 1031 -14388 1065 -14132
rect 1209 -14388 1243 -14132
rect 1387 -14388 1421 -14132
rect 1565 -14388 1599 -14132
rect 1743 -14388 1777 -14132
rect 1921 -14388 1955 -14132
rect 2099 -14388 2133 -14132
rect 2277 -14388 2311 -14132
rect 2455 -14388 2489 -14132
rect 2633 -14388 2667 -14132
rect 2811 -14388 2845 -14132
rect 2989 -14388 3023 -14132
rect 3167 -14388 3201 -14132
rect 3345 -14388 3379 -14132
rect 3523 -14388 3557 -14132
rect 3701 -14388 3735 -14132
rect 3879 -14388 3913 -14132
rect 4057 -14388 4091 -14132
rect 5577 -14388 5611 -14132
rect 5755 -14388 5789 -14132
rect 5933 -14388 5967 -14132
rect 6111 -14388 6145 -14132
rect 6289 -14388 6323 -14132
rect 6467 -14388 6501 -14132
rect 6645 -14388 6679 -14132
rect 6823 -14388 6857 -14132
rect 7001 -14388 7035 -14132
rect 7179 -14388 7213 -14132
rect 7357 -14388 7391 -14132
rect 7535 -14388 7569 -14132
rect 7713 -14388 7747 -14132
rect 7891 -14388 7925 -14132
rect 8069 -14388 8103 -14132
rect 8247 -14388 8281 -14132
rect 8425 -14388 8459 -14132
rect 8603 -14388 8637 -14132
rect 8781 -14388 8815 -14132
rect 8959 -14388 8993 -14132
rect 9137 -14388 9171 -14132
rect 9315 -14388 9349 -14132
rect 9493 -14388 9527 -14132
rect 9671 -14388 9705 -14132
rect 9849 -14388 9883 -14132
rect 10027 -14388 10061 -14132
rect 10205 -14388 10239 -14132
rect 10383 -14388 10417 -14132
rect 10561 -14388 10595 -14132
rect 10739 -14388 10773 -14132
rect 10917 -14388 10951 -14132
rect 11095 -14388 11129 -14132
rect 11273 -14388 11307 -14132
rect 11451 -14388 11485 -14132
rect 11629 -14388 11663 -14132
rect 11807 -14388 11841 -14132
rect 11985 -14388 12019 -14132
rect 12163 -14388 12197 -14132
rect 12341 -14388 12375 -14132
rect 12519 -14388 12553 -14132
rect 12697 -14388 12731 -14132
rect -2089 -14472 -2045 -14438
rect -1911 -14472 -1867 -14438
rect -1733 -14472 -1689 -14438
rect -1555 -14472 -1511 -14438
rect -1377 -14472 -1333 -14438
rect -1199 -14472 -1155 -14438
rect -1021 -14472 -977 -14438
rect -843 -14472 -799 -14438
rect -665 -14472 -621 -14438
rect -487 -14472 -443 -14438
rect -309 -14472 -265 -14438
rect -131 -14472 -87 -14438
rect 47 -14472 91 -14438
rect 225 -14472 269 -14438
rect 403 -14472 447 -14438
rect 581 -14472 625 -14438
rect 759 -14472 803 -14438
rect 937 -14472 981 -14438
rect 1115 -14472 1159 -14438
rect 1293 -14472 1337 -14438
rect 1471 -14472 1515 -14438
rect 1649 -14472 1693 -14438
rect 1827 -14472 1871 -14438
rect 2005 -14472 2049 -14438
rect 2183 -14472 2227 -14438
rect 2361 -14472 2405 -14438
rect 2539 -14472 2583 -14438
rect 2717 -14472 2761 -14438
rect 2895 -14472 2939 -14438
rect 3073 -14472 3117 -14438
rect 3251 -14472 3295 -14438
rect 3429 -14472 3473 -14438
rect 3607 -14472 3651 -14438
rect 3785 -14472 3829 -14438
rect 3963 -14472 4007 -14438
rect 5661 -14472 5705 -14438
rect 5839 -14472 5883 -14438
rect 6017 -14472 6061 -14438
rect 6195 -14472 6239 -14438
rect 6373 -14472 6417 -14438
rect 6551 -14472 6595 -14438
rect 6729 -14472 6773 -14438
rect 6907 -14472 6951 -14438
rect 7085 -14472 7129 -14438
rect 7263 -14472 7307 -14438
rect 7441 -14472 7485 -14438
rect 7619 -14472 7663 -14438
rect 7797 -14472 7841 -14438
rect 7975 -14472 8019 -14438
rect 8153 -14472 8197 -14438
rect 8331 -14472 8375 -14438
rect 8509 -14472 8553 -14438
rect 8687 -14472 8731 -14438
rect 8865 -14472 8909 -14438
rect 9043 -14472 9087 -14438
rect 9221 -14472 9265 -14438
rect 9399 -14472 9443 -14438
rect 9577 -14472 9621 -14438
rect 9755 -14472 9799 -14438
rect 9933 -14472 9977 -14438
rect 10111 -14472 10155 -14438
rect 10289 -14472 10333 -14438
rect 10467 -14472 10511 -14438
rect 10645 -14472 10689 -14438
rect 10823 -14472 10867 -14438
rect 11001 -14472 11045 -14438
rect 11179 -14472 11223 -14438
rect 11357 -14472 11401 -14438
rect 11535 -14472 11579 -14438
rect 11713 -14472 11757 -14438
rect 11891 -14472 11935 -14438
rect 12069 -14472 12113 -14438
rect 12247 -14472 12291 -14438
rect 12425 -14472 12469 -14438
rect 12603 -14472 12647 -14438
rect -5944 -14734 -5900 -14700
rect -5766 -14734 -5722 -14700
rect -5588 -14734 -5544 -14700
rect -5410 -14734 -5366 -14700
rect -5232 -14734 -5188 -14700
rect -5054 -14734 -5010 -14700
rect -4876 -14734 -4832 -14700
rect -4698 -14734 -4654 -14700
rect -4520 -14734 -4476 -14700
rect -4342 -14734 -4298 -14700
rect -4164 -14734 -4120 -14700
rect -5944 -15044 -5900 -15010
rect -5766 -15044 -5722 -15010
rect -5588 -15044 -5544 -15010
rect -5410 -15044 -5366 -15010
rect -5232 -15044 -5188 -15010
rect -5054 -15044 -5010 -15010
rect -4876 -15044 -4832 -15010
rect -4698 -15044 -4654 -15010
rect -4520 -15044 -4476 -15010
rect -4342 -15044 -4298 -15010
rect -4164 -15044 -4120 -15010
rect 4543 -15047 4721 -14869
rect -6028 -15350 -5994 -15094
rect -5850 -15350 -5816 -15094
rect -5672 -15350 -5638 -15094
rect -5494 -15350 -5460 -15094
rect -5316 -15350 -5282 -15094
rect -5138 -15350 -5104 -15094
rect -4960 -15350 -4926 -15094
rect -4782 -15350 -4748 -15094
rect -4604 -15350 -4570 -15094
rect -4426 -15350 -4392 -15094
rect -4248 -15350 -4214 -15094
rect -2089 -15082 -2045 -15048
rect -1911 -15082 -1867 -15048
rect -1733 -15082 -1689 -15048
rect -1555 -15082 -1511 -15048
rect -1377 -15082 -1333 -15048
rect -1199 -15082 -1155 -15048
rect -1021 -15082 -977 -15048
rect -843 -15082 -799 -15048
rect -665 -15082 -621 -15048
rect -487 -15082 -443 -15048
rect -309 -15082 -265 -15048
rect -131 -15082 -87 -15048
rect 47 -15082 91 -15048
rect 225 -15082 269 -15048
rect 403 -15082 447 -15048
rect 581 -15082 625 -15048
rect 759 -15082 803 -15048
rect 937 -15082 981 -15048
rect 1115 -15082 1159 -15048
rect 1293 -15082 1337 -15048
rect 1471 -15082 1515 -15048
rect 1649 -15082 1693 -15048
rect 1827 -15082 1871 -15048
rect 2005 -15082 2049 -15048
rect 2183 -15082 2227 -15048
rect 2361 -15082 2405 -15048
rect 2539 -15082 2583 -15048
rect 2717 -15082 2761 -15048
rect 2895 -15082 2939 -15048
rect 3073 -15082 3117 -15048
rect 3251 -15082 3295 -15048
rect 3429 -15082 3473 -15048
rect 3607 -15082 3651 -15048
rect 3785 -15082 3829 -15048
rect 3963 -15082 4007 -15048
rect 5661 -15082 5705 -15048
rect 5839 -15082 5883 -15048
rect 6017 -15082 6061 -15048
rect 6195 -15082 6239 -15048
rect 6373 -15082 6417 -15048
rect 6551 -15082 6595 -15048
rect 6729 -15082 6773 -15048
rect 6907 -15082 6951 -15048
rect 7085 -15082 7129 -15048
rect 7263 -15082 7307 -15048
rect 7441 -15082 7485 -15048
rect 7619 -15082 7663 -15048
rect 7797 -15082 7841 -15048
rect 7975 -15082 8019 -15048
rect 8153 -15082 8197 -15048
rect 8331 -15082 8375 -15048
rect 8509 -15082 8553 -15048
rect 8687 -15082 8731 -15048
rect 8865 -15082 8909 -15048
rect 9043 -15082 9087 -15048
rect 9221 -15082 9265 -15048
rect 9399 -15082 9443 -15048
rect 9577 -15082 9621 -15048
rect 9755 -15082 9799 -15048
rect 9933 -15082 9977 -15048
rect 10111 -15082 10155 -15048
rect 10289 -15082 10333 -15048
rect 10467 -15082 10511 -15048
rect 10645 -15082 10689 -15048
rect 10823 -15082 10867 -15048
rect 11001 -15082 11045 -15048
rect 11179 -15082 11223 -15048
rect 11357 -15082 11401 -15048
rect 11535 -15082 11579 -15048
rect 11713 -15082 11757 -15048
rect 11891 -15082 11935 -15048
rect 12069 -15082 12113 -15048
rect 12247 -15082 12291 -15048
rect 12425 -15082 12469 -15048
rect 12603 -15082 12647 -15048
rect -4070 -15350 -4036 -15094
rect -5944 -15434 -5900 -15400
rect -5766 -15434 -5722 -15400
rect -5588 -15434 -5544 -15400
rect -5410 -15434 -5366 -15400
rect -5232 -15434 -5188 -15400
rect -5054 -15434 -5010 -15400
rect -4876 -15434 -4832 -15400
rect -4698 -15434 -4654 -15400
rect -4520 -15434 -4476 -15400
rect -4342 -15434 -4298 -15400
rect -4164 -15434 -4120 -15400
rect -2985 -15454 -2807 -15276
rect -2173 -15388 -2139 -15132
rect -1995 -15388 -1961 -15132
rect -1817 -15388 -1783 -15132
rect -1639 -15388 -1605 -15132
rect -1461 -15388 -1427 -15132
rect -1283 -15388 -1249 -15132
rect -1105 -15388 -1071 -15132
rect -927 -15388 -893 -15132
rect -749 -15388 -715 -15132
rect -571 -15388 -537 -15132
rect -393 -15388 -359 -15132
rect -215 -15388 -181 -15132
rect -37 -15388 -3 -15132
rect 141 -15388 175 -15132
rect 319 -15388 353 -15132
rect 497 -15388 531 -15132
rect 675 -15388 709 -15132
rect 853 -15388 887 -15132
rect 1031 -15388 1065 -15132
rect 1209 -15388 1243 -15132
rect 1387 -15388 1421 -15132
rect 1565 -15388 1599 -15132
rect 1743 -15388 1777 -15132
rect 1921 -15388 1955 -15132
rect 2099 -15388 2133 -15132
rect 2277 -15388 2311 -15132
rect 2455 -15388 2489 -15132
rect 2633 -15388 2667 -15132
rect 2811 -15388 2845 -15132
rect 2989 -15388 3023 -15132
rect 3167 -15388 3201 -15132
rect 3345 -15388 3379 -15132
rect 3523 -15388 3557 -15132
rect 3701 -15388 3735 -15132
rect 3879 -15388 3913 -15132
rect 4057 -15388 4091 -15132
rect 5577 -15388 5611 -15132
rect 5755 -15388 5789 -15132
rect 5933 -15388 5967 -15132
rect 6111 -15388 6145 -15132
rect 6289 -15388 6323 -15132
rect 6467 -15388 6501 -15132
rect 6645 -15388 6679 -15132
rect 6823 -15388 6857 -15132
rect 7001 -15388 7035 -15132
rect 7179 -15388 7213 -15132
rect 7357 -15388 7391 -15132
rect 7535 -15388 7569 -15132
rect 7713 -15388 7747 -15132
rect 7891 -15388 7925 -15132
rect 8069 -15388 8103 -15132
rect 8247 -15388 8281 -15132
rect 8425 -15388 8459 -15132
rect 8603 -15388 8637 -15132
rect 8781 -15388 8815 -15132
rect 8959 -15388 8993 -15132
rect 9137 -15388 9171 -15132
rect 9315 -15388 9349 -15132
rect 9493 -15388 9527 -15132
rect 9671 -15388 9705 -15132
rect 9849 -15388 9883 -15132
rect 10027 -15388 10061 -15132
rect 10205 -15388 10239 -15132
rect 10383 -15388 10417 -15132
rect 10561 -15388 10595 -15132
rect 10739 -15388 10773 -15132
rect 10917 -15388 10951 -15132
rect 11095 -15388 11129 -15132
rect 11273 -15388 11307 -15132
rect 11451 -15388 11485 -15132
rect 11629 -15388 11663 -15132
rect 11807 -15388 11841 -15132
rect 11985 -15388 12019 -15132
rect 12163 -15388 12197 -15132
rect 12341 -15388 12375 -15132
rect 12519 -15388 12553 -15132
rect 12697 -15388 12731 -15132
rect -2089 -15472 -2045 -15438
rect -1911 -15472 -1867 -15438
rect -1733 -15472 -1689 -15438
rect -1555 -15472 -1511 -15438
rect -1377 -15472 -1333 -15438
rect -1199 -15472 -1155 -15438
rect -1021 -15472 -977 -15438
rect -843 -15472 -799 -15438
rect -665 -15472 -621 -15438
rect -487 -15472 -443 -15438
rect -309 -15472 -265 -15438
rect -131 -15472 -87 -15438
rect 47 -15472 91 -15438
rect 225 -15472 269 -15438
rect 403 -15472 447 -15438
rect 581 -15472 625 -15438
rect 759 -15472 803 -15438
rect 937 -15472 981 -15438
rect 1115 -15472 1159 -15438
rect 1293 -15472 1337 -15438
rect 1471 -15472 1515 -15438
rect 1649 -15472 1693 -15438
rect 1827 -15472 1871 -15438
rect 2005 -15472 2049 -15438
rect 2183 -15472 2227 -15438
rect 2361 -15472 2405 -15438
rect 2539 -15472 2583 -15438
rect 2717 -15472 2761 -15438
rect 2895 -15472 2939 -15438
rect 3073 -15472 3117 -15438
rect 3251 -15472 3295 -15438
rect 3429 -15472 3473 -15438
rect 3607 -15472 3651 -15438
rect 3785 -15472 3829 -15438
rect 3963 -15472 4007 -15438
rect 5661 -15472 5705 -15438
rect 5839 -15472 5883 -15438
rect 6017 -15472 6061 -15438
rect 6195 -15472 6239 -15438
rect 6373 -15472 6417 -15438
rect 6551 -15472 6595 -15438
rect 6729 -15472 6773 -15438
rect 6907 -15472 6951 -15438
rect 7085 -15472 7129 -15438
rect 7263 -15472 7307 -15438
rect 7441 -15472 7485 -15438
rect 7619 -15472 7663 -15438
rect 7797 -15472 7841 -15438
rect 7975 -15472 8019 -15438
rect 8153 -15472 8197 -15438
rect 8331 -15472 8375 -15438
rect 8509 -15472 8553 -15438
rect 8687 -15472 8731 -15438
rect 8865 -15472 8909 -15438
rect 9043 -15472 9087 -15438
rect 9221 -15472 9265 -15438
rect 9399 -15472 9443 -15438
rect 9577 -15472 9621 -15438
rect 9755 -15472 9799 -15438
rect 9933 -15472 9977 -15438
rect 10111 -15472 10155 -15438
rect 10289 -15472 10333 -15438
rect 10467 -15472 10511 -15438
rect 10645 -15472 10689 -15438
rect 10823 -15472 10867 -15438
rect 11001 -15472 11045 -15438
rect 11179 -15472 11223 -15438
rect 11357 -15472 11401 -15438
rect 11535 -15472 11579 -15438
rect 11713 -15472 11757 -15438
rect 11891 -15472 11935 -15438
rect 12069 -15472 12113 -15438
rect 12247 -15472 12291 -15438
rect 12425 -15472 12469 -15438
rect 12603 -15472 12647 -15438
rect -5944 -15744 -5900 -15710
rect -5766 -15744 -5722 -15710
rect -5588 -15744 -5544 -15710
rect -5410 -15744 -5366 -15710
rect -5232 -15744 -5188 -15710
rect -5054 -15744 -5010 -15710
rect -4876 -15744 -4832 -15710
rect -4698 -15744 -4654 -15710
rect -4520 -15744 -4476 -15710
rect -4342 -15744 -4298 -15710
rect -4164 -15744 -4120 -15710
rect -6028 -16050 -5994 -15794
rect -5850 -16050 -5816 -15794
rect -5672 -16050 -5638 -15794
rect -5494 -16050 -5460 -15794
rect -5316 -16050 -5282 -15794
rect -5138 -16050 -5104 -15794
rect -4960 -16050 -4926 -15794
rect -4782 -16050 -4748 -15794
rect -4604 -16050 -4570 -15794
rect -4426 -16050 -4392 -15794
rect -4248 -16050 -4214 -15794
rect -4070 -16050 -4036 -15794
rect -2089 -16082 -2045 -16048
rect -1911 -16082 -1867 -16048
rect -1733 -16082 -1689 -16048
rect -1555 -16082 -1511 -16048
rect -1377 -16082 -1333 -16048
rect -1199 -16082 -1155 -16048
rect -1021 -16082 -977 -16048
rect -843 -16082 -799 -16048
rect -665 -16082 -621 -16048
rect -487 -16082 -443 -16048
rect -309 -16082 -265 -16048
rect -131 -16082 -87 -16048
rect 47 -16082 91 -16048
rect 225 -16082 269 -16048
rect 403 -16082 447 -16048
rect 581 -16082 625 -16048
rect 759 -16082 803 -16048
rect 937 -16082 981 -16048
rect 1115 -16082 1159 -16048
rect 1293 -16082 1337 -16048
rect 1471 -16082 1515 -16048
rect 1649 -16082 1693 -16048
rect 1827 -16082 1871 -16048
rect 2005 -16082 2049 -16048
rect 2183 -16082 2227 -16048
rect 2361 -16082 2405 -16048
rect 2539 -16082 2583 -16048
rect 2717 -16082 2761 -16048
rect 2895 -16082 2939 -16048
rect 3073 -16082 3117 -16048
rect 3251 -16082 3295 -16048
rect 3429 -16082 3473 -16048
rect 3607 -16082 3651 -16048
rect 3785 -16082 3829 -16048
rect 3963 -16082 4007 -16048
rect 5661 -16082 5705 -16048
rect 5839 -16082 5883 -16048
rect 6017 -16082 6061 -16048
rect 6195 -16082 6239 -16048
rect 6373 -16082 6417 -16048
rect 6551 -16082 6595 -16048
rect 6729 -16082 6773 -16048
rect 6907 -16082 6951 -16048
rect 7085 -16082 7129 -16048
rect 7263 -16082 7307 -16048
rect 7441 -16082 7485 -16048
rect 7619 -16082 7663 -16048
rect 7797 -16082 7841 -16048
rect 7975 -16082 8019 -16048
rect 8153 -16082 8197 -16048
rect 8331 -16082 8375 -16048
rect 8509 -16082 8553 -16048
rect 8687 -16082 8731 -16048
rect 8865 -16082 8909 -16048
rect 9043 -16082 9087 -16048
rect 9221 -16082 9265 -16048
rect 9399 -16082 9443 -16048
rect 9577 -16082 9621 -16048
rect 9755 -16082 9799 -16048
rect 9933 -16082 9977 -16048
rect 10111 -16082 10155 -16048
rect 10289 -16082 10333 -16048
rect 10467 -16082 10511 -16048
rect 10645 -16082 10689 -16048
rect 10823 -16082 10867 -16048
rect 11001 -16082 11045 -16048
rect 11179 -16082 11223 -16048
rect 11357 -16082 11401 -16048
rect 11535 -16082 11579 -16048
rect 11713 -16082 11757 -16048
rect 11891 -16082 11935 -16048
rect 12069 -16082 12113 -16048
rect 12247 -16082 12291 -16048
rect 12425 -16082 12469 -16048
rect 12603 -16082 12647 -16048
rect -5944 -16134 -5900 -16100
rect -5766 -16134 -5722 -16100
rect -5588 -16134 -5544 -16100
rect -5410 -16134 -5366 -16100
rect -5232 -16134 -5188 -16100
rect -5054 -16134 -5010 -16100
rect -4876 -16134 -4832 -16100
rect -4698 -16134 -4654 -16100
rect -4520 -16134 -4476 -16100
rect -4342 -16134 -4298 -16100
rect -4164 -16134 -4120 -16100
rect -2173 -16388 -2139 -16132
rect -1995 -16388 -1961 -16132
rect -1817 -16388 -1783 -16132
rect -1639 -16388 -1605 -16132
rect -1461 -16388 -1427 -16132
rect -1283 -16388 -1249 -16132
rect -1105 -16388 -1071 -16132
rect -927 -16388 -893 -16132
rect -749 -16388 -715 -16132
rect -571 -16388 -537 -16132
rect -393 -16388 -359 -16132
rect -215 -16388 -181 -16132
rect -37 -16388 -3 -16132
rect 141 -16388 175 -16132
rect 319 -16388 353 -16132
rect 497 -16388 531 -16132
rect 675 -16388 709 -16132
rect 853 -16388 887 -16132
rect 1031 -16388 1065 -16132
rect 1209 -16388 1243 -16132
rect 1387 -16388 1421 -16132
rect 1565 -16388 1599 -16132
rect 1743 -16388 1777 -16132
rect 1921 -16388 1955 -16132
rect 2099 -16388 2133 -16132
rect 2277 -16388 2311 -16132
rect 2455 -16388 2489 -16132
rect 2633 -16388 2667 -16132
rect 2811 -16388 2845 -16132
rect 2989 -16388 3023 -16132
rect 3167 -16388 3201 -16132
rect 3345 -16388 3379 -16132
rect 3523 -16388 3557 -16132
rect 3701 -16388 3735 -16132
rect 3879 -16388 3913 -16132
rect 4057 -16388 4091 -16132
rect 5577 -16388 5611 -16132
rect 5755 -16388 5789 -16132
rect 5933 -16388 5967 -16132
rect 6111 -16388 6145 -16132
rect 6289 -16388 6323 -16132
rect 6467 -16388 6501 -16132
rect 6645 -16388 6679 -16132
rect 6823 -16388 6857 -16132
rect 7001 -16388 7035 -16132
rect 7179 -16388 7213 -16132
rect 7357 -16388 7391 -16132
rect 7535 -16388 7569 -16132
rect 7713 -16388 7747 -16132
rect 7891 -16388 7925 -16132
rect 8069 -16388 8103 -16132
rect 8247 -16388 8281 -16132
rect 8425 -16388 8459 -16132
rect 8603 -16388 8637 -16132
rect 8781 -16388 8815 -16132
rect 8959 -16388 8993 -16132
rect 9137 -16388 9171 -16132
rect 9315 -16388 9349 -16132
rect 9493 -16388 9527 -16132
rect 9671 -16388 9705 -16132
rect 9849 -16388 9883 -16132
rect 10027 -16388 10061 -16132
rect 10205 -16388 10239 -16132
rect 10383 -16388 10417 -16132
rect 10561 -16388 10595 -16132
rect 10739 -16388 10773 -16132
rect 10917 -16388 10951 -16132
rect 11095 -16388 11129 -16132
rect 11273 -16388 11307 -16132
rect 11451 -16388 11485 -16132
rect 11629 -16388 11663 -16132
rect 11807 -16388 11841 -16132
rect 11985 -16388 12019 -16132
rect 12163 -16388 12197 -16132
rect 12341 -16388 12375 -16132
rect 12519 -16388 12553 -16132
rect 12697 -16388 12731 -16132
rect -5944 -16444 -5900 -16410
rect -5766 -16444 -5722 -16410
rect -5588 -16444 -5544 -16410
rect -5410 -16444 -5366 -16410
rect -5232 -16444 -5188 -16410
rect -5054 -16444 -5010 -16410
rect -4876 -16444 -4832 -16410
rect -4698 -16444 -4654 -16410
rect -4520 -16444 -4476 -16410
rect -4342 -16444 -4298 -16410
rect -4164 -16444 -4120 -16410
rect -2089 -16472 -2045 -16438
rect -1911 -16472 -1867 -16438
rect -1733 -16472 -1689 -16438
rect -1555 -16472 -1511 -16438
rect -1377 -16472 -1333 -16438
rect -1199 -16472 -1155 -16438
rect -1021 -16472 -977 -16438
rect -843 -16472 -799 -16438
rect -665 -16472 -621 -16438
rect -487 -16472 -443 -16438
rect -309 -16472 -265 -16438
rect -131 -16472 -87 -16438
rect 47 -16472 91 -16438
rect 225 -16472 269 -16438
rect 403 -16472 447 -16438
rect 581 -16472 625 -16438
rect 759 -16472 803 -16438
rect 937 -16472 981 -16438
rect 1115 -16472 1159 -16438
rect 1293 -16472 1337 -16438
rect 1471 -16472 1515 -16438
rect 1649 -16472 1693 -16438
rect 1827 -16472 1871 -16438
rect 2005 -16472 2049 -16438
rect 2183 -16472 2227 -16438
rect 2361 -16472 2405 -16438
rect 2539 -16472 2583 -16438
rect 2717 -16472 2761 -16438
rect 2895 -16472 2939 -16438
rect 3073 -16472 3117 -16438
rect 3251 -16472 3295 -16438
rect 3429 -16472 3473 -16438
rect 3607 -16472 3651 -16438
rect 3785 -16472 3829 -16438
rect 3963 -16472 4007 -16438
rect 5661 -16472 5705 -16438
rect 5839 -16472 5883 -16438
rect 6017 -16472 6061 -16438
rect 6195 -16472 6239 -16438
rect 6373 -16472 6417 -16438
rect 6551 -16472 6595 -16438
rect 6729 -16472 6773 -16438
rect 6907 -16472 6951 -16438
rect 7085 -16472 7129 -16438
rect 7263 -16472 7307 -16438
rect 7441 -16472 7485 -16438
rect 7619 -16472 7663 -16438
rect 7797 -16472 7841 -16438
rect 7975 -16472 8019 -16438
rect 8153 -16472 8197 -16438
rect 8331 -16472 8375 -16438
rect 8509 -16472 8553 -16438
rect 8687 -16472 8731 -16438
rect 8865 -16472 8909 -16438
rect 9043 -16472 9087 -16438
rect 9221 -16472 9265 -16438
rect 9399 -16472 9443 -16438
rect 9577 -16472 9621 -16438
rect 9755 -16472 9799 -16438
rect 9933 -16472 9977 -16438
rect 10111 -16472 10155 -16438
rect 10289 -16472 10333 -16438
rect 10467 -16472 10511 -16438
rect 10645 -16472 10689 -16438
rect 10823 -16472 10867 -16438
rect 11001 -16472 11045 -16438
rect 11179 -16472 11223 -16438
rect 11357 -16472 11401 -16438
rect 11535 -16472 11579 -16438
rect 11713 -16472 11757 -16438
rect 11891 -16472 11935 -16438
rect 12069 -16472 12113 -16438
rect 12247 -16472 12291 -16438
rect 12425 -16472 12469 -16438
rect 12603 -16472 12647 -16438
rect -6028 -16750 -5994 -16494
rect -5850 -16750 -5816 -16494
rect -5672 -16750 -5638 -16494
rect -5494 -16750 -5460 -16494
rect -5316 -16750 -5282 -16494
rect -5138 -16750 -5104 -16494
rect -4960 -16750 -4926 -16494
rect -4782 -16750 -4748 -16494
rect -4604 -16750 -4570 -16494
rect -4426 -16750 -4392 -16494
rect -4248 -16750 -4214 -16494
rect -4070 -16750 -4036 -16494
rect -5944 -16834 -5900 -16800
rect -5766 -16834 -5722 -16800
rect -5588 -16834 -5544 -16800
rect -5410 -16834 -5366 -16800
rect -5232 -16834 -5188 -16800
rect -5054 -16834 -5010 -16800
rect -4876 -16834 -4832 -16800
rect -4698 -16834 -4654 -16800
rect -4520 -16834 -4476 -16800
rect -4342 -16834 -4298 -16800
rect -4164 -16834 -4120 -16800
rect -7323 -17559 13384 -17459
<< metal1 >>
rect 7034 2713 7080 2891
rect 7250 2775 8332 2809
rect 7034 2327 7040 2713
rect 7074 2327 7080 2713
rect 7135 2665 7145 2717
rect 7197 2665 7207 2717
rect 7250 2625 7284 2775
rect 7327 2665 7337 2717
rect 7389 2665 7399 2717
rect 7442 2625 7476 2775
rect 7519 2665 7529 2717
rect 7581 2665 7591 2717
rect 7634 2625 7668 2775
rect 7711 2665 7721 2717
rect 7773 2665 7783 2717
rect 7826 2625 7860 2775
rect 7902 2665 7912 2717
rect 7964 2665 7974 2717
rect 8018 2625 8052 2775
rect 8095 2665 8105 2717
rect 8157 2665 8167 2717
rect 7148 2613 7194 2625
rect 7148 2365 7154 2613
rect 7188 2365 7194 2613
rect 7148 2353 7194 2365
rect 7244 2613 7290 2625
rect 7244 2365 7250 2613
rect 7284 2365 7290 2613
rect 7244 2353 7290 2365
rect 7340 2613 7386 2625
rect 7340 2365 7346 2613
rect 7380 2365 7386 2613
rect 7340 2353 7386 2365
rect 7436 2613 7482 2625
rect 7436 2365 7442 2613
rect 7476 2365 7482 2613
rect 7436 2353 7482 2365
rect 7532 2613 7578 2625
rect 7532 2365 7538 2613
rect 7572 2365 7578 2613
rect 7532 2353 7578 2365
rect 7628 2613 7674 2625
rect 7628 2365 7634 2613
rect 7668 2365 7674 2613
rect 7628 2353 7674 2365
rect 7724 2613 7770 2625
rect 7724 2365 7730 2613
rect 7764 2365 7770 2613
rect 7724 2353 7770 2365
rect 7820 2613 7866 2625
rect 7820 2365 7826 2613
rect 7860 2365 7866 2613
rect 7820 2353 7866 2365
rect 7916 2613 7962 2625
rect 7916 2365 7922 2613
rect 7956 2365 7962 2613
rect 7916 2353 7962 2365
rect 8012 2613 8058 2625
rect 8012 2365 8018 2613
rect 8052 2365 8058 2613
rect 8012 2353 8058 2365
rect 8108 2613 8154 2625
rect 8108 2365 8114 2613
rect 8148 2365 8154 2613
rect 8108 2353 8154 2365
rect 7034 2315 7080 2327
rect 7154 2212 7188 2353
rect 7346 2212 7380 2353
rect 7538 2212 7572 2353
rect 7730 2212 7764 2353
rect 7922 2212 7956 2353
rect 8114 2226 8148 2353
rect 8070 2212 8080 2226
rect 5608 2178 8080 2212
rect -7605 -1260 3704 -1200
rect -7605 -1353 -7379 -1260
rect 3329 -1353 3704 -1260
rect -7605 -1467 3704 -1353
rect -5059 -1807 -5025 -1467
rect -5945 -1808 -3809 -1807
rect -5945 -1841 -3776 -1808
rect -6234 -2039 -6158 -2023
rect -6056 -2039 -5980 -2023
rect -5945 -2039 -5911 -1841
rect -5877 -1963 -5867 -1910
rect -5814 -1963 -5804 -1910
rect -5699 -1963 -5689 -1910
rect -5636 -1963 -5626 -1910
rect -5520 -1963 -5510 -1910
rect -5457 -1963 -5447 -1910
rect -5343 -1963 -5333 -1910
rect -5280 -1963 -5270 -1910
rect -5165 -1963 -5155 -1910
rect -5102 -1963 -5092 -1910
rect -4986 -1963 -4976 -1910
rect -4923 -1963 -4913 -1910
rect -4809 -1963 -4799 -1910
rect -4746 -1963 -4736 -1910
rect -4631 -1963 -4621 -1910
rect -4568 -1963 -4558 -1910
rect -4453 -1963 -4443 -1910
rect -4390 -1963 -4380 -1910
rect -4275 -1963 -4265 -1910
rect -4212 -1963 -4202 -1910
rect -4096 -1963 -4086 -1910
rect -4033 -1963 -4023 -1910
rect -3919 -1963 -3909 -1910
rect -3856 -1963 -3846 -1910
rect -5857 -2023 -5823 -1963
rect -5679 -2023 -5645 -1963
rect -5501 -2023 -5467 -1963
rect -5322 -2023 -5288 -1963
rect -5145 -2023 -5111 -1963
rect -4967 -2023 -4933 -1963
rect -4789 -2023 -4755 -1963
rect -4611 -2023 -4577 -1963
rect -4433 -2023 -4399 -1963
rect -4255 -2023 -4221 -1963
rect -4077 -2023 -4043 -1963
rect -3898 -2023 -3864 -1963
rect -6302 -2073 -6218 -2039
rect -6174 -2073 -6040 -2039
rect -5996 -2073 -5911 -2039
rect -6302 -2120 -6268 -2073
rect -6234 -2079 -6158 -2073
rect -6126 -2120 -6092 -2073
rect -6056 -2079 -5980 -2073
rect -5945 -2120 -5911 -2073
rect -5878 -2039 -5802 -2023
rect -5878 -2073 -5862 -2039
rect -5818 -2073 -5802 -2039
rect -5878 -2079 -5802 -2073
rect -5700 -2039 -5624 -2023
rect -5700 -2073 -5684 -2039
rect -5640 -2073 -5624 -2039
rect -5700 -2079 -5624 -2073
rect -5522 -2039 -5446 -2023
rect -5522 -2073 -5506 -2039
rect -5462 -2073 -5446 -2039
rect -5522 -2079 -5446 -2073
rect -5344 -2039 -5268 -2023
rect -5344 -2073 -5328 -2039
rect -5284 -2073 -5268 -2039
rect -5344 -2079 -5268 -2073
rect -5166 -2039 -5090 -2023
rect -5166 -2073 -5150 -2039
rect -5106 -2073 -5090 -2039
rect -5166 -2079 -5090 -2073
rect -4988 -2039 -4912 -2023
rect -4988 -2073 -4972 -2039
rect -4928 -2073 -4912 -2039
rect -4988 -2079 -4912 -2073
rect -4810 -2039 -4734 -2023
rect -4810 -2073 -4794 -2039
rect -4750 -2073 -4734 -2039
rect -4810 -2079 -4734 -2073
rect -4632 -2039 -4556 -2023
rect -4632 -2073 -4616 -2039
rect -4572 -2073 -4556 -2039
rect -4632 -2079 -4556 -2073
rect -4454 -2039 -4378 -2023
rect -4454 -2073 -4438 -2039
rect -4394 -2073 -4378 -2039
rect -4454 -2079 -4378 -2073
rect -4276 -2039 -4200 -2023
rect -4276 -2073 -4260 -2039
rect -4216 -2073 -4200 -2039
rect -4276 -2079 -4200 -2073
rect -4098 -2039 -4022 -2023
rect -4098 -2073 -4082 -2039
rect -4038 -2073 -4022 -2039
rect -4098 -2079 -4022 -2073
rect -3920 -2039 -3844 -2023
rect -3920 -2073 -3904 -2039
rect -3860 -2073 -3844 -2039
rect -3920 -2079 -3844 -2073
rect -3810 -2120 -3776 -1841
rect -1119 -1963 -1109 -1910
rect -1056 -1963 -1046 -1910
rect -3742 -2039 -3666 -2023
rect -3742 -2073 -3726 -2039
rect -3682 -2073 -3666 -2039
rect -3742 -2079 -3666 -2073
rect -3564 -2039 -3488 -2023
rect -3564 -2073 -3548 -2039
rect -3504 -2073 -3488 -2039
rect -3564 -2079 -3488 -2073
rect -6308 -2132 -6262 -2120
rect -6308 -2388 -6302 -2132
rect -6268 -2388 -6262 -2132
rect -6308 -2400 -6262 -2388
rect -6130 -2132 -6084 -2120
rect -6130 -2388 -6124 -2132
rect -6090 -2388 -6084 -2132
rect -6130 -2400 -6084 -2388
rect -5952 -2132 -5906 -2120
rect -5952 -2388 -5946 -2132
rect -5912 -2388 -5906 -2132
rect -5952 -2400 -5906 -2388
rect -5774 -2132 -5728 -2120
rect -5774 -2388 -5768 -2132
rect -5734 -2388 -5728 -2132
rect -5774 -2400 -5728 -2388
rect -5596 -2132 -5550 -2120
rect -5596 -2388 -5590 -2132
rect -5556 -2388 -5550 -2132
rect -5596 -2400 -5550 -2388
rect -5418 -2132 -5372 -2120
rect -5418 -2388 -5412 -2132
rect -5378 -2388 -5372 -2132
rect -5418 -2400 -5372 -2388
rect -5240 -2132 -5194 -2120
rect -5240 -2388 -5234 -2132
rect -5200 -2388 -5194 -2132
rect -5240 -2400 -5194 -2388
rect -5062 -2132 -5016 -2120
rect -5062 -2388 -5056 -2132
rect -5022 -2388 -5016 -2132
rect -5062 -2400 -5016 -2388
rect -4884 -2132 -4838 -2120
rect -4884 -2388 -4878 -2132
rect -4844 -2388 -4838 -2132
rect -4884 -2400 -4838 -2388
rect -4706 -2132 -4660 -2120
rect -4706 -2388 -4700 -2132
rect -4666 -2388 -4660 -2132
rect -4706 -2400 -4660 -2388
rect -4528 -2132 -4482 -2120
rect -4528 -2388 -4522 -2132
rect -4488 -2388 -4482 -2132
rect -4528 -2400 -4482 -2388
rect -4350 -2132 -4304 -2120
rect -4350 -2388 -4344 -2132
rect -4310 -2388 -4304 -2132
rect -4350 -2400 -4304 -2388
rect -4172 -2132 -4126 -2120
rect -4172 -2388 -4166 -2132
rect -4132 -2388 -4126 -2132
rect -4172 -2400 -4126 -2388
rect -3994 -2132 -3948 -2120
rect -3994 -2388 -3988 -2132
rect -3954 -2388 -3948 -2132
rect -3994 -2400 -3948 -2388
rect -3816 -2132 -3770 -2120
rect -3816 -2388 -3810 -2132
rect -3776 -2388 -3770 -2132
rect -3816 -2400 -3770 -2388
rect -3638 -2132 -3592 -2120
rect -3638 -2388 -3632 -2132
rect -3598 -2388 -3592 -2132
rect -3638 -2400 -3592 -2388
rect -3460 -2132 -3414 -2120
rect -3460 -2388 -3454 -2132
rect -3420 -2388 -3414 -2132
rect -3460 -2400 -3414 -2388
rect -6234 -2447 -6158 -2441
rect -6234 -2481 -6218 -2447
rect -6174 -2481 -6158 -2447
rect -6234 -2497 -6158 -2481
rect -6056 -2447 -5980 -2441
rect -6056 -2481 -6040 -2447
rect -5996 -2481 -5980 -2447
rect -6056 -2497 -5980 -2481
rect -6508 -2582 -6498 -2529
rect -6445 -2582 -6435 -2529
rect -6635 -3454 -6625 -3401
rect -6572 -3454 -6562 -3401
rect -6625 -5322 -6572 -3454
rect -6498 -3640 -6445 -2582
rect -6054 -2833 -6044 -2780
rect -5991 -2833 -5981 -2780
rect -6035 -2893 -6001 -2833
rect -6234 -2909 -6158 -2893
rect -6234 -2911 -6218 -2909
rect -6302 -2943 -6218 -2911
rect -6174 -2911 -6158 -2909
rect -6056 -2909 -5980 -2893
rect -6174 -2943 -6090 -2911
rect -6302 -2945 -6090 -2943
rect -6302 -2990 -6268 -2945
rect -6234 -2949 -6158 -2945
rect -6124 -2990 -6090 -2945
rect -6056 -2943 -6040 -2909
rect -5996 -2943 -5980 -2909
rect -6056 -2949 -5980 -2943
rect -5946 -2990 -5912 -2400
rect -5878 -2447 -5802 -2441
rect -5878 -2481 -5862 -2447
rect -5818 -2481 -5802 -2447
rect -5878 -2497 -5802 -2481
rect -5856 -2780 -5822 -2497
rect -5768 -2530 -5734 -2400
rect -5700 -2447 -5624 -2441
rect -5700 -2481 -5684 -2447
rect -5640 -2481 -5624 -2447
rect -5700 -2497 -5624 -2481
rect -5787 -2583 -5777 -2530
rect -5724 -2583 -5714 -2530
rect -5876 -2833 -5866 -2780
rect -5813 -2833 -5803 -2780
rect -5856 -2893 -5822 -2833
rect -5679 -2893 -5645 -2497
rect -5878 -2909 -5802 -2893
rect -5878 -2943 -5862 -2909
rect -5818 -2943 -5802 -2909
rect -5878 -2949 -5802 -2943
rect -5700 -2909 -5624 -2893
rect -5700 -2943 -5684 -2909
rect -5640 -2943 -5624 -2909
rect -5700 -2949 -5624 -2943
rect -5590 -2990 -5556 -2400
rect -5522 -2447 -5446 -2441
rect -5522 -2481 -5506 -2447
rect -5462 -2481 -5446 -2447
rect -5522 -2497 -5446 -2481
rect -5501 -2893 -5467 -2497
rect -5412 -2668 -5378 -2400
rect -5344 -2447 -5268 -2441
rect -5344 -2481 -5328 -2447
rect -5284 -2481 -5268 -2447
rect -5344 -2497 -5268 -2481
rect -5431 -2721 -5421 -2668
rect -5368 -2721 -5358 -2668
rect -5323 -2893 -5289 -2497
rect -5522 -2909 -5446 -2893
rect -5522 -2943 -5506 -2909
rect -5462 -2943 -5446 -2909
rect -5522 -2949 -5446 -2943
rect -5344 -2909 -5268 -2893
rect -5344 -2943 -5328 -2909
rect -5284 -2943 -5268 -2909
rect -5344 -2949 -5268 -2943
rect -5234 -2990 -5200 -2400
rect -5166 -2447 -5090 -2441
rect -5166 -2481 -5150 -2447
rect -5106 -2481 -5090 -2447
rect -5166 -2497 -5090 -2481
rect -5145 -2893 -5111 -2497
rect -5056 -2530 -5022 -2400
rect -4988 -2447 -4912 -2441
rect -4988 -2481 -4972 -2447
rect -4928 -2481 -4912 -2447
rect -4988 -2497 -4912 -2481
rect -5076 -2583 -5066 -2530
rect -5013 -2583 -5003 -2530
rect -4967 -2893 -4933 -2497
rect -5166 -2909 -5090 -2893
rect -5166 -2943 -5150 -2909
rect -5106 -2943 -5090 -2909
rect -5166 -2949 -5090 -2943
rect -4988 -2909 -4912 -2893
rect -4988 -2943 -4972 -2909
rect -4928 -2943 -4912 -2909
rect -4988 -2949 -4912 -2943
rect -4878 -2990 -4844 -2400
rect -4810 -2447 -4734 -2441
rect -4810 -2481 -4794 -2447
rect -4750 -2481 -4734 -2447
rect -4810 -2497 -4734 -2481
rect -4789 -2893 -4755 -2497
rect -4700 -2668 -4666 -2400
rect -4632 -2447 -4556 -2441
rect -4632 -2481 -4616 -2447
rect -4572 -2481 -4556 -2447
rect -4632 -2497 -4556 -2481
rect -4720 -2721 -4710 -2668
rect -4657 -2721 -4647 -2668
rect -4611 -2893 -4577 -2497
rect -4810 -2909 -4734 -2893
rect -4810 -2943 -4794 -2909
rect -4750 -2943 -4734 -2909
rect -4810 -2949 -4734 -2943
rect -4632 -2909 -4556 -2893
rect -4632 -2943 -4616 -2909
rect -4572 -2943 -4556 -2909
rect -4632 -2949 -4556 -2943
rect -4522 -2990 -4488 -2400
rect -4454 -2447 -4378 -2441
rect -4454 -2481 -4438 -2447
rect -4394 -2481 -4378 -2447
rect -4454 -2497 -4378 -2481
rect -4433 -2893 -4399 -2497
rect -4344 -2530 -4310 -2400
rect -4276 -2447 -4200 -2441
rect -4276 -2481 -4260 -2447
rect -4216 -2481 -4200 -2447
rect -4276 -2497 -4200 -2481
rect -4364 -2583 -4354 -2530
rect -4301 -2583 -4291 -2530
rect -4255 -2893 -4221 -2497
rect -4454 -2909 -4378 -2893
rect -4454 -2943 -4438 -2909
rect -4394 -2943 -4378 -2909
rect -4454 -2949 -4378 -2943
rect -4276 -2909 -4200 -2893
rect -4276 -2943 -4260 -2909
rect -4216 -2943 -4200 -2909
rect -4276 -2949 -4200 -2943
rect -4166 -2990 -4132 -2400
rect -4098 -2447 -4022 -2441
rect -4098 -2481 -4082 -2447
rect -4038 -2481 -4022 -2447
rect -4098 -2497 -4022 -2481
rect -4077 -2893 -4043 -2497
rect -3988 -2668 -3954 -2400
rect -3920 -2447 -3844 -2441
rect -3920 -2481 -3904 -2447
rect -3860 -2481 -3844 -2447
rect -3920 -2497 -3844 -2481
rect -3810 -2446 -3776 -2400
rect -3742 -2446 -3666 -2441
rect -3633 -2446 -3599 -2400
rect -3564 -2446 -3488 -2441
rect -3454 -2446 -3420 -2400
rect -1099 -2425 -1065 -1963
rect -3810 -2447 -3420 -2446
rect -3810 -2480 -3726 -2447
rect -4008 -2721 -3998 -2668
rect -3945 -2721 -3935 -2668
rect -3899 -2780 -3865 -2497
rect -3918 -2833 -3908 -2780
rect -3855 -2833 -3845 -2780
rect -3899 -2893 -3865 -2833
rect -4098 -2909 -4022 -2893
rect -4098 -2943 -4082 -2909
rect -4038 -2943 -4022 -2909
rect -4098 -2949 -4022 -2943
rect -3920 -2909 -3844 -2893
rect -3920 -2943 -3904 -2909
rect -3860 -2943 -3844 -2909
rect -3920 -2949 -3844 -2943
rect -3810 -2990 -3776 -2480
rect -3742 -2481 -3726 -2480
rect -3682 -2480 -3548 -2447
rect -3682 -2481 -3666 -2480
rect -3742 -2497 -3666 -2481
rect -3564 -2481 -3548 -2480
rect -3504 -2480 -3420 -2447
rect -1119 -2478 -1109 -2425
rect -1056 -2478 -1046 -2425
rect -762 -2478 -752 -2425
rect -699 -2478 -689 -2425
rect -3504 -2481 -3488 -2480
rect -3564 -2497 -3488 -2481
rect -2634 -2611 -2624 -2558
rect -2571 -2611 -2561 -2558
rect -1295 -2611 -1285 -2558
rect -1232 -2611 -1222 -2558
rect -3308 -2721 -3298 -2668
rect -3245 -2721 -3235 -2668
rect -3741 -2833 -3731 -2780
rect -3678 -2833 -3668 -2780
rect -3721 -2893 -3687 -2833
rect -3742 -2909 -3666 -2893
rect -3742 -2943 -3726 -2909
rect -3682 -2943 -3666 -2909
rect -3742 -2949 -3666 -2943
rect -3564 -2909 -3488 -2893
rect -3564 -2943 -3548 -2909
rect -3504 -2943 -3488 -2909
rect -3564 -2949 -3488 -2943
rect -6308 -3002 -6262 -2990
rect -6308 -3258 -6302 -3002
rect -6268 -3258 -6262 -3002
rect -6308 -3270 -6262 -3258
rect -6130 -3002 -6084 -2990
rect -6130 -3258 -6124 -3002
rect -6090 -3258 -6084 -3002
rect -6130 -3270 -6084 -3258
rect -5952 -3002 -5906 -2990
rect -5952 -3258 -5946 -3002
rect -5912 -3258 -5906 -3002
rect -5952 -3270 -5906 -3258
rect -5774 -3002 -5728 -2990
rect -5774 -3258 -5768 -3002
rect -5734 -3258 -5728 -3002
rect -5774 -3270 -5728 -3258
rect -5596 -3002 -5550 -2990
rect -5596 -3258 -5590 -3002
rect -5556 -3258 -5550 -3002
rect -5596 -3270 -5550 -3258
rect -5418 -3002 -5372 -2990
rect -5418 -3258 -5412 -3002
rect -5378 -3258 -5372 -3002
rect -5418 -3270 -5372 -3258
rect -5240 -3002 -5194 -2990
rect -5240 -3258 -5234 -3002
rect -5200 -3258 -5194 -3002
rect -5240 -3270 -5194 -3258
rect -5062 -3002 -5016 -2990
rect -5062 -3258 -5056 -3002
rect -5022 -3258 -5016 -3002
rect -5062 -3270 -5016 -3258
rect -4884 -3002 -4838 -2990
rect -4884 -3258 -4878 -3002
rect -4844 -3258 -4838 -3002
rect -4884 -3270 -4838 -3258
rect -4706 -3002 -4660 -2990
rect -4706 -3258 -4700 -3002
rect -4666 -3258 -4660 -3002
rect -4706 -3270 -4660 -3258
rect -4528 -3002 -4482 -2990
rect -4528 -3258 -4522 -3002
rect -4488 -3258 -4482 -3002
rect -4528 -3270 -4482 -3258
rect -4350 -3002 -4304 -2990
rect -4350 -3258 -4344 -3002
rect -4310 -3258 -4304 -3002
rect -4350 -3270 -4304 -3258
rect -4172 -3002 -4126 -2990
rect -4172 -3258 -4166 -3002
rect -4132 -3258 -4126 -3002
rect -4172 -3270 -4126 -3258
rect -3994 -3002 -3948 -2990
rect -3994 -3258 -3988 -3002
rect -3954 -3258 -3948 -3002
rect -3994 -3270 -3948 -3258
rect -3816 -3002 -3770 -2990
rect -3816 -3258 -3810 -3002
rect -3776 -3258 -3770 -3002
rect -3816 -3270 -3770 -3258
rect -3638 -3002 -3592 -2990
rect -3638 -3258 -3632 -3002
rect -3598 -3258 -3592 -3002
rect -3638 -3270 -3592 -3258
rect -3460 -3002 -3414 -2990
rect -3460 -3258 -3454 -3002
rect -3420 -3258 -3414 -3002
rect -3460 -3270 -3414 -3258
rect -6234 -3317 -6158 -3311
rect -6234 -3351 -6218 -3317
rect -6174 -3351 -6158 -3317
rect -6234 -3367 -6158 -3351
rect -6124 -3401 -6090 -3270
rect -6056 -3317 -5980 -3311
rect -6056 -3351 -6040 -3317
rect -5996 -3351 -5980 -3317
rect -6056 -3367 -5980 -3351
rect -6144 -3454 -6134 -3401
rect -6081 -3454 -6071 -3401
rect -6508 -3693 -6498 -3640
rect -6445 -3693 -6435 -3640
rect -6498 -4271 -6445 -3693
rect -6035 -3763 -6001 -3367
rect -6234 -3778 -6158 -3763
rect -6302 -3779 -6090 -3778
rect -6302 -3812 -6218 -3779
rect -6302 -3860 -6268 -3812
rect -6234 -3813 -6218 -3812
rect -6174 -3812 -6090 -3779
rect -6174 -3813 -6158 -3812
rect -6234 -3819 -6158 -3813
rect -6124 -3860 -6090 -3812
rect -6056 -3779 -5980 -3763
rect -6056 -3813 -6040 -3779
rect -5996 -3813 -5980 -3779
rect -6056 -3819 -5980 -3813
rect -5946 -3860 -5912 -3270
rect -5878 -3317 -5802 -3311
rect -5878 -3351 -5862 -3317
rect -5818 -3351 -5802 -3317
rect -5878 -3367 -5802 -3351
rect -5857 -3763 -5823 -3367
rect -5768 -3516 -5734 -3270
rect -5700 -3317 -5624 -3311
rect -5700 -3351 -5684 -3317
rect -5640 -3351 -5624 -3317
rect -5700 -3367 -5624 -3351
rect -5787 -3569 -5777 -3516
rect -5724 -3569 -5714 -3516
rect -5679 -3763 -5645 -3367
rect -5878 -3779 -5802 -3763
rect -5878 -3813 -5862 -3779
rect -5818 -3813 -5802 -3779
rect -5878 -3819 -5802 -3813
rect -5700 -3779 -5624 -3763
rect -5700 -3813 -5684 -3779
rect -5640 -3813 -5624 -3779
rect -5700 -3819 -5624 -3813
rect -5590 -3860 -5556 -3270
rect -5522 -3317 -5446 -3311
rect -5522 -3351 -5506 -3317
rect -5462 -3351 -5446 -3317
rect -5522 -3367 -5446 -3351
rect -5501 -3763 -5467 -3367
rect -5412 -3640 -5378 -3270
rect -5344 -3317 -5268 -3311
rect -5344 -3351 -5328 -3317
rect -5284 -3351 -5268 -3317
rect -5344 -3367 -5268 -3351
rect -5432 -3693 -5422 -3640
rect -5369 -3693 -5359 -3640
rect -5323 -3763 -5289 -3367
rect -5522 -3779 -5446 -3763
rect -5522 -3813 -5506 -3779
rect -5462 -3813 -5446 -3779
rect -5522 -3819 -5446 -3813
rect -5344 -3779 -5268 -3763
rect -5344 -3813 -5328 -3779
rect -5284 -3813 -5268 -3779
rect -5344 -3819 -5268 -3813
rect -5234 -3860 -5200 -3270
rect -5166 -3317 -5090 -3311
rect -5166 -3351 -5150 -3317
rect -5106 -3351 -5090 -3317
rect -5166 -3367 -5090 -3351
rect -5145 -3763 -5111 -3367
rect -5056 -3401 -5022 -3270
rect -4988 -3317 -4912 -3311
rect -4988 -3351 -4972 -3317
rect -4928 -3351 -4912 -3317
rect -4988 -3367 -4912 -3351
rect -5076 -3454 -5066 -3401
rect -5013 -3454 -5003 -3401
rect -4967 -3763 -4933 -3367
rect -5166 -3779 -5090 -3763
rect -5166 -3813 -5150 -3779
rect -5106 -3813 -5090 -3779
rect -5166 -3819 -5090 -3813
rect -4988 -3779 -4912 -3763
rect -4988 -3813 -4972 -3779
rect -4928 -3813 -4912 -3779
rect -4988 -3819 -4912 -3813
rect -4878 -3860 -4844 -3270
rect -4810 -3317 -4734 -3311
rect -4810 -3351 -4794 -3317
rect -4750 -3351 -4734 -3317
rect -4810 -3367 -4734 -3351
rect -4789 -3763 -4755 -3367
rect -4700 -3401 -4666 -3270
rect -4632 -3317 -4556 -3311
rect -4632 -3351 -4616 -3317
rect -4572 -3351 -4556 -3317
rect -4632 -3367 -4556 -3351
rect -4720 -3454 -4710 -3401
rect -4657 -3454 -4647 -3401
rect -4611 -3763 -4577 -3367
rect -4810 -3779 -4734 -3763
rect -4810 -3813 -4794 -3779
rect -4750 -3813 -4734 -3779
rect -4810 -3819 -4734 -3813
rect -4632 -3779 -4556 -3763
rect -4632 -3813 -4616 -3779
rect -4572 -3813 -4556 -3779
rect -4632 -3819 -4556 -3813
rect -4522 -3860 -4488 -3270
rect -4454 -3317 -4378 -3311
rect -4454 -3351 -4438 -3317
rect -4394 -3351 -4378 -3317
rect -4454 -3367 -4378 -3351
rect -4433 -3763 -4399 -3367
rect -4344 -3640 -4310 -3270
rect -4276 -3317 -4200 -3311
rect -4276 -3351 -4260 -3317
rect -4216 -3351 -4200 -3317
rect -4276 -3367 -4200 -3351
rect -4363 -3693 -4353 -3640
rect -4300 -3693 -4290 -3640
rect -4254 -3763 -4220 -3367
rect -4454 -3779 -4378 -3763
rect -4454 -3813 -4438 -3779
rect -4394 -3813 -4378 -3779
rect -4454 -3819 -4378 -3813
rect -4276 -3779 -4200 -3763
rect -4276 -3813 -4260 -3779
rect -4216 -3813 -4200 -3779
rect -4276 -3819 -4200 -3813
rect -4166 -3860 -4132 -3270
rect -4098 -3317 -4022 -3311
rect -4098 -3351 -4082 -3317
rect -4038 -3351 -4022 -3317
rect -4098 -3367 -4022 -3351
rect -4077 -3763 -4043 -3367
rect -3988 -3516 -3954 -3270
rect -3920 -3317 -3844 -3311
rect -3920 -3351 -3904 -3317
rect -3860 -3351 -3844 -3317
rect -3920 -3367 -3844 -3351
rect -4008 -3569 -3998 -3516
rect -3945 -3569 -3935 -3516
rect -3899 -3763 -3865 -3367
rect -4098 -3779 -4022 -3763
rect -4098 -3813 -4082 -3779
rect -4038 -3813 -4022 -3779
rect -4098 -3819 -4022 -3813
rect -3920 -3779 -3844 -3763
rect -3920 -3813 -3904 -3779
rect -3860 -3813 -3844 -3779
rect -3920 -3819 -3844 -3813
rect -3810 -3860 -3776 -3270
rect -3742 -3317 -3666 -3311
rect -3742 -3351 -3726 -3317
rect -3682 -3351 -3666 -3317
rect -3742 -3367 -3666 -3351
rect -3632 -3316 -3598 -3270
rect -3564 -3316 -3488 -3311
rect -3454 -3316 -3420 -3270
rect -3632 -3317 -3420 -3316
rect -3632 -3350 -3548 -3317
rect -3721 -3763 -3687 -3367
rect -3632 -3401 -3598 -3350
rect -3564 -3351 -3548 -3350
rect -3504 -3350 -3420 -3317
rect -3504 -3351 -3488 -3350
rect -3564 -3367 -3488 -3351
rect -3652 -3454 -3642 -3401
rect -3589 -3454 -3579 -3401
rect -3298 -3516 -3245 -2721
rect -3141 -3454 -3131 -3401
rect -3078 -3454 -3068 -3401
rect -3308 -3569 -3298 -3516
rect -3245 -3569 -3235 -3516
rect -3742 -3779 -3666 -3763
rect -3742 -3813 -3726 -3779
rect -3682 -3813 -3666 -3779
rect -3742 -3819 -3666 -3813
rect -3564 -3779 -3488 -3763
rect -3564 -3813 -3548 -3779
rect -3504 -3813 -3488 -3779
rect -3564 -3819 -3488 -3813
rect -6308 -3872 -6262 -3860
rect -6308 -4128 -6302 -3872
rect -6268 -4128 -6262 -3872
rect -6308 -4140 -6262 -4128
rect -6130 -3872 -6084 -3860
rect -6130 -4128 -6124 -3872
rect -6090 -4128 -6084 -3872
rect -6130 -4140 -6084 -4128
rect -5952 -3872 -5906 -3860
rect -5952 -4128 -5946 -3872
rect -5912 -4128 -5906 -3872
rect -5952 -4140 -5906 -4128
rect -5774 -3872 -5728 -3860
rect -5774 -4128 -5768 -3872
rect -5734 -4128 -5728 -3872
rect -5774 -4140 -5728 -4128
rect -5596 -3872 -5550 -3860
rect -5596 -4128 -5590 -3872
rect -5556 -4128 -5550 -3872
rect -5596 -4140 -5550 -4128
rect -5418 -3872 -5372 -3860
rect -5418 -4128 -5412 -3872
rect -5378 -4128 -5372 -3872
rect -5418 -4140 -5372 -4128
rect -5240 -3872 -5194 -3860
rect -5240 -4128 -5234 -3872
rect -5200 -4128 -5194 -3872
rect -5240 -4140 -5194 -4128
rect -5062 -3872 -5016 -3860
rect -5062 -4128 -5056 -3872
rect -5022 -4128 -5016 -3872
rect -5062 -4140 -5016 -4128
rect -4884 -3872 -4838 -3860
rect -4884 -4128 -4878 -3872
rect -4844 -4128 -4838 -3872
rect -4884 -4140 -4838 -4128
rect -4706 -3872 -4660 -3860
rect -4706 -4128 -4700 -3872
rect -4666 -4128 -4660 -3872
rect -4706 -4140 -4660 -4128
rect -4528 -3872 -4482 -3860
rect -4528 -4128 -4522 -3872
rect -4488 -4128 -4482 -3872
rect -4528 -4140 -4482 -4128
rect -4350 -3872 -4304 -3860
rect -4350 -4128 -4344 -3872
rect -4310 -4128 -4304 -3872
rect -4350 -4140 -4304 -4128
rect -4172 -3872 -4126 -3860
rect -4172 -4128 -4166 -3872
rect -4132 -4128 -4126 -3872
rect -4172 -4140 -4126 -4128
rect -3994 -3872 -3948 -3860
rect -3994 -4128 -3988 -3872
rect -3954 -4128 -3948 -3872
rect -3994 -4140 -3948 -4128
rect -3816 -3872 -3770 -3860
rect -3816 -4128 -3810 -3872
rect -3776 -4128 -3770 -3872
rect -3816 -4140 -3770 -4128
rect -3638 -3872 -3592 -3860
rect -3638 -4128 -3632 -3872
rect -3598 -4128 -3592 -3872
rect -3638 -4140 -3592 -4128
rect -3460 -3872 -3414 -3860
rect -3460 -4128 -3454 -3872
rect -3420 -4128 -3414 -3872
rect -3460 -4140 -3414 -4128
rect -6234 -4187 -6158 -4181
rect -6234 -4221 -6218 -4187
rect -6174 -4221 -6158 -4187
rect -6234 -4237 -6158 -4221
rect -6508 -4324 -6498 -4271
rect -6445 -4324 -6435 -4271
rect -6498 -5141 -6445 -4324
rect -6124 -4390 -6090 -4140
rect -6056 -4187 -5980 -4181
rect -6056 -4221 -6040 -4187
rect -5996 -4221 -5980 -4187
rect -6056 -4237 -5980 -4221
rect -6144 -4443 -6134 -4390
rect -6081 -4443 -6071 -4390
rect -6035 -4633 -6001 -4237
rect -6234 -4649 -6158 -4633
rect -6056 -4649 -5980 -4633
rect -6302 -4683 -6218 -4649
rect -6174 -4683 -6090 -4649
rect -6302 -4730 -6268 -4683
rect -6234 -4689 -6158 -4683
rect -6124 -4730 -6090 -4683
rect -6056 -4683 -6040 -4649
rect -5996 -4683 -5980 -4649
rect -6056 -4689 -5980 -4683
rect -5946 -4730 -5912 -4140
rect -5878 -4187 -5802 -4181
rect -5878 -4221 -5862 -4187
rect -5818 -4221 -5802 -4187
rect -5878 -4237 -5802 -4221
rect -5857 -4633 -5823 -4237
rect -5768 -4271 -5734 -4140
rect -5700 -4187 -5624 -4181
rect -5700 -4221 -5684 -4187
rect -5640 -4221 -5624 -4187
rect -5700 -4237 -5624 -4221
rect -5788 -4324 -5778 -4271
rect -5725 -4324 -5715 -4271
rect -5679 -4633 -5645 -4237
rect -5878 -4649 -5802 -4633
rect -5878 -4683 -5862 -4649
rect -5818 -4683 -5802 -4649
rect -5878 -4689 -5802 -4683
rect -5700 -4649 -5624 -4633
rect -5700 -4683 -5684 -4649
rect -5640 -4683 -5624 -4649
rect -5700 -4689 -5624 -4683
rect -5590 -4730 -5556 -4140
rect -5522 -4187 -5446 -4181
rect -5522 -4221 -5506 -4187
rect -5462 -4221 -5446 -4187
rect -5522 -4237 -5446 -4221
rect -5501 -4633 -5467 -4237
rect -5412 -4506 -5378 -4140
rect -5344 -4187 -5268 -4181
rect -5344 -4221 -5328 -4187
rect -5284 -4221 -5268 -4187
rect -5344 -4237 -5268 -4221
rect -5432 -4559 -5422 -4506
rect -5369 -4559 -5359 -4506
rect -5323 -4633 -5289 -4237
rect -5522 -4649 -5446 -4633
rect -5522 -4683 -5506 -4649
rect -5462 -4683 -5446 -4649
rect -5522 -4689 -5446 -4683
rect -5344 -4649 -5268 -4633
rect -5344 -4683 -5328 -4649
rect -5284 -4683 -5268 -4649
rect -5344 -4689 -5268 -4683
rect -5234 -4730 -5200 -4140
rect -5166 -4187 -5090 -4181
rect -5166 -4221 -5150 -4187
rect -5106 -4221 -5090 -4187
rect -5166 -4237 -5090 -4221
rect -5145 -4633 -5111 -4237
rect -5056 -4390 -5022 -4140
rect -4988 -4187 -4912 -4181
rect -4988 -4221 -4972 -4187
rect -4928 -4221 -4912 -4187
rect -4988 -4237 -4912 -4221
rect -5076 -4443 -5066 -4390
rect -5013 -4443 -5003 -4390
rect -4967 -4633 -4933 -4237
rect -5166 -4649 -5090 -4633
rect -5166 -4683 -5150 -4649
rect -5106 -4683 -5090 -4649
rect -5166 -4689 -5090 -4683
rect -4988 -4649 -4912 -4633
rect -4988 -4683 -4972 -4649
rect -4928 -4683 -4912 -4649
rect -4988 -4689 -4912 -4683
rect -4878 -4730 -4844 -4140
rect -4810 -4187 -4734 -4181
rect -4810 -4221 -4794 -4187
rect -4750 -4221 -4734 -4187
rect -4810 -4237 -4734 -4221
rect -4789 -4633 -4755 -4237
rect -4700 -4390 -4666 -4140
rect -4632 -4187 -4556 -4181
rect -4632 -4221 -4616 -4187
rect -4572 -4221 -4556 -4187
rect -4632 -4237 -4556 -4221
rect -4719 -4443 -4709 -4390
rect -4656 -4443 -4646 -4390
rect -4611 -4633 -4577 -4237
rect -4810 -4649 -4734 -4633
rect -4810 -4683 -4794 -4649
rect -4750 -4683 -4734 -4649
rect -4810 -4689 -4734 -4683
rect -4632 -4649 -4556 -4633
rect -4632 -4683 -4616 -4649
rect -4572 -4683 -4556 -4649
rect -4632 -4689 -4556 -4683
rect -4522 -4730 -4488 -4140
rect -4454 -4187 -4378 -4181
rect -4454 -4221 -4438 -4187
rect -4394 -4221 -4378 -4187
rect -4454 -4237 -4378 -4221
rect -4433 -4633 -4399 -4237
rect -4344 -4506 -4310 -4140
rect -4276 -4187 -4200 -4181
rect -4276 -4221 -4260 -4187
rect -4216 -4221 -4200 -4187
rect -4276 -4237 -4200 -4221
rect -4363 -4559 -4353 -4506
rect -4300 -4559 -4290 -4506
rect -4255 -4633 -4221 -4237
rect -4454 -4649 -4378 -4633
rect -4454 -4683 -4438 -4649
rect -4394 -4683 -4378 -4649
rect -4454 -4689 -4378 -4683
rect -4276 -4649 -4200 -4633
rect -4276 -4683 -4260 -4649
rect -4216 -4683 -4200 -4649
rect -4276 -4689 -4200 -4683
rect -4166 -4730 -4132 -4140
rect -4098 -4187 -4022 -4181
rect -4098 -4221 -4082 -4187
rect -4038 -4221 -4022 -4187
rect -4098 -4237 -4022 -4221
rect -4077 -4633 -4043 -4237
rect -3988 -4271 -3954 -4140
rect -3920 -4187 -3844 -4181
rect -3920 -4221 -3904 -4187
rect -3860 -4221 -3844 -4187
rect -3920 -4237 -3844 -4221
rect -4008 -4324 -3998 -4271
rect -3945 -4324 -3935 -4271
rect -3899 -4633 -3865 -4237
rect -4098 -4649 -4022 -4633
rect -4098 -4683 -4082 -4649
rect -4038 -4683 -4022 -4649
rect -4098 -4689 -4022 -4683
rect -3920 -4649 -3844 -4633
rect -3920 -4683 -3904 -4649
rect -3860 -4683 -3844 -4649
rect -3920 -4689 -3844 -4683
rect -3810 -4730 -3776 -4140
rect -3742 -4187 -3666 -4181
rect -3742 -4221 -3726 -4187
rect -3682 -4221 -3666 -4187
rect -3742 -4237 -3666 -4221
rect -3632 -4186 -3598 -4140
rect -3564 -4186 -3488 -4181
rect -3453 -4186 -3419 -4140
rect -3632 -4187 -3419 -4186
rect -3632 -4220 -3548 -4187
rect -3721 -4633 -3687 -4237
rect -3632 -4390 -3598 -4220
rect -3564 -4221 -3548 -4220
rect -3504 -4220 -3419 -4187
rect -3504 -4221 -3488 -4220
rect -3564 -4237 -3488 -4221
rect -3652 -4443 -3642 -4390
rect -3589 -4443 -3579 -4390
rect -3298 -4506 -3245 -3569
rect -3308 -4559 -3298 -4506
rect -3245 -4559 -3235 -4506
rect -3742 -4649 -3666 -4633
rect -3742 -4683 -3726 -4649
rect -3682 -4683 -3666 -4649
rect -3742 -4689 -3666 -4683
rect -3564 -4649 -3488 -4633
rect -3564 -4683 -3548 -4649
rect -3504 -4683 -3488 -4649
rect -3564 -4689 -3488 -4683
rect -6308 -4742 -6262 -4730
rect -6308 -4998 -6302 -4742
rect -6268 -4998 -6262 -4742
rect -6308 -5010 -6262 -4998
rect -6130 -4742 -6084 -4730
rect -6130 -4998 -6124 -4742
rect -6090 -4998 -6084 -4742
rect -6130 -5010 -6084 -4998
rect -5952 -4742 -5906 -4730
rect -5952 -4998 -5946 -4742
rect -5912 -4998 -5906 -4742
rect -5952 -5010 -5906 -4998
rect -5774 -4742 -5728 -4730
rect -5774 -4998 -5768 -4742
rect -5734 -4998 -5728 -4742
rect -5774 -5010 -5728 -4998
rect -5596 -4742 -5550 -4730
rect -5596 -4998 -5590 -4742
rect -5556 -4998 -5550 -4742
rect -5596 -5010 -5550 -4998
rect -5418 -4742 -5372 -4730
rect -5418 -4998 -5412 -4742
rect -5378 -4998 -5372 -4742
rect -5418 -5010 -5372 -4998
rect -5240 -4742 -5194 -4730
rect -5240 -4998 -5234 -4742
rect -5200 -4998 -5194 -4742
rect -5240 -5010 -5194 -4998
rect -5062 -4742 -5016 -4730
rect -5062 -4998 -5056 -4742
rect -5022 -4998 -5016 -4742
rect -5062 -5010 -5016 -4998
rect -4884 -4742 -4838 -4730
rect -4884 -4998 -4878 -4742
rect -4844 -4998 -4838 -4742
rect -4884 -5010 -4838 -4998
rect -4706 -4742 -4660 -4730
rect -4706 -4998 -4700 -4742
rect -4666 -4998 -4660 -4742
rect -4706 -5010 -4660 -4998
rect -4528 -4742 -4482 -4730
rect -4528 -4998 -4522 -4742
rect -4488 -4998 -4482 -4742
rect -4528 -5010 -4482 -4998
rect -4350 -4742 -4304 -4730
rect -4350 -4998 -4344 -4742
rect -4310 -4998 -4304 -4742
rect -4350 -5010 -4304 -4998
rect -4172 -4742 -4126 -4730
rect -4172 -4998 -4166 -4742
rect -4132 -4998 -4126 -4742
rect -4172 -5010 -4126 -4998
rect -3994 -4742 -3948 -4730
rect -3994 -4998 -3988 -4742
rect -3954 -4998 -3948 -4742
rect -3994 -5010 -3948 -4998
rect -3816 -4742 -3770 -4730
rect -3816 -4998 -3810 -4742
rect -3776 -4998 -3770 -4742
rect -3816 -5010 -3770 -4998
rect -3638 -4742 -3592 -4730
rect -3638 -4998 -3632 -4742
rect -3598 -4998 -3592 -4742
rect -3638 -5010 -3592 -4998
rect -3460 -4742 -3414 -4730
rect -3460 -4998 -3454 -4742
rect -3420 -4998 -3414 -4742
rect -3460 -5010 -3414 -4998
rect -6234 -5057 -6158 -5051
rect -6234 -5091 -6218 -5057
rect -6174 -5091 -6158 -5057
rect -6234 -5107 -6158 -5091
rect -6508 -5194 -6498 -5141
rect -6445 -5194 -6435 -5141
rect -6635 -5375 -6625 -5322
rect -6572 -5375 -6562 -5322
rect -6498 -6248 -6445 -5194
rect -6124 -5232 -6090 -5010
rect -6056 -5057 -5980 -5051
rect -6056 -5091 -6040 -5057
rect -5996 -5091 -5980 -5057
rect -6056 -5107 -5980 -5091
rect -6144 -5285 -6134 -5232
rect -6081 -5285 -6071 -5232
rect -6234 -5518 -6158 -5503
rect -6301 -5519 -6091 -5518
rect -6056 -5519 -5980 -5503
rect -5946 -5519 -5912 -5010
rect -5878 -5057 -5802 -5051
rect -5878 -5091 -5862 -5057
rect -5818 -5091 -5802 -5057
rect -5878 -5107 -5802 -5091
rect -5857 -5503 -5823 -5107
rect -5768 -5415 -5734 -5010
rect -5700 -5057 -5624 -5051
rect -5700 -5091 -5684 -5057
rect -5640 -5091 -5624 -5057
rect -5700 -5107 -5624 -5091
rect -5787 -5468 -5777 -5415
rect -5724 -5468 -5714 -5415
rect -5679 -5503 -5645 -5107
rect -6301 -5552 -6218 -5519
rect -6301 -5600 -6267 -5552
rect -6234 -5553 -6218 -5552
rect -6174 -5552 -6040 -5519
rect -6174 -5553 -6158 -5552
rect -6234 -5559 -6158 -5553
rect -6125 -5553 -6040 -5552
rect -5996 -5553 -5912 -5519
rect -6125 -5600 -6091 -5553
rect -6056 -5559 -5980 -5553
rect -5946 -5600 -5912 -5553
rect -5878 -5519 -5802 -5503
rect -5878 -5553 -5862 -5519
rect -5818 -5553 -5802 -5519
rect -5878 -5559 -5802 -5553
rect -5700 -5519 -5624 -5503
rect -5700 -5553 -5684 -5519
rect -5640 -5553 -5624 -5519
rect -5700 -5559 -5624 -5553
rect -5590 -5600 -5556 -5010
rect -5522 -5057 -5446 -5051
rect -5522 -5091 -5506 -5057
rect -5462 -5091 -5446 -5057
rect -5522 -5107 -5446 -5091
rect -5501 -5503 -5467 -5107
rect -5412 -5141 -5378 -5010
rect -5344 -5057 -5268 -5051
rect -5344 -5091 -5328 -5057
rect -5284 -5091 -5268 -5057
rect -5344 -5107 -5268 -5091
rect -5432 -5194 -5422 -5141
rect -5369 -5194 -5359 -5141
rect -5323 -5503 -5289 -5107
rect -5522 -5519 -5446 -5503
rect -5522 -5553 -5506 -5519
rect -5462 -5553 -5446 -5519
rect -5522 -5559 -5446 -5553
rect -5344 -5519 -5268 -5503
rect -5344 -5553 -5328 -5519
rect -5284 -5553 -5268 -5519
rect -5344 -5559 -5268 -5553
rect -5234 -5600 -5200 -5010
rect -5166 -5057 -5090 -5051
rect -5166 -5091 -5150 -5057
rect -5106 -5091 -5090 -5057
rect -5166 -5107 -5090 -5091
rect -5145 -5503 -5111 -5107
rect -5056 -5233 -5022 -5010
rect -4988 -5057 -4912 -5051
rect -4988 -5091 -4972 -5057
rect -4928 -5091 -4912 -5057
rect -4988 -5107 -4912 -5091
rect -5076 -5286 -5066 -5233
rect -5013 -5286 -5003 -5233
rect -4967 -5503 -4933 -5107
rect -5166 -5519 -5090 -5503
rect -5166 -5553 -5150 -5519
rect -5106 -5553 -5090 -5519
rect -5166 -5559 -5090 -5553
rect -4988 -5519 -4912 -5503
rect -4988 -5553 -4972 -5519
rect -4928 -5553 -4912 -5519
rect -4988 -5559 -4912 -5553
rect -4878 -5600 -4844 -5010
rect -4810 -5057 -4734 -5051
rect -4810 -5091 -4794 -5057
rect -4750 -5091 -4734 -5057
rect -4810 -5107 -4734 -5091
rect -4789 -5503 -4755 -5107
rect -4700 -5322 -4666 -5010
rect -4632 -5057 -4556 -5051
rect -4632 -5091 -4616 -5057
rect -4572 -5091 -4556 -5057
rect -4632 -5107 -4556 -5091
rect -4720 -5375 -4710 -5322
rect -4657 -5375 -4647 -5322
rect -4611 -5503 -4577 -5107
rect -4810 -5519 -4734 -5503
rect -4810 -5553 -4794 -5519
rect -4750 -5553 -4734 -5519
rect -4810 -5559 -4734 -5553
rect -4632 -5519 -4556 -5503
rect -4632 -5553 -4616 -5519
rect -4572 -5553 -4556 -5519
rect -4632 -5559 -4556 -5553
rect -4522 -5600 -4488 -5010
rect -4454 -5057 -4378 -5051
rect -4454 -5091 -4438 -5057
rect -4394 -5091 -4378 -5057
rect -4454 -5107 -4378 -5091
rect -4433 -5503 -4399 -5107
rect -4344 -5141 -4310 -5010
rect -4276 -5057 -4200 -5051
rect -4276 -5091 -4260 -5057
rect -4216 -5091 -4200 -5057
rect -4276 -5107 -4200 -5091
rect -4363 -5194 -4353 -5141
rect -4300 -5194 -4290 -5141
rect -4255 -5503 -4221 -5107
rect -4454 -5519 -4378 -5503
rect -4454 -5553 -4438 -5519
rect -4394 -5553 -4378 -5519
rect -4454 -5559 -4378 -5553
rect -4276 -5519 -4200 -5503
rect -4276 -5553 -4260 -5519
rect -4216 -5553 -4200 -5519
rect -4276 -5559 -4200 -5553
rect -4166 -5600 -4132 -5010
rect -4098 -5057 -4022 -5051
rect -4098 -5091 -4082 -5057
rect -4038 -5091 -4022 -5057
rect -4098 -5107 -4022 -5091
rect -4077 -5503 -4043 -5107
rect -3988 -5415 -3954 -5010
rect -3920 -5057 -3844 -5051
rect -3920 -5091 -3904 -5057
rect -3860 -5091 -3844 -5057
rect -3920 -5107 -3844 -5091
rect -4007 -5468 -3997 -5415
rect -3944 -5468 -3934 -5415
rect -3899 -5503 -3865 -5107
rect -4098 -5519 -4022 -5503
rect -4098 -5553 -4082 -5519
rect -4038 -5553 -4022 -5519
rect -4098 -5559 -4022 -5553
rect -3920 -5519 -3844 -5503
rect -3920 -5553 -3904 -5519
rect -3860 -5553 -3844 -5519
rect -3920 -5559 -3844 -5553
rect -3810 -5600 -3776 -5010
rect -3742 -5057 -3666 -5051
rect -3742 -5091 -3726 -5057
rect -3682 -5091 -3666 -5057
rect -3742 -5107 -3666 -5091
rect -3632 -5056 -3598 -5010
rect -3564 -5056 -3488 -5051
rect -3453 -5056 -3419 -5010
rect -3632 -5057 -3419 -5056
rect -3632 -5090 -3548 -5057
rect -3632 -5319 -3598 -5090
rect -3564 -5091 -3548 -5090
rect -3504 -5090 -3419 -5057
rect -3504 -5091 -3488 -5090
rect -3564 -5107 -3488 -5091
rect -3652 -5372 -3642 -5319
rect -3589 -5372 -3579 -5319
rect -3298 -5416 -3245 -4559
rect -3130 -5233 -3077 -3454
rect -3140 -5286 -3130 -5233
rect -3077 -5286 -3067 -5233
rect -2624 -5324 -2571 -2611
rect -1386 -2791 -1310 -2775
rect -1386 -2825 -1370 -2791
rect -1326 -2825 -1310 -2791
rect -1386 -2831 -1310 -2825
rect -1276 -2872 -1242 -2611
rect -1207 -2718 -1197 -2665
rect -1144 -2718 -1134 -2665
rect -1187 -2775 -1153 -2718
rect -1208 -2791 -1132 -2775
rect -1208 -2825 -1192 -2791
rect -1148 -2825 -1132 -2791
rect -1208 -2831 -1132 -2825
rect -1099 -2872 -1065 -2478
rect -940 -2611 -930 -2558
rect -877 -2611 -867 -2558
rect -1029 -2718 -1019 -2665
rect -966 -2718 -956 -2665
rect -1009 -2775 -975 -2718
rect -1030 -2791 -954 -2775
rect -1030 -2825 -1014 -2791
rect -970 -2825 -954 -2791
rect -1030 -2831 -954 -2825
rect -920 -2872 -886 -2611
rect -851 -2718 -841 -2665
rect -788 -2718 -778 -2665
rect -831 -2775 -797 -2718
rect -852 -2791 -776 -2775
rect -852 -2825 -836 -2791
rect -792 -2825 -776 -2791
rect -852 -2831 -776 -2825
rect -742 -2872 -708 -2478
rect -208 -2605 182 -2571
rect -674 -2791 -598 -2775
rect -674 -2825 -658 -2791
rect -614 -2825 -598 -2791
rect -674 -2831 -598 -2825
rect -496 -2791 -420 -2775
rect -496 -2825 -480 -2791
rect -436 -2825 -420 -2791
rect -496 -2831 -420 -2825
rect -318 -2791 -242 -2775
rect -318 -2825 -302 -2791
rect -258 -2825 -242 -2791
rect -318 -2831 -242 -2825
rect -208 -2872 -174 -2605
rect -139 -2718 -129 -2665
rect -76 -2718 -66 -2665
rect 40 -2718 50 -2665
rect 103 -2718 113 -2665
rect -119 -2775 -85 -2718
rect 59 -2775 93 -2718
rect -140 -2791 -64 -2775
rect -140 -2825 -124 -2791
rect -80 -2825 -64 -2791
rect -140 -2831 -64 -2825
rect 38 -2791 114 -2775
rect 38 -2825 54 -2791
rect 98 -2825 114 -2791
rect 38 -2831 114 -2825
rect 148 -2872 182 -2605
rect 217 -2718 227 -2665
rect 280 -2718 290 -2665
rect 237 -2775 271 -2718
rect 594 -2775 628 -1467
rect 5327 -2258 5337 -2205
rect 5390 -2258 5400 -2205
rect 1909 -2479 1919 -2426
rect 1972 -2479 1982 -2426
rect 2265 -2479 2275 -2426
rect 2328 -2479 2338 -2426
rect 1038 -2611 1428 -2577
rect 930 -2718 940 -2665
rect 993 -2718 1003 -2665
rect 949 -2775 983 -2718
rect 216 -2791 292 -2775
rect 216 -2825 232 -2791
rect 276 -2825 292 -2791
rect 216 -2831 292 -2825
rect 394 -2791 470 -2775
rect 394 -2825 410 -2791
rect 454 -2825 470 -2791
rect 394 -2831 470 -2825
rect 572 -2791 648 -2775
rect 572 -2825 588 -2791
rect 632 -2825 648 -2791
rect 572 -2831 648 -2825
rect 750 -2791 826 -2775
rect 750 -2825 766 -2791
rect 810 -2825 826 -2791
rect 750 -2831 826 -2825
rect 928 -2791 1004 -2775
rect 928 -2825 944 -2791
rect 988 -2825 1004 -2791
rect 928 -2831 1004 -2825
rect 1038 -2872 1072 -2611
rect 1107 -2718 1117 -2665
rect 1170 -2718 1180 -2665
rect 1285 -2718 1295 -2665
rect 1348 -2718 1358 -2665
rect 1127 -2775 1161 -2718
rect 1305 -2775 1339 -2718
rect 1106 -2791 1182 -2775
rect 1106 -2825 1122 -2791
rect 1166 -2825 1182 -2791
rect 1106 -2831 1182 -2825
rect 1284 -2791 1360 -2775
rect 1284 -2825 1300 -2791
rect 1344 -2825 1360 -2791
rect 1284 -2831 1360 -2825
rect 1394 -2872 1428 -2611
rect 1462 -2791 1538 -2775
rect 1462 -2825 1478 -2791
rect 1522 -2825 1538 -2791
rect 1462 -2831 1538 -2825
rect 1640 -2791 1716 -2775
rect 1640 -2825 1656 -2791
rect 1700 -2825 1716 -2791
rect 1640 -2831 1716 -2825
rect 1818 -2791 1894 -2775
rect 1818 -2825 1834 -2791
rect 1878 -2825 1894 -2791
rect 1818 -2831 1894 -2825
rect 1928 -2872 1962 -2479
rect 2087 -2607 2097 -2554
rect 2150 -2607 2160 -2554
rect 1997 -2718 2007 -2665
rect 2060 -2718 2070 -2665
rect 2017 -2775 2051 -2718
rect 1996 -2791 2072 -2775
rect 1996 -2825 2012 -2791
rect 2056 -2825 2072 -2791
rect 1996 -2831 2072 -2825
rect 2105 -2872 2139 -2607
rect 2176 -2718 2186 -2665
rect 2239 -2718 2249 -2665
rect 2195 -2775 2229 -2718
rect 2174 -2791 2250 -2775
rect 2174 -2825 2190 -2791
rect 2234 -2825 2250 -2791
rect 2174 -2831 2250 -2825
rect 2285 -2872 2319 -2479
rect 3183 -2480 3193 -2427
rect 3246 -2480 3256 -2427
rect 2443 -2607 2453 -2554
rect 2506 -2606 2931 -2554
rect 2506 -2607 2516 -2606
rect 2353 -2718 2363 -2665
rect 2416 -2718 2426 -2665
rect 2373 -2775 2407 -2718
rect 2352 -2791 2428 -2775
rect 2352 -2825 2368 -2791
rect 2412 -2825 2428 -2791
rect 2352 -2831 2428 -2825
rect 2462 -2872 2496 -2607
rect 2530 -2791 2606 -2775
rect 2530 -2825 2546 -2791
rect 2590 -2825 2606 -2791
rect 2530 -2831 2606 -2825
rect -1460 -2884 -1414 -2872
rect -2198 -3043 -1996 -3037
rect -2198 -3221 -2186 -3043
rect -2008 -3221 -1996 -3043
rect -1460 -3140 -1454 -2884
rect -1420 -3140 -1414 -2884
rect -1460 -3152 -1414 -3140
rect -1282 -2884 -1236 -2872
rect -1282 -3140 -1276 -2884
rect -1242 -3140 -1236 -2884
rect -1282 -3152 -1236 -3140
rect -1104 -2884 -1058 -2872
rect -1104 -3140 -1098 -2884
rect -1064 -3140 -1058 -2884
rect -1104 -3152 -1058 -3140
rect -926 -2884 -880 -2872
rect -926 -3140 -920 -2884
rect -886 -3140 -880 -2884
rect -926 -3152 -880 -3140
rect -748 -2884 -702 -2872
rect -748 -3140 -742 -2884
rect -708 -3140 -702 -2884
rect -748 -3152 -702 -3140
rect -570 -2884 -524 -2872
rect -570 -3140 -564 -2884
rect -530 -3140 -524 -2884
rect -570 -3152 -524 -3140
rect -392 -2884 -346 -2872
rect -392 -3140 -386 -2884
rect -352 -3140 -346 -2884
rect -392 -3152 -346 -3140
rect -214 -2884 -168 -2872
rect -214 -3140 -208 -2884
rect -174 -3140 -168 -2884
rect -214 -3152 -168 -3140
rect -36 -2884 10 -2872
rect -36 -3140 -30 -2884
rect 4 -3140 10 -2884
rect -36 -3152 10 -3140
rect 142 -2884 188 -2872
rect 142 -3140 148 -2884
rect 182 -3140 188 -2884
rect 142 -3152 188 -3140
rect 320 -2884 366 -2872
rect 320 -3140 326 -2884
rect 360 -3140 366 -2884
rect 320 -3152 366 -3140
rect 498 -2884 544 -2872
rect 498 -3140 504 -2884
rect 538 -3140 544 -2884
rect 498 -3152 544 -3140
rect 676 -2884 722 -2872
rect 676 -3140 682 -2884
rect 716 -3140 722 -2884
rect 676 -3152 722 -3140
rect 854 -2884 900 -2872
rect 854 -3140 860 -2884
rect 894 -3140 900 -2884
rect 854 -3152 900 -3140
rect 1032 -2884 1078 -2872
rect 1032 -3140 1038 -2884
rect 1072 -3140 1078 -2884
rect 1032 -3152 1078 -3140
rect 1210 -2884 1256 -2872
rect 1210 -3140 1216 -2884
rect 1250 -3140 1256 -2884
rect 1210 -3152 1256 -3140
rect 1388 -2884 1434 -2872
rect 1388 -3140 1394 -2884
rect 1428 -3140 1434 -2884
rect 1388 -3152 1434 -3140
rect 1566 -2884 1612 -2872
rect 1566 -3140 1572 -2884
rect 1606 -3140 1612 -2884
rect 1566 -3152 1612 -3140
rect 1744 -2884 1790 -2872
rect 1744 -3140 1750 -2884
rect 1784 -3140 1790 -2884
rect 1744 -3152 1790 -3140
rect 1922 -2884 1968 -2872
rect 1922 -3140 1928 -2884
rect 1962 -3140 1968 -2884
rect 1922 -3152 1968 -3140
rect 2100 -2884 2146 -2872
rect 2100 -3140 2106 -2884
rect 2140 -3140 2146 -2884
rect 2100 -3152 2146 -3140
rect 2278 -2884 2324 -2872
rect 2278 -3140 2284 -2884
rect 2318 -3140 2324 -2884
rect 2278 -3152 2324 -3140
rect 2456 -2884 2502 -2872
rect 2456 -3140 2462 -2884
rect 2496 -3140 2502 -2884
rect 2456 -3152 2502 -3140
rect 2634 -2884 2680 -2872
rect 2634 -3140 2640 -2884
rect 2674 -3140 2680 -2884
rect 2634 -3152 2680 -3140
rect -2198 -3227 -1996 -3221
rect -1454 -3282 -1420 -3152
rect -1386 -3199 -1310 -3193
rect -1386 -3233 -1370 -3199
rect -1326 -3233 -1310 -3199
rect -1386 -3249 -1310 -3233
rect -1365 -3282 -1331 -3249
rect -1276 -3282 -1242 -3152
rect -1208 -3199 -1132 -3193
rect -1208 -3233 -1192 -3199
rect -1148 -3233 -1132 -3199
rect -1208 -3249 -1132 -3233
rect -1030 -3199 -954 -3193
rect -1030 -3233 -1014 -3199
rect -970 -3233 -954 -3199
rect -1030 -3249 -954 -3233
rect -852 -3199 -776 -3193
rect -852 -3233 -836 -3199
rect -792 -3233 -776 -3199
rect -852 -3249 -776 -3233
rect -674 -3199 -598 -3193
rect -674 -3233 -658 -3199
rect -614 -3233 -598 -3199
rect -674 -3249 -598 -3233
rect -1454 -3316 -1242 -3282
rect -1454 -3317 -1420 -3316
rect -1655 -3510 -1645 -3449
rect -1584 -3510 -1574 -3449
rect -2014 -4465 -2004 -4412
rect -1951 -4465 -1941 -4412
rect -2003 -4517 -1950 -4465
rect -2634 -5377 -2624 -5324
rect -2571 -5377 -2561 -5324
rect -3308 -5469 -3298 -5416
rect -3245 -5469 -3235 -5416
rect -3742 -5519 -3666 -5503
rect -3742 -5553 -3726 -5519
rect -3682 -5553 -3666 -5519
rect -3742 -5559 -3666 -5553
rect -3564 -5519 -3488 -5503
rect -3564 -5553 -3548 -5519
rect -3504 -5553 -3488 -5519
rect -3564 -5559 -3488 -5553
rect -6308 -5612 -6262 -5600
rect -6308 -5868 -6302 -5612
rect -6268 -5868 -6262 -5612
rect -6308 -5880 -6262 -5868
rect -6130 -5612 -6084 -5600
rect -6130 -5868 -6124 -5612
rect -6090 -5868 -6084 -5612
rect -6130 -5880 -6084 -5868
rect -5952 -5612 -5906 -5600
rect -5952 -5868 -5946 -5612
rect -5912 -5868 -5906 -5612
rect -5952 -5880 -5906 -5868
rect -5774 -5612 -5728 -5600
rect -5774 -5868 -5768 -5612
rect -5734 -5868 -5728 -5612
rect -5774 -5880 -5728 -5868
rect -5596 -5612 -5550 -5600
rect -5596 -5868 -5590 -5612
rect -5556 -5868 -5550 -5612
rect -5596 -5880 -5550 -5868
rect -5418 -5612 -5372 -5600
rect -5418 -5868 -5412 -5612
rect -5378 -5868 -5372 -5612
rect -5418 -5880 -5372 -5868
rect -5240 -5612 -5194 -5600
rect -5240 -5868 -5234 -5612
rect -5200 -5868 -5194 -5612
rect -5240 -5880 -5194 -5868
rect -5062 -5612 -5016 -5600
rect -5062 -5868 -5056 -5612
rect -5022 -5868 -5016 -5612
rect -5062 -5880 -5016 -5868
rect -4884 -5612 -4838 -5600
rect -4884 -5868 -4878 -5612
rect -4844 -5868 -4838 -5612
rect -4884 -5880 -4838 -5868
rect -4706 -5612 -4660 -5600
rect -4706 -5868 -4700 -5612
rect -4666 -5868 -4660 -5612
rect -4706 -5880 -4660 -5868
rect -4528 -5612 -4482 -5600
rect -4528 -5868 -4522 -5612
rect -4488 -5868 -4482 -5612
rect -4528 -5880 -4482 -5868
rect -4350 -5612 -4304 -5600
rect -4350 -5868 -4344 -5612
rect -4310 -5868 -4304 -5612
rect -4350 -5880 -4304 -5868
rect -4172 -5612 -4126 -5600
rect -4172 -5868 -4166 -5612
rect -4132 -5868 -4126 -5612
rect -4172 -5880 -4126 -5868
rect -3994 -5612 -3948 -5600
rect -3994 -5868 -3988 -5612
rect -3954 -5868 -3948 -5612
rect -3994 -5880 -3948 -5868
rect -3816 -5612 -3770 -5600
rect -3816 -5868 -3810 -5612
rect -3776 -5868 -3770 -5612
rect -3816 -5880 -3770 -5868
rect -3638 -5612 -3592 -5600
rect -3638 -5868 -3632 -5612
rect -3598 -5868 -3592 -5612
rect -3638 -5880 -3592 -5868
rect -3460 -5612 -3414 -5600
rect -3460 -5868 -3454 -5612
rect -3420 -5868 -3414 -5612
rect -3460 -5880 -3414 -5868
rect -6234 -5927 -6158 -5921
rect -6234 -5961 -6218 -5927
rect -6174 -5961 -6158 -5927
rect -6234 -5977 -6158 -5961
rect -6056 -5927 -5980 -5921
rect -6056 -5961 -6040 -5927
rect -5996 -5961 -5980 -5927
rect -6056 -5977 -5980 -5961
rect -5946 -6016 -5912 -5880
rect -5878 -5927 -5802 -5921
rect -5878 -5961 -5862 -5927
rect -5818 -5961 -5802 -5927
rect -5878 -5977 -5802 -5961
rect -5966 -6069 -5956 -6016
rect -5903 -6069 -5893 -6016
rect -5768 -6131 -5734 -5880
rect -5700 -5927 -5624 -5921
rect -5700 -5961 -5684 -5927
rect -5640 -5961 -5624 -5927
rect -5700 -5977 -5624 -5961
rect -5590 -6016 -5556 -5880
rect -5522 -5927 -5446 -5921
rect -5522 -5961 -5506 -5927
rect -5462 -5961 -5446 -5927
rect -5522 -5977 -5446 -5961
rect -5611 -6069 -5601 -6016
rect -5548 -6069 -5538 -6016
rect -5788 -6184 -5778 -6131
rect -5725 -6184 -5715 -6131
rect -5412 -6248 -5378 -5880
rect -5344 -5927 -5268 -5921
rect -5344 -5961 -5328 -5927
rect -5284 -5961 -5268 -5927
rect -5344 -5977 -5268 -5961
rect -5234 -6016 -5200 -5880
rect -5166 -5927 -5090 -5921
rect -5166 -5961 -5150 -5927
rect -5106 -5961 -5090 -5927
rect -5166 -5977 -5090 -5961
rect -5254 -6069 -5244 -6016
rect -5191 -6069 -5181 -6016
rect -5056 -6131 -5022 -5880
rect -4988 -5927 -4912 -5921
rect -4988 -5961 -4972 -5927
rect -4928 -5961 -4912 -5927
rect -4988 -5977 -4912 -5961
rect -5075 -6184 -5065 -6131
rect -5012 -6184 -5002 -6131
rect -6508 -6301 -6498 -6248
rect -6445 -6301 -6435 -6248
rect -5431 -6301 -5421 -6248
rect -5368 -6301 -5358 -6248
rect -4967 -6376 -4933 -5977
rect -4878 -6016 -4844 -5880
rect -4810 -5927 -4734 -5921
rect -4810 -5961 -4794 -5927
rect -4750 -5961 -4734 -5927
rect -4810 -5977 -4734 -5961
rect -4898 -6069 -4888 -6016
rect -4835 -6069 -4825 -6016
rect -4700 -6248 -4666 -5880
rect -4632 -5927 -4556 -5921
rect -4632 -5961 -4616 -5927
rect -4572 -5961 -4556 -5927
rect -4632 -5977 -4556 -5961
rect -4720 -6301 -4710 -6248
rect -4657 -6301 -4647 -6248
rect -4613 -6376 -4579 -5977
rect -4522 -6016 -4488 -5880
rect -4454 -5927 -4378 -5921
rect -4454 -5961 -4438 -5927
rect -4394 -5961 -4378 -5927
rect -4454 -5977 -4378 -5961
rect -4542 -6069 -4532 -6016
rect -4479 -6069 -4469 -6016
rect -4344 -6131 -4310 -5880
rect -4276 -5927 -4200 -5921
rect -4276 -5961 -4260 -5927
rect -4216 -5961 -4200 -5927
rect -4276 -5977 -4200 -5961
rect -4166 -6016 -4132 -5880
rect -4098 -5927 -4022 -5921
rect -4098 -5961 -4082 -5927
rect -4038 -5961 -4022 -5927
rect -4098 -5977 -4022 -5961
rect -4185 -6069 -4175 -6016
rect -4122 -6069 -4112 -6016
rect -4364 -6184 -4354 -6131
rect -4301 -6184 -4291 -6131
rect -3988 -6247 -3954 -5880
rect -3920 -5927 -3844 -5921
rect -3920 -5961 -3904 -5927
rect -3860 -5961 -3844 -5927
rect -3920 -5977 -3844 -5961
rect -3810 -5928 -3776 -5880
rect -3742 -5927 -3666 -5921
rect -3742 -5928 -3726 -5927
rect -3810 -5961 -3726 -5928
rect -3682 -5928 -3666 -5927
rect -3632 -5928 -3598 -5880
rect -3564 -5927 -3488 -5921
rect -3564 -5928 -3548 -5927
rect -3682 -5961 -3548 -5928
rect -3504 -5928 -3488 -5927
rect -3455 -5928 -3421 -5880
rect -3504 -5961 -3421 -5928
rect -3810 -5962 -3421 -5961
rect -3810 -6016 -3776 -5962
rect -3742 -5977 -3666 -5962
rect -3564 -5977 -3488 -5962
rect -3830 -6069 -3820 -6016
rect -3767 -6069 -3757 -6016
rect -3298 -6131 -3245 -5469
rect -3046 -5662 -2844 -5656
rect -3046 -5840 -3034 -5662
rect -2856 -5840 -2844 -5662
rect -3046 -5846 -2844 -5840
rect -2624 -6007 -2571 -5377
rect -2634 -6060 -2624 -6007
rect -2571 -6060 -2561 -6007
rect -3308 -6184 -3298 -6131
rect -3245 -6184 -3235 -6131
rect -4008 -6300 -3998 -6247
rect -3945 -6300 -3935 -6247
rect -3988 -6301 -3954 -6300
rect -4967 -6378 -4579 -6376
rect -4967 -6410 -4786 -6378
rect -4796 -6431 -4786 -6410
rect -4733 -6410 -4579 -6378
rect -4733 -6431 -4723 -6410
rect -2002 -6714 -1950 -4517
rect -1886 -5285 -1876 -5232
rect -1823 -5285 -1813 -5232
rect -1646 -5278 -1585 -3510
rect -1296 -3624 -1286 -3571
rect -1233 -3624 -1223 -3571
rect -1386 -3691 -1310 -3675
rect -1386 -3725 -1370 -3691
rect -1326 -3725 -1310 -3691
rect -1386 -3731 -1310 -3725
rect -1276 -3772 -1242 -3624
rect -1186 -3675 -1152 -3249
rect -1118 -3509 -1108 -3456
rect -1055 -3509 -1045 -3456
rect -1208 -3691 -1132 -3675
rect -1208 -3725 -1192 -3691
rect -1148 -3725 -1132 -3691
rect -1208 -3731 -1132 -3725
rect -1098 -3772 -1064 -3509
rect -1009 -3675 -975 -3249
rect -939 -3624 -929 -3571
rect -876 -3624 -866 -3571
rect -1030 -3691 -954 -3675
rect -1030 -3725 -1014 -3691
rect -970 -3725 -954 -3691
rect -1030 -3731 -954 -3725
rect -919 -3772 -885 -3624
rect -831 -3675 -797 -3249
rect -653 -3282 -619 -3249
rect -563 -3282 -529 -3152
rect -496 -3199 -420 -3193
rect -496 -3233 -480 -3199
rect -436 -3233 -420 -3199
rect -496 -3249 -420 -3233
rect -474 -3282 -440 -3249
rect -385 -3282 -351 -3152
rect -318 -3199 -242 -3193
rect -318 -3233 -302 -3199
rect -258 -3233 -242 -3199
rect -318 -3249 -242 -3233
rect -295 -3282 -261 -3249
rect -653 -3301 -261 -3282
rect -653 -3316 -484 -3301
rect -494 -3354 -484 -3316
rect -431 -3316 -261 -3301
rect -431 -3354 -421 -3316
rect -760 -3509 -750 -3456
rect -697 -3509 -687 -3456
rect -406 -3509 -396 -3456
rect -343 -3509 -333 -3456
rect -852 -3691 -776 -3675
rect -852 -3725 -836 -3691
rect -792 -3725 -776 -3691
rect -852 -3731 -776 -3725
rect -742 -3772 -708 -3509
rect -583 -3624 -573 -3571
rect -520 -3624 -510 -3571
rect -674 -3691 -598 -3675
rect -674 -3725 -658 -3691
rect -614 -3725 -598 -3691
rect -674 -3731 -598 -3725
rect -564 -3772 -530 -3624
rect -496 -3691 -420 -3675
rect -496 -3725 -480 -3691
rect -436 -3725 -420 -3691
rect -496 -3731 -420 -3725
rect -386 -3772 -352 -3509
rect -208 -3571 -174 -3152
rect -140 -3199 -64 -3193
rect -140 -3233 -124 -3199
rect -80 -3233 -64 -3199
rect -140 -3249 -64 -3233
rect -227 -3624 -217 -3571
rect -164 -3624 -154 -3571
rect -318 -3691 -242 -3675
rect -318 -3725 -302 -3691
rect -258 -3725 -242 -3691
rect -318 -3731 -242 -3725
rect -208 -3772 -174 -3624
rect -119 -3675 -85 -3249
rect -30 -3456 4 -3152
rect 38 -3199 114 -3193
rect 38 -3233 54 -3199
rect 98 -3233 114 -3199
rect 38 -3249 114 -3233
rect 216 -3199 292 -3193
rect 216 -3233 232 -3199
rect 276 -3233 292 -3199
rect 216 -3249 292 -3233
rect 327 -3456 361 -3152
rect 394 -3199 470 -3193
rect 394 -3233 410 -3199
rect 454 -3233 470 -3199
rect 394 -3249 470 -3233
rect 414 -3283 448 -3249
rect 504 -3283 538 -3152
rect 572 -3199 648 -3193
rect 572 -3233 588 -3199
rect 632 -3233 648 -3199
rect 572 -3249 648 -3233
rect 592 -3283 626 -3249
rect 682 -3283 716 -3152
rect 750 -3199 826 -3193
rect 750 -3233 766 -3199
rect 810 -3233 826 -3199
rect 750 -3249 826 -3233
rect 771 -3283 805 -3249
rect 414 -3301 805 -3283
rect 414 -3317 583 -3301
rect 573 -3354 583 -3317
rect 636 -3317 805 -3301
rect 636 -3354 646 -3317
rect -49 -3509 -39 -3456
rect 14 -3509 24 -3456
rect 307 -3509 317 -3456
rect 370 -3509 380 -3456
rect -140 -3691 -64 -3675
rect -140 -3725 -124 -3691
rect -80 -3725 -64 -3691
rect -140 -3731 -64 -3725
rect -30 -3772 4 -3509
rect 589 -3598 623 -3354
rect 860 -3456 894 -3152
rect 928 -3199 1004 -3193
rect 928 -3233 944 -3199
rect 988 -3233 1004 -3199
rect 928 -3249 1004 -3233
rect 1106 -3199 1182 -3193
rect 1106 -3233 1122 -3199
rect 1166 -3233 1182 -3199
rect 1106 -3249 1182 -3233
rect 1216 -3456 1250 -3152
rect 1284 -3199 1360 -3193
rect 1284 -3233 1300 -3199
rect 1344 -3233 1360 -3199
rect 1284 -3249 1360 -3233
rect 840 -3509 850 -3456
rect 903 -3509 913 -3456
rect 1196 -3509 1206 -3456
rect 1259 -3509 1269 -3456
rect 59 -3632 1160 -3598
rect 59 -3675 93 -3632
rect 149 -3633 271 -3632
rect 38 -3691 114 -3675
rect 38 -3725 54 -3691
rect 98 -3725 114 -3691
rect 38 -3731 114 -3725
rect 149 -3772 183 -3633
rect 237 -3675 271 -3633
rect 948 -3675 982 -3632
rect 216 -3691 292 -3675
rect 216 -3725 232 -3691
rect 276 -3725 292 -3691
rect 216 -3731 292 -3725
rect 394 -3691 470 -3675
rect 394 -3725 410 -3691
rect 454 -3725 470 -3691
rect 394 -3731 470 -3725
rect 572 -3691 648 -3675
rect 572 -3725 588 -3691
rect 632 -3725 648 -3691
rect 572 -3731 648 -3725
rect 750 -3691 826 -3675
rect 750 -3725 766 -3691
rect 810 -3725 826 -3691
rect 750 -3731 826 -3725
rect 928 -3691 1004 -3675
rect 928 -3725 944 -3691
rect 988 -3725 1004 -3691
rect 928 -3731 1004 -3725
rect 1038 -3772 1072 -3632
rect 1126 -3675 1160 -3632
rect 1106 -3691 1182 -3675
rect 1106 -3725 1122 -3691
rect 1166 -3725 1182 -3691
rect 1106 -3731 1182 -3725
rect 1216 -3772 1250 -3509
rect 1306 -3675 1340 -3249
rect 1394 -3564 1428 -3152
rect 1462 -3199 1538 -3193
rect 1462 -3233 1478 -3199
rect 1522 -3233 1538 -3199
rect 1462 -3249 1538 -3233
rect 1482 -3283 1516 -3249
rect 1572 -3283 1606 -3152
rect 1640 -3199 1716 -3193
rect 1640 -3233 1656 -3199
rect 1700 -3233 1716 -3199
rect 1640 -3249 1716 -3233
rect 1662 -3283 1696 -3249
rect 1750 -3283 1784 -3152
rect 1818 -3199 1894 -3193
rect 1818 -3233 1834 -3199
rect 1878 -3233 1894 -3199
rect 1818 -3249 1894 -3233
rect 1996 -3199 2072 -3193
rect 1996 -3233 2012 -3199
rect 2056 -3233 2072 -3199
rect 1996 -3249 2072 -3233
rect 2174 -3199 2250 -3193
rect 2174 -3233 2190 -3199
rect 2234 -3233 2250 -3199
rect 2174 -3249 2250 -3233
rect 2352 -3199 2428 -3193
rect 2352 -3233 2368 -3199
rect 2412 -3233 2428 -3199
rect 2352 -3249 2428 -3233
rect 1840 -3283 1874 -3249
rect 1482 -3301 1874 -3283
rect 1482 -3317 1654 -3301
rect 1644 -3354 1654 -3317
rect 1707 -3317 1874 -3301
rect 1707 -3354 1717 -3317
rect 1552 -3509 1562 -3456
rect 1615 -3509 1625 -3456
rect 1909 -3509 1919 -3456
rect 1972 -3509 1982 -3456
rect 1374 -3617 1384 -3564
rect 1437 -3617 1447 -3564
rect 1284 -3691 1360 -3675
rect 1284 -3725 1300 -3691
rect 1344 -3725 1360 -3691
rect 1284 -3731 1360 -3725
rect 1394 -3772 1428 -3617
rect 1462 -3691 1538 -3675
rect 1462 -3725 1478 -3691
rect 1522 -3725 1538 -3691
rect 1462 -3731 1538 -3725
rect 1572 -3772 1606 -3509
rect 1731 -3617 1741 -3564
rect 1794 -3617 1804 -3564
rect 1640 -3691 1716 -3675
rect 1640 -3725 1656 -3691
rect 1700 -3725 1716 -3691
rect 1640 -3731 1716 -3725
rect 1750 -3772 1784 -3617
rect 1818 -3691 1894 -3675
rect 1818 -3725 1834 -3691
rect 1878 -3725 1894 -3691
rect 1818 -3731 1894 -3725
rect 1929 -3772 1963 -3509
rect 2017 -3675 2051 -3249
rect 2087 -3617 2097 -3564
rect 2150 -3617 2160 -3564
rect 1996 -3691 2072 -3675
rect 1996 -3725 2012 -3691
rect 2056 -3725 2072 -3691
rect 1996 -3731 2072 -3725
rect 2106 -3772 2140 -3617
rect 2196 -3675 2230 -3249
rect 2265 -3509 2275 -3456
rect 2328 -3509 2338 -3456
rect 2174 -3691 2250 -3675
rect 2174 -3725 2190 -3691
rect 2234 -3725 2250 -3691
rect 2174 -3731 2250 -3725
rect 2284 -3772 2318 -3509
rect 2373 -3675 2407 -3249
rect 2462 -3284 2496 -3152
rect 2530 -3199 2606 -3193
rect 2530 -3233 2546 -3199
rect 2590 -3233 2606 -3199
rect 2530 -3249 2606 -3233
rect 2551 -3284 2585 -3249
rect 2641 -3284 2675 -3152
rect 2462 -3318 2675 -3284
rect 2441 -3617 2451 -3564
rect 2504 -3617 2514 -3564
rect 2352 -3691 2428 -3675
rect 2352 -3725 2368 -3691
rect 2412 -3725 2428 -3691
rect 2352 -3731 2428 -3725
rect 2462 -3772 2496 -3617
rect 2530 -3691 2606 -3675
rect 2530 -3725 2546 -3691
rect 2590 -3725 2606 -3691
rect 2530 -3731 2606 -3725
rect -1460 -3784 -1414 -3772
rect -1460 -4040 -1454 -3784
rect -1420 -4040 -1414 -3784
rect -1460 -4052 -1414 -4040
rect -1282 -3784 -1236 -3772
rect -1282 -4040 -1276 -3784
rect -1242 -4040 -1236 -3784
rect -1282 -4052 -1236 -4040
rect -1104 -3784 -1058 -3772
rect -1104 -4040 -1098 -3784
rect -1064 -4040 -1058 -3784
rect -1104 -4052 -1058 -4040
rect -926 -3784 -880 -3772
rect -926 -4040 -920 -3784
rect -886 -4040 -880 -3784
rect -926 -4052 -880 -4040
rect -748 -3784 -702 -3772
rect -748 -4040 -742 -3784
rect -708 -4040 -702 -3784
rect -748 -4052 -702 -4040
rect -570 -3784 -524 -3772
rect -570 -4040 -564 -3784
rect -530 -4040 -524 -3784
rect -570 -4052 -524 -4040
rect -392 -3784 -346 -3772
rect -392 -4040 -386 -3784
rect -352 -4040 -346 -3784
rect -392 -4052 -346 -4040
rect -214 -3784 -168 -3772
rect -214 -4040 -208 -3784
rect -174 -4040 -168 -3784
rect -214 -4052 -168 -4040
rect -36 -3784 10 -3772
rect -36 -4040 -30 -3784
rect 4 -4040 10 -3784
rect -36 -4052 10 -4040
rect 142 -3784 188 -3772
rect 142 -4040 148 -3784
rect 182 -4040 188 -3784
rect 142 -4052 188 -4040
rect 320 -3784 366 -3772
rect 320 -4040 326 -3784
rect 360 -4040 366 -3784
rect 320 -4052 366 -4040
rect 498 -3784 544 -3772
rect 498 -4040 504 -3784
rect 538 -4040 544 -3784
rect 498 -4052 544 -4040
rect 676 -3784 722 -3772
rect 676 -4040 682 -3784
rect 716 -4040 722 -3784
rect 676 -4052 722 -4040
rect 854 -3784 900 -3772
rect 854 -4040 860 -3784
rect 894 -4040 900 -3784
rect 854 -4052 900 -4040
rect 1032 -3784 1078 -3772
rect 1032 -4040 1038 -3784
rect 1072 -4040 1078 -3784
rect 1032 -4052 1078 -4040
rect 1210 -3784 1256 -3772
rect 1210 -4040 1216 -3784
rect 1250 -4040 1256 -3784
rect 1210 -4052 1256 -4040
rect 1388 -3784 1434 -3772
rect 1388 -4040 1394 -3784
rect 1428 -4040 1434 -3784
rect 1388 -4052 1434 -4040
rect 1566 -3784 1612 -3772
rect 1566 -4040 1572 -3784
rect 1606 -4040 1612 -3784
rect 1566 -4052 1612 -4040
rect 1744 -3784 1790 -3772
rect 1744 -4040 1750 -3784
rect 1784 -4040 1790 -3784
rect 1744 -4052 1790 -4040
rect 1922 -3784 1968 -3772
rect 1922 -4040 1928 -3784
rect 1962 -4040 1968 -3784
rect 1922 -4052 1968 -4040
rect 2100 -3784 2146 -3772
rect 2100 -4040 2106 -3784
rect 2140 -4040 2146 -3784
rect 2100 -4052 2146 -4040
rect 2278 -3784 2324 -3772
rect 2278 -4040 2284 -3784
rect 2318 -4040 2324 -3784
rect 2278 -4052 2324 -4040
rect 2456 -3784 2502 -3772
rect 2456 -4040 2462 -3784
rect 2496 -4040 2502 -3784
rect 2456 -4052 2502 -4040
rect 2634 -3784 2680 -3772
rect 2634 -4040 2640 -3784
rect 2674 -4040 2680 -3784
rect 2634 -4052 2680 -4040
rect -1454 -4184 -1420 -4052
rect -1386 -4099 -1310 -4093
rect -1386 -4133 -1370 -4099
rect -1326 -4133 -1310 -4099
rect -1386 -4149 -1310 -4133
rect -1366 -4184 -1332 -4149
rect -1276 -4184 -1242 -4052
rect -1208 -4099 -1132 -4093
rect -1208 -4133 -1192 -4099
rect -1148 -4133 -1132 -4099
rect -1208 -4149 -1132 -4133
rect -1030 -4099 -954 -4093
rect -1030 -4133 -1014 -4099
rect -970 -4133 -954 -4099
rect -1030 -4149 -954 -4133
rect -852 -4099 -776 -4093
rect -852 -4133 -836 -4099
rect -792 -4133 -776 -4099
rect -852 -4149 -776 -4133
rect -674 -4099 -598 -4093
rect -674 -4133 -658 -4099
rect -614 -4133 -598 -4099
rect -674 -4149 -598 -4133
rect -496 -4099 -420 -4093
rect -496 -4133 -480 -4099
rect -436 -4133 -420 -4099
rect -496 -4149 -420 -4133
rect -318 -4099 -242 -4093
rect -318 -4133 -302 -4099
rect -258 -4133 -242 -4099
rect -318 -4149 -242 -4133
rect -140 -4099 -64 -4093
rect -140 -4133 -124 -4099
rect -80 -4133 -64 -4099
rect -140 -4149 -64 -4133
rect 38 -4099 114 -4093
rect 38 -4133 54 -4099
rect 98 -4133 114 -4099
rect 38 -4149 114 -4133
rect -1454 -4218 -1242 -4184
rect -1454 -4541 -1242 -4507
rect -1454 -4672 -1420 -4541
rect -1365 -4575 -1331 -4541
rect -1386 -4591 -1310 -4575
rect -1386 -4625 -1370 -4591
rect -1326 -4625 -1310 -4591
rect -1386 -4631 -1310 -4625
rect -1276 -4672 -1242 -4541
rect -1187 -4575 -1153 -4149
rect -1009 -4575 -975 -4149
rect -831 -4192 -797 -4149
rect -653 -4192 -619 -4149
rect -474 -4192 -440 -4149
rect -297 -4192 -263 -4149
rect -851 -4245 -841 -4192
rect -788 -4245 -778 -4192
rect -672 -4245 -662 -4192
rect -609 -4245 -599 -4192
rect -493 -4245 -483 -4192
rect -430 -4245 -420 -4192
rect -316 -4245 -306 -4192
rect -253 -4245 -243 -4192
rect -831 -4575 -797 -4245
rect -653 -4575 -619 -4245
rect -474 -4575 -440 -4245
rect -297 -4575 -263 -4245
rect -119 -4575 -85 -4149
rect -1208 -4591 -1132 -4575
rect -1208 -4625 -1192 -4591
rect -1148 -4625 -1132 -4591
rect -1208 -4631 -1132 -4625
rect -1030 -4591 -954 -4575
rect -1030 -4625 -1014 -4591
rect -970 -4625 -954 -4591
rect -1030 -4631 -954 -4625
rect -852 -4591 -776 -4575
rect -852 -4625 -836 -4591
rect -792 -4625 -776 -4591
rect -852 -4631 -776 -4625
rect -674 -4591 -598 -4575
rect -674 -4625 -658 -4591
rect -614 -4625 -598 -4591
rect -674 -4631 -598 -4625
rect -496 -4591 -420 -4575
rect -496 -4625 -480 -4591
rect -436 -4625 -420 -4591
rect -496 -4631 -420 -4625
rect -318 -4591 -242 -4575
rect -318 -4625 -302 -4591
rect -258 -4625 -242 -4591
rect -318 -4631 -242 -4625
rect -140 -4591 -64 -4575
rect -140 -4625 -124 -4591
rect -80 -4625 -64 -4591
rect -140 -4631 -64 -4625
rect 38 -4591 114 -4575
rect 38 -4625 54 -4591
rect 98 -4625 114 -4591
rect 38 -4631 114 -4625
rect 148 -4672 182 -4052
rect 216 -4099 292 -4093
rect 216 -4133 232 -4099
rect 276 -4133 292 -4099
rect 216 -4149 292 -4133
rect 326 -4304 360 -4052
rect 394 -4099 470 -4093
rect 394 -4133 410 -4099
rect 454 -4133 470 -4099
rect 394 -4149 470 -4133
rect 416 -4192 450 -4149
rect 397 -4245 407 -4192
rect 460 -4245 470 -4192
rect 307 -4357 317 -4304
rect 370 -4357 380 -4304
rect 216 -4591 292 -4575
rect 216 -4625 232 -4591
rect 276 -4625 292 -4591
rect 216 -4631 292 -4625
rect 326 -4672 360 -4357
rect 416 -4575 450 -4245
rect 504 -4412 538 -4052
rect 572 -4099 648 -4093
rect 572 -4133 588 -4099
rect 632 -4133 648 -4099
rect 572 -4149 648 -4133
rect 593 -4192 627 -4149
rect 573 -4245 583 -4192
rect 636 -4245 646 -4192
rect 485 -4465 495 -4412
rect 548 -4465 558 -4412
rect 394 -4591 470 -4575
rect 394 -4625 410 -4591
rect 454 -4625 470 -4591
rect 394 -4631 470 -4625
rect 504 -4672 538 -4465
rect 593 -4575 627 -4245
rect 682 -4304 716 -4052
rect 750 -4099 826 -4093
rect 750 -4133 766 -4099
rect 810 -4133 826 -4099
rect 750 -4149 826 -4133
rect 771 -4192 805 -4149
rect 751 -4245 761 -4192
rect 814 -4245 824 -4192
rect 663 -4357 673 -4304
rect 726 -4357 736 -4304
rect 572 -4591 648 -4575
rect 572 -4625 588 -4591
rect 632 -4625 648 -4591
rect 572 -4631 648 -4625
rect 682 -4672 716 -4357
rect 771 -4575 805 -4245
rect 860 -4412 894 -4052
rect 928 -4099 1004 -4093
rect 928 -4133 944 -4099
rect 988 -4133 1004 -4099
rect 928 -4149 1004 -4133
rect 840 -4465 850 -4412
rect 903 -4465 913 -4412
rect 750 -4591 826 -4575
rect 750 -4625 766 -4591
rect 810 -4625 826 -4591
rect 750 -4631 826 -4625
rect 860 -4672 894 -4465
rect 928 -4591 1004 -4575
rect 928 -4625 944 -4591
rect 988 -4625 1004 -4591
rect 928 -4631 1004 -4625
rect 1039 -4672 1073 -4052
rect 1106 -4099 1182 -4093
rect 1106 -4133 1122 -4099
rect 1166 -4133 1182 -4099
rect 1106 -4149 1182 -4133
rect 1284 -4099 1360 -4093
rect 1284 -4133 1300 -4099
rect 1344 -4133 1360 -4099
rect 1284 -4149 1360 -4133
rect 1462 -4099 1538 -4093
rect 1462 -4133 1478 -4099
rect 1522 -4133 1538 -4099
rect 1462 -4149 1538 -4133
rect 1640 -4099 1716 -4093
rect 1640 -4133 1656 -4099
rect 1700 -4133 1716 -4099
rect 1640 -4149 1716 -4133
rect 1818 -4099 1894 -4093
rect 1818 -4133 1834 -4099
rect 1878 -4133 1894 -4099
rect 1818 -4149 1894 -4133
rect 1996 -4099 2072 -4093
rect 1996 -4133 2012 -4099
rect 2056 -4133 2072 -4099
rect 1996 -4149 2072 -4133
rect 2174 -4099 2250 -4093
rect 2174 -4133 2190 -4099
rect 2234 -4133 2250 -4099
rect 2174 -4149 2250 -4133
rect 2352 -4099 2428 -4093
rect 2352 -4133 2368 -4099
rect 2412 -4133 2428 -4099
rect 2352 -4149 2428 -4133
rect 1305 -4575 1339 -4149
rect 1484 -4192 1518 -4149
rect 1661 -4192 1695 -4149
rect 1839 -4192 1873 -4149
rect 2017 -4192 2051 -4149
rect 1464 -4245 1474 -4192
rect 1527 -4245 1537 -4192
rect 1642 -4245 1652 -4192
rect 1705 -4245 1715 -4192
rect 1820 -4245 1830 -4192
rect 1883 -4245 1893 -4192
rect 1998 -4245 2008 -4192
rect 2061 -4245 2071 -4192
rect 1484 -4575 1518 -4245
rect 1661 -4575 1695 -4245
rect 1839 -4575 1873 -4245
rect 2017 -4575 2051 -4245
rect 2195 -4575 2229 -4149
rect 2373 -4575 2407 -4149
rect 2463 -4182 2497 -4052
rect 2530 -4099 2606 -4093
rect 2530 -4133 2546 -4099
rect 2590 -4133 2606 -4099
rect 2530 -4149 2606 -4133
rect 2552 -4182 2586 -4149
rect 2640 -4180 2674 -4052
rect 2640 -4182 2792 -4180
rect 2463 -4214 2792 -4182
rect 2463 -4216 2674 -4214
rect 2528 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect 2550 -4506 2584 -4327
rect 2758 -4446 2792 -4214
rect 2462 -4540 2674 -4506
rect 2736 -4507 2746 -4446
rect 2807 -4507 2817 -4446
rect 2758 -4508 2792 -4507
rect 1106 -4591 1182 -4575
rect 1106 -4625 1122 -4591
rect 1166 -4625 1182 -4591
rect 1106 -4631 1182 -4625
rect 1284 -4591 1360 -4575
rect 1284 -4625 1300 -4591
rect 1344 -4625 1360 -4591
rect 1284 -4631 1360 -4625
rect 1462 -4591 1538 -4575
rect 1462 -4625 1478 -4591
rect 1522 -4625 1538 -4591
rect 1462 -4631 1538 -4625
rect 1640 -4591 1716 -4575
rect 1640 -4625 1656 -4591
rect 1700 -4625 1716 -4591
rect 1640 -4631 1716 -4625
rect 1818 -4591 1894 -4575
rect 1818 -4625 1834 -4591
rect 1878 -4625 1894 -4591
rect 1818 -4631 1894 -4625
rect 1996 -4591 2072 -4575
rect 1996 -4625 2012 -4591
rect 2056 -4625 2072 -4591
rect 1996 -4631 2072 -4625
rect 2174 -4591 2250 -4575
rect 2174 -4625 2190 -4591
rect 2234 -4625 2250 -4591
rect 2174 -4631 2250 -4625
rect 2352 -4591 2428 -4575
rect 2352 -4625 2368 -4591
rect 2412 -4625 2428 -4591
rect 2352 -4631 2428 -4625
rect 2462 -4672 2496 -4540
rect 2550 -4575 2584 -4540
rect 2530 -4591 2606 -4575
rect 2530 -4625 2546 -4591
rect 2590 -4625 2606 -4591
rect 2530 -4631 2606 -4625
rect 2640 -4672 2674 -4540
rect -1460 -4684 -1414 -4672
rect -1460 -4940 -1454 -4684
rect -1420 -4940 -1414 -4684
rect -1460 -4952 -1414 -4940
rect -1282 -4684 -1236 -4672
rect -1282 -4940 -1276 -4684
rect -1242 -4940 -1236 -4684
rect -1282 -4952 -1236 -4940
rect -1104 -4684 -1058 -4672
rect -1104 -4940 -1098 -4684
rect -1064 -4940 -1058 -4684
rect -1104 -4952 -1058 -4940
rect -926 -4684 -880 -4672
rect -926 -4940 -920 -4684
rect -886 -4940 -880 -4684
rect -926 -4952 -880 -4940
rect -748 -4684 -702 -4672
rect -748 -4940 -742 -4684
rect -708 -4940 -702 -4684
rect -748 -4952 -702 -4940
rect -570 -4684 -524 -4672
rect -570 -4940 -564 -4684
rect -530 -4940 -524 -4684
rect -570 -4952 -524 -4940
rect -392 -4684 -346 -4672
rect -392 -4940 -386 -4684
rect -352 -4940 -346 -4684
rect -392 -4952 -346 -4940
rect -214 -4684 -168 -4672
rect -214 -4940 -208 -4684
rect -174 -4940 -168 -4684
rect -214 -4952 -168 -4940
rect -36 -4684 10 -4672
rect -36 -4940 -30 -4684
rect 4 -4940 10 -4684
rect -36 -4952 10 -4940
rect 142 -4684 188 -4672
rect 142 -4940 148 -4684
rect 182 -4940 188 -4684
rect 142 -4952 188 -4940
rect 320 -4684 366 -4672
rect 320 -4940 326 -4684
rect 360 -4940 366 -4684
rect 320 -4952 366 -4940
rect 498 -4684 544 -4672
rect 498 -4940 504 -4684
rect 538 -4940 544 -4684
rect 498 -4952 544 -4940
rect 676 -4684 722 -4672
rect 676 -4940 682 -4684
rect 716 -4940 722 -4684
rect 676 -4952 722 -4940
rect 854 -4684 900 -4672
rect 854 -4940 860 -4684
rect 894 -4940 900 -4684
rect 854 -4952 900 -4940
rect 1032 -4684 1078 -4672
rect 1032 -4940 1038 -4684
rect 1072 -4940 1078 -4684
rect 1032 -4952 1078 -4940
rect 1210 -4684 1256 -4672
rect 1210 -4940 1216 -4684
rect 1250 -4940 1256 -4684
rect 1210 -4952 1256 -4940
rect 1388 -4684 1434 -4672
rect 1388 -4940 1394 -4684
rect 1428 -4940 1434 -4684
rect 1388 -4952 1434 -4940
rect 1566 -4684 1612 -4672
rect 1566 -4940 1572 -4684
rect 1606 -4940 1612 -4684
rect 1566 -4952 1612 -4940
rect 1744 -4684 1790 -4672
rect 1744 -4940 1750 -4684
rect 1784 -4940 1790 -4684
rect 1744 -4952 1790 -4940
rect 1922 -4684 1968 -4672
rect 1922 -4940 1928 -4684
rect 1962 -4940 1968 -4684
rect 1922 -4952 1968 -4940
rect 2100 -4684 2146 -4672
rect 2100 -4940 2106 -4684
rect 2140 -4940 2146 -4684
rect 2100 -4952 2146 -4940
rect 2278 -4684 2324 -4672
rect 2278 -4940 2284 -4684
rect 2318 -4940 2324 -4684
rect 2278 -4952 2324 -4940
rect 2456 -4684 2502 -4672
rect 2456 -4940 2462 -4684
rect 2496 -4940 2502 -4684
rect 2456 -4952 2502 -4940
rect 2634 -4684 2680 -4672
rect 2634 -4940 2640 -4684
rect 2674 -4940 2680 -4684
rect 2634 -4952 2680 -4940
rect -1386 -4999 -1310 -4993
rect -1386 -5033 -1370 -4999
rect -1326 -5033 -1310 -4999
rect -1386 -5049 -1310 -5033
rect -1277 -5097 -1243 -4952
rect -1208 -4999 -1132 -4993
rect -1208 -5033 -1192 -4999
rect -1148 -5033 -1132 -4999
rect -1208 -5049 -1132 -5033
rect -1297 -5150 -1287 -5097
rect -1234 -5150 -1224 -5097
rect -1876 -5337 -1823 -5285
rect -1875 -6364 -1823 -5337
rect -1656 -5339 -1646 -5278
rect -1585 -5339 -1575 -5278
rect -1454 -5442 -1242 -5408
rect -1454 -5572 -1420 -5442
rect -1363 -5475 -1329 -5442
rect -1386 -5491 -1310 -5475
rect -1386 -5525 -1370 -5491
rect -1326 -5525 -1310 -5491
rect -1386 -5531 -1310 -5525
rect -1276 -5572 -1242 -5442
rect -1187 -5475 -1153 -5049
rect -1097 -5213 -1063 -4952
rect -1030 -4999 -954 -4993
rect -1030 -5033 -1014 -4999
rect -970 -5033 -954 -4999
rect -1030 -5049 -954 -5033
rect -1115 -5266 -1105 -5213
rect -1052 -5266 -1042 -5213
rect -1009 -5475 -975 -5049
rect -919 -5097 -885 -4952
rect -852 -4999 -776 -4993
rect -852 -5033 -836 -4999
rect -792 -5033 -776 -4999
rect -852 -5049 -776 -5033
rect -939 -5150 -929 -5097
rect -876 -5150 -866 -5097
rect -830 -5475 -796 -5049
rect -741 -5213 -707 -4952
rect -674 -4999 -598 -4993
rect -674 -5033 -658 -4999
rect -614 -5033 -598 -4999
rect -674 -5049 -598 -5033
rect -563 -5097 -529 -4952
rect -496 -4999 -420 -4993
rect -496 -5033 -480 -4999
rect -436 -5033 -420 -4999
rect -496 -5049 -420 -5033
rect -582 -5150 -572 -5097
rect -519 -5150 -509 -5097
rect -386 -5213 -352 -4952
rect -318 -4999 -242 -4993
rect -318 -5033 -302 -4999
rect -258 -5033 -242 -4999
rect -318 -5049 -242 -5033
rect -208 -5097 -174 -4952
rect -140 -4999 -64 -4993
rect -140 -5033 -124 -4999
rect -80 -5033 -64 -4999
rect -140 -5049 -64 -5033
rect -228 -5150 -218 -5097
rect -165 -5150 -155 -5097
rect -761 -5266 -751 -5213
rect -698 -5266 -688 -5213
rect -406 -5266 -396 -5213
rect -343 -5266 -333 -5213
rect -654 -5434 -262 -5400
rect -654 -5475 -620 -5434
rect -1208 -5491 -1132 -5475
rect -1208 -5525 -1192 -5491
rect -1148 -5525 -1132 -5491
rect -1208 -5531 -1132 -5525
rect -1030 -5491 -954 -5475
rect -1030 -5525 -1014 -5491
rect -970 -5525 -954 -5491
rect -1030 -5531 -954 -5525
rect -852 -5491 -776 -5475
rect -852 -5525 -836 -5491
rect -792 -5525 -776 -5491
rect -852 -5531 -776 -5525
rect -674 -5491 -598 -5475
rect -674 -5525 -658 -5491
rect -614 -5525 -598 -5491
rect -674 -5531 -598 -5525
rect -563 -5572 -529 -5434
rect -474 -5475 -440 -5434
rect -496 -5491 -420 -5475
rect -496 -5525 -480 -5491
rect -436 -5525 -420 -5491
rect -496 -5531 -420 -5525
rect -385 -5572 -351 -5434
rect -296 -5475 -262 -5434
rect -318 -5491 -242 -5475
rect -318 -5525 -302 -5491
rect -258 -5525 -242 -5491
rect -318 -5531 -242 -5525
rect -208 -5572 -174 -5150
rect -119 -5380 -85 -5049
rect -30 -5213 4 -4952
rect 59 -4993 93 -4992
rect 38 -4999 114 -4993
rect 38 -5033 54 -4999
rect 98 -5033 114 -4999
rect 38 -5049 114 -5033
rect 59 -5091 93 -5049
rect 148 -5091 182 -4952
rect 216 -4999 292 -4993
rect 216 -5033 232 -4999
rect 276 -5033 292 -4999
rect 216 -5049 292 -5033
rect 394 -4999 470 -4993
rect 394 -5033 410 -4999
rect 454 -5033 470 -4999
rect 394 -5049 470 -5033
rect 572 -4999 648 -4993
rect 572 -5033 588 -4999
rect 632 -5033 648 -4999
rect 572 -5049 648 -5033
rect 750 -4999 826 -4993
rect 750 -5033 766 -4999
rect 810 -5033 826 -4999
rect 750 -5049 826 -5033
rect 928 -4999 1004 -4993
rect 928 -5033 944 -4999
rect 988 -5033 1004 -4999
rect 928 -5049 1004 -5033
rect 236 -5091 270 -5049
rect 948 -5091 982 -5049
rect 1039 -5091 1073 -4952
rect 1106 -4999 1182 -4993
rect 1106 -5033 1122 -4999
rect 1166 -5033 1182 -4999
rect 1106 -5049 1182 -5033
rect 1128 -5091 1162 -5049
rect 59 -5125 1162 -5091
rect -51 -5266 -41 -5213
rect 12 -5266 22 -5213
rect 306 -5266 316 -5213
rect 369 -5266 379 -5213
rect -138 -5433 -128 -5380
rect -75 -5433 -65 -5380
rect -119 -5475 -85 -5433
rect -140 -5491 -64 -5475
rect -140 -5525 -124 -5491
rect -80 -5525 -64 -5491
rect -140 -5531 -64 -5525
rect -30 -5572 4 -5266
rect 40 -5433 50 -5380
rect 103 -5433 113 -5380
rect 218 -5433 228 -5380
rect 281 -5433 291 -5380
rect 59 -5475 93 -5433
rect 238 -5475 272 -5433
rect 38 -5491 114 -5475
rect 38 -5525 54 -5491
rect 98 -5525 114 -5491
rect 38 -5531 114 -5525
rect 216 -5491 292 -5475
rect 216 -5525 232 -5491
rect 276 -5525 292 -5491
rect 216 -5531 292 -5525
rect 326 -5572 360 -5266
rect 593 -5315 627 -5125
rect 1216 -5213 1250 -4952
rect 1284 -4999 1360 -4993
rect 1284 -5033 1300 -4999
rect 1344 -5033 1360 -4999
rect 1284 -5049 1360 -5033
rect 840 -5266 850 -5213
rect 903 -5266 913 -5213
rect 1197 -5266 1207 -5213
rect 1260 -5266 1270 -5213
rect 415 -5349 804 -5315
rect 415 -5475 449 -5349
rect 394 -5491 470 -5475
rect 394 -5525 410 -5491
rect 454 -5525 470 -5491
rect 394 -5531 470 -5525
rect 505 -5572 539 -5349
rect 592 -5475 626 -5349
rect 572 -5491 648 -5475
rect 572 -5525 588 -5491
rect 632 -5525 648 -5491
rect 572 -5531 648 -5525
rect 681 -5572 715 -5349
rect 770 -5475 804 -5349
rect 750 -5491 826 -5475
rect 750 -5525 766 -5491
rect 810 -5525 826 -5491
rect 750 -5531 826 -5525
rect 860 -5572 894 -5266
rect 930 -5434 940 -5381
rect 993 -5434 1003 -5381
rect 1109 -5433 1119 -5380
rect 1172 -5433 1182 -5380
rect 949 -5475 983 -5434
rect 1128 -5475 1162 -5433
rect 928 -5491 1004 -5475
rect 928 -5525 944 -5491
rect 988 -5525 1004 -5491
rect 928 -5531 1004 -5525
rect 1106 -5491 1182 -5475
rect 1106 -5525 1122 -5491
rect 1166 -5525 1182 -5491
rect 1106 -5531 1182 -5525
rect 1216 -5572 1250 -5266
rect 1306 -5380 1340 -5049
rect 1394 -5093 1428 -4952
rect 1462 -4999 1538 -4993
rect 1462 -5033 1478 -4999
rect 1522 -5033 1538 -4999
rect 1462 -5049 1538 -5033
rect 1375 -5146 1385 -5093
rect 1438 -5146 1448 -5093
rect 1286 -5433 1296 -5380
rect 1349 -5433 1359 -5380
rect 1306 -5475 1340 -5433
rect 1284 -5491 1360 -5475
rect 1284 -5525 1300 -5491
rect 1344 -5525 1360 -5491
rect 1284 -5531 1360 -5525
rect 1394 -5572 1428 -5146
rect 1572 -5213 1606 -4952
rect 1640 -4999 1716 -4993
rect 1640 -5033 1656 -4999
rect 1700 -5033 1716 -4999
rect 1640 -5049 1716 -5033
rect 1750 -5093 1784 -4952
rect 1818 -4999 1894 -4993
rect 1818 -5033 1834 -4999
rect 1878 -5033 1894 -4999
rect 1818 -5049 1894 -5033
rect 1730 -5146 1740 -5093
rect 1793 -5146 1803 -5093
rect 1927 -5213 1961 -4952
rect 1996 -4999 2072 -4993
rect 1996 -5033 2012 -4999
rect 2056 -5033 2072 -4999
rect 1996 -5049 2072 -5033
rect 1553 -5266 1563 -5213
rect 1616 -5266 1626 -5213
rect 1907 -5266 1917 -5213
rect 1970 -5266 1980 -5213
rect 1482 -5433 1874 -5399
rect 1482 -5475 1516 -5433
rect 1462 -5491 1538 -5475
rect 1462 -5525 1478 -5491
rect 1522 -5525 1538 -5491
rect 1462 -5531 1538 -5525
rect 1573 -5572 1607 -5433
rect 1661 -5475 1695 -5433
rect 1640 -5491 1716 -5475
rect 1640 -5525 1656 -5491
rect 1700 -5525 1716 -5491
rect 1640 -5531 1716 -5525
rect 1749 -5572 1783 -5433
rect 1840 -5475 1874 -5433
rect 2018 -5475 2052 -5049
rect 2106 -5093 2140 -4952
rect 2174 -4999 2250 -4993
rect 2174 -5033 2190 -4999
rect 2234 -5033 2250 -4999
rect 2174 -5049 2250 -5033
rect 2086 -5146 2096 -5093
rect 2149 -5146 2159 -5093
rect 2195 -5475 2229 -5049
rect 2284 -5213 2318 -4952
rect 2352 -4999 2428 -4993
rect 2352 -5033 2368 -4999
rect 2412 -5033 2428 -4999
rect 2352 -5049 2428 -5033
rect 2264 -5266 2274 -5213
rect 2327 -5266 2337 -5213
rect 2373 -5475 2407 -5049
rect 2462 -5093 2496 -4952
rect 2530 -4999 2606 -4993
rect 2530 -5033 2546 -4999
rect 2590 -5033 2606 -4999
rect 2530 -5049 2606 -5033
rect 2443 -5146 2453 -5093
rect 2506 -5146 2516 -5093
rect 2463 -5442 2674 -5408
rect 1818 -5491 1894 -5475
rect 1818 -5525 1834 -5491
rect 1878 -5525 1894 -5491
rect 1818 -5531 1894 -5525
rect 1996 -5491 2072 -5475
rect 1996 -5525 2012 -5491
rect 2056 -5525 2072 -5491
rect 1996 -5531 2072 -5525
rect 2174 -5491 2250 -5475
rect 2174 -5525 2190 -5491
rect 2234 -5525 2250 -5491
rect 2174 -5531 2250 -5525
rect 2352 -5491 2428 -5475
rect 2352 -5525 2368 -5491
rect 2412 -5525 2428 -5491
rect 2352 -5531 2428 -5525
rect 2463 -5572 2497 -5442
rect 2550 -5475 2584 -5442
rect 2530 -5491 2606 -5475
rect 2530 -5525 2546 -5491
rect 2590 -5525 2606 -5491
rect 2530 -5531 2606 -5525
rect 2640 -5572 2674 -5442
rect -1460 -5584 -1414 -5572
rect -1460 -5840 -1454 -5584
rect -1420 -5840 -1414 -5584
rect -1460 -5852 -1414 -5840
rect -1282 -5584 -1236 -5572
rect -1282 -5840 -1276 -5584
rect -1242 -5840 -1236 -5584
rect -1282 -5852 -1236 -5840
rect -1104 -5584 -1058 -5572
rect -1104 -5840 -1098 -5584
rect -1064 -5840 -1058 -5584
rect -1104 -5852 -1058 -5840
rect -926 -5584 -880 -5572
rect -926 -5840 -920 -5584
rect -886 -5840 -880 -5584
rect -926 -5852 -880 -5840
rect -748 -5584 -702 -5572
rect -748 -5840 -742 -5584
rect -708 -5840 -702 -5584
rect -748 -5852 -702 -5840
rect -570 -5584 -524 -5572
rect -570 -5840 -564 -5584
rect -530 -5840 -524 -5584
rect -570 -5852 -524 -5840
rect -392 -5584 -346 -5572
rect -392 -5840 -386 -5584
rect -352 -5840 -346 -5584
rect -392 -5852 -346 -5840
rect -214 -5584 -168 -5572
rect -214 -5840 -208 -5584
rect -174 -5840 -168 -5584
rect -214 -5852 -168 -5840
rect -36 -5584 10 -5572
rect -36 -5840 -30 -5584
rect 4 -5840 10 -5584
rect -36 -5852 10 -5840
rect 142 -5584 188 -5572
rect 142 -5840 148 -5584
rect 182 -5840 188 -5584
rect 142 -5852 188 -5840
rect 320 -5584 366 -5572
rect 320 -5840 326 -5584
rect 360 -5840 366 -5584
rect 320 -5852 366 -5840
rect 498 -5584 544 -5572
rect 498 -5840 504 -5584
rect 538 -5840 544 -5584
rect 498 -5852 544 -5840
rect 676 -5584 722 -5572
rect 676 -5840 682 -5584
rect 716 -5840 722 -5584
rect 676 -5852 722 -5840
rect 854 -5584 900 -5572
rect 854 -5840 860 -5584
rect 894 -5840 900 -5584
rect 854 -5852 900 -5840
rect 1032 -5584 1078 -5572
rect 1032 -5840 1038 -5584
rect 1072 -5840 1078 -5584
rect 1032 -5852 1078 -5840
rect 1210 -5584 1256 -5572
rect 1210 -5840 1216 -5584
rect 1250 -5840 1256 -5584
rect 1210 -5852 1256 -5840
rect 1388 -5584 1434 -5572
rect 1388 -5840 1394 -5584
rect 1428 -5840 1434 -5584
rect 1388 -5852 1434 -5840
rect 1566 -5584 1612 -5572
rect 1566 -5840 1572 -5584
rect 1606 -5840 1612 -5584
rect 1566 -5852 1612 -5840
rect 1744 -5584 1790 -5572
rect 1744 -5840 1750 -5584
rect 1784 -5840 1790 -5584
rect 1744 -5852 1790 -5840
rect 1922 -5584 1968 -5572
rect 1922 -5840 1928 -5584
rect 1962 -5840 1968 -5584
rect 1922 -5852 1968 -5840
rect 2100 -5584 2146 -5572
rect 2100 -5840 2106 -5584
rect 2140 -5840 2146 -5584
rect 2100 -5852 2146 -5840
rect 2278 -5584 2324 -5572
rect 2278 -5840 2284 -5584
rect 2318 -5840 2324 -5584
rect 2278 -5852 2324 -5840
rect 2456 -5584 2502 -5572
rect 2456 -5840 2462 -5584
rect 2496 -5840 2502 -5584
rect 2456 -5852 2502 -5840
rect 2634 -5584 2680 -5572
rect 2634 -5840 2640 -5584
rect 2674 -5840 2680 -5584
rect 2634 -5852 2680 -5840
rect -1386 -5899 -1310 -5893
rect -1386 -5933 -1370 -5899
rect -1326 -5933 -1310 -5899
rect -1386 -5949 -1310 -5933
rect -1274 -6364 -1240 -5852
rect -1208 -5899 -1132 -5893
rect -1208 -5933 -1192 -5899
rect -1148 -5933 -1132 -5899
rect -1208 -5949 -1132 -5933
rect -1886 -6417 -1876 -6364
rect -1823 -6417 -1813 -6364
rect -1292 -6417 -1282 -6364
rect -1229 -6417 -1219 -6364
rect -1099 -6479 -1065 -5852
rect -1030 -5899 -954 -5893
rect -1030 -5933 -1014 -5899
rect -970 -5933 -954 -5899
rect -1030 -5949 -954 -5933
rect -919 -6365 -885 -5852
rect -852 -5899 -776 -5893
rect -852 -5933 -836 -5899
rect -792 -5933 -776 -5899
rect -852 -5949 -776 -5933
rect -938 -6417 -928 -6365
rect -876 -6417 -866 -6365
rect -742 -6479 -708 -5852
rect -674 -5899 -598 -5893
rect -674 -5933 -658 -5899
rect -614 -5933 -598 -5899
rect -674 -5949 -598 -5933
rect -496 -5899 -420 -5893
rect -496 -5933 -480 -5899
rect -436 -5933 -420 -5899
rect -496 -5949 -420 -5933
rect -318 -5899 -242 -5893
rect -318 -5933 -302 -5899
rect -258 -5933 -242 -5899
rect -318 -5949 -242 -5933
rect -1120 -6532 -1110 -6479
rect -1057 -6532 -1047 -6479
rect -762 -6532 -752 -6479
rect -699 -6532 -689 -6479
rect -476 -6493 -442 -5949
rect -208 -6077 -174 -5852
rect -140 -5899 -64 -5893
rect -140 -5933 -124 -5899
rect -80 -5933 -64 -5899
rect -140 -5949 -64 -5933
rect 38 -5899 114 -5893
rect 38 -5933 54 -5899
rect 98 -5933 114 -5899
rect 38 -5949 114 -5933
rect 149 -6077 183 -5852
rect 216 -5899 292 -5893
rect 216 -5933 232 -5899
rect 276 -5933 292 -5899
rect 216 -5949 292 -5933
rect 394 -5899 470 -5893
rect 394 -5933 410 -5899
rect 454 -5933 470 -5899
rect 394 -5949 470 -5933
rect 572 -5899 648 -5893
rect 572 -5933 588 -5899
rect 632 -5933 648 -5899
rect 572 -5949 648 -5933
rect 750 -5899 826 -5893
rect 750 -5933 766 -5899
rect 810 -5933 826 -5899
rect 750 -5949 826 -5933
rect 928 -5899 1004 -5893
rect 928 -5933 944 -5899
rect 988 -5933 1004 -5899
rect 928 -5949 1004 -5933
rect -208 -6111 183 -6077
rect 237 -6250 271 -5949
rect 217 -6303 227 -6250
rect 280 -6303 290 -6250
rect 594 -6493 628 -5949
rect 951 -6250 985 -5949
rect 1038 -6081 1072 -5852
rect 1106 -5899 1182 -5893
rect 1106 -5933 1122 -5899
rect 1166 -5933 1182 -5899
rect 1106 -5949 1182 -5933
rect 1284 -5899 1360 -5893
rect 1284 -5933 1300 -5899
rect 1344 -5933 1360 -5899
rect 1284 -5949 1360 -5933
rect 1394 -6081 1428 -5852
rect 1462 -5899 1538 -5893
rect 1462 -5933 1478 -5899
rect 1522 -5933 1538 -5899
rect 1462 -5949 1538 -5933
rect 1640 -5899 1716 -5893
rect 1640 -5933 1656 -5899
rect 1700 -5933 1716 -5899
rect 1640 -5949 1716 -5933
rect 1818 -5899 1894 -5893
rect 1818 -5933 1834 -5899
rect 1878 -5933 1894 -5899
rect 1818 -5949 1894 -5933
rect 1038 -6115 1428 -6081
rect 932 -6303 942 -6250
rect 995 -6303 1005 -6250
rect 1662 -6493 1696 -5949
rect 1928 -6124 1962 -5852
rect 1996 -5899 2072 -5893
rect 1996 -5933 2012 -5899
rect 2056 -5933 2072 -5899
rect 1996 -5949 2072 -5933
rect 2106 -6007 2140 -5852
rect 2174 -5899 2250 -5893
rect 2174 -5933 2190 -5899
rect 2234 -5933 2250 -5899
rect 2174 -5949 2250 -5933
rect 2086 -6060 2096 -6007
rect 2149 -6060 2159 -6007
rect 2284 -6124 2318 -5852
rect 2352 -5899 2428 -5893
rect 2352 -5933 2368 -5899
rect 2412 -5933 2428 -5899
rect 2352 -5949 2428 -5933
rect 2462 -6007 2496 -5852
rect 2530 -5899 2606 -5893
rect 2530 -5933 2546 -5899
rect 2590 -5933 2606 -5899
rect 2530 -5949 2606 -5933
rect 2442 -6060 2452 -6007
rect 2505 -6060 2515 -6007
rect 1908 -6177 1918 -6124
rect 1971 -6177 1981 -6124
rect 2265 -6177 2275 -6124
rect 2328 -6177 2338 -6124
rect 2879 -6365 2931 -2606
rect 3194 -4805 3246 -2480
rect 3184 -4857 3194 -4805
rect 3246 -4857 3256 -4805
rect 4761 -4857 4771 -4805
rect 4823 -4857 4833 -4805
rect 2869 -6417 2879 -6365
rect 2931 -6417 2941 -6365
rect -476 -6527 1696 -6493
rect -742 -6598 -708 -6532
rect 4771 -6597 4823 -4857
rect 5027 -5059 5037 -5006
rect 5090 -5059 5100 -5006
rect 4895 -5265 4905 -5212
rect 4958 -5265 4968 -5212
rect -763 -6651 -753 -6598
rect -700 -6651 -690 -6598
rect 4762 -6650 4772 -6597
rect 4825 -6650 4835 -6597
rect -2013 -6767 -2003 -6714
rect -1950 -6767 -1940 -6714
rect 4771 -6891 4823 -6650
rect 4905 -6889 4958 -5265
rect 5037 -6887 5090 -5059
rect 5337 -5527 5390 -2258
rect 5608 -5207 5683 2178
rect 7034 2063 7080 2075
rect 7034 1863 7040 2063
rect 7074 1863 7080 2063
rect 7154 2045 7188 2178
rect 7346 2045 7380 2178
rect 7538 2045 7572 2178
rect 7730 2045 7764 2178
rect 7922 2045 7956 2178
rect 8070 2162 8080 2178
rect 8144 2162 8154 2226
rect 8298 2212 8332 2775
rect 8372 2665 8382 2717
rect 8434 2665 8461 2717
rect 16034 2713 16080 2891
rect 16250 2775 17332 2809
rect 16034 2327 16040 2713
rect 16074 2327 16080 2713
rect 16135 2665 16145 2717
rect 16197 2665 16207 2717
rect 16250 2625 16284 2775
rect 16327 2665 16337 2717
rect 16389 2665 16399 2717
rect 16442 2625 16476 2775
rect 16519 2665 16529 2717
rect 16581 2665 16591 2717
rect 16634 2625 16668 2775
rect 16711 2665 16721 2717
rect 16773 2665 16783 2717
rect 16826 2625 16860 2775
rect 16902 2665 16912 2717
rect 16964 2665 16974 2717
rect 17018 2625 17052 2775
rect 17095 2665 17105 2717
rect 17157 2665 17167 2717
rect 16148 2613 16194 2625
rect 16148 2365 16154 2613
rect 16188 2365 16194 2613
rect 16148 2353 16194 2365
rect 16244 2613 16290 2625
rect 16244 2365 16250 2613
rect 16284 2365 16290 2613
rect 16244 2353 16290 2365
rect 16340 2613 16386 2625
rect 16340 2365 16346 2613
rect 16380 2365 16386 2613
rect 16340 2353 16386 2365
rect 16436 2613 16482 2625
rect 16436 2365 16442 2613
rect 16476 2365 16482 2613
rect 16436 2353 16482 2365
rect 16532 2613 16578 2625
rect 16532 2365 16538 2613
rect 16572 2365 16578 2613
rect 16532 2353 16578 2365
rect 16628 2613 16674 2625
rect 16628 2365 16634 2613
rect 16668 2365 16674 2613
rect 16628 2353 16674 2365
rect 16724 2613 16770 2625
rect 16724 2365 16730 2613
rect 16764 2365 16770 2613
rect 16724 2353 16770 2365
rect 16820 2613 16866 2625
rect 16820 2365 16826 2613
rect 16860 2365 16866 2613
rect 16820 2353 16866 2365
rect 16916 2613 16962 2625
rect 16916 2365 16922 2613
rect 16956 2365 16962 2613
rect 16916 2353 16962 2365
rect 17012 2613 17058 2625
rect 17012 2365 17018 2613
rect 17052 2365 17058 2613
rect 17012 2353 17058 2365
rect 17108 2613 17154 2625
rect 17108 2365 17114 2613
rect 17148 2365 17154 2613
rect 17108 2353 17154 2365
rect 16034 2315 16080 2327
rect 8617 2212 11513 2228
rect 8298 2178 11513 2212
rect 8114 2045 8148 2162
rect 7148 2033 7194 2045
rect 7148 1953 7154 2033
rect 7188 1953 7194 2033
rect 7148 1941 7194 1953
rect 7244 2033 7290 2045
rect 7244 1953 7250 2033
rect 7284 1953 7290 2033
rect 7244 1941 7290 1953
rect 7340 2033 7386 2045
rect 7340 1953 7346 2033
rect 7380 1953 7386 2033
rect 7340 1941 7386 1953
rect 7436 2033 7482 2045
rect 7436 1953 7442 2033
rect 7476 1953 7482 2033
rect 7436 1941 7482 1953
rect 7532 2033 7578 2045
rect 7532 1953 7538 2033
rect 7572 1953 7578 2033
rect 7532 1941 7578 1953
rect 7628 2033 7674 2045
rect 7628 1953 7634 2033
rect 7668 1953 7674 2033
rect 7628 1941 7674 1953
rect 7724 2033 7770 2045
rect 7724 1953 7730 2033
rect 7764 1953 7770 2033
rect 7724 1941 7770 1953
rect 7820 2033 7866 2045
rect 7820 1953 7826 2033
rect 7860 1953 7866 2033
rect 7820 1941 7866 1953
rect 7916 2033 7962 2045
rect 7916 1953 7922 2033
rect 7956 1953 7962 2033
rect 7916 1941 7962 1953
rect 8012 2033 8058 2045
rect 8012 1953 8018 2033
rect 8052 1953 8058 2033
rect 8012 1941 8058 1953
rect 8108 2033 8154 2045
rect 8108 1953 8114 2033
rect 8148 1953 8154 2033
rect 8108 1941 8154 1953
rect 7138 1909 7204 1913
rect 7034 1691 7080 1863
rect 7135 1857 7145 1909
rect 7197 1857 7207 1909
rect 7138 1853 7204 1857
rect 7250 1801 7284 1941
rect 7330 1909 7396 1913
rect 7327 1857 7337 1909
rect 7389 1857 7399 1909
rect 7330 1853 7396 1857
rect 7442 1801 7476 1941
rect 7522 1910 7588 1913
rect 7520 1858 7530 1910
rect 7582 1858 7592 1910
rect 7522 1853 7588 1858
rect 7634 1801 7668 1941
rect 7714 1910 7780 1913
rect 7712 1858 7722 1910
rect 7774 1858 7784 1910
rect 7714 1853 7780 1858
rect 7826 1801 7860 1941
rect 7906 1910 7972 1913
rect 7904 1858 7914 1910
rect 7966 1858 7976 1910
rect 7906 1853 7972 1858
rect 8018 1801 8052 1941
rect 8098 1910 8164 1913
rect 8095 1858 8105 1910
rect 8157 1858 8167 1910
rect 8098 1853 8164 1858
rect 8298 1801 8332 2178
rect 8617 2164 11513 2178
rect 15783 2164 15793 2228
rect 15857 2212 15867 2228
rect 16154 2212 16188 2353
rect 16346 2212 16380 2353
rect 16538 2212 16572 2353
rect 16730 2212 16764 2353
rect 16922 2212 16956 2353
rect 17114 2212 17148 2353
rect 15857 2178 17148 2212
rect 15857 2164 15867 2178
rect 8372 1858 8382 1910
rect 8434 1858 8461 1910
rect 7250 1767 8332 1801
rect 7034 913 7080 1091
rect 7250 975 8332 1009
rect 7034 527 7040 913
rect 7074 527 7080 913
rect 7135 865 7145 917
rect 7197 865 7207 917
rect 7250 825 7284 975
rect 7327 865 7337 917
rect 7389 865 7399 917
rect 7442 825 7476 975
rect 7519 865 7529 917
rect 7581 865 7591 917
rect 7634 825 7668 975
rect 7711 865 7721 917
rect 7773 865 7783 917
rect 7826 825 7860 975
rect 7902 865 7912 917
rect 7964 865 7974 917
rect 8018 825 8052 975
rect 8095 865 8105 917
rect 8157 865 8167 917
rect 7148 813 7194 825
rect 7148 565 7154 813
rect 7188 565 7194 813
rect 7148 553 7194 565
rect 7244 813 7290 825
rect 7244 565 7250 813
rect 7284 565 7290 813
rect 7244 553 7290 565
rect 7340 813 7386 825
rect 7340 565 7346 813
rect 7380 565 7386 813
rect 7340 553 7386 565
rect 7436 813 7482 825
rect 7436 565 7442 813
rect 7476 565 7482 813
rect 7436 553 7482 565
rect 7532 813 7578 825
rect 7532 565 7538 813
rect 7572 565 7578 813
rect 7532 553 7578 565
rect 7628 813 7674 825
rect 7628 565 7634 813
rect 7668 565 7674 813
rect 7628 553 7674 565
rect 7724 813 7770 825
rect 7724 565 7730 813
rect 7764 565 7770 813
rect 7724 553 7770 565
rect 7820 813 7866 825
rect 7820 565 7826 813
rect 7860 565 7866 813
rect 7820 553 7866 565
rect 7916 813 7962 825
rect 7916 565 7922 813
rect 7956 565 7962 813
rect 7916 553 7962 565
rect 8012 813 8058 825
rect 8012 565 8018 813
rect 8052 565 8058 813
rect 8012 553 8058 565
rect 8108 813 8154 825
rect 8108 565 8114 813
rect 8148 565 8154 813
rect 8108 553 8154 565
rect 7034 515 7080 527
rect 7154 412 7188 553
rect 7346 412 7380 553
rect 7538 412 7572 553
rect 7730 412 7764 553
rect 7922 412 7956 553
rect 8114 426 8148 553
rect 8064 412 8074 426
rect 6216 378 8074 412
rect 6216 -3451 6291 378
rect 7034 263 7080 275
rect 7034 63 7040 263
rect 7074 63 7080 263
rect 7154 245 7188 378
rect 7346 245 7380 378
rect 7538 245 7572 378
rect 7730 245 7764 378
rect 7922 245 7956 378
rect 8064 362 8074 378
rect 8138 362 8148 426
rect 8114 245 8148 362
rect 8298 412 8332 975
rect 10720 943 10730 1007
rect 10794 943 10804 1007
rect 8372 865 8382 917
rect 8434 865 8461 917
rect 8615 412 8625 424
rect 8298 378 8625 412
rect 7148 233 7194 245
rect 7148 153 7154 233
rect 7188 153 7194 233
rect 7148 141 7194 153
rect 7244 233 7290 245
rect 7244 153 7250 233
rect 7284 153 7290 233
rect 7244 141 7290 153
rect 7340 233 7386 245
rect 7340 153 7346 233
rect 7380 153 7386 233
rect 7340 141 7386 153
rect 7436 233 7482 245
rect 7436 153 7442 233
rect 7476 153 7482 233
rect 7436 141 7482 153
rect 7532 233 7578 245
rect 7532 153 7538 233
rect 7572 153 7578 233
rect 7532 141 7578 153
rect 7628 233 7674 245
rect 7628 153 7634 233
rect 7668 153 7674 233
rect 7628 141 7674 153
rect 7724 233 7770 245
rect 7724 153 7730 233
rect 7764 153 7770 233
rect 7724 141 7770 153
rect 7820 233 7866 245
rect 7820 153 7826 233
rect 7860 153 7866 233
rect 7820 141 7866 153
rect 7916 233 7962 245
rect 7916 153 7922 233
rect 7956 153 7962 233
rect 7916 141 7962 153
rect 8012 233 8058 245
rect 8012 153 8018 233
rect 8052 153 8058 233
rect 8012 141 8058 153
rect 8108 233 8154 245
rect 8108 153 8114 233
rect 8148 153 8154 233
rect 8108 141 8154 153
rect 7138 109 7204 113
rect 7034 -109 7080 63
rect 7135 57 7145 109
rect 7197 57 7207 109
rect 7138 53 7204 57
rect 7250 1 7284 141
rect 7330 109 7396 113
rect 7327 57 7337 109
rect 7389 57 7399 109
rect 7330 53 7396 57
rect 7442 1 7476 141
rect 7522 110 7588 113
rect 7520 58 7530 110
rect 7582 58 7592 110
rect 7522 53 7588 58
rect 7634 1 7668 141
rect 7714 110 7780 113
rect 7712 58 7722 110
rect 7774 58 7784 110
rect 7714 53 7780 58
rect 7826 1 7860 141
rect 7906 110 7972 113
rect 7904 58 7914 110
rect 7966 58 7976 110
rect 7906 53 7972 58
rect 8018 1 8052 141
rect 8098 110 8164 113
rect 8095 58 8105 110
rect 8157 58 8167 110
rect 8098 53 8164 58
rect 8298 1 8332 378
rect 8615 360 8625 378
rect 8689 360 8699 424
rect 8372 58 8382 110
rect 8434 58 8461 110
rect 7250 -33 8332 1
rect 7034 -887 7080 -709
rect 7250 -825 8332 -791
rect 7034 -1273 7040 -887
rect 7074 -1273 7080 -887
rect 7135 -935 7145 -883
rect 7197 -935 7207 -883
rect 7250 -975 7284 -825
rect 7327 -935 7337 -883
rect 7389 -935 7399 -883
rect 7442 -975 7476 -825
rect 7519 -935 7529 -883
rect 7581 -935 7591 -883
rect 7634 -975 7668 -825
rect 7711 -935 7721 -883
rect 7773 -935 7783 -883
rect 7826 -975 7860 -825
rect 7902 -935 7912 -883
rect 7964 -935 7974 -883
rect 8018 -975 8052 -825
rect 8095 -935 8105 -883
rect 8157 -935 8167 -883
rect 7148 -987 7194 -975
rect 7148 -1235 7154 -987
rect 7188 -1235 7194 -987
rect 7148 -1247 7194 -1235
rect 7244 -987 7290 -975
rect 7244 -1235 7250 -987
rect 7284 -1235 7290 -987
rect 7244 -1247 7290 -1235
rect 7340 -987 7386 -975
rect 7340 -1235 7346 -987
rect 7380 -1235 7386 -987
rect 7340 -1247 7386 -1235
rect 7436 -987 7482 -975
rect 7436 -1235 7442 -987
rect 7476 -1235 7482 -987
rect 7436 -1247 7482 -1235
rect 7532 -987 7578 -975
rect 7532 -1235 7538 -987
rect 7572 -1235 7578 -987
rect 7532 -1247 7578 -1235
rect 7628 -987 7674 -975
rect 7628 -1235 7634 -987
rect 7668 -1235 7674 -987
rect 7628 -1247 7674 -1235
rect 7724 -987 7770 -975
rect 7724 -1235 7730 -987
rect 7764 -1235 7770 -987
rect 7724 -1247 7770 -1235
rect 7820 -987 7866 -975
rect 7820 -1235 7826 -987
rect 7860 -1235 7866 -987
rect 7820 -1247 7866 -1235
rect 7916 -987 7962 -975
rect 7916 -1235 7922 -987
rect 7956 -1235 7962 -987
rect 7916 -1247 7962 -1235
rect 8012 -987 8058 -975
rect 8012 -1235 8018 -987
rect 8052 -1235 8058 -987
rect 8012 -1247 8058 -1235
rect 8108 -987 8154 -975
rect 8108 -1235 8114 -987
rect 8148 -1235 8154 -987
rect 8108 -1247 8154 -1235
rect 7034 -1285 7080 -1273
rect 7154 -1388 7188 -1247
rect 7346 -1388 7380 -1247
rect 7538 -1388 7572 -1247
rect 7730 -1388 7764 -1247
rect 7922 -1388 7956 -1247
rect 8114 -1374 8148 -1247
rect 8068 -1388 8078 -1374
rect 6674 -1422 8078 -1388
rect 6674 -2199 6749 -1422
rect 7034 -1537 7080 -1525
rect 7034 -1737 7040 -1537
rect 7074 -1737 7080 -1537
rect 7154 -1555 7188 -1422
rect 7346 -1555 7380 -1422
rect 7538 -1555 7572 -1422
rect 7730 -1555 7764 -1422
rect 7922 -1555 7956 -1422
rect 8068 -1438 8078 -1422
rect 8142 -1438 8152 -1374
rect 8298 -1388 8332 -825
rect 8372 -935 8382 -883
rect 8434 -935 8461 -883
rect 8658 -1388 8668 -1375
rect 8298 -1422 8668 -1388
rect 8114 -1555 8148 -1438
rect 7148 -1567 7194 -1555
rect 7148 -1647 7154 -1567
rect 7188 -1647 7194 -1567
rect 7148 -1659 7194 -1647
rect 7244 -1567 7290 -1555
rect 7244 -1647 7250 -1567
rect 7284 -1647 7290 -1567
rect 7244 -1659 7290 -1647
rect 7340 -1567 7386 -1555
rect 7340 -1647 7346 -1567
rect 7380 -1647 7386 -1567
rect 7340 -1659 7386 -1647
rect 7436 -1567 7482 -1555
rect 7436 -1647 7442 -1567
rect 7476 -1647 7482 -1567
rect 7436 -1659 7482 -1647
rect 7532 -1567 7578 -1555
rect 7532 -1647 7538 -1567
rect 7572 -1647 7578 -1567
rect 7532 -1659 7578 -1647
rect 7628 -1567 7674 -1555
rect 7628 -1647 7634 -1567
rect 7668 -1647 7674 -1567
rect 7628 -1659 7674 -1647
rect 7724 -1567 7770 -1555
rect 7724 -1647 7730 -1567
rect 7764 -1647 7770 -1567
rect 7724 -1659 7770 -1647
rect 7820 -1567 7866 -1555
rect 7820 -1647 7826 -1567
rect 7860 -1647 7866 -1567
rect 7820 -1659 7866 -1647
rect 7916 -1567 7962 -1555
rect 7916 -1647 7922 -1567
rect 7956 -1647 7962 -1567
rect 7916 -1659 7962 -1647
rect 8012 -1567 8058 -1555
rect 8012 -1647 8018 -1567
rect 8052 -1647 8058 -1567
rect 8012 -1659 8058 -1647
rect 8108 -1567 8154 -1555
rect 8108 -1647 8114 -1567
rect 8148 -1647 8154 -1567
rect 8108 -1659 8154 -1647
rect 7138 -1691 7204 -1687
rect 7034 -1909 7080 -1737
rect 7135 -1743 7145 -1691
rect 7197 -1743 7207 -1691
rect 7138 -1747 7204 -1743
rect 7250 -1799 7284 -1659
rect 7330 -1691 7396 -1687
rect 7327 -1743 7337 -1691
rect 7389 -1743 7399 -1691
rect 7330 -1747 7396 -1743
rect 7442 -1799 7476 -1659
rect 7522 -1690 7588 -1687
rect 7520 -1742 7530 -1690
rect 7582 -1742 7592 -1690
rect 7522 -1747 7588 -1742
rect 7634 -1799 7668 -1659
rect 7714 -1690 7780 -1687
rect 7712 -1742 7722 -1690
rect 7774 -1742 7784 -1690
rect 7714 -1747 7780 -1742
rect 7826 -1799 7860 -1659
rect 7906 -1690 7972 -1687
rect 7904 -1742 7914 -1690
rect 7966 -1742 7976 -1690
rect 7906 -1747 7972 -1742
rect 8018 -1799 8052 -1659
rect 8098 -1690 8164 -1687
rect 8095 -1742 8105 -1690
rect 8157 -1742 8167 -1690
rect 8098 -1747 8164 -1742
rect 8298 -1799 8332 -1422
rect 8658 -1439 8668 -1422
rect 8732 -1439 8742 -1375
rect 10730 -1623 10794 943
rect 11449 -906 11513 2164
rect 16034 2063 16080 2075
rect 16034 1863 16040 2063
rect 16074 1863 16080 2063
rect 16154 2045 16188 2178
rect 16346 2045 16380 2178
rect 16538 2045 16572 2178
rect 16730 2045 16764 2178
rect 16922 2045 16956 2178
rect 17114 2045 17148 2178
rect 17298 2212 17332 2775
rect 17372 2665 17382 2717
rect 17434 2665 17461 2717
rect 17298 2178 18412 2212
rect 16148 2033 16194 2045
rect 16148 1953 16154 2033
rect 16188 1953 16194 2033
rect 16148 1941 16194 1953
rect 16244 2033 16290 2045
rect 16244 1953 16250 2033
rect 16284 1953 16290 2033
rect 16244 1941 16290 1953
rect 16340 2033 16386 2045
rect 16340 1953 16346 2033
rect 16380 1953 16386 2033
rect 16340 1941 16386 1953
rect 16436 2033 16482 2045
rect 16436 1953 16442 2033
rect 16476 1953 16482 2033
rect 16436 1941 16482 1953
rect 16532 2033 16578 2045
rect 16532 1953 16538 2033
rect 16572 1953 16578 2033
rect 16532 1941 16578 1953
rect 16628 2033 16674 2045
rect 16628 1953 16634 2033
rect 16668 1953 16674 2033
rect 16628 1941 16674 1953
rect 16724 2033 16770 2045
rect 16724 1953 16730 2033
rect 16764 1953 16770 2033
rect 16724 1941 16770 1953
rect 16820 2033 16866 2045
rect 16820 1953 16826 2033
rect 16860 1953 16866 2033
rect 16820 1941 16866 1953
rect 16916 2033 16962 2045
rect 16916 1953 16922 2033
rect 16956 1953 16962 2033
rect 16916 1941 16962 1953
rect 17012 2033 17058 2045
rect 17012 1953 17018 2033
rect 17052 1953 17058 2033
rect 17012 1941 17058 1953
rect 17108 2033 17154 2045
rect 17108 1953 17114 2033
rect 17148 1953 17154 2033
rect 17108 1941 17154 1953
rect 16138 1909 16204 1913
rect 16034 1691 16080 1863
rect 16135 1857 16145 1909
rect 16197 1857 16207 1909
rect 16138 1853 16204 1857
rect 16250 1801 16284 1941
rect 16330 1909 16396 1913
rect 16327 1857 16337 1909
rect 16389 1857 16399 1909
rect 16330 1853 16396 1857
rect 16442 1801 16476 1941
rect 16522 1910 16588 1913
rect 16520 1858 16530 1910
rect 16582 1858 16592 1910
rect 16522 1853 16588 1858
rect 16634 1801 16668 1941
rect 16714 1910 16780 1913
rect 16712 1858 16722 1910
rect 16774 1858 16784 1910
rect 16714 1853 16780 1858
rect 16826 1801 16860 1941
rect 16906 1910 16972 1913
rect 16904 1858 16914 1910
rect 16966 1858 16976 1910
rect 16906 1853 16972 1858
rect 17018 1801 17052 1941
rect 17098 1910 17164 1913
rect 17095 1858 17105 1910
rect 17157 1858 17167 1910
rect 17098 1853 17164 1858
rect 17298 1801 17332 2178
rect 17372 1858 17382 1910
rect 17434 1858 17461 1910
rect 16250 1767 17332 1801
rect 16034 913 16080 1091
rect 16250 975 17332 1009
rect 16034 527 16040 913
rect 16074 527 16080 913
rect 16135 865 16145 917
rect 16197 865 16207 917
rect 16250 825 16284 975
rect 16327 865 16337 917
rect 16389 865 16399 917
rect 16442 825 16476 975
rect 16519 865 16529 917
rect 16581 865 16591 917
rect 16634 825 16668 975
rect 16711 865 16721 917
rect 16773 865 16783 917
rect 16826 825 16860 975
rect 16902 865 16912 917
rect 16964 865 16974 917
rect 17018 825 17052 975
rect 17095 865 17105 917
rect 17157 865 17167 917
rect 16148 813 16194 825
rect 16148 565 16154 813
rect 16188 565 16194 813
rect 16148 553 16194 565
rect 16244 813 16290 825
rect 16244 565 16250 813
rect 16284 565 16290 813
rect 16244 553 16290 565
rect 16340 813 16386 825
rect 16340 565 16346 813
rect 16380 565 16386 813
rect 16340 553 16386 565
rect 16436 813 16482 825
rect 16436 565 16442 813
rect 16476 565 16482 813
rect 16436 553 16482 565
rect 16532 813 16578 825
rect 16532 565 16538 813
rect 16572 565 16578 813
rect 16532 553 16578 565
rect 16628 813 16674 825
rect 16628 565 16634 813
rect 16668 565 16674 813
rect 16628 553 16674 565
rect 16724 813 16770 825
rect 16724 565 16730 813
rect 16764 565 16770 813
rect 16724 553 16770 565
rect 16820 813 16866 825
rect 16820 565 16826 813
rect 16860 565 16866 813
rect 16820 553 16866 565
rect 16916 813 16962 825
rect 16916 565 16922 813
rect 16956 565 16962 813
rect 16916 553 16962 565
rect 17012 813 17058 825
rect 17012 565 17018 813
rect 17052 565 17058 813
rect 17012 553 17058 565
rect 17108 813 17154 825
rect 17108 565 17114 813
rect 17148 565 17154 813
rect 17108 553 17154 565
rect 16034 515 16080 527
rect 15796 362 15806 426
rect 15870 412 15880 426
rect 16154 412 16188 553
rect 16346 412 16380 553
rect 16538 412 16572 553
rect 16730 412 16764 553
rect 16922 412 16956 553
rect 17114 412 17148 553
rect 15870 378 17148 412
rect 15870 362 15880 378
rect 16034 263 16080 275
rect 12249 25 12259 89
rect 12323 25 12333 89
rect 16034 63 16040 263
rect 16074 63 16080 263
rect 16154 245 16188 378
rect 16346 245 16380 378
rect 16538 245 16572 378
rect 16730 245 16764 378
rect 16922 245 16956 378
rect 17114 245 17148 378
rect 17298 412 17332 975
rect 17372 865 17382 917
rect 17434 865 17461 917
rect 17298 378 17901 412
rect 16148 233 16194 245
rect 16148 153 16154 233
rect 16188 153 16194 233
rect 16148 141 16194 153
rect 16244 233 16290 245
rect 16244 153 16250 233
rect 16284 153 16290 233
rect 16244 141 16290 153
rect 16340 233 16386 245
rect 16340 153 16346 233
rect 16380 153 16386 233
rect 16340 141 16386 153
rect 16436 233 16482 245
rect 16436 153 16442 233
rect 16476 153 16482 233
rect 16436 141 16482 153
rect 16532 233 16578 245
rect 16532 153 16538 233
rect 16572 153 16578 233
rect 16532 141 16578 153
rect 16628 233 16674 245
rect 16628 153 16634 233
rect 16668 153 16674 233
rect 16628 141 16674 153
rect 16724 233 16770 245
rect 16724 153 16730 233
rect 16764 153 16770 233
rect 16724 141 16770 153
rect 16820 233 16866 245
rect 16820 153 16826 233
rect 16860 153 16866 233
rect 16820 141 16866 153
rect 16916 233 16962 245
rect 16916 153 16922 233
rect 16956 153 16962 233
rect 16916 141 16962 153
rect 17012 233 17058 245
rect 17012 153 17018 233
rect 17052 153 17058 233
rect 17012 141 17058 153
rect 17108 233 17154 245
rect 17108 153 17114 233
rect 17148 153 17154 233
rect 17108 141 17154 153
rect 16138 109 16204 113
rect 12259 -385 12323 25
rect 16034 -109 16080 63
rect 16135 57 16145 109
rect 16197 57 16207 109
rect 16138 53 16204 57
rect 16250 1 16284 141
rect 16330 109 16396 113
rect 16327 57 16337 109
rect 16389 57 16399 109
rect 16330 53 16396 57
rect 16442 1 16476 141
rect 16522 110 16588 113
rect 16520 58 16530 110
rect 16582 58 16592 110
rect 16522 53 16588 58
rect 16634 1 16668 141
rect 16714 110 16780 113
rect 16712 58 16722 110
rect 16774 58 16784 110
rect 16714 53 16780 58
rect 16826 1 16860 141
rect 16906 110 16972 113
rect 16904 58 16914 110
rect 16966 58 16976 110
rect 16906 53 16972 58
rect 17018 1 17052 141
rect 17098 110 17164 113
rect 17095 58 17105 110
rect 17157 58 17167 110
rect 17098 53 17164 58
rect 17298 1 17332 378
rect 17372 58 17382 110
rect 17434 58 17461 110
rect 16250 -33 17332 1
rect 12249 -449 12259 -385
rect 12323 -449 12333 -385
rect 12933 -541 15268 -537
rect 12860 -605 12870 -541
rect 12934 -601 15268 -541
rect 15332 -601 15342 -537
rect 12934 -605 12944 -601
rect 16034 -887 16080 -709
rect 16250 -825 17332 -791
rect 11449 -970 12208 -906
rect 12272 -970 12282 -906
rect 13976 -1143 14309 -1079
rect 14373 -1143 14383 -1079
rect 12400 -1321 12410 -1257
rect 12474 -1321 12484 -1257
rect 12410 -1384 12474 -1321
rect 10730 -1687 10968 -1623
rect 8372 -1742 8382 -1690
rect 8434 -1742 8461 -1690
rect 7250 -1833 8332 -1799
rect 9425 -2050 9435 -1986
rect 9499 -2050 10733 -1986
rect 10797 -2050 10807 -1986
rect 6670 -2263 6680 -2199
rect 6744 -2263 6754 -2199
rect 6674 -3188 6749 -2263
rect 10904 -2315 10968 -1687
rect 9425 -2379 9435 -2315
rect 9499 -2379 10968 -2315
rect 7034 -2687 7080 -2509
rect 7250 -2625 8332 -2591
rect 7034 -3073 7040 -2687
rect 7074 -3073 7080 -2687
rect 7135 -2735 7145 -2683
rect 7197 -2735 7207 -2683
rect 7250 -2775 7284 -2625
rect 7327 -2735 7337 -2683
rect 7389 -2735 7399 -2683
rect 7442 -2775 7476 -2625
rect 7519 -2735 7529 -2683
rect 7581 -2735 7591 -2683
rect 7634 -2775 7668 -2625
rect 7711 -2735 7721 -2683
rect 7773 -2735 7783 -2683
rect 7826 -2775 7860 -2625
rect 7902 -2735 7912 -2683
rect 7964 -2735 7974 -2683
rect 8018 -2775 8052 -2625
rect 8095 -2735 8105 -2683
rect 8157 -2735 8167 -2683
rect 7148 -2787 7194 -2775
rect 7148 -3035 7154 -2787
rect 7188 -3035 7194 -2787
rect 7148 -3047 7194 -3035
rect 7244 -2787 7290 -2775
rect 7244 -3035 7250 -2787
rect 7284 -3035 7290 -2787
rect 7244 -3047 7290 -3035
rect 7340 -2787 7386 -2775
rect 7340 -3035 7346 -2787
rect 7380 -3035 7386 -2787
rect 7340 -3047 7386 -3035
rect 7436 -2787 7482 -2775
rect 7436 -3035 7442 -2787
rect 7476 -3035 7482 -2787
rect 7436 -3047 7482 -3035
rect 7532 -2787 7578 -2775
rect 7532 -3035 7538 -2787
rect 7572 -3035 7578 -2787
rect 7532 -3047 7578 -3035
rect 7628 -2787 7674 -2775
rect 7628 -3035 7634 -2787
rect 7668 -3035 7674 -2787
rect 7628 -3047 7674 -3035
rect 7724 -2787 7770 -2775
rect 7724 -3035 7730 -2787
rect 7764 -3035 7770 -2787
rect 7724 -3047 7770 -3035
rect 7820 -2787 7866 -2775
rect 7820 -3035 7826 -2787
rect 7860 -3035 7866 -2787
rect 7820 -3047 7866 -3035
rect 7916 -2787 7962 -2775
rect 7916 -3035 7922 -2787
rect 7956 -3035 7962 -2787
rect 7916 -3047 7962 -3035
rect 8012 -2787 8058 -2775
rect 8012 -3035 8018 -2787
rect 8052 -3035 8058 -2787
rect 8012 -3047 8058 -3035
rect 8108 -2787 8154 -2775
rect 8108 -3035 8114 -2787
rect 8148 -3035 8154 -2787
rect 8108 -3047 8154 -3035
rect 7034 -3085 7080 -3073
rect 7154 -3188 7188 -3047
rect 7346 -3188 7380 -3047
rect 7538 -3188 7572 -3047
rect 7730 -3188 7764 -3047
rect 7922 -3188 7956 -3047
rect 8114 -3174 8148 -3047
rect 8065 -3188 8075 -3174
rect 6674 -3222 8075 -3188
rect 7034 -3337 7080 -3325
rect 6212 -3515 6222 -3451
rect 6286 -3515 6296 -3451
rect 6216 -4988 6291 -3515
rect 7034 -3537 7040 -3337
rect 7074 -3537 7080 -3337
rect 7154 -3355 7188 -3222
rect 7346 -3355 7380 -3222
rect 7538 -3355 7572 -3222
rect 7730 -3355 7764 -3222
rect 7922 -3355 7956 -3222
rect 8065 -3238 8075 -3222
rect 8139 -3238 8149 -3174
rect 8298 -3188 8332 -2625
rect 8372 -2735 8382 -2683
rect 8434 -2735 8461 -2683
rect 8658 -3188 8668 -3178
rect 8298 -3222 8668 -3188
rect 8114 -3355 8148 -3238
rect 7148 -3367 7194 -3355
rect 7148 -3447 7154 -3367
rect 7188 -3447 7194 -3367
rect 7148 -3459 7194 -3447
rect 7244 -3367 7290 -3355
rect 7244 -3447 7250 -3367
rect 7284 -3447 7290 -3367
rect 7244 -3459 7290 -3447
rect 7340 -3367 7386 -3355
rect 7340 -3447 7346 -3367
rect 7380 -3447 7386 -3367
rect 7340 -3459 7386 -3447
rect 7436 -3367 7482 -3355
rect 7436 -3447 7442 -3367
rect 7476 -3447 7482 -3367
rect 7436 -3459 7482 -3447
rect 7532 -3367 7578 -3355
rect 7532 -3447 7538 -3367
rect 7572 -3447 7578 -3367
rect 7532 -3459 7578 -3447
rect 7628 -3367 7674 -3355
rect 7628 -3447 7634 -3367
rect 7668 -3447 7674 -3367
rect 7628 -3459 7674 -3447
rect 7724 -3367 7770 -3355
rect 7724 -3447 7730 -3367
rect 7764 -3447 7770 -3367
rect 7724 -3459 7770 -3447
rect 7820 -3367 7866 -3355
rect 7820 -3447 7826 -3367
rect 7860 -3447 7866 -3367
rect 7820 -3459 7866 -3447
rect 7916 -3367 7962 -3355
rect 7916 -3447 7922 -3367
rect 7956 -3447 7962 -3367
rect 7916 -3459 7962 -3447
rect 8012 -3367 8058 -3355
rect 8012 -3447 8018 -3367
rect 8052 -3447 8058 -3367
rect 8012 -3459 8058 -3447
rect 8108 -3367 8154 -3355
rect 8108 -3447 8114 -3367
rect 8148 -3447 8154 -3367
rect 8108 -3459 8154 -3447
rect 7138 -3491 7204 -3487
rect 7034 -3709 7080 -3537
rect 7135 -3543 7145 -3491
rect 7197 -3543 7207 -3491
rect 7138 -3547 7204 -3543
rect 7250 -3599 7284 -3459
rect 7330 -3491 7396 -3487
rect 7327 -3543 7337 -3491
rect 7389 -3543 7399 -3491
rect 7330 -3547 7396 -3543
rect 7442 -3599 7476 -3459
rect 7522 -3490 7588 -3487
rect 7520 -3542 7530 -3490
rect 7582 -3542 7592 -3490
rect 7522 -3547 7588 -3542
rect 7634 -3599 7668 -3459
rect 7714 -3490 7780 -3487
rect 7712 -3542 7722 -3490
rect 7774 -3542 7784 -3490
rect 7714 -3547 7780 -3542
rect 7826 -3599 7860 -3459
rect 7906 -3490 7972 -3487
rect 7904 -3542 7914 -3490
rect 7966 -3542 7976 -3490
rect 7906 -3547 7972 -3542
rect 8018 -3599 8052 -3459
rect 8098 -3490 8164 -3487
rect 8095 -3542 8105 -3490
rect 8157 -3542 8167 -3490
rect 8098 -3547 8164 -3542
rect 8298 -3599 8332 -3222
rect 8658 -3242 8668 -3222
rect 8732 -3242 8742 -3178
rect 12410 -3246 12473 -1384
rect 13976 -1827 14040 -1143
rect 16034 -1273 16040 -887
rect 16074 -1273 16080 -887
rect 16135 -935 16145 -883
rect 16197 -935 16207 -883
rect 16250 -975 16284 -825
rect 16327 -935 16337 -883
rect 16389 -935 16399 -883
rect 16442 -975 16476 -825
rect 16519 -935 16529 -883
rect 16581 -935 16591 -883
rect 16634 -975 16668 -825
rect 16711 -935 16721 -883
rect 16773 -935 16783 -883
rect 16826 -975 16860 -825
rect 16902 -935 16912 -883
rect 16964 -935 16974 -883
rect 17018 -975 17052 -825
rect 17095 -935 17105 -883
rect 17157 -935 17167 -883
rect 16148 -987 16194 -975
rect 16148 -1235 16154 -987
rect 16188 -1235 16194 -987
rect 16148 -1247 16194 -1235
rect 16244 -987 16290 -975
rect 16244 -1235 16250 -987
rect 16284 -1235 16290 -987
rect 16244 -1247 16290 -1235
rect 16340 -987 16386 -975
rect 16340 -1235 16346 -987
rect 16380 -1235 16386 -987
rect 16340 -1247 16386 -1235
rect 16436 -987 16482 -975
rect 16436 -1235 16442 -987
rect 16476 -1235 16482 -987
rect 16436 -1247 16482 -1235
rect 16532 -987 16578 -975
rect 16532 -1235 16538 -987
rect 16572 -1235 16578 -987
rect 16532 -1247 16578 -1235
rect 16628 -987 16674 -975
rect 16628 -1235 16634 -987
rect 16668 -1235 16674 -987
rect 16628 -1247 16674 -1235
rect 16724 -987 16770 -975
rect 16724 -1235 16730 -987
rect 16764 -1235 16770 -987
rect 16724 -1247 16770 -1235
rect 16820 -987 16866 -975
rect 16820 -1235 16826 -987
rect 16860 -1235 16866 -987
rect 16820 -1247 16866 -1235
rect 16916 -987 16962 -975
rect 16916 -1235 16922 -987
rect 16956 -1235 16962 -987
rect 16916 -1247 16962 -1235
rect 17012 -987 17058 -975
rect 17012 -1235 17018 -987
rect 17052 -1235 17058 -987
rect 17012 -1247 17058 -1235
rect 17108 -987 17154 -975
rect 17108 -1235 17114 -987
rect 17148 -1235 17154 -987
rect 17108 -1247 17154 -1235
rect 16034 -1285 16080 -1273
rect 15851 -1438 15861 -1374
rect 15925 -1388 15935 -1374
rect 16154 -1388 16188 -1247
rect 16346 -1388 16380 -1247
rect 16538 -1388 16572 -1247
rect 16730 -1388 16764 -1247
rect 16922 -1388 16956 -1247
rect 17114 -1388 17148 -1247
rect 15925 -1422 17148 -1388
rect 15925 -1438 15935 -1422
rect 16034 -1537 16080 -1525
rect 16034 -1737 16040 -1537
rect 16074 -1737 16080 -1537
rect 16154 -1555 16188 -1422
rect 16346 -1555 16380 -1422
rect 16538 -1555 16572 -1422
rect 16730 -1555 16764 -1422
rect 16922 -1555 16956 -1422
rect 17114 -1555 17148 -1422
rect 17298 -1388 17332 -825
rect 17372 -935 17382 -883
rect 17434 -935 17461 -883
rect 17826 -1388 17901 378
rect 17298 -1422 17901 -1388
rect 16148 -1567 16194 -1555
rect 16148 -1647 16154 -1567
rect 16188 -1647 16194 -1567
rect 16148 -1659 16194 -1647
rect 16244 -1567 16290 -1555
rect 16244 -1647 16250 -1567
rect 16284 -1647 16290 -1567
rect 16244 -1659 16290 -1647
rect 16340 -1567 16386 -1555
rect 16340 -1647 16346 -1567
rect 16380 -1647 16386 -1567
rect 16340 -1659 16386 -1647
rect 16436 -1567 16482 -1555
rect 16436 -1647 16442 -1567
rect 16476 -1647 16482 -1567
rect 16436 -1659 16482 -1647
rect 16532 -1567 16578 -1555
rect 16532 -1647 16538 -1567
rect 16572 -1647 16578 -1567
rect 16532 -1659 16578 -1647
rect 16628 -1567 16674 -1555
rect 16628 -1647 16634 -1567
rect 16668 -1647 16674 -1567
rect 16628 -1659 16674 -1647
rect 16724 -1567 16770 -1555
rect 16724 -1647 16730 -1567
rect 16764 -1647 16770 -1567
rect 16724 -1659 16770 -1647
rect 16820 -1567 16866 -1555
rect 16820 -1647 16826 -1567
rect 16860 -1647 16866 -1567
rect 16820 -1659 16866 -1647
rect 16916 -1567 16962 -1555
rect 16916 -1647 16922 -1567
rect 16956 -1647 16962 -1567
rect 16916 -1659 16962 -1647
rect 17012 -1567 17058 -1555
rect 17012 -1647 17018 -1567
rect 17052 -1647 17058 -1567
rect 17012 -1659 17058 -1647
rect 17108 -1567 17154 -1555
rect 17108 -1647 17114 -1567
rect 17148 -1647 17154 -1567
rect 17108 -1659 17154 -1647
rect 16138 -1691 16204 -1687
rect 13966 -1891 13976 -1827
rect 14040 -1891 14050 -1827
rect 16034 -1909 16080 -1737
rect 16135 -1743 16145 -1691
rect 16197 -1743 16207 -1691
rect 16138 -1747 16204 -1743
rect 16250 -1799 16284 -1659
rect 16330 -1691 16396 -1687
rect 16327 -1743 16337 -1691
rect 16389 -1743 16399 -1691
rect 16330 -1747 16396 -1743
rect 16442 -1799 16476 -1659
rect 16522 -1690 16588 -1687
rect 16520 -1742 16530 -1690
rect 16582 -1742 16592 -1690
rect 16522 -1747 16588 -1742
rect 16634 -1799 16668 -1659
rect 16714 -1690 16780 -1687
rect 16712 -1742 16722 -1690
rect 16774 -1742 16784 -1690
rect 16714 -1747 16780 -1742
rect 16826 -1799 16860 -1659
rect 16906 -1690 16972 -1687
rect 16904 -1742 16914 -1690
rect 16966 -1742 16976 -1690
rect 16906 -1747 16972 -1742
rect 17018 -1799 17052 -1659
rect 17098 -1690 17164 -1687
rect 17095 -1742 17105 -1690
rect 17157 -1742 17167 -1690
rect 17098 -1747 17164 -1742
rect 17298 -1799 17332 -1422
rect 17372 -1742 17382 -1690
rect 17434 -1742 17461 -1690
rect 16250 -1833 17332 -1799
rect 16034 -2687 16080 -2509
rect 16250 -2625 17332 -2591
rect 16034 -3073 16040 -2687
rect 16074 -3073 16080 -2687
rect 16135 -2735 16145 -2683
rect 16197 -2735 16207 -2683
rect 16250 -2775 16284 -2625
rect 16327 -2735 16337 -2683
rect 16389 -2735 16399 -2683
rect 16442 -2775 16476 -2625
rect 16519 -2735 16529 -2683
rect 16581 -2735 16591 -2683
rect 16634 -2775 16668 -2625
rect 16711 -2735 16721 -2683
rect 16773 -2735 16783 -2683
rect 16826 -2775 16860 -2625
rect 16902 -2735 16912 -2683
rect 16964 -2735 16974 -2683
rect 17018 -2775 17052 -2625
rect 17095 -2735 17105 -2683
rect 17157 -2735 17167 -2683
rect 16148 -2787 16194 -2775
rect 16148 -3035 16154 -2787
rect 16188 -3035 16194 -2787
rect 16148 -3047 16194 -3035
rect 16244 -2787 16290 -2775
rect 16244 -3035 16250 -2787
rect 16284 -3035 16290 -2787
rect 16244 -3047 16290 -3035
rect 16340 -2787 16386 -2775
rect 16340 -3035 16346 -2787
rect 16380 -3035 16386 -2787
rect 16340 -3047 16386 -3035
rect 16436 -2787 16482 -2775
rect 16436 -3035 16442 -2787
rect 16476 -3035 16482 -2787
rect 16436 -3047 16482 -3035
rect 16532 -2787 16578 -2775
rect 16532 -3035 16538 -2787
rect 16572 -3035 16578 -2787
rect 16532 -3047 16578 -3035
rect 16628 -2787 16674 -2775
rect 16628 -3035 16634 -2787
rect 16668 -3035 16674 -2787
rect 16628 -3047 16674 -3035
rect 16724 -2787 16770 -2775
rect 16724 -3035 16730 -2787
rect 16764 -3035 16770 -2787
rect 16724 -3047 16770 -3035
rect 16820 -2787 16866 -2775
rect 16820 -3035 16826 -2787
rect 16860 -3035 16866 -2787
rect 16820 -3047 16866 -3035
rect 16916 -2787 16962 -2775
rect 16916 -3035 16922 -2787
rect 16956 -3035 16962 -2787
rect 16916 -3047 16962 -3035
rect 17012 -2787 17058 -2775
rect 17012 -3035 17018 -2787
rect 17052 -3035 17058 -2787
rect 17012 -3047 17058 -3035
rect 17108 -2787 17154 -2775
rect 17108 -3035 17114 -2787
rect 17148 -3035 17154 -2787
rect 17108 -3047 17154 -3035
rect 16034 -3085 16080 -3073
rect 15856 -3236 15866 -3172
rect 15930 -3188 15940 -3172
rect 16154 -3188 16188 -3047
rect 16346 -3188 16380 -3047
rect 16538 -3188 16572 -3047
rect 16730 -3188 16764 -3047
rect 16922 -3188 16956 -3047
rect 17114 -3188 17148 -3047
rect 15930 -3222 17148 -3188
rect 15930 -3236 15940 -3222
rect 12400 -3310 12410 -3246
rect 12474 -3310 12484 -3246
rect 16034 -3337 16080 -3325
rect 8372 -3542 8382 -3490
rect 8434 -3542 8461 -3490
rect 16034 -3537 16040 -3337
rect 16074 -3537 16080 -3337
rect 16154 -3355 16188 -3222
rect 16346 -3355 16380 -3222
rect 16538 -3355 16572 -3222
rect 16730 -3355 16764 -3222
rect 16922 -3355 16956 -3222
rect 17114 -3355 17148 -3222
rect 17298 -3188 17332 -2625
rect 17372 -2735 17382 -2683
rect 17434 -2735 17461 -2683
rect 17826 -3188 17901 -1422
rect 17298 -3222 17901 -3188
rect 16148 -3367 16194 -3355
rect 16148 -3447 16154 -3367
rect 16188 -3447 16194 -3367
rect 16148 -3459 16194 -3447
rect 16244 -3367 16290 -3355
rect 16244 -3447 16250 -3367
rect 16284 -3447 16290 -3367
rect 16244 -3459 16290 -3447
rect 16340 -3367 16386 -3355
rect 16340 -3447 16346 -3367
rect 16380 -3447 16386 -3367
rect 16340 -3459 16386 -3447
rect 16436 -3367 16482 -3355
rect 16436 -3447 16442 -3367
rect 16476 -3447 16482 -3367
rect 16436 -3459 16482 -3447
rect 16532 -3367 16578 -3355
rect 16532 -3447 16538 -3367
rect 16572 -3447 16578 -3367
rect 16532 -3459 16578 -3447
rect 16628 -3367 16674 -3355
rect 16628 -3447 16634 -3367
rect 16668 -3447 16674 -3367
rect 16628 -3459 16674 -3447
rect 16724 -3367 16770 -3355
rect 16724 -3447 16730 -3367
rect 16764 -3447 16770 -3367
rect 16724 -3459 16770 -3447
rect 16820 -3367 16866 -3355
rect 16820 -3447 16826 -3367
rect 16860 -3447 16866 -3367
rect 16820 -3459 16866 -3447
rect 16916 -3367 16962 -3355
rect 16916 -3447 16922 -3367
rect 16956 -3447 16962 -3367
rect 16916 -3459 16962 -3447
rect 17012 -3367 17058 -3355
rect 17012 -3447 17018 -3367
rect 17052 -3447 17058 -3367
rect 17012 -3459 17058 -3447
rect 17108 -3367 17154 -3355
rect 17108 -3447 17114 -3367
rect 17148 -3447 17154 -3367
rect 17108 -3459 17154 -3447
rect 16138 -3491 16204 -3487
rect 7250 -3633 8332 -3599
rect 16034 -3709 16080 -3537
rect 16135 -3543 16145 -3491
rect 16197 -3543 16207 -3491
rect 16138 -3547 16204 -3543
rect 16250 -3599 16284 -3459
rect 16330 -3491 16396 -3487
rect 16327 -3543 16337 -3491
rect 16389 -3543 16399 -3491
rect 16330 -3547 16396 -3543
rect 16442 -3599 16476 -3459
rect 16522 -3490 16588 -3487
rect 16520 -3542 16530 -3490
rect 16582 -3542 16592 -3490
rect 16522 -3547 16588 -3542
rect 16634 -3599 16668 -3459
rect 16714 -3490 16780 -3487
rect 16712 -3542 16722 -3490
rect 16774 -3542 16784 -3490
rect 16714 -3547 16780 -3542
rect 16826 -3599 16860 -3459
rect 16906 -3490 16972 -3487
rect 16904 -3542 16914 -3490
rect 16966 -3542 16976 -3490
rect 16906 -3547 16972 -3542
rect 17018 -3599 17052 -3459
rect 17098 -3490 17164 -3487
rect 17095 -3542 17105 -3490
rect 17157 -3542 17167 -3490
rect 17098 -3547 17164 -3542
rect 17298 -3599 17332 -3222
rect 17372 -3542 17382 -3490
rect 17434 -3542 17461 -3490
rect 16250 -3633 17332 -3599
rect 8738 -3893 11432 -3829
rect 11496 -3893 11506 -3829
rect 7034 -4487 7080 -4309
rect 7250 -4425 8332 -4391
rect 7034 -4873 7040 -4487
rect 7074 -4873 7080 -4487
rect 7135 -4535 7145 -4483
rect 7197 -4535 7207 -4483
rect 7250 -4575 7284 -4425
rect 7327 -4535 7337 -4483
rect 7389 -4535 7399 -4483
rect 7442 -4575 7476 -4425
rect 7519 -4535 7529 -4483
rect 7581 -4535 7591 -4483
rect 7634 -4575 7668 -4425
rect 7711 -4535 7721 -4483
rect 7773 -4535 7783 -4483
rect 7826 -4575 7860 -4425
rect 7902 -4535 7912 -4483
rect 7964 -4535 7974 -4483
rect 8018 -4575 8052 -4425
rect 8095 -4535 8105 -4483
rect 8157 -4535 8167 -4483
rect 7148 -4587 7194 -4575
rect 7148 -4835 7154 -4587
rect 7188 -4835 7194 -4587
rect 7148 -4847 7194 -4835
rect 7244 -4587 7290 -4575
rect 7244 -4835 7250 -4587
rect 7284 -4835 7290 -4587
rect 7244 -4847 7290 -4835
rect 7340 -4587 7386 -4575
rect 7340 -4835 7346 -4587
rect 7380 -4835 7386 -4587
rect 7340 -4847 7386 -4835
rect 7436 -4587 7482 -4575
rect 7436 -4835 7442 -4587
rect 7476 -4835 7482 -4587
rect 7436 -4847 7482 -4835
rect 7532 -4587 7578 -4575
rect 7532 -4835 7538 -4587
rect 7572 -4835 7578 -4587
rect 7532 -4847 7578 -4835
rect 7628 -4587 7674 -4575
rect 7628 -4835 7634 -4587
rect 7668 -4835 7674 -4587
rect 7628 -4847 7674 -4835
rect 7724 -4587 7770 -4575
rect 7724 -4835 7730 -4587
rect 7764 -4835 7770 -4587
rect 7724 -4847 7770 -4835
rect 7820 -4587 7866 -4575
rect 7820 -4835 7826 -4587
rect 7860 -4835 7866 -4587
rect 7820 -4847 7866 -4835
rect 7916 -4587 7962 -4575
rect 7916 -4835 7922 -4587
rect 7956 -4835 7962 -4587
rect 7916 -4847 7962 -4835
rect 8012 -4587 8058 -4575
rect 8012 -4835 8018 -4587
rect 8052 -4835 8058 -4587
rect 8012 -4847 8058 -4835
rect 8108 -4587 8154 -4575
rect 8108 -4835 8114 -4587
rect 8148 -4835 8154 -4587
rect 8108 -4847 8154 -4835
rect 7034 -4885 7080 -4873
rect 7154 -4988 7188 -4847
rect 7346 -4988 7380 -4847
rect 7538 -4988 7572 -4847
rect 7730 -4988 7764 -4847
rect 7922 -4988 7956 -4847
rect 8114 -4972 8148 -4847
rect 8072 -4988 8082 -4972
rect 6216 -5022 8082 -4988
rect 7034 -5137 7080 -5125
rect 5604 -5271 5614 -5207
rect 5678 -5271 5688 -5207
rect 5327 -5580 5337 -5527
rect 5390 -5580 5400 -5527
rect 5608 -6788 5683 -5271
rect 7034 -5337 7040 -5137
rect 7074 -5337 7080 -5137
rect 7154 -5155 7188 -5022
rect 7346 -5155 7380 -5022
rect 7538 -5155 7572 -5022
rect 7730 -5155 7764 -5022
rect 7922 -5155 7956 -5022
rect 8072 -5036 8082 -5022
rect 8146 -5036 8156 -4972
rect 8298 -4988 8332 -4425
rect 8372 -4535 8382 -4483
rect 8434 -4535 8461 -4483
rect 8738 -4988 8802 -3893
rect 12694 -4007 12704 -3943
rect 12768 -4007 15254 -3943
rect 15318 -4007 15328 -3943
rect 9262 -4192 9272 -4128
rect 9336 -4192 13428 -4128
rect 13492 -4192 13502 -4128
rect 16034 -4487 16080 -4309
rect 16250 -4425 17332 -4391
rect 16034 -4873 16040 -4487
rect 16074 -4873 16080 -4487
rect 16135 -4535 16145 -4483
rect 16197 -4535 16207 -4483
rect 16250 -4575 16284 -4425
rect 16327 -4535 16337 -4483
rect 16389 -4535 16399 -4483
rect 16442 -4575 16476 -4425
rect 16519 -4535 16529 -4483
rect 16581 -4535 16591 -4483
rect 16634 -4575 16668 -4425
rect 16711 -4535 16721 -4483
rect 16773 -4535 16783 -4483
rect 16826 -4575 16860 -4425
rect 16902 -4535 16912 -4483
rect 16964 -4535 16974 -4483
rect 17018 -4575 17052 -4425
rect 17095 -4535 17105 -4483
rect 17157 -4535 17167 -4483
rect 16148 -4587 16194 -4575
rect 16148 -4835 16154 -4587
rect 16188 -4835 16194 -4587
rect 16148 -4847 16194 -4835
rect 16244 -4587 16290 -4575
rect 16244 -4835 16250 -4587
rect 16284 -4835 16290 -4587
rect 16244 -4847 16290 -4835
rect 16340 -4587 16386 -4575
rect 16340 -4835 16346 -4587
rect 16380 -4835 16386 -4587
rect 16340 -4847 16386 -4835
rect 16436 -4587 16482 -4575
rect 16436 -4835 16442 -4587
rect 16476 -4835 16482 -4587
rect 16436 -4847 16482 -4835
rect 16532 -4587 16578 -4575
rect 16532 -4835 16538 -4587
rect 16572 -4835 16578 -4587
rect 16532 -4847 16578 -4835
rect 16628 -4587 16674 -4575
rect 16628 -4835 16634 -4587
rect 16668 -4835 16674 -4587
rect 16628 -4847 16674 -4835
rect 16724 -4587 16770 -4575
rect 16724 -4835 16730 -4587
rect 16764 -4835 16770 -4587
rect 16724 -4847 16770 -4835
rect 16820 -4587 16866 -4575
rect 16820 -4835 16826 -4587
rect 16860 -4835 16866 -4587
rect 16820 -4847 16866 -4835
rect 16916 -4587 16962 -4575
rect 16916 -4835 16922 -4587
rect 16956 -4835 16962 -4587
rect 16916 -4847 16962 -4835
rect 17012 -4587 17058 -4575
rect 17012 -4835 17018 -4587
rect 17052 -4835 17058 -4587
rect 17012 -4847 17058 -4835
rect 17108 -4587 17154 -4575
rect 17108 -4835 17114 -4587
rect 17148 -4835 17154 -4587
rect 17108 -4847 17154 -4835
rect 16034 -4885 16080 -4873
rect 8298 -5022 8802 -4988
rect 8114 -5155 8148 -5036
rect 7148 -5167 7194 -5155
rect 7148 -5247 7154 -5167
rect 7188 -5247 7194 -5167
rect 7148 -5259 7194 -5247
rect 7244 -5167 7290 -5155
rect 7244 -5247 7250 -5167
rect 7284 -5247 7290 -5167
rect 7244 -5259 7290 -5247
rect 7340 -5167 7386 -5155
rect 7340 -5247 7346 -5167
rect 7380 -5247 7386 -5167
rect 7340 -5259 7386 -5247
rect 7436 -5167 7482 -5155
rect 7436 -5247 7442 -5167
rect 7476 -5247 7482 -5167
rect 7436 -5259 7482 -5247
rect 7532 -5167 7578 -5155
rect 7532 -5247 7538 -5167
rect 7572 -5247 7578 -5167
rect 7532 -5259 7578 -5247
rect 7628 -5167 7674 -5155
rect 7628 -5247 7634 -5167
rect 7668 -5247 7674 -5167
rect 7628 -5259 7674 -5247
rect 7724 -5167 7770 -5155
rect 7724 -5247 7730 -5167
rect 7764 -5247 7770 -5167
rect 7724 -5259 7770 -5247
rect 7820 -5167 7866 -5155
rect 7820 -5247 7826 -5167
rect 7860 -5247 7866 -5167
rect 7820 -5259 7866 -5247
rect 7916 -5167 7962 -5155
rect 7916 -5247 7922 -5167
rect 7956 -5247 7962 -5167
rect 7916 -5259 7962 -5247
rect 8012 -5167 8058 -5155
rect 8012 -5247 8018 -5167
rect 8052 -5247 8058 -5167
rect 8012 -5259 8058 -5247
rect 8108 -5167 8154 -5155
rect 8108 -5247 8114 -5167
rect 8148 -5247 8154 -5167
rect 8108 -5259 8154 -5247
rect 7138 -5291 7204 -5287
rect 7034 -5509 7080 -5337
rect 7135 -5343 7145 -5291
rect 7197 -5343 7207 -5291
rect 7138 -5347 7204 -5343
rect 7250 -5399 7284 -5259
rect 7330 -5291 7396 -5287
rect 7327 -5343 7337 -5291
rect 7389 -5343 7399 -5291
rect 7330 -5347 7396 -5343
rect 7442 -5399 7476 -5259
rect 7522 -5290 7588 -5287
rect 7520 -5342 7530 -5290
rect 7582 -5342 7592 -5290
rect 7522 -5347 7588 -5342
rect 7634 -5399 7668 -5259
rect 7714 -5290 7780 -5287
rect 7712 -5342 7722 -5290
rect 7774 -5342 7784 -5290
rect 7714 -5347 7780 -5342
rect 7826 -5399 7860 -5259
rect 7906 -5290 7972 -5287
rect 7904 -5342 7914 -5290
rect 7966 -5342 7976 -5290
rect 7906 -5347 7972 -5342
rect 8018 -5399 8052 -5259
rect 8098 -5290 8164 -5287
rect 8095 -5342 8105 -5290
rect 8157 -5342 8167 -5290
rect 8098 -5347 8164 -5342
rect 8298 -5399 8332 -5022
rect 8738 -5023 8802 -5022
rect 15792 -5040 15802 -4976
rect 15866 -4988 15876 -4976
rect 16154 -4988 16188 -4847
rect 16346 -4988 16380 -4847
rect 16538 -4988 16572 -4847
rect 16730 -4988 16764 -4847
rect 16922 -4988 16956 -4847
rect 17114 -4988 17148 -4847
rect 15866 -5022 17148 -4988
rect 15866 -5040 15876 -5022
rect 16034 -5137 16080 -5125
rect 8372 -5342 8382 -5290
rect 8434 -5342 8461 -5290
rect 16034 -5337 16040 -5137
rect 16074 -5337 16080 -5137
rect 16154 -5155 16188 -5022
rect 16346 -5155 16380 -5022
rect 16538 -5155 16572 -5022
rect 16730 -5155 16764 -5022
rect 16922 -5155 16956 -5022
rect 17114 -5155 17148 -5022
rect 17298 -4988 17332 -4425
rect 17372 -4535 17382 -4483
rect 17434 -4535 17461 -4483
rect 17826 -4988 17901 -3222
rect 17298 -5022 17901 -4988
rect 16148 -5167 16194 -5155
rect 16148 -5247 16154 -5167
rect 16188 -5247 16194 -5167
rect 16148 -5259 16194 -5247
rect 16244 -5167 16290 -5155
rect 16244 -5247 16250 -5167
rect 16284 -5247 16290 -5167
rect 16244 -5259 16290 -5247
rect 16340 -5167 16386 -5155
rect 16340 -5247 16346 -5167
rect 16380 -5247 16386 -5167
rect 16340 -5259 16386 -5247
rect 16436 -5167 16482 -5155
rect 16436 -5247 16442 -5167
rect 16476 -5247 16482 -5167
rect 16436 -5259 16482 -5247
rect 16532 -5167 16578 -5155
rect 16532 -5247 16538 -5167
rect 16572 -5247 16578 -5167
rect 16532 -5259 16578 -5247
rect 16628 -5167 16674 -5155
rect 16628 -5247 16634 -5167
rect 16668 -5247 16674 -5167
rect 16628 -5259 16674 -5247
rect 16724 -5167 16770 -5155
rect 16724 -5247 16730 -5167
rect 16764 -5247 16770 -5167
rect 16724 -5259 16770 -5247
rect 16820 -5167 16866 -5155
rect 16820 -5247 16826 -5167
rect 16860 -5247 16866 -5167
rect 16820 -5259 16866 -5247
rect 16916 -5167 16962 -5155
rect 16916 -5247 16922 -5167
rect 16956 -5247 16962 -5167
rect 16916 -5259 16962 -5247
rect 17012 -5167 17058 -5155
rect 17012 -5247 17018 -5167
rect 17052 -5247 17058 -5167
rect 17012 -5259 17058 -5247
rect 17108 -5167 17154 -5155
rect 17108 -5247 17114 -5167
rect 17148 -5247 17154 -5167
rect 17108 -5259 17154 -5247
rect 16138 -5291 16204 -5287
rect 7250 -5433 8332 -5399
rect 16034 -5509 16080 -5337
rect 16135 -5343 16145 -5291
rect 16197 -5343 16207 -5291
rect 16138 -5347 16204 -5343
rect 16250 -5399 16284 -5259
rect 16330 -5291 16396 -5287
rect 16327 -5343 16337 -5291
rect 16389 -5343 16399 -5291
rect 16330 -5347 16396 -5343
rect 16442 -5399 16476 -5259
rect 16522 -5290 16588 -5287
rect 16520 -5342 16530 -5290
rect 16582 -5342 16592 -5290
rect 16522 -5347 16588 -5342
rect 16634 -5399 16668 -5259
rect 16714 -5290 16780 -5287
rect 16712 -5342 16722 -5290
rect 16774 -5342 16784 -5290
rect 16714 -5347 16780 -5342
rect 16826 -5399 16860 -5259
rect 16906 -5290 16972 -5287
rect 16904 -5342 16914 -5290
rect 16966 -5342 16976 -5290
rect 16906 -5347 16972 -5342
rect 17018 -5399 17052 -5259
rect 17098 -5290 17164 -5287
rect 17095 -5342 17105 -5290
rect 17157 -5342 17167 -5290
rect 17098 -5347 17164 -5342
rect 17298 -5399 17332 -5022
rect 17372 -5342 17382 -5290
rect 17434 -5342 17461 -5290
rect 16250 -5433 17332 -5399
rect 7034 -6287 7080 -6109
rect 7250 -6225 8332 -6191
rect 7034 -6673 7040 -6287
rect 7074 -6673 7080 -6287
rect 7135 -6335 7145 -6283
rect 7197 -6335 7207 -6283
rect 7250 -6375 7284 -6225
rect 7327 -6335 7337 -6283
rect 7389 -6335 7399 -6283
rect 7442 -6375 7476 -6225
rect 7519 -6335 7529 -6283
rect 7581 -6335 7591 -6283
rect 7634 -6375 7668 -6225
rect 7711 -6335 7721 -6283
rect 7773 -6335 7783 -6283
rect 7826 -6375 7860 -6225
rect 7902 -6335 7912 -6283
rect 7964 -6335 7974 -6283
rect 8018 -6375 8052 -6225
rect 8095 -6335 8105 -6283
rect 8157 -6335 8167 -6283
rect 7148 -6387 7194 -6375
rect 7148 -6635 7154 -6387
rect 7188 -6635 7194 -6387
rect 7148 -6647 7194 -6635
rect 7244 -6387 7290 -6375
rect 7244 -6635 7250 -6387
rect 7284 -6635 7290 -6387
rect 7244 -6647 7290 -6635
rect 7340 -6387 7386 -6375
rect 7340 -6635 7346 -6387
rect 7380 -6635 7386 -6387
rect 7340 -6647 7386 -6635
rect 7436 -6387 7482 -6375
rect 7436 -6635 7442 -6387
rect 7476 -6635 7482 -6387
rect 7436 -6647 7482 -6635
rect 7532 -6387 7578 -6375
rect 7532 -6635 7538 -6387
rect 7572 -6635 7578 -6387
rect 7532 -6647 7578 -6635
rect 7628 -6387 7674 -6375
rect 7628 -6635 7634 -6387
rect 7668 -6635 7674 -6387
rect 7628 -6647 7674 -6635
rect 7724 -6387 7770 -6375
rect 7724 -6635 7730 -6387
rect 7764 -6635 7770 -6387
rect 7724 -6647 7770 -6635
rect 7820 -6387 7866 -6375
rect 7820 -6635 7826 -6387
rect 7860 -6635 7866 -6387
rect 7820 -6647 7866 -6635
rect 7916 -6387 7962 -6375
rect 7916 -6635 7922 -6387
rect 7956 -6635 7962 -6387
rect 7916 -6647 7962 -6635
rect 8012 -6387 8058 -6375
rect 8012 -6635 8018 -6387
rect 8052 -6635 8058 -6387
rect 8012 -6647 8058 -6635
rect 8108 -6387 8154 -6375
rect 8108 -6635 8114 -6387
rect 8148 -6635 8154 -6387
rect 8108 -6647 8154 -6635
rect 7034 -6685 7080 -6673
rect 7154 -6788 7188 -6647
rect 7346 -6788 7380 -6647
rect 7538 -6788 7572 -6647
rect 7730 -6788 7764 -6647
rect 7922 -6788 7956 -6647
rect 8114 -6773 8148 -6647
rect 8073 -6788 8083 -6773
rect 5608 -6822 8083 -6788
rect 4760 -6944 4770 -6891
rect 4823 -6944 4833 -6891
rect 4896 -6942 4906 -6889
rect 4959 -6942 4969 -6889
rect 5028 -6940 5038 -6887
rect 5091 -6940 5101 -6887
rect 7034 -6937 7080 -6925
rect 7034 -7137 7040 -6937
rect 7074 -7137 7080 -6937
rect 7154 -6955 7188 -6822
rect 7346 -6955 7380 -6822
rect 7538 -6955 7572 -6822
rect 7730 -6955 7764 -6822
rect 7922 -6955 7956 -6822
rect 8073 -6837 8083 -6822
rect 8147 -6837 8157 -6773
rect 8298 -6788 8332 -6225
rect 8372 -6335 8382 -6283
rect 8434 -6335 8461 -6283
rect 16034 -6287 16080 -6109
rect 16250 -6225 17332 -6191
rect 16034 -6673 16040 -6287
rect 16074 -6673 16080 -6287
rect 16135 -6335 16145 -6283
rect 16197 -6335 16207 -6283
rect 16250 -6375 16284 -6225
rect 16327 -6335 16337 -6283
rect 16389 -6335 16399 -6283
rect 16442 -6375 16476 -6225
rect 16519 -6335 16529 -6283
rect 16581 -6335 16591 -6283
rect 16634 -6375 16668 -6225
rect 16711 -6335 16721 -6283
rect 16773 -6335 16783 -6283
rect 16826 -6375 16860 -6225
rect 16902 -6335 16912 -6283
rect 16964 -6335 16974 -6283
rect 17018 -6375 17052 -6225
rect 17095 -6335 17105 -6283
rect 17157 -6335 17167 -6283
rect 16148 -6387 16194 -6375
rect 16148 -6635 16154 -6387
rect 16188 -6635 16194 -6387
rect 16148 -6647 16194 -6635
rect 16244 -6387 16290 -6375
rect 16244 -6635 16250 -6387
rect 16284 -6635 16290 -6387
rect 16244 -6647 16290 -6635
rect 16340 -6387 16386 -6375
rect 16340 -6635 16346 -6387
rect 16380 -6635 16386 -6387
rect 16340 -6647 16386 -6635
rect 16436 -6387 16482 -6375
rect 16436 -6635 16442 -6387
rect 16476 -6635 16482 -6387
rect 16436 -6647 16482 -6635
rect 16532 -6387 16578 -6375
rect 16532 -6635 16538 -6387
rect 16572 -6635 16578 -6387
rect 16532 -6647 16578 -6635
rect 16628 -6387 16674 -6375
rect 16628 -6635 16634 -6387
rect 16668 -6635 16674 -6387
rect 16628 -6647 16674 -6635
rect 16724 -6387 16770 -6375
rect 16724 -6635 16730 -6387
rect 16764 -6635 16770 -6387
rect 16724 -6647 16770 -6635
rect 16820 -6387 16866 -6375
rect 16820 -6635 16826 -6387
rect 16860 -6635 16866 -6387
rect 16820 -6647 16866 -6635
rect 16916 -6387 16962 -6375
rect 16916 -6635 16922 -6387
rect 16956 -6635 16962 -6387
rect 16916 -6647 16962 -6635
rect 17012 -6387 17058 -6375
rect 17012 -6635 17018 -6387
rect 17052 -6635 17058 -6387
rect 17012 -6647 17058 -6635
rect 17108 -6387 17154 -6375
rect 17108 -6635 17114 -6387
rect 17148 -6635 17154 -6387
rect 17108 -6647 17154 -6635
rect 16034 -6685 16080 -6673
rect 8590 -6788 8600 -6770
rect 8298 -6822 8600 -6788
rect 8114 -6955 8148 -6837
rect 7148 -6967 7194 -6955
rect 7148 -7047 7154 -6967
rect 7188 -7047 7194 -6967
rect 7148 -7059 7194 -7047
rect 7244 -6967 7290 -6955
rect 7244 -7047 7250 -6967
rect 7284 -7047 7290 -6967
rect 7244 -7059 7290 -7047
rect 7340 -6967 7386 -6955
rect 7340 -7047 7346 -6967
rect 7380 -7047 7386 -6967
rect 7340 -7059 7386 -7047
rect 7436 -6967 7482 -6955
rect 7436 -7047 7442 -6967
rect 7476 -7047 7482 -6967
rect 7436 -7059 7482 -7047
rect 7532 -6967 7578 -6955
rect 7532 -7047 7538 -6967
rect 7572 -7047 7578 -6967
rect 7532 -7059 7578 -7047
rect 7628 -6967 7674 -6955
rect 7628 -7047 7634 -6967
rect 7668 -7047 7674 -6967
rect 7628 -7059 7674 -7047
rect 7724 -6967 7770 -6955
rect 7724 -7047 7730 -6967
rect 7764 -7047 7770 -6967
rect 7724 -7059 7770 -7047
rect 7820 -6967 7866 -6955
rect 7820 -7047 7826 -6967
rect 7860 -7047 7866 -6967
rect 7820 -7059 7866 -7047
rect 7916 -6967 7962 -6955
rect 7916 -7047 7922 -6967
rect 7956 -7047 7962 -6967
rect 7916 -7059 7962 -7047
rect 8012 -6967 8058 -6955
rect 8012 -7047 8018 -6967
rect 8052 -7047 8058 -6967
rect 8012 -7059 8058 -7047
rect 8108 -6967 8154 -6955
rect 8108 -7047 8114 -6967
rect 8148 -7047 8154 -6967
rect 8108 -7059 8154 -7047
rect 7138 -7091 7204 -7087
rect 7034 -7309 7080 -7137
rect 7135 -7143 7145 -7091
rect 7197 -7143 7207 -7091
rect 7138 -7147 7204 -7143
rect 7250 -7199 7284 -7059
rect 7330 -7091 7396 -7087
rect 7327 -7143 7337 -7091
rect 7389 -7143 7399 -7091
rect 7330 -7147 7396 -7143
rect 7442 -7199 7476 -7059
rect 7522 -7090 7588 -7087
rect 7520 -7142 7530 -7090
rect 7582 -7142 7592 -7090
rect 7522 -7147 7588 -7142
rect 7634 -7199 7668 -7059
rect 7714 -7090 7780 -7087
rect 7712 -7142 7722 -7090
rect 7774 -7142 7784 -7090
rect 7714 -7147 7780 -7142
rect 7826 -7199 7860 -7059
rect 7906 -7090 7972 -7087
rect 7904 -7142 7914 -7090
rect 7966 -7142 7976 -7090
rect 7906 -7147 7972 -7142
rect 8018 -7199 8052 -7059
rect 8098 -7090 8164 -7087
rect 8095 -7142 8105 -7090
rect 8157 -7142 8167 -7090
rect 8098 -7147 8164 -7142
rect 8298 -7199 8332 -6822
rect 8590 -6834 8600 -6822
rect 8664 -6834 8674 -6770
rect 15810 -6832 15820 -6768
rect 15884 -6788 15894 -6768
rect 16154 -6788 16188 -6647
rect 16346 -6788 16380 -6647
rect 16538 -6788 16572 -6647
rect 16730 -6788 16764 -6647
rect 16922 -6788 16956 -6647
rect 17114 -6788 17148 -6647
rect 15884 -6822 17148 -6788
rect 15884 -6832 15894 -6822
rect 16034 -6937 16080 -6925
rect 8372 -7142 8382 -7090
rect 8434 -7142 8461 -7090
rect 16034 -7137 16040 -6937
rect 16074 -7137 16080 -6937
rect 16154 -6955 16188 -6822
rect 16346 -6955 16380 -6822
rect 16538 -6955 16572 -6822
rect 16730 -6955 16764 -6822
rect 16922 -6955 16956 -6822
rect 17114 -6955 17148 -6822
rect 17298 -6788 17332 -6225
rect 17372 -6335 17382 -6283
rect 17434 -6335 17461 -6283
rect 17826 -6521 17901 -5022
rect 17821 -6585 17831 -6521
rect 17895 -6585 17905 -6521
rect 18337 -6788 18412 2178
rect 17298 -6822 18412 -6788
rect 16148 -6967 16194 -6955
rect 16148 -7047 16154 -6967
rect 16188 -7047 16194 -6967
rect 16148 -7059 16194 -7047
rect 16244 -6967 16290 -6955
rect 16244 -7047 16250 -6967
rect 16284 -7047 16290 -6967
rect 16244 -7059 16290 -7047
rect 16340 -6967 16386 -6955
rect 16340 -7047 16346 -6967
rect 16380 -7047 16386 -6967
rect 16340 -7059 16386 -7047
rect 16436 -6967 16482 -6955
rect 16436 -7047 16442 -6967
rect 16476 -7047 16482 -6967
rect 16436 -7059 16482 -7047
rect 16532 -6967 16578 -6955
rect 16532 -7047 16538 -6967
rect 16572 -7047 16578 -6967
rect 16532 -7059 16578 -7047
rect 16628 -6967 16674 -6955
rect 16628 -7047 16634 -6967
rect 16668 -7047 16674 -6967
rect 16628 -7059 16674 -7047
rect 16724 -6967 16770 -6955
rect 16724 -7047 16730 -6967
rect 16764 -7047 16770 -6967
rect 16724 -7059 16770 -7047
rect 16820 -6967 16866 -6955
rect 16820 -7047 16826 -6967
rect 16860 -7047 16866 -6967
rect 16820 -7059 16866 -7047
rect 16916 -6967 16962 -6955
rect 16916 -7047 16922 -6967
rect 16956 -7047 16962 -6967
rect 16916 -7059 16962 -7047
rect 17012 -6967 17058 -6955
rect 17012 -7047 17018 -6967
rect 17052 -7047 17058 -6967
rect 17012 -7059 17058 -7047
rect 17108 -6967 17154 -6955
rect 17108 -7047 17114 -6967
rect 17148 -7047 17154 -6967
rect 17108 -7059 17154 -7047
rect 16138 -7091 16204 -7087
rect 7250 -7233 8332 -7199
rect 16034 -7309 16080 -7137
rect 16135 -7143 16145 -7091
rect 16197 -7143 16207 -7091
rect 16138 -7147 16204 -7143
rect 16250 -7199 16284 -7059
rect 16330 -7091 16396 -7087
rect 16327 -7143 16337 -7091
rect 16389 -7143 16399 -7091
rect 16330 -7147 16396 -7143
rect 16442 -7199 16476 -7059
rect 16522 -7090 16588 -7087
rect 16520 -7142 16530 -7090
rect 16582 -7142 16592 -7090
rect 16522 -7147 16588 -7142
rect 16634 -7199 16668 -7059
rect 16714 -7090 16780 -7087
rect 16712 -7142 16722 -7090
rect 16774 -7142 16784 -7090
rect 16714 -7147 16780 -7142
rect 16826 -7199 16860 -7059
rect 16906 -7090 16972 -7087
rect 16904 -7142 16914 -7090
rect 16966 -7142 16976 -7090
rect 16906 -7147 16972 -7142
rect 17018 -7199 17052 -7059
rect 17098 -7090 17164 -7087
rect 17095 -7142 17105 -7090
rect 17157 -7142 17167 -7090
rect 17098 -7147 17164 -7142
rect 17298 -7199 17332 -6822
rect 17372 -7142 17382 -7090
rect 17434 -7142 17461 -7090
rect 16250 -7233 17332 -7199
rect -3883 -7697 -3873 -7691
rect -5629 -7731 -3873 -7697
rect -5628 -7862 -5594 -7731
rect -5544 -7774 -5500 -7731
rect -5560 -7790 -5484 -7774
rect -5560 -7824 -5544 -7790
rect -5500 -7824 -5484 -7790
rect -5560 -7830 -5484 -7824
rect -5450 -7862 -5416 -7731
rect -5366 -7774 -5322 -7731
rect -5188 -7774 -5144 -7731
rect -5382 -7790 -5306 -7774
rect -5382 -7824 -5366 -7790
rect -5322 -7824 -5306 -7790
rect -5382 -7830 -5306 -7824
rect -5204 -7790 -5128 -7774
rect -5204 -7824 -5188 -7790
rect -5144 -7824 -5128 -7790
rect -5204 -7830 -5128 -7824
rect -5094 -7862 -5060 -7731
rect -5010 -7774 -4966 -7731
rect -4832 -7774 -4788 -7731
rect -5026 -7790 -4950 -7774
rect -5026 -7824 -5010 -7790
rect -4966 -7824 -4950 -7790
rect -5026 -7830 -4950 -7824
rect -4848 -7790 -4772 -7774
rect -4848 -7824 -4832 -7790
rect -4788 -7824 -4772 -7790
rect -4848 -7830 -4772 -7824
rect -4738 -7862 -4704 -7731
rect -4654 -7774 -4610 -7731
rect -4476 -7774 -4432 -7731
rect -4670 -7790 -4594 -7774
rect -4670 -7824 -4654 -7790
rect -4610 -7824 -4594 -7790
rect -4670 -7830 -4594 -7824
rect -4492 -7790 -4416 -7774
rect -4492 -7824 -4476 -7790
rect -4432 -7824 -4416 -7790
rect -4492 -7830 -4416 -7824
rect -4382 -7862 -4348 -7731
rect -4298 -7774 -4254 -7731
rect -3883 -7743 -3873 -7731
rect -3821 -7743 -3811 -7691
rect -4314 -7790 -4238 -7774
rect -4314 -7824 -4298 -7790
rect -4254 -7824 -4238 -7790
rect -4314 -7830 -4238 -7824
rect -4136 -7790 -4060 -7774
rect -3741 -7790 -3731 -7785
rect -4136 -7824 -4120 -7790
rect -4076 -7824 -4060 -7790
rect -4136 -7830 -4060 -7824
rect -4026 -7824 -3731 -7790
rect -4026 -7862 -3992 -7824
rect -3741 -7837 -3731 -7824
rect -3679 -7837 -3669 -7785
rect -3551 -7840 -3541 -7788
rect -3489 -7840 -3479 -7788
rect -5634 -7874 -5588 -7862
rect -5634 -8130 -5628 -7874
rect -5594 -8130 -5588 -7874
rect -5634 -8142 -5588 -8130
rect -5456 -7874 -5410 -7862
rect -5456 -8130 -5450 -7874
rect -5416 -8130 -5410 -7874
rect -5456 -8142 -5410 -8130
rect -5278 -7874 -5232 -7862
rect -5278 -8130 -5272 -7874
rect -5238 -8130 -5232 -7874
rect -5278 -8142 -5232 -8130
rect -5100 -7874 -5054 -7862
rect -5100 -8130 -5094 -7874
rect -5060 -8130 -5054 -7874
rect -5100 -8142 -5054 -8130
rect -4922 -7874 -4876 -7862
rect -4922 -8130 -4916 -7874
rect -4882 -8130 -4876 -7874
rect -4922 -8142 -4876 -8130
rect -4744 -7874 -4698 -7862
rect -4744 -8130 -4738 -7874
rect -4704 -8130 -4698 -7874
rect -4744 -8142 -4698 -8130
rect -4566 -7874 -4520 -7862
rect -4566 -8130 -4560 -7874
rect -4526 -8130 -4520 -7874
rect -4566 -8142 -4520 -8130
rect -4388 -7874 -4342 -7862
rect -4388 -8130 -4382 -7874
rect -4348 -8130 -4342 -7874
rect -4388 -8142 -4342 -8130
rect -4210 -7874 -4164 -7862
rect -4210 -8130 -4204 -7874
rect -4170 -8130 -4164 -7874
rect -4210 -8142 -4164 -8130
rect -4032 -7874 -3986 -7862
rect -4032 -8130 -4026 -7874
rect -3992 -8130 -3986 -7874
rect -4032 -8142 -3986 -8130
rect -5628 -8412 -5594 -8142
rect -5560 -8180 -5484 -8174
rect -5560 -8214 -5544 -8180
rect -5500 -8214 -5484 -8180
rect -5560 -8230 -5484 -8214
rect -5544 -8324 -5500 -8230
rect -5560 -8340 -5484 -8324
rect -5560 -8374 -5544 -8340
rect -5500 -8374 -5484 -8340
rect -5560 -8380 -5484 -8374
rect -5450 -8412 -5416 -8142
rect -5382 -8180 -5306 -8174
rect -5382 -8214 -5366 -8180
rect -5322 -8214 -5306 -8180
rect -5382 -8230 -5306 -8214
rect -5366 -8324 -5322 -8230
rect -5382 -8340 -5306 -8324
rect -5382 -8374 -5366 -8340
rect -5322 -8374 -5306 -8340
rect -5382 -8380 -5306 -8374
rect -5272 -8412 -5238 -8142
rect -5204 -8180 -5128 -8174
rect -5204 -8214 -5188 -8180
rect -5144 -8214 -5128 -8180
rect -5204 -8230 -5128 -8214
rect -5188 -8324 -5144 -8230
rect -5204 -8340 -5128 -8324
rect -5204 -8374 -5188 -8340
rect -5144 -8374 -5128 -8340
rect -5204 -8380 -5128 -8374
rect -5094 -8412 -5060 -8142
rect -5026 -8180 -4950 -8174
rect -5026 -8214 -5010 -8180
rect -4966 -8214 -4950 -8180
rect -5026 -8230 -4950 -8214
rect -5010 -8324 -4966 -8230
rect -5026 -8340 -4950 -8324
rect -5026 -8374 -5010 -8340
rect -4966 -8374 -4950 -8340
rect -5026 -8380 -4950 -8374
rect -4916 -8412 -4882 -8142
rect -4848 -8180 -4772 -8174
rect -4848 -8214 -4832 -8180
rect -4788 -8214 -4772 -8180
rect -4848 -8230 -4772 -8214
rect -4832 -8324 -4788 -8230
rect -4848 -8340 -4772 -8324
rect -4848 -8374 -4832 -8340
rect -4788 -8374 -4772 -8340
rect -4848 -8380 -4772 -8374
rect -4738 -8412 -4704 -8142
rect -4670 -8180 -4594 -8174
rect -4670 -8214 -4654 -8180
rect -4610 -8214 -4594 -8180
rect -4670 -8230 -4594 -8214
rect -4654 -8324 -4610 -8230
rect -4670 -8340 -4594 -8324
rect -4670 -8374 -4654 -8340
rect -4610 -8374 -4594 -8340
rect -4670 -8380 -4594 -8374
rect -4560 -8412 -4526 -8142
rect -4492 -8180 -4416 -8174
rect -4492 -8214 -4476 -8180
rect -4432 -8214 -4416 -8180
rect -4492 -8230 -4416 -8214
rect -4476 -8324 -4432 -8230
rect -4492 -8340 -4416 -8324
rect -4492 -8374 -4476 -8340
rect -4432 -8374 -4416 -8340
rect -4492 -8380 -4416 -8374
rect -4382 -8412 -4348 -8142
rect -4314 -8180 -4238 -8174
rect -4314 -8214 -4298 -8180
rect -4254 -8214 -4238 -8180
rect -4314 -8230 -4238 -8214
rect -4298 -8324 -4254 -8230
rect -4314 -8340 -4238 -8324
rect -4314 -8374 -4298 -8340
rect -4254 -8374 -4238 -8340
rect -4314 -8380 -4238 -8374
rect -4204 -8412 -4170 -8142
rect -4136 -8180 -4060 -8174
rect -4136 -8214 -4120 -8180
rect -4076 -8214 -4060 -8180
rect -4136 -8230 -4060 -8214
rect -4120 -8324 -4076 -8230
rect -4136 -8340 -4060 -8324
rect -4136 -8374 -4120 -8340
rect -4076 -8374 -4060 -8340
rect -4136 -8380 -4060 -8374
rect -4026 -8412 -3992 -8142
rect -5634 -8424 -5588 -8412
rect -5634 -8680 -5628 -8424
rect -5594 -8680 -5588 -8424
rect -5634 -8692 -5588 -8680
rect -5456 -8424 -5410 -8412
rect -5456 -8680 -5450 -8424
rect -5416 -8680 -5410 -8424
rect -5456 -8692 -5410 -8680
rect -5278 -8424 -5232 -8412
rect -5278 -8680 -5272 -8424
rect -5238 -8680 -5232 -8424
rect -5278 -8692 -5232 -8680
rect -5100 -8424 -5054 -8412
rect -5100 -8680 -5094 -8424
rect -5060 -8680 -5054 -8424
rect -5100 -8692 -5054 -8680
rect -4922 -8424 -4876 -8412
rect -4922 -8680 -4916 -8424
rect -4882 -8680 -4876 -8424
rect -4922 -8692 -4876 -8680
rect -4744 -8424 -4698 -8412
rect -4744 -8680 -4738 -8424
rect -4704 -8680 -4698 -8424
rect -4744 -8692 -4698 -8680
rect -4566 -8424 -4520 -8412
rect -4566 -8680 -4560 -8424
rect -4526 -8680 -4520 -8424
rect -4566 -8692 -4520 -8680
rect -4388 -8424 -4342 -8412
rect -4388 -8680 -4382 -8424
rect -4348 -8680 -4342 -8424
rect -4388 -8692 -4342 -8680
rect -4210 -8424 -4164 -8412
rect -4210 -8680 -4204 -8424
rect -4170 -8680 -4164 -8424
rect -4210 -8692 -4164 -8680
rect -4032 -8424 -3986 -8412
rect -4032 -8680 -4026 -8424
rect -3992 -8680 -3986 -8424
rect -4032 -8692 -3986 -8680
rect -5628 -8962 -5594 -8692
rect -5560 -8730 -5484 -8724
rect -5560 -8764 -5544 -8730
rect -5500 -8764 -5484 -8730
rect -5560 -8780 -5484 -8764
rect -5544 -8874 -5500 -8780
rect -5560 -8890 -5484 -8874
rect -5560 -8924 -5544 -8890
rect -5500 -8924 -5484 -8890
rect -5560 -8930 -5484 -8924
rect -5450 -8962 -5416 -8692
rect -5382 -8730 -5306 -8724
rect -5382 -8764 -5366 -8730
rect -5322 -8764 -5306 -8730
rect -5382 -8780 -5306 -8764
rect -5366 -8874 -5322 -8780
rect -5382 -8890 -5306 -8874
rect -5382 -8924 -5366 -8890
rect -5322 -8924 -5306 -8890
rect -5382 -8930 -5306 -8924
rect -5272 -8962 -5238 -8692
rect -5204 -8730 -5128 -8724
rect -5204 -8764 -5188 -8730
rect -5144 -8764 -5128 -8730
rect -5204 -8780 -5128 -8764
rect -5188 -8874 -5144 -8780
rect -5204 -8890 -5128 -8874
rect -5204 -8924 -5188 -8890
rect -5144 -8924 -5128 -8890
rect -5204 -8930 -5128 -8924
rect -5094 -8962 -5060 -8692
rect -5026 -8730 -4950 -8724
rect -5026 -8764 -5010 -8730
rect -4966 -8764 -4950 -8730
rect -5026 -8780 -4950 -8764
rect -5010 -8874 -4966 -8780
rect -5026 -8890 -4950 -8874
rect -5026 -8924 -5010 -8890
rect -4966 -8924 -4950 -8890
rect -5026 -8930 -4950 -8924
rect -4916 -8962 -4882 -8692
rect -4848 -8730 -4772 -8724
rect -4848 -8764 -4832 -8730
rect -4788 -8764 -4772 -8730
rect -4848 -8780 -4772 -8764
rect -4832 -8874 -4788 -8780
rect -4848 -8890 -4772 -8874
rect -4848 -8924 -4832 -8890
rect -4788 -8924 -4772 -8890
rect -4848 -8930 -4772 -8924
rect -4738 -8962 -4704 -8692
rect -4670 -8730 -4594 -8724
rect -4670 -8764 -4654 -8730
rect -4610 -8764 -4594 -8730
rect -4670 -8780 -4594 -8764
rect -4654 -8874 -4610 -8780
rect -4670 -8890 -4594 -8874
rect -4670 -8924 -4654 -8890
rect -4610 -8924 -4594 -8890
rect -4670 -8930 -4594 -8924
rect -4560 -8962 -4526 -8692
rect -4492 -8730 -4416 -8724
rect -4492 -8764 -4476 -8730
rect -4432 -8764 -4416 -8730
rect -4492 -8780 -4416 -8764
rect -4476 -8874 -4432 -8780
rect -4492 -8890 -4416 -8874
rect -4492 -8924 -4476 -8890
rect -4432 -8924 -4416 -8890
rect -4492 -8930 -4416 -8924
rect -4382 -8962 -4348 -8692
rect -4314 -8730 -4238 -8724
rect -4314 -8764 -4298 -8730
rect -4254 -8764 -4238 -8730
rect -4314 -8780 -4238 -8764
rect -4298 -8874 -4254 -8780
rect -4314 -8890 -4238 -8874
rect -4314 -8924 -4298 -8890
rect -4254 -8924 -4238 -8890
rect -4314 -8930 -4238 -8924
rect -4204 -8962 -4170 -8692
rect -4136 -8730 -4060 -8724
rect -4136 -8764 -4120 -8730
rect -4076 -8764 -4060 -8730
rect -4136 -8780 -4060 -8764
rect -4120 -8874 -4076 -8780
rect -4136 -8890 -4060 -8874
rect -4136 -8924 -4120 -8890
rect -4076 -8924 -4060 -8890
rect -4136 -8930 -4060 -8924
rect -4026 -8962 -3992 -8692
rect -5634 -8974 -5588 -8962
rect -5634 -9230 -5628 -8974
rect -5594 -9230 -5588 -8974
rect -5634 -9242 -5588 -9230
rect -5456 -8974 -5410 -8962
rect -5456 -9230 -5450 -8974
rect -5416 -9230 -5410 -8974
rect -5456 -9242 -5410 -9230
rect -5278 -8974 -5232 -8962
rect -5278 -9230 -5272 -8974
rect -5238 -9230 -5232 -8974
rect -5278 -9242 -5232 -9230
rect -5100 -8974 -5054 -8962
rect -5100 -9230 -5094 -8974
rect -5060 -9230 -5054 -8974
rect -5100 -9242 -5054 -9230
rect -4922 -8974 -4876 -8962
rect -4922 -9230 -4916 -8974
rect -4882 -9230 -4876 -8974
rect -4922 -9242 -4876 -9230
rect -4744 -8974 -4698 -8962
rect -4744 -9230 -4738 -8974
rect -4704 -9230 -4698 -8974
rect -4744 -9242 -4698 -9230
rect -4566 -8974 -4520 -8962
rect -4566 -9230 -4560 -8974
rect -4526 -9230 -4520 -8974
rect -4566 -9242 -4520 -9230
rect -4388 -8974 -4342 -8962
rect -4388 -9230 -4382 -8974
rect -4348 -9230 -4342 -8974
rect -4388 -9242 -4342 -9230
rect -4210 -8974 -4164 -8962
rect -4210 -9230 -4204 -8974
rect -4170 -9230 -4164 -8974
rect -4210 -9242 -4164 -9230
rect -4032 -8974 -3986 -8962
rect -4032 -9230 -4026 -8974
rect -3992 -9230 -3986 -8974
rect -4032 -9242 -3986 -9230
rect -5628 -9512 -5594 -9242
rect -5560 -9280 -5484 -9274
rect -5560 -9314 -5544 -9280
rect -5500 -9314 -5484 -9280
rect -5560 -9330 -5484 -9314
rect -5544 -9424 -5500 -9330
rect -5560 -9440 -5484 -9424
rect -5560 -9474 -5544 -9440
rect -5500 -9474 -5484 -9440
rect -5560 -9480 -5484 -9474
rect -5450 -9512 -5416 -9242
rect -5382 -9280 -5306 -9274
rect -5382 -9314 -5366 -9280
rect -5322 -9314 -5306 -9280
rect -5382 -9330 -5306 -9314
rect -5366 -9424 -5322 -9330
rect -5382 -9440 -5306 -9424
rect -5382 -9474 -5366 -9440
rect -5322 -9474 -5306 -9440
rect -5382 -9480 -5306 -9474
rect -5272 -9512 -5238 -9242
rect -5204 -9280 -5128 -9274
rect -5204 -9314 -5188 -9280
rect -5144 -9314 -5128 -9280
rect -5204 -9330 -5128 -9314
rect -5188 -9424 -5144 -9330
rect -5204 -9440 -5128 -9424
rect -5204 -9474 -5188 -9440
rect -5144 -9474 -5128 -9440
rect -5204 -9480 -5128 -9474
rect -5094 -9512 -5060 -9242
rect -5026 -9280 -4950 -9274
rect -5026 -9314 -5010 -9280
rect -4966 -9314 -4950 -9280
rect -5026 -9330 -4950 -9314
rect -5010 -9424 -4966 -9330
rect -5026 -9440 -4950 -9424
rect -5026 -9474 -5010 -9440
rect -4966 -9474 -4950 -9440
rect -5026 -9480 -4950 -9474
rect -4916 -9512 -4882 -9242
rect -4848 -9280 -4772 -9274
rect -4848 -9314 -4832 -9280
rect -4788 -9314 -4772 -9280
rect -4848 -9330 -4772 -9314
rect -4832 -9424 -4788 -9330
rect -4848 -9440 -4772 -9424
rect -4848 -9474 -4832 -9440
rect -4788 -9474 -4772 -9440
rect -4848 -9480 -4772 -9474
rect -4738 -9512 -4704 -9242
rect -4670 -9280 -4594 -9274
rect -4670 -9314 -4654 -9280
rect -4610 -9314 -4594 -9280
rect -4670 -9330 -4594 -9314
rect -4654 -9424 -4610 -9330
rect -4670 -9440 -4594 -9424
rect -4670 -9474 -4654 -9440
rect -4610 -9474 -4594 -9440
rect -4670 -9480 -4594 -9474
rect -4560 -9512 -4526 -9242
rect -4492 -9280 -4416 -9274
rect -4492 -9314 -4476 -9280
rect -4432 -9314 -4416 -9280
rect -4492 -9330 -4416 -9314
rect -4476 -9424 -4432 -9330
rect -4492 -9440 -4416 -9424
rect -4492 -9474 -4476 -9440
rect -4432 -9474 -4416 -9440
rect -4492 -9480 -4416 -9474
rect -4382 -9512 -4348 -9242
rect -4314 -9280 -4238 -9274
rect -4314 -9314 -4298 -9280
rect -4254 -9314 -4238 -9280
rect -4314 -9330 -4238 -9314
rect -4298 -9424 -4254 -9330
rect -4314 -9440 -4238 -9424
rect -4314 -9474 -4298 -9440
rect -4254 -9474 -4238 -9440
rect -4314 -9480 -4238 -9474
rect -4204 -9512 -4170 -9242
rect -4136 -9280 -4060 -9274
rect -4136 -9314 -4120 -9280
rect -4076 -9314 -4060 -9280
rect -4136 -9330 -4060 -9314
rect -4120 -9424 -4076 -9330
rect -4136 -9440 -4060 -9424
rect -4136 -9474 -4120 -9440
rect -4076 -9474 -4060 -9440
rect -4136 -9480 -4060 -9474
rect -4026 -9512 -3992 -9242
rect -5634 -9524 -5588 -9512
rect -5634 -9780 -5628 -9524
rect -5594 -9780 -5588 -9524
rect -5634 -9792 -5588 -9780
rect -5456 -9524 -5410 -9512
rect -5456 -9780 -5450 -9524
rect -5416 -9780 -5410 -9524
rect -5456 -9792 -5410 -9780
rect -5278 -9524 -5232 -9512
rect -5278 -9780 -5272 -9524
rect -5238 -9780 -5232 -9524
rect -5278 -9792 -5232 -9780
rect -5100 -9524 -5054 -9512
rect -5100 -9780 -5094 -9524
rect -5060 -9780 -5054 -9524
rect -5100 -9792 -5054 -9780
rect -4922 -9524 -4876 -9512
rect -4922 -9780 -4916 -9524
rect -4882 -9780 -4876 -9524
rect -4922 -9792 -4876 -9780
rect -4744 -9524 -4698 -9512
rect -4744 -9780 -4738 -9524
rect -4704 -9780 -4698 -9524
rect -4744 -9792 -4698 -9780
rect -4566 -9524 -4520 -9512
rect -4566 -9780 -4560 -9524
rect -4526 -9780 -4520 -9524
rect -4566 -9792 -4520 -9780
rect -4388 -9524 -4342 -9512
rect -4388 -9780 -4382 -9524
rect -4348 -9780 -4342 -9524
rect -4388 -9792 -4342 -9780
rect -4210 -9524 -4164 -9512
rect -4210 -9780 -4204 -9524
rect -4170 -9780 -4164 -9524
rect -4210 -9792 -4164 -9780
rect -4032 -9524 -3986 -9512
rect -4032 -9780 -4026 -9524
rect -3992 -9780 -3986 -9524
rect -4032 -9792 -3986 -9780
rect -5628 -10062 -5594 -9792
rect -5560 -9830 -5484 -9824
rect -5560 -9864 -5544 -9830
rect -5500 -9864 -5484 -9830
rect -5560 -9880 -5484 -9864
rect -5544 -9974 -5500 -9880
rect -5560 -9990 -5484 -9974
rect -5560 -10024 -5544 -9990
rect -5500 -10024 -5484 -9990
rect -5560 -10030 -5484 -10024
rect -5450 -10062 -5416 -9792
rect -5382 -9830 -5306 -9824
rect -5382 -9864 -5366 -9830
rect -5322 -9864 -5306 -9830
rect -5382 -9880 -5306 -9864
rect -5366 -9974 -5322 -9880
rect -5382 -9990 -5306 -9974
rect -5382 -10024 -5366 -9990
rect -5322 -10024 -5306 -9990
rect -5382 -10030 -5306 -10024
rect -5272 -10062 -5238 -9792
rect -5204 -9830 -5128 -9824
rect -5204 -9864 -5188 -9830
rect -5144 -9864 -5128 -9830
rect -5204 -9880 -5128 -9864
rect -5188 -9974 -5144 -9880
rect -5204 -9990 -5128 -9974
rect -5204 -10024 -5188 -9990
rect -5144 -10024 -5128 -9990
rect -5204 -10030 -5128 -10024
rect -5094 -10062 -5060 -9792
rect -5026 -9830 -4950 -9824
rect -5026 -9864 -5010 -9830
rect -4966 -9864 -4950 -9830
rect -5026 -9880 -4950 -9864
rect -5010 -9974 -4966 -9880
rect -5026 -9990 -4950 -9974
rect -5026 -10024 -5010 -9990
rect -4966 -10024 -4950 -9990
rect -5026 -10030 -4950 -10024
rect -4916 -10062 -4882 -9792
rect -4848 -9830 -4772 -9824
rect -4848 -9864 -4832 -9830
rect -4788 -9864 -4772 -9830
rect -4848 -9880 -4772 -9864
rect -4832 -9974 -4788 -9880
rect -4848 -9990 -4772 -9974
rect -4848 -10024 -4832 -9990
rect -4788 -10024 -4772 -9990
rect -4848 -10030 -4772 -10024
rect -4738 -10062 -4704 -9792
rect -4670 -9830 -4594 -9824
rect -4670 -9864 -4654 -9830
rect -4610 -9864 -4594 -9830
rect -4670 -9880 -4594 -9864
rect -4654 -9974 -4610 -9880
rect -4670 -9990 -4594 -9974
rect -4670 -10024 -4654 -9990
rect -4610 -10024 -4594 -9990
rect -4670 -10030 -4594 -10024
rect -4560 -10062 -4526 -9792
rect -4492 -9830 -4416 -9824
rect -4492 -9864 -4476 -9830
rect -4432 -9864 -4416 -9830
rect -4492 -9880 -4416 -9864
rect -4476 -9974 -4432 -9880
rect -4492 -9990 -4416 -9974
rect -4492 -10024 -4476 -9990
rect -4432 -10024 -4416 -9990
rect -4492 -10030 -4416 -10024
rect -4382 -10062 -4348 -9792
rect -4314 -9830 -4238 -9824
rect -4314 -9864 -4298 -9830
rect -4254 -9864 -4238 -9830
rect -4314 -9880 -4238 -9864
rect -4298 -9974 -4254 -9880
rect -4314 -9990 -4238 -9974
rect -4314 -10024 -4298 -9990
rect -4254 -10024 -4238 -9990
rect -4314 -10030 -4238 -10024
rect -4204 -10062 -4170 -9792
rect -4136 -9830 -4060 -9824
rect -4136 -9864 -4120 -9830
rect -4076 -9864 -4060 -9830
rect -4136 -9880 -4060 -9864
rect -4120 -9974 -4076 -9880
rect -4136 -9990 -4060 -9974
rect -4136 -10024 -4120 -9990
rect -4076 -10024 -4060 -9990
rect -4136 -10030 -4060 -10024
rect -4026 -10062 -3992 -9792
rect -5634 -10074 -5588 -10062
rect -5634 -10330 -5628 -10074
rect -5594 -10330 -5588 -10074
rect -5634 -10342 -5588 -10330
rect -5456 -10074 -5410 -10062
rect -5456 -10330 -5450 -10074
rect -5416 -10330 -5410 -10074
rect -5456 -10342 -5410 -10330
rect -5278 -10074 -5232 -10062
rect -5278 -10330 -5272 -10074
rect -5238 -10330 -5232 -10074
rect -5278 -10342 -5232 -10330
rect -5100 -10074 -5054 -10062
rect -5100 -10330 -5094 -10074
rect -5060 -10330 -5054 -10074
rect -5100 -10342 -5054 -10330
rect -4922 -10074 -4876 -10062
rect -4922 -10330 -4916 -10074
rect -4882 -10330 -4876 -10074
rect -4922 -10342 -4876 -10330
rect -4744 -10074 -4698 -10062
rect -4744 -10330 -4738 -10074
rect -4704 -10330 -4698 -10074
rect -4744 -10342 -4698 -10330
rect -4566 -10074 -4520 -10062
rect -4566 -10330 -4560 -10074
rect -4526 -10330 -4520 -10074
rect -4566 -10342 -4520 -10330
rect -4388 -10074 -4342 -10062
rect -4388 -10330 -4382 -10074
rect -4348 -10330 -4342 -10074
rect -4388 -10342 -4342 -10330
rect -4210 -10074 -4164 -10062
rect -4210 -10330 -4204 -10074
rect -4170 -10330 -4164 -10074
rect -4210 -10342 -4164 -10330
rect -4032 -10074 -3986 -10062
rect -4032 -10330 -4026 -10074
rect -3992 -10330 -3986 -10074
rect -4032 -10342 -3986 -10330
rect -5628 -10612 -5594 -10342
rect -5560 -10380 -5484 -10374
rect -5560 -10414 -5544 -10380
rect -5500 -10414 -5484 -10380
rect -5560 -10430 -5484 -10414
rect -5544 -10524 -5500 -10430
rect -5560 -10540 -5484 -10524
rect -5560 -10574 -5544 -10540
rect -5500 -10574 -5484 -10540
rect -5560 -10580 -5484 -10574
rect -5450 -10612 -5416 -10342
rect -5382 -10380 -5306 -10374
rect -5382 -10414 -5366 -10380
rect -5322 -10414 -5306 -10380
rect -5382 -10430 -5306 -10414
rect -5366 -10524 -5322 -10430
rect -5382 -10540 -5306 -10524
rect -5382 -10574 -5366 -10540
rect -5322 -10574 -5306 -10540
rect -5382 -10580 -5306 -10574
rect -5272 -10612 -5238 -10342
rect -5204 -10380 -5128 -10374
rect -5204 -10414 -5188 -10380
rect -5144 -10414 -5128 -10380
rect -5204 -10430 -5128 -10414
rect -5188 -10524 -5144 -10430
rect -5204 -10540 -5128 -10524
rect -5204 -10574 -5188 -10540
rect -5144 -10574 -5128 -10540
rect -5204 -10580 -5128 -10574
rect -5094 -10612 -5060 -10342
rect -5026 -10380 -4950 -10374
rect -5026 -10414 -5010 -10380
rect -4966 -10414 -4950 -10380
rect -5026 -10430 -4950 -10414
rect -5010 -10524 -4966 -10430
rect -5026 -10540 -4950 -10524
rect -5026 -10574 -5010 -10540
rect -4966 -10574 -4950 -10540
rect -5026 -10580 -4950 -10574
rect -4916 -10612 -4882 -10342
rect -4848 -10380 -4772 -10374
rect -4848 -10414 -4832 -10380
rect -4788 -10414 -4772 -10380
rect -4848 -10430 -4772 -10414
rect -4832 -10524 -4788 -10430
rect -4848 -10540 -4772 -10524
rect -4848 -10574 -4832 -10540
rect -4788 -10574 -4772 -10540
rect -4848 -10580 -4772 -10574
rect -4738 -10612 -4704 -10342
rect -4670 -10380 -4594 -10374
rect -4670 -10414 -4654 -10380
rect -4610 -10414 -4594 -10380
rect -4670 -10430 -4594 -10414
rect -4654 -10524 -4610 -10430
rect -4670 -10540 -4594 -10524
rect -4670 -10574 -4654 -10540
rect -4610 -10574 -4594 -10540
rect -4670 -10580 -4594 -10574
rect -4560 -10612 -4526 -10342
rect -4492 -10380 -4416 -10374
rect -4492 -10414 -4476 -10380
rect -4432 -10414 -4416 -10380
rect -4492 -10430 -4416 -10414
rect -4476 -10524 -4432 -10430
rect -4492 -10540 -4416 -10524
rect -4492 -10574 -4476 -10540
rect -4432 -10574 -4416 -10540
rect -4492 -10580 -4416 -10574
rect -4382 -10612 -4348 -10342
rect -4314 -10380 -4238 -10374
rect -4314 -10414 -4298 -10380
rect -4254 -10414 -4238 -10380
rect -4314 -10430 -4238 -10414
rect -4298 -10524 -4254 -10430
rect -4314 -10540 -4238 -10524
rect -4314 -10574 -4298 -10540
rect -4254 -10574 -4238 -10540
rect -4314 -10580 -4238 -10574
rect -4204 -10612 -4170 -10342
rect -4136 -10380 -4060 -10374
rect -4136 -10414 -4120 -10380
rect -4076 -10414 -4060 -10380
rect -4136 -10430 -4060 -10414
rect -4120 -10524 -4076 -10430
rect -4136 -10540 -4060 -10524
rect -4136 -10574 -4120 -10540
rect -4076 -10574 -4060 -10540
rect -4136 -10580 -4060 -10574
rect -4026 -10612 -3992 -10342
rect -5634 -10624 -5588 -10612
rect -5634 -10880 -5628 -10624
rect -5594 -10880 -5588 -10624
rect -5634 -10892 -5588 -10880
rect -5456 -10624 -5410 -10612
rect -5456 -10880 -5450 -10624
rect -5416 -10880 -5410 -10624
rect -5456 -10892 -5410 -10880
rect -5278 -10624 -5232 -10612
rect -5278 -10880 -5272 -10624
rect -5238 -10880 -5232 -10624
rect -5278 -10892 -5232 -10880
rect -5100 -10624 -5054 -10612
rect -5100 -10880 -5094 -10624
rect -5060 -10880 -5054 -10624
rect -5100 -10892 -5054 -10880
rect -4922 -10624 -4876 -10612
rect -4922 -10880 -4916 -10624
rect -4882 -10880 -4876 -10624
rect -4922 -10892 -4876 -10880
rect -4744 -10624 -4698 -10612
rect -4744 -10880 -4738 -10624
rect -4704 -10880 -4698 -10624
rect -4744 -10892 -4698 -10880
rect -4566 -10624 -4520 -10612
rect -4566 -10880 -4560 -10624
rect -4526 -10880 -4520 -10624
rect -4566 -10892 -4520 -10880
rect -4388 -10624 -4342 -10612
rect -4388 -10880 -4382 -10624
rect -4348 -10880 -4342 -10624
rect -4388 -10892 -4342 -10880
rect -4210 -10624 -4164 -10612
rect -4210 -10880 -4204 -10624
rect -4170 -10880 -4164 -10624
rect -4210 -10892 -4164 -10880
rect -4032 -10624 -3986 -10612
rect -4032 -10880 -4026 -10624
rect -3992 -10880 -3986 -10624
rect -4032 -10892 -3986 -10880
rect -5628 -11162 -5594 -10892
rect -5560 -10930 -5484 -10924
rect -5560 -10964 -5544 -10930
rect -5500 -10964 -5484 -10930
rect -5560 -10980 -5484 -10964
rect -5544 -11074 -5500 -10980
rect -5560 -11090 -5484 -11074
rect -5560 -11124 -5544 -11090
rect -5500 -11124 -5484 -11090
rect -5560 -11130 -5484 -11124
rect -5450 -11162 -5416 -10892
rect -5382 -10930 -5306 -10924
rect -5382 -10964 -5366 -10930
rect -5322 -10964 -5306 -10930
rect -5382 -10980 -5306 -10964
rect -5366 -11074 -5322 -10980
rect -5382 -11090 -5306 -11074
rect -5382 -11124 -5366 -11090
rect -5322 -11124 -5306 -11090
rect -5382 -11130 -5306 -11124
rect -5272 -11162 -5238 -10892
rect -5204 -10930 -5128 -10924
rect -5204 -10964 -5188 -10930
rect -5144 -10964 -5128 -10930
rect -5204 -10980 -5128 -10964
rect -5188 -11074 -5144 -10980
rect -5204 -11090 -5128 -11074
rect -5204 -11124 -5188 -11090
rect -5144 -11124 -5128 -11090
rect -5204 -11130 -5128 -11124
rect -5094 -11162 -5060 -10892
rect -5026 -10930 -4950 -10924
rect -5026 -10964 -5010 -10930
rect -4966 -10964 -4950 -10930
rect -5026 -10980 -4950 -10964
rect -5010 -11074 -4966 -10980
rect -5026 -11090 -4950 -11074
rect -5026 -11124 -5010 -11090
rect -4966 -11124 -4950 -11090
rect -5026 -11130 -4950 -11124
rect -4916 -11162 -4882 -10892
rect -4848 -10930 -4772 -10924
rect -4848 -10964 -4832 -10930
rect -4788 -10964 -4772 -10930
rect -4848 -10980 -4772 -10964
rect -4832 -11074 -4788 -10980
rect -4848 -11090 -4772 -11074
rect -4848 -11124 -4832 -11090
rect -4788 -11124 -4772 -11090
rect -4848 -11130 -4772 -11124
rect -4738 -11162 -4704 -10892
rect -4670 -10930 -4594 -10924
rect -4670 -10964 -4654 -10930
rect -4610 -10964 -4594 -10930
rect -4670 -10980 -4594 -10964
rect -4654 -11074 -4610 -10980
rect -4670 -11090 -4594 -11074
rect -4670 -11124 -4654 -11090
rect -4610 -11124 -4594 -11090
rect -4670 -11130 -4594 -11124
rect -4560 -11162 -4526 -10892
rect -4492 -10930 -4416 -10924
rect -4492 -10964 -4476 -10930
rect -4432 -10964 -4416 -10930
rect -4492 -10980 -4416 -10964
rect -4476 -11074 -4432 -10980
rect -4492 -11090 -4416 -11074
rect -4492 -11124 -4476 -11090
rect -4432 -11124 -4416 -11090
rect -4492 -11130 -4416 -11124
rect -4382 -11162 -4348 -10892
rect -4314 -10930 -4238 -10924
rect -4314 -10964 -4298 -10930
rect -4254 -10964 -4238 -10930
rect -4314 -10980 -4238 -10964
rect -4298 -11074 -4254 -10980
rect -4314 -11090 -4238 -11074
rect -4314 -11124 -4298 -11090
rect -4254 -11124 -4238 -11090
rect -4314 -11130 -4238 -11124
rect -4204 -11162 -4170 -10892
rect -4136 -10930 -4060 -10924
rect -4136 -10964 -4120 -10930
rect -4076 -10964 -4060 -10930
rect -4136 -10980 -4060 -10964
rect -4120 -11074 -4076 -10980
rect -4136 -11090 -4060 -11074
rect -4136 -11124 -4120 -11090
rect -4076 -11124 -4060 -11090
rect -4136 -11130 -4060 -11124
rect -4026 -11162 -3992 -10892
rect -5634 -11174 -5588 -11162
rect -5634 -11430 -5628 -11174
rect -5594 -11430 -5588 -11174
rect -5634 -11442 -5588 -11430
rect -5456 -11174 -5410 -11162
rect -5456 -11430 -5450 -11174
rect -5416 -11430 -5410 -11174
rect -5456 -11442 -5410 -11430
rect -5278 -11174 -5232 -11162
rect -5278 -11430 -5272 -11174
rect -5238 -11430 -5232 -11174
rect -5278 -11442 -5232 -11430
rect -5100 -11174 -5054 -11162
rect -5100 -11430 -5094 -11174
rect -5060 -11430 -5054 -11174
rect -5100 -11442 -5054 -11430
rect -4922 -11174 -4876 -11162
rect -4922 -11430 -4916 -11174
rect -4882 -11430 -4876 -11174
rect -4922 -11442 -4876 -11430
rect -4744 -11174 -4698 -11162
rect -4744 -11430 -4738 -11174
rect -4704 -11430 -4698 -11174
rect -4744 -11442 -4698 -11430
rect -4566 -11174 -4520 -11162
rect -4566 -11430 -4560 -11174
rect -4526 -11430 -4520 -11174
rect -4566 -11442 -4520 -11430
rect -4388 -11174 -4342 -11162
rect -4388 -11430 -4382 -11174
rect -4348 -11430 -4342 -11174
rect -4388 -11442 -4342 -11430
rect -4210 -11174 -4164 -11162
rect -4210 -11430 -4204 -11174
rect -4170 -11430 -4164 -11174
rect -4210 -11442 -4164 -11430
rect -4032 -11174 -3986 -11162
rect -4032 -11430 -4026 -11174
rect -3992 -11430 -3986 -11174
rect -4032 -11442 -3986 -11430
rect -5628 -11712 -5594 -11442
rect -5560 -11480 -5484 -11474
rect -5560 -11514 -5544 -11480
rect -5500 -11514 -5484 -11480
rect -5560 -11530 -5484 -11514
rect -5544 -11624 -5500 -11530
rect -5560 -11640 -5484 -11624
rect -5560 -11674 -5544 -11640
rect -5500 -11674 -5484 -11640
rect -5560 -11680 -5484 -11674
rect -5450 -11712 -5416 -11442
rect -5382 -11480 -5306 -11474
rect -5382 -11514 -5366 -11480
rect -5322 -11514 -5306 -11480
rect -5382 -11530 -5306 -11514
rect -5364 -11624 -5320 -11530
rect -5382 -11640 -5306 -11624
rect -5382 -11674 -5366 -11640
rect -5322 -11674 -5306 -11640
rect -5382 -11680 -5306 -11674
rect -5272 -11712 -5238 -11442
rect -5204 -11480 -5128 -11474
rect -5204 -11514 -5188 -11480
rect -5144 -11514 -5128 -11480
rect -5204 -11530 -5128 -11514
rect -5188 -11624 -5144 -11530
rect -5204 -11640 -5128 -11624
rect -5204 -11674 -5188 -11640
rect -5144 -11674 -5128 -11640
rect -5204 -11680 -5128 -11674
rect -5094 -11712 -5060 -11442
rect -5026 -11480 -4950 -11474
rect -5026 -11514 -5010 -11480
rect -4966 -11514 -4950 -11480
rect -5026 -11530 -4950 -11514
rect -5010 -11624 -4966 -11530
rect -5026 -11640 -4950 -11624
rect -5026 -11674 -5010 -11640
rect -4966 -11674 -4950 -11640
rect -5026 -11680 -4950 -11674
rect -4916 -11712 -4882 -11442
rect -4848 -11480 -4772 -11474
rect -4848 -11514 -4832 -11480
rect -4788 -11514 -4772 -11480
rect -4848 -11530 -4772 -11514
rect -4832 -11624 -4788 -11530
rect -4848 -11640 -4772 -11624
rect -4848 -11674 -4832 -11640
rect -4788 -11674 -4772 -11640
rect -4848 -11680 -4772 -11674
rect -4738 -11712 -4704 -11442
rect -4670 -11480 -4594 -11474
rect -4670 -11514 -4654 -11480
rect -4610 -11514 -4594 -11480
rect -4670 -11530 -4594 -11514
rect -4654 -11624 -4610 -11530
rect -4670 -11640 -4594 -11624
rect -4670 -11674 -4654 -11640
rect -4610 -11674 -4594 -11640
rect -4670 -11680 -4594 -11674
rect -4560 -11712 -4526 -11442
rect -4492 -11480 -4416 -11474
rect -4492 -11514 -4476 -11480
rect -4432 -11514 -4416 -11480
rect -4492 -11530 -4416 -11514
rect -4476 -11624 -4432 -11530
rect -4492 -11640 -4416 -11624
rect -4492 -11674 -4476 -11640
rect -4432 -11674 -4416 -11640
rect -4492 -11680 -4416 -11674
rect -4382 -11712 -4348 -11442
rect -4314 -11480 -4238 -11474
rect -4314 -11514 -4298 -11480
rect -4254 -11514 -4238 -11480
rect -4314 -11530 -4238 -11514
rect -4298 -11624 -4254 -11530
rect -4314 -11640 -4238 -11624
rect -4314 -11674 -4298 -11640
rect -4254 -11674 -4238 -11640
rect -4314 -11680 -4238 -11674
rect -4204 -11712 -4170 -11442
rect -4136 -11480 -4060 -11474
rect -4136 -11514 -4120 -11480
rect -4076 -11514 -4060 -11480
rect -4136 -11530 -4060 -11514
rect -4120 -11624 -4076 -11530
rect -4136 -11640 -4060 -11624
rect -4136 -11674 -4120 -11640
rect -4076 -11674 -4060 -11640
rect -4136 -11680 -4060 -11674
rect -4026 -11712 -3992 -11442
rect -5634 -11724 -5588 -11712
rect -5634 -11980 -5628 -11724
rect -5594 -11980 -5588 -11724
rect -5634 -11992 -5588 -11980
rect -5456 -11724 -5410 -11712
rect -5456 -11980 -5450 -11724
rect -5416 -11980 -5410 -11724
rect -5456 -11992 -5410 -11980
rect -5278 -11724 -5232 -11712
rect -5278 -11980 -5272 -11724
rect -5238 -11980 -5232 -11724
rect -5278 -11992 -5232 -11980
rect -5100 -11724 -5054 -11712
rect -5100 -11980 -5094 -11724
rect -5060 -11980 -5054 -11724
rect -5100 -11992 -5054 -11980
rect -4922 -11724 -4876 -11712
rect -4922 -11980 -4916 -11724
rect -4882 -11980 -4876 -11724
rect -4922 -11992 -4876 -11980
rect -4744 -11724 -4698 -11712
rect -4744 -11980 -4738 -11724
rect -4704 -11980 -4698 -11724
rect -4744 -11992 -4698 -11980
rect -4566 -11724 -4520 -11712
rect -4566 -11980 -4560 -11724
rect -4526 -11980 -4520 -11724
rect -4566 -11992 -4520 -11980
rect -4388 -11724 -4342 -11712
rect -4388 -11980 -4382 -11724
rect -4348 -11980 -4342 -11724
rect -4388 -11992 -4342 -11980
rect -4210 -11724 -4164 -11712
rect -4210 -11980 -4204 -11724
rect -4170 -11980 -4164 -11724
rect -4210 -11992 -4164 -11980
rect -4032 -11724 -3986 -11712
rect -4032 -11980 -4026 -11724
rect -3992 -11980 -3986 -11724
rect -4032 -11992 -3986 -11980
rect -5560 -12030 -5484 -12024
rect -5560 -12064 -5544 -12030
rect -5500 -12064 -5484 -12030
rect -5560 -12080 -5484 -12064
rect -5382 -12030 -5306 -12024
rect -5382 -12064 -5366 -12030
rect -5322 -12064 -5306 -12030
rect -5382 -12080 -5306 -12064
rect -5272 -12119 -5238 -11992
rect -5204 -12030 -5128 -12024
rect -5204 -12064 -5188 -12030
rect -5144 -12064 -5128 -12030
rect -5204 -12080 -5128 -12064
rect -5026 -12030 -4950 -12024
rect -5026 -12064 -5010 -12030
rect -4966 -12064 -4950 -12030
rect -5026 -12080 -4950 -12064
rect -4916 -12119 -4882 -11992
rect -4848 -12030 -4772 -12024
rect -4848 -12064 -4832 -12030
rect -4788 -12064 -4772 -12030
rect -4848 -12080 -4772 -12064
rect -4670 -12030 -4594 -12024
rect -4670 -12064 -4654 -12030
rect -4610 -12064 -4594 -12030
rect -4670 -12080 -4594 -12064
rect -4560 -12119 -4526 -11992
rect -4492 -12030 -4416 -12024
rect -4492 -12064 -4476 -12030
rect -4432 -12064 -4416 -12030
rect -4492 -12080 -4416 -12064
rect -4314 -12030 -4238 -12024
rect -4314 -12064 -4298 -12030
rect -4254 -12064 -4238 -12030
rect -4314 -12080 -4238 -12064
rect -4204 -12119 -4170 -11992
rect -4136 -12030 -4060 -12024
rect -4136 -12064 -4120 -12030
rect -4076 -12064 -4060 -12030
rect -4136 -12080 -4060 -12064
rect -4113 -12119 -4079 -12080
rect -4026 -12119 -3992 -11992
rect -5272 -12153 -3611 -12119
rect -5512 -12324 -5502 -12271
rect -5449 -12324 -5439 -12271
rect -6976 -12565 -6077 -12512
rect -6024 -12565 -6014 -12512
rect -5636 -12565 -5626 -12512
rect -5573 -12565 -5563 -12512
rect -6233 -13115 -6223 -13062
rect -6170 -13115 -6160 -13062
rect -6976 -13905 -6426 -13852
rect -6373 -13905 -6363 -13852
rect -6223 -14055 -6170 -13115
rect -6077 -13745 -6024 -12565
rect -5617 -12612 -5583 -12565
rect -5922 -12628 -5778 -12612
rect -5922 -12662 -5867 -12628
rect -5833 -12662 -5778 -12628
rect -5922 -12668 -5778 -12662
rect -5633 -12628 -5567 -12612
rect -5633 -12662 -5617 -12628
rect -5583 -12662 -5567 -12628
rect -5633 -12668 -5567 -12662
rect -5922 -12700 -5876 -12668
rect -5824 -12700 -5778 -12668
rect -5492 -12700 -5458 -12324
rect -5010 -12325 -5000 -12272
rect -4947 -12325 -4937 -12272
rect -4512 -12324 -4502 -12271
rect -4449 -12324 -4439 -12271
rect -5386 -12441 -5376 -12388
rect -5323 -12441 -5313 -12388
rect -5137 -12441 -5127 -12388
rect -5074 -12441 -5064 -12388
rect -5367 -12612 -5333 -12441
rect -5117 -12612 -5083 -12441
rect -5383 -12628 -5317 -12612
rect -5383 -12662 -5367 -12628
rect -5333 -12662 -5317 -12628
rect -5383 -12668 -5317 -12662
rect -5133 -12628 -5067 -12612
rect -5133 -12662 -5117 -12628
rect -5083 -12662 -5067 -12628
rect -5133 -12668 -5067 -12662
rect -4992 -12700 -4958 -12325
rect -4887 -12565 -4877 -12512
rect -4824 -12565 -4814 -12512
rect -4637 -12565 -4627 -12512
rect -4574 -12565 -4564 -12512
rect -4867 -12612 -4833 -12565
rect -4617 -12612 -4583 -12565
rect -4883 -12628 -4817 -12612
rect -4883 -12662 -4867 -12628
rect -4833 -12662 -4817 -12628
rect -4883 -12668 -4817 -12662
rect -4633 -12628 -4567 -12612
rect -4633 -12662 -4617 -12628
rect -4583 -12662 -4567 -12628
rect -4633 -12668 -4567 -12662
rect -4492 -12700 -4458 -12324
rect -4387 -12441 -4377 -12388
rect -4324 -12441 -4314 -12388
rect -4367 -12612 -4333 -12441
rect -3938 -12442 -3928 -12389
rect -3875 -12442 -3865 -12389
rect -4383 -12628 -4317 -12612
rect -4383 -12662 -4367 -12628
rect -4333 -12662 -4317 -12628
rect -4383 -12668 -4317 -12662
rect -4172 -12628 -4028 -12612
rect -4172 -12662 -4117 -12628
rect -4083 -12662 -4028 -12628
rect -4172 -12668 -4028 -12662
rect -4172 -12700 -4126 -12668
rect -5923 -12712 -5877 -12700
rect -5923 -12928 -5917 -12712
rect -5883 -12928 -5877 -12712
rect -5824 -12712 -5626 -12700
rect -5824 -12740 -5817 -12712
rect -5923 -12940 -5877 -12928
rect -5823 -12928 -5817 -12740
rect -5783 -12740 -5667 -12712
rect -5783 -12900 -5777 -12740
rect -5673 -12900 -5667 -12740
rect -5783 -12928 -5667 -12900
rect -5633 -12740 -5626 -12712
rect -5574 -12712 -5376 -12700
rect -5574 -12740 -5567 -12712
rect -5633 -12928 -5627 -12740
rect -5573 -12900 -5567 -12740
rect -5823 -12940 -5627 -12928
rect -5574 -12928 -5567 -12900
rect -5533 -12740 -5417 -12712
rect -5533 -12900 -5527 -12740
rect -5423 -12900 -5417 -12740
rect -5533 -12928 -5417 -12900
rect -5383 -12740 -5376 -12712
rect -5324 -12712 -5126 -12700
rect -5324 -12740 -5317 -12712
rect -5383 -12900 -5377 -12740
rect -5323 -12900 -5317 -12740
rect -5383 -12928 -5376 -12900
rect -5574 -12940 -5376 -12928
rect -5324 -12928 -5317 -12900
rect -5283 -12740 -5167 -12712
rect -5283 -12900 -5277 -12740
rect -5173 -12900 -5167 -12740
rect -5283 -12928 -5167 -12900
rect -5133 -12740 -5126 -12712
rect -5074 -12712 -4876 -12700
rect -5074 -12740 -5067 -12712
rect -5133 -12900 -5127 -12740
rect -5073 -12900 -5067 -12740
rect -5133 -12928 -5126 -12900
rect -5324 -12940 -5126 -12928
rect -5074 -12928 -5067 -12900
rect -5033 -12740 -4917 -12712
rect -5033 -12900 -5027 -12740
rect -4923 -12900 -4917 -12740
rect -5033 -12928 -4917 -12900
rect -4883 -12740 -4876 -12712
rect -4823 -12712 -4625 -12700
rect -4883 -12900 -4877 -12740
rect -4823 -12900 -4817 -12712
rect -4883 -12928 -4876 -12900
rect -5074 -12940 -4876 -12928
rect -4825 -12928 -4817 -12900
rect -4783 -12740 -4667 -12712
rect -4783 -12900 -4777 -12740
rect -4673 -12900 -4667 -12740
rect -4783 -12928 -4667 -12900
rect -4633 -12740 -4625 -12712
rect -4574 -12712 -4376 -12700
rect -4574 -12740 -4567 -12712
rect -4633 -12928 -4627 -12740
rect -4573 -12900 -4567 -12740
rect -4825 -12940 -4627 -12928
rect -4574 -12928 -4567 -12900
rect -4533 -12740 -4417 -12712
rect -4533 -12900 -4527 -12740
rect -4423 -12900 -4417 -12740
rect -4533 -12928 -4417 -12900
rect -4383 -12740 -4376 -12712
rect -4324 -12712 -4126 -12700
rect -4074 -12700 -4028 -12668
rect -4074 -12712 -4027 -12700
rect -4324 -12740 -4317 -12712
rect -4383 -12900 -4377 -12740
rect -4323 -12900 -4317 -12740
rect -4383 -12928 -4376 -12900
rect -4574 -12940 -4376 -12928
rect -4324 -12928 -4317 -12900
rect -4283 -12740 -4167 -12712
rect -4283 -12900 -4277 -12740
rect -4173 -12900 -4167 -12740
rect -4283 -12928 -4167 -12900
rect -4133 -12740 -4126 -12712
rect -4133 -12900 -4127 -12740
rect -4133 -12928 -4126 -12900
rect -4324 -12940 -4126 -12928
rect -4073 -12928 -4067 -12712
rect -4033 -12928 -4027 -12712
rect -4073 -12940 -4027 -12928
rect -5883 -12978 -5817 -12972
rect -5883 -13012 -5867 -12978
rect -5833 -13012 -5817 -12978
rect -5883 -13028 -5817 -13012
rect -5744 -13062 -5704 -12940
rect -5633 -12978 -5567 -12972
rect -5633 -13012 -5617 -12978
rect -5583 -13012 -5567 -12978
rect -5633 -13028 -5567 -13012
rect -5761 -13115 -5751 -13062
rect -5698 -13115 -5688 -13062
rect -5883 -13308 -5817 -13292
rect -5883 -13342 -5867 -13308
rect -5833 -13342 -5817 -13308
rect -5883 -13348 -5817 -13342
rect -5633 -13308 -5567 -13292
rect -5633 -13342 -5617 -13308
rect -5583 -13342 -5567 -13308
rect -5633 -13348 -5567 -13342
rect -5495 -13380 -5455 -12940
rect -5383 -12978 -5317 -12972
rect -5383 -13012 -5367 -12978
rect -5333 -13012 -5317 -12978
rect -5383 -13028 -5317 -13012
rect -5245 -13189 -5205 -12940
rect -5133 -12978 -5067 -12972
rect -5133 -13012 -5117 -12978
rect -5083 -13012 -5067 -12978
rect -5133 -13028 -5067 -13012
rect -5261 -13242 -5251 -13189
rect -5198 -13242 -5188 -13189
rect -5383 -13308 -5317 -13292
rect -5383 -13342 -5367 -13308
rect -5333 -13342 -5317 -13308
rect -5383 -13348 -5317 -13342
rect -5133 -13308 -5067 -13292
rect -5133 -13342 -5117 -13308
rect -5083 -13342 -5067 -13308
rect -5133 -13348 -5067 -13342
rect -4995 -13380 -4955 -12940
rect -4883 -12978 -4817 -12972
rect -4883 -13012 -4867 -12978
rect -4833 -13012 -4817 -12978
rect -4883 -13028 -4817 -13012
rect -4746 -13062 -4706 -12940
rect -4633 -12978 -4567 -12972
rect -4633 -13012 -4617 -12978
rect -4583 -13012 -4567 -12978
rect -4633 -13028 -4567 -13012
rect -4762 -13115 -4752 -13062
rect -4699 -13115 -4689 -13062
rect -4883 -13308 -4817 -13292
rect -4883 -13342 -4867 -13308
rect -4833 -13342 -4817 -13308
rect -4883 -13348 -4817 -13342
rect -4633 -13308 -4567 -13292
rect -4633 -13342 -4617 -13308
rect -4583 -13342 -4567 -13308
rect -4633 -13348 -4567 -13342
rect -4495 -13380 -4455 -12940
rect -4383 -12978 -4317 -12972
rect -4383 -13012 -4367 -12978
rect -4333 -13012 -4317 -12978
rect -4383 -13028 -4317 -13012
rect -4244 -13189 -4204 -12940
rect -4133 -12978 -4067 -12972
rect -4133 -13012 -4117 -12978
rect -4083 -13012 -4067 -12978
rect -4133 -13028 -4067 -13012
rect -4261 -13242 -4251 -13189
rect -4198 -13242 -4188 -13189
rect -4383 -13308 -4317 -13292
rect -4383 -13342 -4367 -13308
rect -4333 -13342 -4317 -13308
rect -4383 -13348 -4317 -13342
rect -4133 -13308 -4067 -13292
rect -4133 -13342 -4117 -13308
rect -4083 -13342 -4067 -13308
rect -4133 -13348 -4067 -13342
rect -5923 -13392 -5877 -13380
rect -5923 -13608 -5917 -13392
rect -5883 -13608 -5877 -13392
rect -5824 -13392 -5626 -13380
rect -5824 -13420 -5817 -13392
rect -5823 -13580 -5817 -13420
rect -5824 -13608 -5817 -13580
rect -5783 -13420 -5667 -13392
rect -5783 -13580 -5777 -13420
rect -5673 -13580 -5667 -13420
rect -5783 -13608 -5667 -13580
rect -5633 -13420 -5626 -13392
rect -5574 -13392 -5376 -13380
rect -5574 -13420 -5567 -13392
rect -5633 -13580 -5627 -13420
rect -5573 -13580 -5567 -13420
rect -5633 -13608 -5626 -13580
rect -5923 -13620 -5876 -13608
rect -5922 -13652 -5876 -13620
rect -5824 -13620 -5626 -13608
rect -5574 -13608 -5567 -13580
rect -5533 -13420 -5417 -13392
rect -5533 -13580 -5527 -13420
rect -5423 -13580 -5417 -13420
rect -5533 -13608 -5417 -13580
rect -5383 -13420 -5376 -13392
rect -5324 -13392 -5126 -13380
rect -5324 -13420 -5317 -13392
rect -5383 -13580 -5377 -13420
rect -5323 -13580 -5317 -13420
rect -5383 -13608 -5376 -13580
rect -5574 -13620 -5376 -13608
rect -5324 -13608 -5317 -13580
rect -5283 -13420 -5167 -13392
rect -5283 -13580 -5277 -13420
rect -5173 -13580 -5167 -13420
rect -5283 -13608 -5167 -13580
rect -5133 -13420 -5126 -13392
rect -5074 -13392 -4876 -13380
rect -5074 -13420 -5067 -13392
rect -5133 -13580 -5127 -13420
rect -5073 -13580 -5067 -13420
rect -5133 -13608 -5126 -13580
rect -5324 -13620 -5126 -13608
rect -5074 -13608 -5067 -13580
rect -5033 -13420 -4917 -13392
rect -5033 -13580 -5027 -13420
rect -4923 -13580 -4917 -13420
rect -5033 -13608 -4917 -13580
rect -4883 -13420 -4876 -13392
rect -4824 -13392 -4626 -13380
rect -4824 -13420 -4817 -13392
rect -4883 -13580 -4877 -13420
rect -4823 -13580 -4817 -13420
rect -4883 -13608 -4876 -13580
rect -5074 -13620 -4876 -13608
rect -4824 -13608 -4817 -13580
rect -4783 -13420 -4667 -13392
rect -4783 -13580 -4777 -13420
rect -4673 -13580 -4667 -13420
rect -4783 -13608 -4667 -13580
rect -4633 -13420 -4626 -13392
rect -4574 -13392 -4376 -13380
rect -4574 -13420 -4567 -13392
rect -4633 -13580 -4627 -13420
rect -4573 -13580 -4567 -13420
rect -4633 -13608 -4626 -13580
rect -4824 -13620 -4626 -13608
rect -4574 -13608 -4567 -13580
rect -4533 -13420 -4417 -13392
rect -4533 -13580 -4527 -13420
rect -4423 -13580 -4417 -13420
rect -4533 -13608 -4417 -13580
rect -4383 -13420 -4376 -13392
rect -4324 -13392 -4126 -13380
rect -4324 -13420 -4317 -13392
rect -4383 -13580 -4377 -13420
rect -4323 -13580 -4317 -13420
rect -4383 -13608 -4376 -13580
rect -4574 -13620 -4376 -13608
rect -4324 -13608 -4317 -13580
rect -4283 -13420 -4167 -13392
rect -4283 -13580 -4277 -13420
rect -4173 -13580 -4167 -13420
rect -4283 -13608 -4167 -13580
rect -4133 -13420 -4126 -13392
rect -4073 -13392 -4027 -13380
rect -4133 -13580 -4127 -13420
rect -4133 -13608 -4126 -13580
rect -4073 -13608 -4067 -13392
rect -4033 -13608 -4027 -13392
rect -4324 -13620 -4126 -13608
rect -5824 -13652 -5778 -13620
rect -5922 -13658 -5778 -13652
rect -5922 -13692 -5867 -13658
rect -5833 -13692 -5778 -13658
rect -5922 -13708 -5778 -13692
rect -6087 -13798 -6077 -13745
rect -6024 -13798 -6014 -13745
rect -5720 -13957 -5686 -13620
rect -5633 -13658 -5567 -13652
rect -5633 -13692 -5617 -13658
rect -5583 -13692 -5567 -13658
rect -5633 -13708 -5567 -13692
rect -5383 -13658 -5317 -13652
rect -5383 -13692 -5367 -13658
rect -5333 -13692 -5317 -13658
rect -5383 -13708 -5317 -13692
rect -5617 -13852 -5583 -13708
rect -5367 -13745 -5333 -13708
rect -5386 -13798 -5376 -13745
rect -5323 -13798 -5313 -13745
rect -5636 -13905 -5626 -13852
rect -5573 -13905 -5563 -13852
rect -5740 -14010 -5730 -13957
rect -5677 -14010 -5667 -13957
rect -5240 -14055 -5206 -13620
rect -5133 -13658 -5067 -13652
rect -5133 -13692 -5117 -13658
rect -5083 -13692 -5067 -13658
rect -5133 -13708 -5067 -13692
rect -4883 -13658 -4817 -13652
rect -4883 -13692 -4867 -13658
rect -4833 -13692 -4817 -13658
rect -4883 -13708 -4817 -13692
rect -5117 -13745 -5083 -13708
rect -5136 -13798 -5126 -13745
rect -5073 -13798 -5063 -13745
rect -4867 -13852 -4833 -13708
rect -4887 -13905 -4877 -13852
rect -4824 -13905 -4814 -13852
rect -4742 -13957 -4708 -13620
rect -4633 -13658 -4567 -13652
rect -4633 -13692 -4617 -13658
rect -4583 -13692 -4567 -13658
rect -4633 -13708 -4567 -13692
rect -4383 -13658 -4317 -13652
rect -4383 -13692 -4367 -13658
rect -4333 -13692 -4317 -13658
rect -4383 -13708 -4317 -13692
rect -4617 -13852 -4583 -13708
rect -4367 -13745 -4333 -13708
rect -4386 -13798 -4376 -13745
rect -4323 -13798 -4313 -13745
rect -4637 -13905 -4627 -13852
rect -4574 -13905 -4564 -13852
rect -4762 -14010 -4752 -13957
rect -4699 -14010 -4689 -13957
rect -4240 -14055 -4206 -13620
rect -4172 -13652 -4126 -13620
rect -4074 -13620 -4027 -13608
rect -4074 -13652 -4028 -13620
rect -4172 -13658 -4028 -13652
rect -4172 -13692 -4117 -13658
rect -4083 -13692 -4028 -13658
rect -4172 -13708 -4028 -13692
rect -3928 -13852 -3875 -12442
rect -3798 -13242 -3788 -13189
rect -3735 -13242 -3725 -13189
rect -3938 -13905 -3928 -13852
rect -3875 -13905 -3865 -13852
rect -3928 -13906 -3875 -13905
rect -3788 -13957 -3735 -13242
rect -3798 -14010 -3788 -13957
rect -3735 -14010 -3725 -13957
rect -6233 -14108 -6223 -14055
rect -6170 -14108 -6160 -14055
rect -5260 -14108 -5250 -14055
rect -5197 -14108 -5187 -14055
rect -4260 -14108 -4250 -14055
rect -4197 -14108 -4187 -14055
rect -6965 -14260 -4303 -14226
rect -6028 -14382 -5994 -14260
rect -5939 -14294 -5905 -14260
rect -5960 -14310 -5884 -14294
rect -5960 -14344 -5944 -14310
rect -5900 -14344 -5884 -14310
rect -5960 -14350 -5884 -14344
rect -5850 -14382 -5816 -14260
rect -5761 -14294 -5727 -14260
rect -5583 -14294 -5549 -14260
rect -5405 -14294 -5371 -14260
rect -5227 -14294 -5193 -14260
rect -5049 -14294 -5015 -14260
rect -4871 -14294 -4837 -14260
rect -4693 -14294 -4659 -14260
rect -4515 -14294 -4481 -14260
rect -4337 -14294 -4303 -14260
rect -4248 -14260 -4036 -14226
rect -5782 -14310 -5706 -14294
rect -5782 -14344 -5766 -14310
rect -5722 -14344 -5706 -14310
rect -5782 -14350 -5706 -14344
rect -5604 -14310 -5528 -14294
rect -5604 -14344 -5588 -14310
rect -5544 -14344 -5528 -14310
rect -5604 -14350 -5528 -14344
rect -5426 -14310 -5350 -14294
rect -5426 -14344 -5410 -14310
rect -5366 -14344 -5350 -14310
rect -5426 -14350 -5350 -14344
rect -5248 -14310 -5172 -14294
rect -5248 -14344 -5232 -14310
rect -5188 -14344 -5172 -14310
rect -5248 -14350 -5172 -14344
rect -5070 -14310 -4994 -14294
rect -5070 -14344 -5054 -14310
rect -5010 -14344 -4994 -14310
rect -5070 -14350 -4994 -14344
rect -4892 -14310 -4816 -14294
rect -4892 -14344 -4876 -14310
rect -4832 -14344 -4816 -14310
rect -4892 -14350 -4816 -14344
rect -4714 -14310 -4638 -14294
rect -4714 -14344 -4698 -14310
rect -4654 -14344 -4638 -14310
rect -4714 -14350 -4638 -14344
rect -4536 -14310 -4460 -14294
rect -4536 -14344 -4520 -14310
rect -4476 -14344 -4460 -14310
rect -4536 -14350 -4460 -14344
rect -4358 -14310 -4282 -14294
rect -4358 -14344 -4342 -14310
rect -4298 -14344 -4282 -14310
rect -4358 -14350 -4282 -14344
rect -4248 -14382 -4214 -14260
rect -4159 -14294 -4125 -14260
rect -4180 -14310 -4104 -14294
rect -4180 -14344 -4164 -14310
rect -4120 -14344 -4104 -14310
rect -4180 -14350 -4104 -14344
rect -4070 -14382 -4036 -14260
rect -6034 -14394 -5988 -14382
rect -6034 -14650 -6028 -14394
rect -5994 -14650 -5988 -14394
rect -6034 -14662 -5988 -14650
rect -5856 -14394 -5810 -14382
rect -5856 -14650 -5850 -14394
rect -5816 -14650 -5810 -14394
rect -5856 -14662 -5810 -14650
rect -5678 -14394 -5632 -14382
rect -5678 -14650 -5672 -14394
rect -5638 -14650 -5632 -14394
rect -5678 -14662 -5632 -14650
rect -5500 -14394 -5454 -14382
rect -5500 -14650 -5494 -14394
rect -5460 -14650 -5454 -14394
rect -5500 -14662 -5454 -14650
rect -5322 -14394 -5276 -14382
rect -5322 -14650 -5316 -14394
rect -5282 -14650 -5276 -14394
rect -5322 -14662 -5276 -14650
rect -5144 -14394 -5098 -14382
rect -5144 -14650 -5138 -14394
rect -5104 -14650 -5098 -14394
rect -5144 -14662 -5098 -14650
rect -4966 -14394 -4920 -14382
rect -4966 -14650 -4960 -14394
rect -4926 -14650 -4920 -14394
rect -4966 -14662 -4920 -14650
rect -4788 -14394 -4742 -14382
rect -4788 -14650 -4782 -14394
rect -4748 -14650 -4742 -14394
rect -4788 -14662 -4742 -14650
rect -4610 -14394 -4564 -14382
rect -4610 -14650 -4604 -14394
rect -4570 -14650 -4564 -14394
rect -4610 -14662 -4564 -14650
rect -4432 -14394 -4386 -14382
rect -4432 -14650 -4426 -14394
rect -4392 -14650 -4386 -14394
rect -4432 -14662 -4386 -14650
rect -4254 -14394 -4208 -14382
rect -4254 -14650 -4248 -14394
rect -4214 -14650 -4208 -14394
rect -4254 -14662 -4208 -14650
rect -4076 -14394 -4030 -14382
rect -4076 -14650 -4070 -14394
rect -4036 -14650 -4030 -14394
rect -4076 -14662 -4030 -14650
rect -5960 -14700 -5884 -14694
rect -5960 -14734 -5944 -14700
rect -5900 -14734 -5884 -14700
rect -5960 -14750 -5884 -14734
rect -5850 -14795 -5816 -14662
rect -5782 -14700 -5706 -14694
rect -5782 -14734 -5766 -14700
rect -5722 -14734 -5706 -14700
rect -5782 -14750 -5706 -14734
rect -6169 -14848 -6159 -14795
rect -6106 -14848 -6096 -14795
rect -5870 -14848 -5860 -14795
rect -5807 -14848 -5797 -14795
rect -6159 -15482 -6106 -14848
rect -6028 -14959 -5816 -14925
rect -6027 -15082 -5993 -14959
rect -5939 -14994 -5905 -14959
rect -5960 -15010 -5884 -14994
rect -5960 -15044 -5944 -15010
rect -5900 -15044 -5884 -15010
rect -5960 -15050 -5884 -15044
rect -5850 -15082 -5816 -14959
rect -5761 -14994 -5727 -14750
rect -5782 -15010 -5706 -14994
rect -5782 -15044 -5766 -15010
rect -5722 -15044 -5706 -15010
rect -5782 -15050 -5706 -15044
rect -5672 -15082 -5638 -14662
rect -5604 -14700 -5528 -14694
rect -5604 -14734 -5588 -14700
rect -5544 -14734 -5528 -14700
rect -5604 -14750 -5528 -14734
rect -5583 -14994 -5549 -14750
rect -5494 -14901 -5460 -14662
rect -5426 -14700 -5350 -14694
rect -5426 -14734 -5410 -14700
rect -5366 -14734 -5350 -14700
rect -5426 -14750 -5350 -14734
rect -5514 -14954 -5504 -14901
rect -5451 -14954 -5441 -14901
rect -5405 -14994 -5371 -14750
rect -5604 -15010 -5528 -14994
rect -5604 -15044 -5588 -15010
rect -5544 -15044 -5528 -15010
rect -5604 -15050 -5528 -15044
rect -5426 -15010 -5350 -14994
rect -5426 -15044 -5410 -15010
rect -5366 -15044 -5350 -15010
rect -5426 -15050 -5350 -15044
rect -5316 -15082 -5282 -14662
rect -5248 -14700 -5172 -14694
rect -5248 -14734 -5232 -14700
rect -5188 -14734 -5172 -14700
rect -5248 -14750 -5172 -14734
rect -5227 -14994 -5193 -14750
rect -5138 -14795 -5104 -14662
rect -5070 -14700 -4994 -14694
rect -5070 -14734 -5054 -14700
rect -5010 -14734 -4994 -14700
rect -5070 -14750 -4994 -14734
rect -5157 -14848 -5147 -14795
rect -5094 -14848 -5084 -14795
rect -5049 -14994 -5015 -14750
rect -5248 -15010 -5172 -14994
rect -5248 -15044 -5232 -15010
rect -5188 -15044 -5172 -15010
rect -5248 -15050 -5172 -15044
rect -5070 -15010 -4994 -14994
rect -5070 -15044 -5054 -15010
rect -5010 -15044 -4994 -15010
rect -5070 -15050 -4994 -15044
rect -4960 -15082 -4926 -14662
rect -4892 -14700 -4816 -14694
rect -4892 -14734 -4876 -14700
rect -4832 -14734 -4816 -14700
rect -4892 -14750 -4816 -14734
rect -4871 -14994 -4837 -14750
rect -4782 -14901 -4748 -14662
rect -4714 -14700 -4638 -14694
rect -4714 -14734 -4698 -14700
rect -4654 -14734 -4638 -14700
rect -4714 -14750 -4638 -14734
rect -4801 -14954 -4791 -14901
rect -4738 -14954 -4728 -14901
rect -4693 -14994 -4659 -14750
rect -4892 -15010 -4816 -14994
rect -4892 -15044 -4876 -15010
rect -4832 -15044 -4816 -15010
rect -4892 -15050 -4816 -15044
rect -4714 -15010 -4638 -14994
rect -4714 -15044 -4698 -15010
rect -4654 -15044 -4638 -15010
rect -4714 -15050 -4638 -15044
rect -4604 -15082 -4570 -14662
rect -4536 -14700 -4460 -14694
rect -4536 -14734 -4520 -14700
rect -4476 -14734 -4460 -14700
rect -4536 -14750 -4460 -14734
rect -4515 -14994 -4481 -14750
rect -4426 -14795 -4392 -14662
rect -4358 -14700 -4282 -14694
rect -4358 -14734 -4342 -14700
rect -4298 -14734 -4282 -14700
rect -4358 -14750 -4282 -14734
rect -4446 -14848 -4436 -14795
rect -4383 -14848 -4373 -14795
rect -4337 -14994 -4303 -14750
rect -4248 -14925 -4214 -14662
rect -4180 -14700 -4104 -14694
rect -4180 -14734 -4164 -14700
rect -4120 -14734 -4104 -14700
rect -4180 -14750 -4104 -14734
rect -3664 -14901 -3611 -12153
rect -3541 -13137 -3489 -7840
rect 4761 -7907 4771 -7854
rect 4824 -7907 4834 -7854
rect 4896 -7905 4906 -7852
rect 4959 -7905 4969 -7852
rect 5027 -7903 5037 -7850
rect 5090 -7903 5100 -7850
rect -3392 -7986 -3382 -7933
rect -3329 -7986 -3319 -7933
rect -1392 -7975 -1382 -7922
rect -1329 -7975 -1319 -7922
rect -3542 -13189 -3489 -13137
rect -3552 -13242 -3542 -13189
rect -3489 -13242 -3479 -13189
rect -3382 -14055 -3329 -7986
rect -1372 -8032 -1338 -7975
rect -1213 -7976 -1203 -7923
rect -1150 -7976 -1140 -7923
rect -1035 -7975 -1025 -7922
rect -972 -7975 -962 -7922
rect -858 -7975 -848 -7922
rect -795 -7975 -785 -7922
rect -680 -7975 -670 -7922
rect -617 -7975 -607 -7922
rect -500 -7975 -490 -7922
rect -437 -7975 -427 -7922
rect 745 -7975 755 -7922
rect 808 -7975 818 -7922
rect 922 -7975 932 -7922
rect 985 -7975 995 -7922
rect 1102 -7975 1112 -7922
rect 1165 -7975 1175 -7922
rect -1194 -8032 -1160 -7976
rect -1016 -8032 -982 -7975
rect -838 -8032 -804 -7975
rect -660 -8032 -626 -7975
rect -481 -8032 -447 -7975
rect 765 -8032 799 -7975
rect 942 -8032 976 -7975
rect 1121 -8032 1155 -7975
rect 1279 -7976 1289 -7923
rect 1342 -7976 1352 -7923
rect 1457 -7975 1467 -7922
rect 1520 -7975 1530 -7922
rect 1634 -7975 1644 -7922
rect 1697 -7975 1707 -7922
rect 2880 -7975 2890 -7922
rect 2943 -7975 2953 -7922
rect 3059 -7975 3069 -7922
rect 3122 -7975 3132 -7922
rect 3237 -7975 3247 -7922
rect 3300 -7975 3310 -7922
rect 3414 -7975 3424 -7922
rect 3477 -7975 3487 -7922
rect 1298 -8032 1332 -7976
rect 1476 -8032 1510 -7975
rect 1654 -8032 1688 -7975
rect 2900 -8032 2934 -7975
rect 3078 -8032 3112 -7975
rect 3256 -8032 3290 -7975
rect 3434 -8032 3468 -7975
rect 3593 -7976 3603 -7923
rect 3656 -7976 3666 -7923
rect 3768 -7975 3778 -7922
rect 3831 -7975 3841 -7922
rect 3612 -8032 3646 -7976
rect 3790 -8032 3824 -7975
rect 4198 -7976 4208 -7923
rect 4261 -7976 4271 -7923
rect -2105 -8048 -2029 -8032
rect -2105 -8082 -2089 -8048
rect -2045 -8082 -2029 -8048
rect -2105 -8088 -2029 -8082
rect -1927 -8048 -1851 -8032
rect -1927 -8082 -1911 -8048
rect -1867 -8082 -1851 -8048
rect -1927 -8088 -1851 -8082
rect -1749 -8048 -1673 -8032
rect -1749 -8082 -1733 -8048
rect -1689 -8082 -1673 -8048
rect -1749 -8088 -1673 -8082
rect -1571 -8048 -1495 -8032
rect -1571 -8082 -1555 -8048
rect -1511 -8082 -1495 -8048
rect -1571 -8088 -1495 -8082
rect -1393 -8048 -1317 -8032
rect -1393 -8082 -1377 -8048
rect -1333 -8082 -1317 -8048
rect -1393 -8088 -1317 -8082
rect -1215 -8048 -1139 -8032
rect -1215 -8082 -1199 -8048
rect -1155 -8082 -1139 -8048
rect -1215 -8088 -1139 -8082
rect -1037 -8048 -961 -8032
rect -1037 -8082 -1021 -8048
rect -977 -8082 -961 -8048
rect -1037 -8088 -961 -8082
rect -859 -8048 -783 -8032
rect -859 -8082 -843 -8048
rect -799 -8082 -783 -8048
rect -859 -8088 -783 -8082
rect -681 -8048 -605 -8032
rect -681 -8082 -665 -8048
rect -621 -8082 -605 -8048
rect -681 -8088 -605 -8082
rect -503 -8048 -427 -8032
rect -503 -8082 -487 -8048
rect -443 -8082 -427 -8048
rect -503 -8088 -427 -8082
rect -325 -8048 -249 -8032
rect -325 -8082 -309 -8048
rect -265 -8082 -249 -8048
rect -325 -8088 -249 -8082
rect -147 -8048 -71 -8032
rect -147 -8082 -131 -8048
rect -87 -8082 -71 -8048
rect -147 -8088 -71 -8082
rect 31 -8048 107 -8032
rect 31 -8082 47 -8048
rect 91 -8082 107 -8048
rect 31 -8088 107 -8082
rect 209 -8048 285 -8032
rect 209 -8082 225 -8048
rect 269 -8082 285 -8048
rect 209 -8088 285 -8082
rect 387 -8048 463 -8032
rect 387 -8082 403 -8048
rect 447 -8082 463 -8048
rect 387 -8088 463 -8082
rect 565 -8048 641 -8032
rect 565 -8082 581 -8048
rect 625 -8082 641 -8048
rect 565 -8088 641 -8082
rect 743 -8048 819 -8032
rect 743 -8082 759 -8048
rect 803 -8082 819 -8048
rect 743 -8088 819 -8082
rect 921 -8048 997 -8032
rect 921 -8082 937 -8048
rect 981 -8082 997 -8048
rect 921 -8088 997 -8082
rect 1099 -8048 1175 -8032
rect 1099 -8082 1115 -8048
rect 1159 -8082 1175 -8048
rect 1099 -8088 1175 -8082
rect 1277 -8048 1353 -8032
rect 1277 -8082 1293 -8048
rect 1337 -8082 1353 -8048
rect 1277 -8088 1353 -8082
rect 1455 -8048 1531 -8032
rect 1455 -8082 1471 -8048
rect 1515 -8082 1531 -8048
rect 1455 -8088 1531 -8082
rect 1633 -8048 1709 -8032
rect 1633 -8082 1649 -8048
rect 1693 -8082 1709 -8048
rect 1633 -8088 1709 -8082
rect 1811 -8048 1887 -8032
rect 1811 -8082 1827 -8048
rect 1871 -8082 1887 -8048
rect 1811 -8088 1887 -8082
rect 1989 -8048 2065 -8032
rect 1989 -8082 2005 -8048
rect 2049 -8082 2065 -8048
rect 1989 -8088 2065 -8082
rect 2167 -8048 2243 -8032
rect 2167 -8082 2183 -8048
rect 2227 -8082 2243 -8048
rect 2167 -8088 2243 -8082
rect 2345 -8048 2421 -8032
rect 2345 -8082 2361 -8048
rect 2405 -8082 2421 -8048
rect 2345 -8088 2421 -8082
rect 2523 -8048 2599 -8032
rect 2523 -8082 2539 -8048
rect 2583 -8082 2599 -8048
rect 2523 -8088 2599 -8082
rect 2701 -8048 2777 -8032
rect 2701 -8082 2717 -8048
rect 2761 -8082 2777 -8048
rect 2701 -8088 2777 -8082
rect 2879 -8048 2955 -8032
rect 2879 -8082 2895 -8048
rect 2939 -8082 2955 -8048
rect 2879 -8088 2955 -8082
rect 3057 -8048 3133 -8032
rect 3057 -8082 3073 -8048
rect 3117 -8082 3133 -8048
rect 3057 -8088 3133 -8082
rect 3235 -8048 3311 -8032
rect 3235 -8082 3251 -8048
rect 3295 -8082 3311 -8048
rect 3235 -8088 3311 -8082
rect 3413 -8048 3489 -8032
rect 3413 -8082 3429 -8048
rect 3473 -8082 3489 -8048
rect 3413 -8088 3489 -8082
rect 3591 -8048 3667 -8032
rect 3591 -8082 3607 -8048
rect 3651 -8082 3667 -8048
rect 3591 -8088 3667 -8082
rect 3769 -8048 3845 -8032
rect 3769 -8082 3785 -8048
rect 3829 -8082 3845 -8048
rect 3769 -8088 3845 -8082
rect 3947 -8048 4023 -8032
rect 3947 -8082 3963 -8048
rect 4007 -8082 4023 -8048
rect 3947 -8088 4023 -8082
rect -2179 -8132 -2133 -8120
rect -2179 -8388 -2173 -8132
rect -2139 -8388 -2133 -8132
rect -2179 -8400 -2133 -8388
rect -2001 -8132 -1955 -8120
rect -2001 -8388 -1995 -8132
rect -1961 -8388 -1955 -8132
rect -2001 -8400 -1955 -8388
rect -1823 -8132 -1777 -8120
rect -1823 -8388 -1817 -8132
rect -1783 -8388 -1777 -8132
rect -1823 -8400 -1777 -8388
rect -1645 -8132 -1599 -8120
rect -1645 -8388 -1639 -8132
rect -1605 -8388 -1599 -8132
rect -1645 -8400 -1599 -8388
rect -1467 -8132 -1421 -8120
rect -1467 -8388 -1461 -8132
rect -1427 -8388 -1421 -8132
rect -1467 -8400 -1421 -8388
rect -1289 -8132 -1243 -8120
rect -1289 -8388 -1283 -8132
rect -1249 -8388 -1243 -8132
rect -1289 -8400 -1243 -8388
rect -1111 -8132 -1065 -8120
rect -1111 -8388 -1105 -8132
rect -1071 -8388 -1065 -8132
rect -1111 -8400 -1065 -8388
rect -933 -8132 -887 -8120
rect -933 -8388 -927 -8132
rect -893 -8388 -887 -8132
rect -933 -8400 -887 -8388
rect -755 -8132 -709 -8120
rect -755 -8388 -749 -8132
rect -715 -8388 -709 -8132
rect -755 -8400 -709 -8388
rect -577 -8132 -531 -8120
rect -577 -8388 -571 -8132
rect -537 -8388 -531 -8132
rect -577 -8400 -531 -8388
rect -399 -8132 -353 -8120
rect -399 -8388 -393 -8132
rect -359 -8388 -353 -8132
rect -399 -8400 -353 -8388
rect -221 -8132 -175 -8120
rect -221 -8388 -215 -8132
rect -181 -8388 -175 -8132
rect -221 -8400 -175 -8388
rect -43 -8132 3 -8120
rect -43 -8388 -37 -8132
rect -3 -8388 3 -8132
rect -43 -8400 3 -8388
rect 135 -8132 181 -8120
rect 135 -8388 141 -8132
rect 175 -8388 181 -8132
rect 135 -8400 181 -8388
rect 313 -8132 359 -8120
rect 313 -8388 319 -8132
rect 353 -8388 359 -8132
rect 313 -8400 359 -8388
rect 491 -8132 537 -8120
rect 491 -8388 497 -8132
rect 531 -8388 537 -8132
rect 491 -8400 537 -8388
rect 669 -8132 715 -8120
rect 669 -8388 675 -8132
rect 709 -8388 715 -8132
rect 669 -8400 715 -8388
rect 847 -8132 893 -8120
rect 847 -8388 853 -8132
rect 887 -8388 893 -8132
rect 847 -8400 893 -8388
rect 1025 -8132 1071 -8120
rect 1025 -8388 1031 -8132
rect 1065 -8388 1071 -8132
rect 1025 -8400 1071 -8388
rect 1203 -8132 1249 -8120
rect 1203 -8388 1209 -8132
rect 1243 -8388 1249 -8132
rect 1203 -8400 1249 -8388
rect 1381 -8132 1427 -8120
rect 1381 -8388 1387 -8132
rect 1421 -8388 1427 -8132
rect 1381 -8400 1427 -8388
rect 1559 -8132 1605 -8120
rect 1559 -8388 1565 -8132
rect 1599 -8388 1605 -8132
rect 1559 -8400 1605 -8388
rect 1737 -8132 1783 -8120
rect 1737 -8388 1743 -8132
rect 1777 -8388 1783 -8132
rect 1737 -8400 1783 -8388
rect 1915 -8132 1961 -8120
rect 1915 -8388 1921 -8132
rect 1955 -8388 1961 -8132
rect 1915 -8400 1961 -8388
rect 2093 -8132 2139 -8120
rect 2093 -8388 2099 -8132
rect 2133 -8388 2139 -8132
rect 2093 -8400 2139 -8388
rect 2271 -8132 2317 -8120
rect 2271 -8388 2277 -8132
rect 2311 -8388 2317 -8132
rect 2271 -8400 2317 -8388
rect 2449 -8132 2495 -8120
rect 2449 -8388 2455 -8132
rect 2489 -8388 2495 -8132
rect 2449 -8400 2495 -8388
rect 2627 -8132 2673 -8120
rect 2627 -8388 2633 -8132
rect 2667 -8388 2673 -8132
rect 2627 -8400 2673 -8388
rect 2805 -8132 2851 -8120
rect 2805 -8388 2811 -8132
rect 2845 -8388 2851 -8132
rect 2805 -8400 2851 -8388
rect 2983 -8132 3029 -8120
rect 2983 -8388 2989 -8132
rect 3023 -8388 3029 -8132
rect 2983 -8400 3029 -8388
rect 3161 -8132 3207 -8120
rect 3161 -8388 3167 -8132
rect 3201 -8388 3207 -8132
rect 3161 -8400 3207 -8388
rect 3339 -8132 3385 -8120
rect 3339 -8388 3345 -8132
rect 3379 -8388 3385 -8132
rect 3339 -8400 3385 -8388
rect 3517 -8132 3563 -8120
rect 3517 -8388 3523 -8132
rect 3557 -8388 3563 -8132
rect 3517 -8400 3563 -8388
rect 3695 -8132 3741 -8120
rect 3695 -8388 3701 -8132
rect 3735 -8388 3741 -8132
rect 3695 -8400 3741 -8388
rect 3873 -8132 3919 -8120
rect 3873 -8388 3879 -8132
rect 3913 -8388 3919 -8132
rect 3873 -8400 3919 -8388
rect 4051 -8132 4097 -8120
rect 4051 -8388 4057 -8132
rect 4091 -8388 4097 -8132
rect 4051 -8400 4097 -8388
rect -2171 -8440 -2137 -8400
rect -2105 -8438 -2029 -8432
rect -2105 -8440 -2089 -8438
rect -2171 -8472 -2089 -8440
rect -2045 -8440 -2029 -8438
rect -1995 -8440 -1961 -8400
rect -2045 -8472 -1961 -8440
rect -2171 -8474 -1961 -8472
rect -2105 -8488 -2029 -8474
rect -1995 -8767 -1961 -8474
rect -1927 -8438 -1851 -8432
rect -1927 -8472 -1911 -8438
rect -1867 -8472 -1851 -8438
rect -1927 -8488 -1851 -8472
rect -1906 -8534 -1872 -8488
rect -1926 -8587 -1916 -8534
rect -1863 -8587 -1853 -8534
rect -1817 -8653 -1783 -8400
rect -1749 -8438 -1673 -8432
rect -1749 -8472 -1733 -8438
rect -1689 -8472 -1673 -8438
rect -1749 -8488 -1673 -8472
rect -1729 -8534 -1695 -8488
rect -1749 -8587 -1739 -8534
rect -1686 -8587 -1676 -8534
rect -1836 -8706 -1826 -8653
rect -1773 -8706 -1763 -8653
rect -2457 -8820 -2447 -8767
rect -2394 -8820 -2384 -8767
rect -2015 -8820 -2005 -8767
rect -1952 -8820 -1942 -8767
rect -2997 -9276 -2795 -9270
rect -2997 -9454 -2985 -9276
rect -2807 -9454 -2795 -9276
rect -2997 -9460 -2795 -9454
rect -2997 -11276 -2795 -11270
rect -2997 -11454 -2985 -11276
rect -2807 -11454 -2795 -11276
rect -2997 -11460 -2795 -11454
rect -2447 -12272 -2394 -8820
rect -2105 -9048 -2029 -9032
rect -2105 -9082 -2089 -9048
rect -2045 -9082 -2029 -9048
rect -2105 -9088 -2029 -9082
rect -1995 -9120 -1961 -8820
rect -1927 -9048 -1851 -9032
rect -1927 -9082 -1911 -9048
rect -1867 -9082 -1851 -9048
rect -1927 -9088 -1851 -9082
rect -1817 -9120 -1783 -8706
rect -1639 -8767 -1605 -8400
rect -1571 -8438 -1495 -8432
rect -1571 -8472 -1555 -8438
rect -1511 -8472 -1495 -8438
rect -1571 -8488 -1495 -8472
rect -1549 -8534 -1515 -8488
rect -1568 -8587 -1558 -8534
rect -1505 -8587 -1495 -8534
rect -1461 -8653 -1427 -8400
rect -1393 -8438 -1317 -8432
rect -1393 -8472 -1377 -8438
rect -1333 -8472 -1317 -8438
rect -1393 -8488 -1317 -8472
rect -1392 -8587 -1382 -8534
rect -1329 -8587 -1319 -8534
rect -1480 -8706 -1470 -8653
rect -1417 -8706 -1407 -8653
rect -1658 -8820 -1648 -8767
rect -1595 -8820 -1585 -8767
rect -1749 -9048 -1673 -9032
rect -1749 -9082 -1733 -9048
rect -1689 -9082 -1673 -9048
rect -1749 -9088 -1673 -9082
rect -1639 -9120 -1605 -8820
rect -1571 -9048 -1495 -9032
rect -1571 -9082 -1555 -9048
rect -1511 -9082 -1495 -9048
rect -1571 -9088 -1495 -9082
rect -1461 -9120 -1427 -8706
rect -1372 -9032 -1338 -8587
rect -1283 -8767 -1249 -8400
rect -1215 -8438 -1139 -8432
rect -1215 -8472 -1199 -8438
rect -1155 -8472 -1139 -8438
rect -1215 -8488 -1139 -8472
rect -1213 -8587 -1203 -8534
rect -1150 -8587 -1140 -8534
rect -1303 -8820 -1293 -8767
rect -1240 -8820 -1230 -8767
rect -1393 -9048 -1317 -9032
rect -1393 -9082 -1377 -9048
rect -1333 -9082 -1317 -9048
rect -1393 -9088 -1317 -9082
rect -1283 -9120 -1249 -8820
rect -1193 -9032 -1159 -8587
rect -1105 -8653 -1071 -8400
rect -1037 -8438 -961 -8432
rect -1037 -8472 -1021 -8438
rect -977 -8472 -961 -8438
rect -1037 -8488 -961 -8472
rect -1036 -8587 -1026 -8534
rect -973 -8587 -963 -8534
rect -1125 -8706 -1115 -8653
rect -1062 -8706 -1052 -8653
rect -1215 -9048 -1139 -9032
rect -1215 -9082 -1199 -9048
rect -1155 -9082 -1139 -9048
rect -1215 -9088 -1139 -9082
rect -1105 -9120 -1071 -8706
rect -1016 -9032 -982 -8587
rect -927 -8767 -893 -8400
rect -859 -8438 -783 -8432
rect -859 -8472 -843 -8438
rect -799 -8472 -783 -8438
rect -859 -8488 -783 -8472
rect -858 -8587 -848 -8534
rect -795 -8587 -785 -8534
rect -946 -8820 -936 -8767
rect -883 -8820 -873 -8767
rect -1037 -9048 -961 -9032
rect -1037 -9082 -1021 -9048
rect -977 -9082 -961 -9048
rect -1037 -9088 -961 -9082
rect -927 -9120 -893 -8820
rect -838 -9032 -804 -8587
rect -749 -8653 -715 -8400
rect -681 -8438 -605 -8432
rect -681 -8472 -665 -8438
rect -621 -8472 -605 -8438
rect -681 -8488 -605 -8472
rect -680 -8587 -670 -8534
rect -617 -8587 -607 -8534
rect -768 -8706 -758 -8653
rect -705 -8706 -695 -8653
rect -859 -9048 -783 -9032
rect -859 -9082 -843 -9048
rect -799 -9082 -783 -9048
rect -859 -9088 -783 -9082
rect -749 -9120 -715 -8706
rect -660 -9032 -626 -8587
rect -571 -8766 -537 -8400
rect -503 -8438 -427 -8432
rect -503 -8472 -487 -8438
rect -443 -8472 -427 -8438
rect -503 -8488 -427 -8472
rect -501 -8587 -491 -8534
rect -438 -8587 -428 -8534
rect -590 -8819 -580 -8766
rect -527 -8819 -517 -8766
rect -681 -9048 -605 -9032
rect -681 -9082 -665 -9048
rect -621 -9082 -605 -9048
rect -681 -9088 -605 -9082
rect -571 -9120 -537 -8819
rect -482 -9032 -448 -8587
rect -393 -8653 -359 -8400
rect -325 -8438 -249 -8432
rect -325 -8472 -309 -8438
rect -265 -8472 -249 -8438
rect -325 -8488 -249 -8472
rect -304 -8534 -270 -8488
rect -324 -8587 -314 -8534
rect -261 -8587 -251 -8534
rect -412 -8706 -402 -8653
rect -349 -8706 -339 -8653
rect -503 -9048 -427 -9032
rect -503 -9082 -487 -9048
rect -443 -9082 -427 -9048
rect -503 -9088 -427 -9082
rect -393 -9120 -359 -8706
rect -215 -8767 -181 -8400
rect -147 -8438 -71 -8432
rect -147 -8472 -131 -8438
rect -87 -8472 -71 -8438
rect -147 -8488 -71 -8472
rect -126 -8534 -92 -8488
rect -146 -8587 -136 -8534
rect -83 -8587 -73 -8534
rect -37 -8653 -3 -8400
rect 31 -8438 107 -8432
rect 31 -8472 47 -8438
rect 91 -8472 107 -8438
rect 31 -8488 107 -8472
rect 52 -8534 86 -8488
rect 32 -8587 42 -8534
rect 95 -8587 105 -8534
rect -57 -8706 -47 -8653
rect 6 -8706 16 -8653
rect -235 -8820 -225 -8767
rect -172 -8820 -162 -8767
rect -325 -9048 -249 -9032
rect -325 -9082 -309 -9048
rect -265 -9082 -249 -9048
rect -325 -9088 -249 -9082
rect -215 -9120 -181 -8820
rect -147 -9048 -71 -9032
rect -147 -9082 -131 -9048
rect -87 -9082 -71 -9048
rect -147 -9088 -71 -9082
rect -37 -9120 -3 -8706
rect 141 -8768 175 -8400
rect 209 -8438 285 -8432
rect 209 -8472 225 -8438
rect 269 -8472 285 -8438
rect 209 -8488 285 -8472
rect 230 -8534 264 -8488
rect 211 -8587 221 -8534
rect 274 -8587 284 -8534
rect 319 -8653 353 -8400
rect 387 -8438 463 -8432
rect 387 -8472 403 -8438
rect 447 -8472 463 -8438
rect 387 -8488 463 -8472
rect 408 -8534 442 -8488
rect 388 -8587 398 -8534
rect 451 -8587 461 -8534
rect 300 -8706 310 -8653
rect 363 -8706 373 -8653
rect 122 -8821 132 -8768
rect 185 -8821 195 -8768
rect 31 -9048 107 -9032
rect 31 -9082 47 -9048
rect 91 -9082 107 -9048
rect 31 -9088 107 -9082
rect 141 -9120 175 -8821
rect 209 -9048 285 -9032
rect 209 -9082 225 -9048
rect 269 -9082 285 -9048
rect 209 -9088 285 -9082
rect 319 -9120 353 -8706
rect 497 -8766 531 -8400
rect 565 -8438 641 -8432
rect 565 -8472 581 -8438
rect 625 -8472 641 -8438
rect 565 -8488 641 -8472
rect 586 -8534 620 -8488
rect 567 -8587 577 -8534
rect 630 -8587 640 -8534
rect 675 -8653 709 -8400
rect 743 -8438 819 -8432
rect 743 -8472 759 -8438
rect 803 -8472 819 -8438
rect 743 -8488 819 -8472
rect 744 -8587 754 -8534
rect 807 -8587 817 -8534
rect 656 -8706 666 -8653
rect 719 -8706 729 -8653
rect 479 -8819 489 -8766
rect 542 -8819 552 -8766
rect 387 -9048 463 -9032
rect 387 -9082 403 -9048
rect 447 -9082 463 -9048
rect 387 -9088 463 -9082
rect 497 -9120 531 -8819
rect 565 -9048 641 -9032
rect 565 -9082 581 -9048
rect 625 -9082 641 -9048
rect 565 -9088 641 -9082
rect 675 -9120 709 -8706
rect 764 -9032 798 -8587
rect 853 -8766 887 -8400
rect 921 -8438 997 -8432
rect 921 -8472 937 -8438
rect 981 -8472 997 -8438
rect 921 -8488 997 -8472
rect 922 -8587 932 -8534
rect 985 -8587 995 -8534
rect 833 -8819 843 -8766
rect 896 -8819 906 -8766
rect 743 -9048 819 -9032
rect 743 -9082 759 -9048
rect 803 -9082 819 -9048
rect 743 -9088 819 -9082
rect 853 -9120 887 -8819
rect 942 -9032 976 -8587
rect 1031 -8653 1065 -8400
rect 1099 -8438 1175 -8432
rect 1099 -8472 1115 -8438
rect 1159 -8472 1175 -8438
rect 1099 -8488 1175 -8472
rect 1101 -8587 1111 -8534
rect 1164 -8587 1174 -8534
rect 1012 -8706 1022 -8653
rect 1075 -8706 1085 -8653
rect 921 -9048 997 -9032
rect 921 -9082 937 -9048
rect 981 -9082 997 -9048
rect 921 -9088 997 -9082
rect 1031 -9120 1065 -8706
rect 1120 -9032 1154 -8587
rect 1209 -8767 1243 -8400
rect 1277 -8438 1353 -8432
rect 1277 -8472 1293 -8438
rect 1337 -8472 1353 -8438
rect 1277 -8488 1353 -8472
rect 1279 -8587 1289 -8534
rect 1342 -8587 1352 -8534
rect 1191 -8820 1201 -8767
rect 1254 -8820 1264 -8767
rect 1099 -9048 1175 -9032
rect 1099 -9082 1115 -9048
rect 1159 -9082 1175 -9048
rect 1099 -9088 1175 -9082
rect 1209 -9120 1243 -8820
rect 1298 -9032 1332 -8587
rect 1387 -8653 1421 -8400
rect 1455 -8438 1531 -8432
rect 1455 -8472 1471 -8438
rect 1515 -8472 1531 -8438
rect 1455 -8488 1531 -8472
rect 1456 -8587 1466 -8534
rect 1519 -8587 1529 -8534
rect 1367 -8706 1377 -8653
rect 1430 -8706 1440 -8653
rect 1277 -9048 1353 -9032
rect 1277 -9082 1293 -9048
rect 1337 -9082 1353 -9048
rect 1277 -9088 1353 -9082
rect 1387 -9120 1421 -8706
rect 1476 -9032 1510 -8587
rect 1565 -8767 1599 -8400
rect 1633 -8438 1709 -8432
rect 1633 -8472 1649 -8438
rect 1693 -8472 1709 -8438
rect 1633 -8488 1709 -8472
rect 1634 -8587 1644 -8534
rect 1697 -8587 1707 -8534
rect 1546 -8820 1556 -8767
rect 1609 -8820 1619 -8767
rect 1455 -9048 1531 -9032
rect 1455 -9082 1471 -9048
rect 1515 -9082 1531 -9048
rect 1455 -9088 1531 -9082
rect 1565 -9120 1599 -8820
rect 1654 -9032 1688 -8587
rect 1743 -8653 1777 -8400
rect 1811 -8438 1887 -8432
rect 1811 -8472 1827 -8438
rect 1871 -8472 1887 -8438
rect 1811 -8488 1887 -8472
rect 1832 -8534 1866 -8488
rect 1812 -8587 1822 -8534
rect 1875 -8587 1885 -8534
rect 1723 -8706 1733 -8653
rect 1786 -8706 1796 -8653
rect 1633 -9048 1709 -9032
rect 1633 -9082 1649 -9048
rect 1693 -9082 1709 -9048
rect 1633 -9088 1709 -9082
rect 1743 -9120 1777 -8706
rect 1921 -8767 1955 -8400
rect 1989 -8438 2065 -8432
rect 1989 -8472 2005 -8438
rect 2049 -8472 2065 -8438
rect 1989 -8488 2065 -8472
rect 2010 -8534 2044 -8488
rect 1990 -8587 2000 -8534
rect 2053 -8587 2063 -8534
rect 2099 -8653 2133 -8400
rect 2167 -8438 2243 -8432
rect 2167 -8472 2183 -8438
rect 2227 -8472 2243 -8438
rect 2167 -8488 2243 -8472
rect 2188 -8534 2222 -8488
rect 2168 -8587 2178 -8534
rect 2231 -8587 2241 -8534
rect 2080 -8706 2090 -8653
rect 2143 -8706 2153 -8653
rect 1901 -8820 1911 -8767
rect 1964 -8820 1974 -8767
rect 1811 -9048 1887 -9032
rect 1811 -9082 1827 -9048
rect 1871 -9082 1887 -9048
rect 1811 -9088 1887 -9082
rect 1921 -9120 1955 -8820
rect 1989 -9048 2065 -9032
rect 1989 -9082 2005 -9048
rect 2049 -9082 2065 -9048
rect 1989 -9088 2065 -9082
rect 2099 -9120 2133 -8706
rect 2277 -8767 2311 -8400
rect 2345 -8438 2421 -8432
rect 2345 -8472 2361 -8438
rect 2405 -8472 2421 -8438
rect 2345 -8488 2421 -8472
rect 2367 -8534 2401 -8488
rect 2347 -8587 2357 -8534
rect 2410 -8587 2420 -8534
rect 2455 -8653 2489 -8400
rect 2523 -8438 2599 -8432
rect 2523 -8472 2539 -8438
rect 2583 -8472 2599 -8438
rect 2523 -8488 2599 -8472
rect 2544 -8534 2578 -8488
rect 2524 -8587 2534 -8534
rect 2587 -8587 2597 -8534
rect 2436 -8706 2446 -8653
rect 2499 -8706 2509 -8653
rect 2257 -8820 2267 -8767
rect 2320 -8820 2330 -8767
rect 2167 -9048 2243 -9032
rect 2167 -9082 2183 -9048
rect 2227 -9082 2243 -9048
rect 2167 -9088 2243 -9082
rect 2277 -9120 2311 -8820
rect 2345 -9048 2421 -9032
rect 2345 -9082 2361 -9048
rect 2405 -9082 2421 -9048
rect 2345 -9088 2421 -9082
rect 2455 -9120 2489 -8706
rect 2633 -8767 2667 -8400
rect 2701 -8438 2777 -8432
rect 2701 -8472 2717 -8438
rect 2761 -8472 2777 -8438
rect 2701 -8488 2777 -8472
rect 2722 -8534 2756 -8488
rect 2702 -8587 2712 -8534
rect 2765 -8587 2775 -8534
rect 2811 -8653 2845 -8400
rect 2879 -8438 2955 -8432
rect 2879 -8472 2895 -8438
rect 2939 -8472 2955 -8438
rect 2879 -8488 2955 -8472
rect 2880 -8587 2890 -8534
rect 2943 -8587 2953 -8534
rect 2792 -8706 2802 -8653
rect 2855 -8706 2865 -8653
rect 2614 -8820 2624 -8767
rect 2677 -8820 2687 -8767
rect 2523 -9048 2599 -9032
rect 2523 -9082 2539 -9048
rect 2583 -9082 2599 -9048
rect 2523 -9088 2599 -9082
rect 2633 -9120 2667 -8820
rect 2701 -9048 2777 -9032
rect 2701 -9082 2717 -9048
rect 2761 -9082 2777 -9048
rect 2701 -9088 2777 -9082
rect 2811 -9120 2845 -8706
rect 2900 -9032 2934 -8587
rect 2989 -8767 3023 -8400
rect 3057 -8438 3133 -8432
rect 3057 -8472 3073 -8438
rect 3117 -8472 3133 -8438
rect 3057 -8488 3133 -8472
rect 3058 -8587 3068 -8534
rect 3121 -8587 3131 -8534
rect 2970 -8820 2980 -8767
rect 3033 -8820 3043 -8767
rect 2879 -9048 2955 -9032
rect 2879 -9082 2895 -9048
rect 2939 -9082 2955 -9048
rect 2879 -9088 2955 -9082
rect 2989 -9120 3023 -8820
rect 3078 -9032 3112 -8587
rect 3167 -8653 3201 -8400
rect 3235 -8438 3311 -8432
rect 3235 -8472 3251 -8438
rect 3295 -8472 3311 -8438
rect 3235 -8488 3311 -8472
rect 3236 -8587 3246 -8534
rect 3299 -8587 3309 -8534
rect 3148 -8706 3158 -8653
rect 3211 -8706 3221 -8653
rect 3057 -9048 3133 -9032
rect 3057 -9082 3073 -9048
rect 3117 -9082 3133 -9048
rect 3057 -9088 3133 -9082
rect 3167 -9120 3201 -8706
rect 3256 -9032 3290 -8587
rect 3345 -8767 3379 -8400
rect 3413 -8438 3489 -8432
rect 3413 -8472 3429 -8438
rect 3473 -8472 3489 -8438
rect 3413 -8488 3489 -8472
rect 3414 -8587 3424 -8534
rect 3477 -8587 3487 -8534
rect 3326 -8820 3336 -8767
rect 3389 -8820 3399 -8767
rect 3235 -9048 3311 -9032
rect 3235 -9082 3251 -9048
rect 3295 -9082 3311 -9048
rect 3235 -9088 3311 -9082
rect 3345 -9120 3379 -8820
rect 3434 -9032 3468 -8587
rect 3523 -8653 3557 -8400
rect 3591 -8438 3667 -8432
rect 3591 -8472 3607 -8438
rect 3651 -8472 3667 -8438
rect 3591 -8488 3667 -8472
rect 3592 -8587 3602 -8534
rect 3655 -8587 3665 -8534
rect 3503 -8706 3513 -8653
rect 3566 -8706 3576 -8653
rect 3413 -9048 3489 -9032
rect 3413 -9082 3429 -9048
rect 3473 -9082 3489 -9048
rect 3413 -9088 3489 -9082
rect 3523 -9120 3557 -8706
rect 3612 -9032 3646 -8587
rect 3701 -8767 3735 -8400
rect 3769 -8438 3845 -8432
rect 3769 -8472 3785 -8438
rect 3829 -8472 3845 -8438
rect 3769 -8488 3845 -8472
rect 3879 -8440 3913 -8400
rect 3947 -8438 4023 -8432
rect 3947 -8440 3963 -8438
rect 3879 -8472 3963 -8440
rect 4007 -8440 4023 -8438
rect 4056 -8440 4090 -8400
rect 4007 -8472 4090 -8440
rect 3879 -8474 4090 -8472
rect 3771 -8587 3781 -8534
rect 3834 -8587 3844 -8534
rect 3682 -8820 3692 -8767
rect 3745 -8820 3755 -8767
rect 3591 -9048 3667 -9032
rect 3591 -9082 3607 -9048
rect 3651 -9082 3667 -9048
rect 3591 -9088 3667 -9082
rect 3701 -9120 3735 -8820
rect 3790 -9032 3824 -8587
rect 3879 -8653 3913 -8474
rect 3947 -8488 4023 -8474
rect 3859 -8706 3869 -8653
rect 3922 -8706 3932 -8653
rect 3769 -9048 3845 -9032
rect 3769 -9082 3785 -9048
rect 3829 -9082 3845 -9048
rect 3769 -9088 3845 -9082
rect 3879 -9120 3913 -8706
rect 3947 -9048 4023 -9032
rect 3947 -9082 3963 -9048
rect 4007 -9082 4023 -9048
rect 3947 -9088 4023 -9082
rect -2179 -9132 -2133 -9120
rect -2179 -9388 -2173 -9132
rect -2139 -9388 -2133 -9132
rect -2179 -9400 -2133 -9388
rect -2001 -9132 -1955 -9120
rect -2001 -9388 -1995 -9132
rect -1961 -9388 -1955 -9132
rect -2001 -9400 -1955 -9388
rect -1823 -9132 -1777 -9120
rect -1823 -9388 -1817 -9132
rect -1783 -9388 -1777 -9132
rect -1823 -9400 -1777 -9388
rect -1645 -9132 -1599 -9120
rect -1645 -9388 -1639 -9132
rect -1605 -9388 -1599 -9132
rect -1645 -9400 -1599 -9388
rect -1467 -9132 -1421 -9120
rect -1467 -9388 -1461 -9132
rect -1427 -9388 -1421 -9132
rect -1467 -9400 -1421 -9388
rect -1289 -9132 -1243 -9120
rect -1289 -9388 -1283 -9132
rect -1249 -9388 -1243 -9132
rect -1289 -9400 -1243 -9388
rect -1111 -9132 -1065 -9120
rect -1111 -9388 -1105 -9132
rect -1071 -9388 -1065 -9132
rect -1111 -9400 -1065 -9388
rect -933 -9132 -887 -9120
rect -933 -9388 -927 -9132
rect -893 -9388 -887 -9132
rect -933 -9400 -887 -9388
rect -755 -9132 -709 -9120
rect -755 -9388 -749 -9132
rect -715 -9388 -709 -9132
rect -755 -9400 -709 -9388
rect -577 -9132 -531 -9120
rect -577 -9388 -571 -9132
rect -537 -9388 -531 -9132
rect -577 -9400 -531 -9388
rect -399 -9132 -353 -9120
rect -399 -9388 -393 -9132
rect -359 -9388 -353 -9132
rect -399 -9400 -353 -9388
rect -221 -9132 -175 -9120
rect -221 -9388 -215 -9132
rect -181 -9388 -175 -9132
rect -221 -9400 -175 -9388
rect -43 -9132 3 -9120
rect -43 -9388 -37 -9132
rect -3 -9388 3 -9132
rect -43 -9400 3 -9388
rect 135 -9132 181 -9120
rect 135 -9388 141 -9132
rect 175 -9388 181 -9132
rect 135 -9400 181 -9388
rect 313 -9132 359 -9120
rect 313 -9388 319 -9132
rect 353 -9388 359 -9132
rect 313 -9400 359 -9388
rect 491 -9132 537 -9120
rect 491 -9388 497 -9132
rect 531 -9388 537 -9132
rect 491 -9400 537 -9388
rect 669 -9132 715 -9120
rect 669 -9388 675 -9132
rect 709 -9388 715 -9132
rect 669 -9400 715 -9388
rect 847 -9132 893 -9120
rect 847 -9388 853 -9132
rect 887 -9388 893 -9132
rect 847 -9400 893 -9388
rect 1025 -9132 1071 -9120
rect 1025 -9388 1031 -9132
rect 1065 -9388 1071 -9132
rect 1025 -9400 1071 -9388
rect 1203 -9132 1249 -9120
rect 1203 -9388 1209 -9132
rect 1243 -9388 1249 -9132
rect 1203 -9400 1249 -9388
rect 1381 -9132 1427 -9120
rect 1381 -9388 1387 -9132
rect 1421 -9388 1427 -9132
rect 1381 -9400 1427 -9388
rect 1559 -9132 1605 -9120
rect 1559 -9388 1565 -9132
rect 1599 -9388 1605 -9132
rect 1559 -9400 1605 -9388
rect 1737 -9132 1783 -9120
rect 1737 -9388 1743 -9132
rect 1777 -9388 1783 -9132
rect 1737 -9400 1783 -9388
rect 1915 -9132 1961 -9120
rect 1915 -9388 1921 -9132
rect 1955 -9388 1961 -9132
rect 1915 -9400 1961 -9388
rect 2093 -9132 2139 -9120
rect 2093 -9388 2099 -9132
rect 2133 -9388 2139 -9132
rect 2093 -9400 2139 -9388
rect 2271 -9132 2317 -9120
rect 2271 -9388 2277 -9132
rect 2311 -9388 2317 -9132
rect 2271 -9400 2317 -9388
rect 2449 -9132 2495 -9120
rect 2449 -9388 2455 -9132
rect 2489 -9388 2495 -9132
rect 2449 -9400 2495 -9388
rect 2627 -9132 2673 -9120
rect 2627 -9388 2633 -9132
rect 2667 -9388 2673 -9132
rect 2627 -9400 2673 -9388
rect 2805 -9132 2851 -9120
rect 2805 -9388 2811 -9132
rect 2845 -9388 2851 -9132
rect 2805 -9400 2851 -9388
rect 2983 -9132 3029 -9120
rect 2983 -9388 2989 -9132
rect 3023 -9388 3029 -9132
rect 2983 -9400 3029 -9388
rect 3161 -9132 3207 -9120
rect 3161 -9388 3167 -9132
rect 3201 -9388 3207 -9132
rect 3161 -9400 3207 -9388
rect 3339 -9132 3385 -9120
rect 3339 -9388 3345 -9132
rect 3379 -9388 3385 -9132
rect 3339 -9400 3385 -9388
rect 3517 -9132 3563 -9120
rect 3517 -9388 3523 -9132
rect 3557 -9388 3563 -9132
rect 3517 -9400 3563 -9388
rect 3695 -9132 3741 -9120
rect 3695 -9388 3701 -9132
rect 3735 -9388 3741 -9132
rect 3695 -9400 3741 -9388
rect 3873 -9132 3919 -9120
rect 3873 -9388 3879 -9132
rect 3913 -9388 3919 -9132
rect 3873 -9400 3919 -9388
rect 4051 -9132 4097 -9120
rect 4051 -9388 4057 -9132
rect 4091 -9388 4097 -9132
rect 4051 -9400 4097 -9388
rect -2174 -9439 -2140 -9400
rect -2105 -9438 -2029 -9432
rect -2105 -9439 -2089 -9438
rect -2174 -9472 -2089 -9439
rect -2045 -9439 -2029 -9438
rect -1995 -9439 -1961 -9400
rect -2045 -9472 -1961 -9439
rect -2174 -9473 -1961 -9472
rect -2105 -9488 -2029 -9473
rect -2325 -9978 -2315 -9925
rect -2262 -9978 -2252 -9925
rect -2457 -12325 -2447 -12272
rect -2394 -12325 -2384 -12272
rect -2997 -13276 -2795 -13270
rect -2997 -13454 -2985 -13276
rect -2807 -13454 -2795 -13276
rect -2997 -13460 -2795 -13454
rect -3392 -14108 -3382 -14055
rect -3329 -14108 -3319 -14055
rect -4248 -14959 -4036 -14925
rect -3946 -14954 -3936 -14901
rect -3883 -14954 -3611 -14901
rect -4536 -15010 -4460 -14994
rect -4536 -15044 -4520 -15010
rect -4476 -15044 -4460 -15010
rect -4536 -15050 -4460 -15044
rect -4358 -15010 -4282 -14994
rect -4358 -15044 -4342 -15010
rect -4298 -15044 -4282 -15010
rect -4358 -15050 -4282 -15044
rect -4248 -15082 -4214 -14959
rect -4159 -14994 -4125 -14959
rect -4180 -15010 -4104 -14994
rect -4180 -15044 -4164 -15010
rect -4120 -15044 -4104 -15010
rect -4180 -15050 -4104 -15044
rect -4070 -15082 -4036 -14959
rect -3936 -15006 -3883 -14954
rect -6034 -15094 -5988 -15082
rect -6034 -15350 -6028 -15094
rect -5994 -15350 -5988 -15094
rect -6034 -15362 -5988 -15350
rect -5856 -15094 -5810 -15082
rect -5856 -15350 -5850 -15094
rect -5816 -15350 -5810 -15094
rect -5856 -15362 -5810 -15350
rect -5678 -15094 -5632 -15082
rect -5678 -15350 -5672 -15094
rect -5638 -15350 -5632 -15094
rect -5678 -15362 -5632 -15350
rect -5500 -15094 -5454 -15082
rect -5500 -15350 -5494 -15094
rect -5460 -15350 -5454 -15094
rect -5500 -15362 -5454 -15350
rect -5322 -15094 -5276 -15082
rect -5322 -15350 -5316 -15094
rect -5282 -15350 -5276 -15094
rect -5322 -15362 -5276 -15350
rect -5144 -15094 -5098 -15082
rect -5144 -15350 -5138 -15094
rect -5104 -15350 -5098 -15094
rect -5144 -15362 -5098 -15350
rect -4966 -15094 -4920 -15082
rect -4966 -15350 -4960 -15094
rect -4926 -15350 -4920 -15094
rect -4966 -15362 -4920 -15350
rect -4788 -15094 -4742 -15082
rect -4788 -15350 -4782 -15094
rect -4748 -15350 -4742 -15094
rect -4788 -15362 -4742 -15350
rect -4610 -15094 -4564 -15082
rect -4610 -15350 -4604 -15094
rect -4570 -15350 -4564 -15094
rect -4610 -15362 -4564 -15350
rect -4432 -15094 -4386 -15082
rect -4432 -15350 -4426 -15094
rect -4392 -15350 -4386 -15094
rect -4432 -15362 -4386 -15350
rect -4254 -15094 -4208 -15082
rect -4254 -15350 -4248 -15094
rect -4214 -15350 -4208 -15094
rect -4254 -15362 -4208 -15350
rect -4076 -15094 -4030 -15082
rect -4076 -15350 -4070 -15094
rect -4036 -15350 -4030 -15094
rect -4076 -15362 -4030 -15350
rect -5960 -15400 -5884 -15394
rect -5960 -15434 -5944 -15400
rect -5900 -15434 -5884 -15400
rect -5960 -15450 -5884 -15434
rect -6169 -15535 -6159 -15482
rect -6106 -15535 -6096 -15482
rect -6159 -16193 -6106 -15535
rect -5850 -15588 -5816 -15362
rect -5782 -15400 -5706 -15394
rect -5782 -15434 -5766 -15400
rect -5722 -15434 -5706 -15400
rect -5782 -15450 -5706 -15434
rect -5870 -15641 -5860 -15588
rect -5807 -15641 -5797 -15588
rect -5761 -15694 -5727 -15450
rect -5960 -15710 -5884 -15694
rect -5960 -15744 -5944 -15710
rect -5900 -15744 -5884 -15710
rect -5960 -15750 -5884 -15744
rect -5782 -15710 -5706 -15694
rect -5782 -15744 -5766 -15710
rect -5722 -15744 -5706 -15710
rect -5782 -15750 -5706 -15744
rect -5672 -15782 -5638 -15362
rect -5604 -15400 -5528 -15394
rect -5604 -15434 -5588 -15400
rect -5544 -15434 -5528 -15400
rect -5604 -15450 -5528 -15434
rect -5583 -15694 -5549 -15450
rect -5494 -15481 -5460 -15362
rect -5426 -15400 -5350 -15394
rect -5426 -15434 -5410 -15400
rect -5366 -15434 -5350 -15400
rect -5426 -15450 -5350 -15434
rect -5514 -15534 -5504 -15481
rect -5451 -15534 -5441 -15481
rect -5405 -15694 -5371 -15450
rect -5604 -15710 -5528 -15694
rect -5604 -15744 -5588 -15710
rect -5544 -15744 -5528 -15710
rect -5604 -15750 -5528 -15744
rect -5426 -15710 -5350 -15694
rect -5426 -15744 -5410 -15710
rect -5366 -15744 -5350 -15710
rect -5426 -15750 -5350 -15744
rect -5316 -15782 -5282 -15362
rect -5248 -15400 -5172 -15394
rect -5248 -15434 -5232 -15400
rect -5188 -15434 -5172 -15400
rect -5248 -15450 -5172 -15434
rect -5227 -15694 -5193 -15450
rect -5138 -15589 -5104 -15362
rect -5070 -15400 -4994 -15394
rect -5070 -15434 -5054 -15400
rect -5010 -15434 -4994 -15400
rect -5070 -15450 -4994 -15434
rect -5158 -15642 -5148 -15589
rect -5095 -15642 -5085 -15589
rect -5049 -15694 -5015 -15450
rect -5248 -15710 -5172 -15694
rect -5248 -15744 -5232 -15710
rect -5188 -15744 -5172 -15710
rect -5248 -15750 -5172 -15744
rect -5070 -15710 -4994 -15694
rect -5070 -15744 -5054 -15710
rect -5010 -15744 -4994 -15710
rect -5070 -15750 -4994 -15744
rect -4960 -15782 -4926 -15362
rect -4892 -15400 -4816 -15394
rect -4892 -15434 -4876 -15400
rect -4832 -15434 -4816 -15400
rect -4892 -15450 -4816 -15434
rect -4871 -15694 -4837 -15450
rect -4782 -15481 -4748 -15362
rect -4714 -15400 -4638 -15394
rect -4714 -15434 -4698 -15400
rect -4654 -15434 -4638 -15400
rect -4714 -15450 -4638 -15434
rect -4802 -15534 -4792 -15481
rect -4739 -15534 -4729 -15481
rect -4693 -15694 -4659 -15450
rect -4892 -15710 -4816 -15694
rect -4892 -15744 -4876 -15710
rect -4832 -15744 -4816 -15710
rect -4892 -15750 -4816 -15744
rect -4714 -15710 -4638 -15694
rect -4714 -15744 -4698 -15710
rect -4654 -15744 -4638 -15710
rect -4714 -15750 -4638 -15744
rect -4604 -15782 -4570 -15362
rect -4536 -15400 -4460 -15394
rect -4536 -15434 -4520 -15400
rect -4476 -15434 -4460 -15400
rect -4536 -15450 -4460 -15434
rect -4515 -15694 -4481 -15450
rect -4426 -15589 -4392 -15362
rect -4358 -15400 -4282 -15394
rect -4358 -15434 -4342 -15400
rect -4298 -15434 -4282 -15400
rect -4358 -15450 -4282 -15434
rect -4445 -15641 -4435 -15589
rect -4383 -15641 -4373 -15589
rect -4337 -15694 -4303 -15450
rect -4536 -15710 -4460 -15694
rect -4536 -15744 -4520 -15710
rect -4476 -15744 -4460 -15710
rect -4536 -15750 -4460 -15744
rect -4358 -15710 -4282 -15694
rect -4358 -15744 -4342 -15710
rect -4298 -15744 -4282 -15710
rect -4358 -15750 -4282 -15744
rect -4248 -15782 -4214 -15362
rect -4180 -15400 -4104 -15394
rect -4180 -15434 -4164 -15400
rect -4120 -15434 -4104 -15400
rect -4180 -15450 -4104 -15434
rect -3935 -15589 -3883 -15006
rect -2997 -15276 -2795 -15270
rect -2997 -15454 -2985 -15276
rect -2807 -15454 -2795 -15276
rect -2997 -15460 -2795 -15454
rect -3945 -15641 -3935 -15589
rect -3883 -15641 -3873 -15589
rect -4180 -15710 -4104 -15694
rect -4180 -15744 -4164 -15710
rect -4120 -15744 -4104 -15710
rect -4180 -15750 -4104 -15744
rect -6034 -15794 -5988 -15782
rect -6034 -16050 -6028 -15794
rect -5994 -16050 -5988 -15794
rect -6034 -16062 -5988 -16050
rect -5856 -15794 -5810 -15782
rect -5856 -16050 -5850 -15794
rect -5816 -16050 -5810 -15794
rect -5856 -16062 -5810 -16050
rect -5678 -15794 -5632 -15782
rect -5678 -16050 -5672 -15794
rect -5638 -16050 -5632 -15794
rect -5678 -16062 -5632 -16050
rect -5500 -15794 -5454 -15782
rect -5500 -16050 -5494 -15794
rect -5460 -16050 -5454 -15794
rect -5500 -16062 -5454 -16050
rect -5322 -15794 -5276 -15782
rect -5322 -16050 -5316 -15794
rect -5282 -16050 -5276 -15794
rect -5322 -16062 -5276 -16050
rect -5144 -15794 -5098 -15782
rect -5144 -16050 -5138 -15794
rect -5104 -16050 -5098 -15794
rect -5144 -16062 -5098 -16050
rect -4966 -15794 -4920 -15782
rect -4966 -16050 -4960 -15794
rect -4926 -16050 -4920 -15794
rect -4966 -16062 -4920 -16050
rect -4788 -15794 -4742 -15782
rect -4788 -16050 -4782 -15794
rect -4748 -16050 -4742 -15794
rect -4788 -16062 -4742 -16050
rect -4610 -15794 -4564 -15782
rect -4610 -16050 -4604 -15794
rect -4570 -16050 -4564 -15794
rect -4610 -16062 -4564 -16050
rect -4432 -15794 -4386 -15782
rect -4432 -16050 -4426 -15794
rect -4392 -16050 -4386 -15794
rect -4432 -16062 -4386 -16050
rect -4254 -15794 -4208 -15782
rect -4254 -16050 -4248 -15794
rect -4214 -16050 -4208 -15794
rect -4254 -16062 -4208 -16050
rect -4076 -15794 -4030 -15782
rect -4076 -16050 -4070 -15794
rect -4036 -16050 -4030 -15794
rect -4076 -16062 -4030 -16050
rect -6028 -16185 -5994 -16062
rect -5960 -16100 -5884 -16094
rect -5960 -16134 -5944 -16100
rect -5900 -16134 -5884 -16100
rect -5960 -16150 -5884 -16134
rect -5939 -16185 -5905 -16150
rect -5850 -16185 -5816 -16062
rect -5782 -16100 -5706 -16094
rect -5782 -16134 -5766 -16100
rect -5722 -16134 -5706 -16100
rect -5782 -16150 -5706 -16134
rect -6169 -16246 -6159 -16193
rect -6106 -16246 -6096 -16193
rect -6028 -16219 -5816 -16185
rect -6159 -17007 -6106 -16246
rect -5850 -16294 -5816 -16219
rect -5870 -16347 -5860 -16294
rect -5807 -16347 -5797 -16294
rect -5761 -16394 -5727 -16150
rect -5960 -16410 -5884 -16394
rect -5960 -16444 -5944 -16410
rect -5900 -16444 -5884 -16410
rect -5960 -16450 -5884 -16444
rect -5782 -16410 -5706 -16394
rect -5782 -16444 -5766 -16410
rect -5722 -16444 -5706 -16410
rect -5782 -16450 -5706 -16444
rect -5672 -16482 -5638 -16062
rect -5604 -16100 -5528 -16094
rect -5604 -16134 -5588 -16100
rect -5544 -16134 -5528 -16100
rect -5604 -16150 -5528 -16134
rect -5583 -16394 -5549 -16150
rect -5494 -16193 -5460 -16062
rect -5426 -16100 -5350 -16094
rect -5426 -16134 -5410 -16100
rect -5366 -16134 -5350 -16100
rect -5426 -16150 -5350 -16134
rect -5514 -16246 -5504 -16193
rect -5451 -16246 -5441 -16193
rect -5405 -16394 -5371 -16150
rect -5604 -16410 -5528 -16394
rect -5604 -16444 -5588 -16410
rect -5544 -16444 -5528 -16410
rect -5604 -16450 -5528 -16444
rect -5426 -16410 -5350 -16394
rect -5426 -16444 -5410 -16410
rect -5366 -16444 -5350 -16410
rect -5426 -16450 -5350 -16444
rect -5316 -16482 -5282 -16062
rect -5248 -16100 -5172 -16094
rect -5248 -16134 -5232 -16100
rect -5188 -16134 -5172 -16100
rect -5248 -16150 -5172 -16134
rect -5227 -16394 -5193 -16150
rect -5138 -16294 -5104 -16062
rect -5070 -16100 -4994 -16094
rect -5070 -16134 -5054 -16100
rect -5010 -16134 -4994 -16100
rect -5070 -16150 -4994 -16134
rect -5158 -16347 -5148 -16294
rect -5095 -16347 -5085 -16294
rect -5049 -16394 -5015 -16150
rect -5248 -16410 -5172 -16394
rect -5248 -16444 -5232 -16410
rect -5188 -16444 -5172 -16410
rect -5248 -16450 -5172 -16444
rect -5070 -16410 -4994 -16394
rect -5070 -16444 -5054 -16410
rect -5010 -16444 -4994 -16410
rect -5070 -16450 -4994 -16444
rect -4960 -16482 -4926 -16062
rect -4892 -16100 -4816 -16094
rect -4892 -16134 -4876 -16100
rect -4832 -16134 -4816 -16100
rect -4892 -16150 -4816 -16134
rect -4871 -16394 -4837 -16150
rect -4782 -16193 -4748 -16062
rect -4714 -16100 -4638 -16094
rect -4714 -16134 -4698 -16100
rect -4654 -16134 -4638 -16100
rect -4714 -16150 -4638 -16134
rect -4802 -16246 -4792 -16193
rect -4739 -16246 -4729 -16193
rect -4693 -16394 -4659 -16150
rect -4892 -16410 -4816 -16394
rect -4892 -16444 -4876 -16410
rect -4832 -16444 -4816 -16410
rect -4892 -16450 -4816 -16444
rect -4714 -16410 -4638 -16394
rect -4714 -16444 -4698 -16410
rect -4654 -16444 -4638 -16410
rect -4714 -16450 -4638 -16444
rect -4604 -16482 -4570 -16062
rect -4536 -16100 -4460 -16094
rect -4536 -16134 -4520 -16100
rect -4476 -16134 -4460 -16100
rect -4536 -16150 -4460 -16134
rect -4515 -16394 -4481 -16150
rect -4426 -16294 -4392 -16062
rect -4358 -16100 -4282 -16094
rect -4358 -16134 -4342 -16100
rect -4298 -16134 -4282 -16100
rect -4358 -16150 -4282 -16134
rect -4446 -16347 -4436 -16294
rect -4383 -16347 -4373 -16294
rect -4337 -16394 -4303 -16150
rect -4248 -16185 -4214 -16062
rect -4180 -16100 -4104 -16094
rect -4180 -16134 -4164 -16100
rect -4120 -16134 -4104 -16100
rect -4180 -16150 -4104 -16134
rect -4159 -16185 -4125 -16150
rect -4070 -16185 -4036 -16062
rect -4248 -16219 -4036 -16185
rect -4536 -16410 -4460 -16394
rect -4536 -16444 -4520 -16410
rect -4476 -16444 -4460 -16410
rect -4536 -16450 -4460 -16444
rect -4358 -16410 -4282 -16394
rect -4358 -16444 -4342 -16410
rect -4298 -16444 -4282 -16410
rect -4358 -16450 -4282 -16444
rect -4248 -16482 -4214 -16219
rect -3935 -16295 -3883 -15641
rect -2447 -15821 -2394 -12325
rect -2315 -14543 -2262 -9978
rect -2105 -10048 -2029 -10032
rect -2105 -10049 -2089 -10048
rect -2175 -10082 -2089 -10049
rect -2045 -10049 -2029 -10048
rect -1995 -10049 -1961 -9473
rect -1927 -9438 -1851 -9432
rect -1927 -9472 -1911 -9438
rect -1867 -9472 -1851 -9438
rect -1927 -9488 -1851 -9472
rect -1906 -9546 -1872 -9488
rect -1926 -9599 -1916 -9546
rect -1863 -9599 -1853 -9546
rect -1926 -9978 -1916 -9925
rect -1863 -9978 -1853 -9925
rect -1906 -10032 -1872 -9978
rect -2045 -10082 -1961 -10049
rect -2175 -10083 -1961 -10082
rect -2175 -10120 -2141 -10083
rect -2105 -10088 -2029 -10083
rect -1995 -10120 -1961 -10083
rect -1927 -10048 -1851 -10032
rect -1927 -10082 -1911 -10048
rect -1867 -10082 -1851 -10048
rect -1927 -10088 -1851 -10082
rect -1817 -10120 -1783 -9400
rect -1749 -9438 -1673 -9432
rect -1749 -9472 -1733 -9438
rect -1689 -9472 -1673 -9438
rect -1749 -9488 -1673 -9472
rect -1728 -9546 -1694 -9488
rect -1748 -9599 -1738 -9546
rect -1685 -9599 -1675 -9546
rect -1748 -9979 -1738 -9926
rect -1685 -9979 -1675 -9926
rect -1728 -10032 -1694 -9979
rect -1749 -10048 -1673 -10032
rect -1749 -10082 -1733 -10048
rect -1689 -10082 -1673 -10048
rect -1749 -10088 -1673 -10082
rect -1639 -10120 -1605 -9400
rect -1571 -9438 -1495 -9432
rect -1571 -9472 -1555 -9438
rect -1511 -9472 -1495 -9438
rect -1571 -9488 -1495 -9472
rect -1549 -9546 -1515 -9488
rect -1568 -9599 -1558 -9546
rect -1505 -9599 -1495 -9546
rect -1570 -9978 -1560 -9925
rect -1507 -9978 -1497 -9925
rect -1550 -10032 -1516 -9978
rect -1571 -10048 -1495 -10032
rect -1571 -10082 -1555 -10048
rect -1511 -10082 -1495 -10048
rect -1571 -10088 -1495 -10082
rect -1461 -10120 -1427 -9400
rect -1393 -9438 -1317 -9432
rect -1393 -9472 -1377 -9438
rect -1333 -9472 -1317 -9438
rect -1393 -9488 -1317 -9472
rect -1372 -9924 -1338 -9488
rect -1392 -9977 -1382 -9924
rect -1329 -9977 -1319 -9924
rect -1393 -10048 -1317 -10032
rect -1393 -10082 -1377 -10048
rect -1333 -10082 -1317 -10048
rect -1393 -10088 -1317 -10082
rect -1283 -10120 -1249 -9400
rect -1215 -9438 -1139 -9432
rect -1215 -9472 -1199 -9438
rect -1155 -9472 -1139 -9438
rect -1215 -9488 -1139 -9472
rect -1215 -10048 -1139 -10032
rect -1215 -10082 -1199 -10048
rect -1155 -10082 -1139 -10048
rect -1215 -10088 -1139 -10082
rect -1105 -10120 -1071 -9400
rect -1037 -9438 -961 -9432
rect -1037 -9472 -1021 -9438
rect -977 -9472 -961 -9438
rect -1037 -9488 -961 -9472
rect -1037 -10048 -961 -10032
rect -1037 -10082 -1021 -10048
rect -977 -10082 -961 -10048
rect -1037 -10088 -961 -10082
rect -927 -10120 -893 -9400
rect -859 -9438 -783 -9432
rect -859 -9472 -843 -9438
rect -799 -9472 -783 -9438
rect -859 -9488 -783 -9472
rect -859 -10048 -783 -10032
rect -859 -10082 -843 -10048
rect -799 -10082 -783 -10048
rect -859 -10088 -783 -10082
rect -749 -10120 -715 -9400
rect -681 -9438 -605 -9432
rect -681 -9472 -665 -9438
rect -621 -9472 -605 -9438
rect -681 -9488 -605 -9472
rect -681 -10048 -605 -10032
rect -681 -10082 -665 -10048
rect -621 -10082 -605 -10048
rect -681 -10088 -605 -10082
rect -571 -10120 -537 -9400
rect -503 -9438 -427 -9432
rect -503 -9472 -487 -9438
rect -443 -9472 -427 -9438
rect -503 -9488 -427 -9472
rect -503 -10048 -427 -10032
rect -503 -10082 -487 -10048
rect -443 -10082 -427 -10048
rect -503 -10088 -427 -10082
rect -393 -10120 -359 -9400
rect -325 -9438 -249 -9432
rect -325 -9472 -309 -9438
rect -265 -9472 -249 -9438
rect -325 -9488 -249 -9472
rect -303 -9546 -269 -9488
rect -322 -9599 -312 -9546
rect -259 -9599 -249 -9546
rect -324 -9978 -314 -9925
rect -261 -9978 -251 -9925
rect -304 -10032 -270 -9978
rect -325 -10048 -249 -10032
rect -325 -10082 -309 -10048
rect -265 -10082 -249 -10048
rect -325 -10088 -249 -10082
rect -215 -10120 -181 -9400
rect -147 -9438 -71 -9432
rect -147 -9472 -131 -9438
rect -87 -9472 -71 -9438
rect -147 -9488 -71 -9472
rect -126 -9545 -92 -9488
rect -146 -9598 -136 -9545
rect -83 -9598 -73 -9545
rect -146 -9979 -136 -9926
rect -83 -9979 -73 -9926
rect -126 -10032 -92 -9979
rect -147 -10048 -71 -10032
rect -147 -10082 -131 -10048
rect -87 -10082 -71 -10048
rect -147 -10088 -71 -10082
rect -37 -10120 -3 -9400
rect 31 -9438 107 -9432
rect 31 -9472 47 -9438
rect 91 -9472 107 -9438
rect 31 -9488 107 -9472
rect 52 -9546 86 -9488
rect 32 -9599 42 -9546
rect 95 -9599 105 -9546
rect 33 -9978 43 -9925
rect 96 -9978 106 -9925
rect 52 -10032 86 -9978
rect 31 -10048 107 -10032
rect 31 -10082 47 -10048
rect 91 -10082 107 -10048
rect 31 -10088 107 -10082
rect 141 -10120 175 -9400
rect 209 -9438 285 -9432
rect 209 -9472 225 -9438
rect 269 -9472 285 -9438
rect 209 -9488 285 -9472
rect 231 -9545 265 -9488
rect 212 -9598 222 -9545
rect 275 -9598 285 -9545
rect 210 -9978 220 -9925
rect 273 -9978 283 -9925
rect 230 -10032 264 -9978
rect 209 -10048 285 -10032
rect 209 -10082 225 -10048
rect 269 -10082 285 -10048
rect 209 -10088 285 -10082
rect 319 -10120 353 -9400
rect 387 -9438 463 -9432
rect 387 -9472 403 -9438
rect 447 -9472 463 -9438
rect 387 -9488 463 -9472
rect 408 -9546 442 -9488
rect 389 -9599 399 -9546
rect 452 -9599 462 -9546
rect 388 -9978 398 -9925
rect 451 -9978 461 -9925
rect 408 -10032 442 -9978
rect 387 -10048 463 -10032
rect 387 -10082 403 -10048
rect 447 -10082 463 -10048
rect 387 -10088 463 -10082
rect 497 -10120 531 -9400
rect 565 -9438 641 -9432
rect 565 -9472 581 -9438
rect 625 -9472 641 -9438
rect 565 -9488 641 -9472
rect 587 -9546 621 -9488
rect 567 -9599 577 -9546
rect 630 -9599 640 -9546
rect 566 -9978 576 -9925
rect 629 -9978 639 -9925
rect 586 -10032 620 -9978
rect 565 -10048 641 -10032
rect 565 -10082 581 -10048
rect 625 -10082 641 -10048
rect 565 -10088 641 -10082
rect 675 -10120 709 -9400
rect 743 -9438 819 -9432
rect 743 -9472 759 -9438
rect 803 -9472 819 -9438
rect 743 -9488 819 -9472
rect 921 -9438 997 -9432
rect 921 -9472 937 -9438
rect 981 -9472 997 -9438
rect 921 -9488 997 -9472
rect 743 -10048 819 -10032
rect 743 -10082 759 -10048
rect 803 -10082 819 -10048
rect 743 -10088 819 -10082
rect 921 -10048 997 -10032
rect 921 -10082 937 -10048
rect 981 -10082 997 -10048
rect 921 -10088 997 -10082
rect 1031 -10120 1065 -9400
rect 1099 -9438 1175 -9432
rect 1099 -9472 1115 -9438
rect 1159 -9472 1175 -9438
rect 1099 -9488 1175 -9472
rect 1099 -10048 1175 -10032
rect 1099 -10082 1115 -10048
rect 1159 -10082 1175 -10048
rect 1099 -10088 1175 -10082
rect 1209 -10120 1243 -9400
rect 1277 -9438 1353 -9432
rect 1277 -9472 1293 -9438
rect 1337 -9472 1353 -9438
rect 1277 -9488 1353 -9472
rect 1277 -10048 1353 -10032
rect 1277 -10082 1293 -10048
rect 1337 -10082 1353 -10048
rect 1277 -10088 1353 -10082
rect 1387 -10120 1421 -9400
rect 1455 -9438 1531 -9432
rect 1455 -9472 1471 -9438
rect 1515 -9472 1531 -9438
rect 1455 -9488 1531 -9472
rect 1455 -10048 1531 -10032
rect 1455 -10082 1471 -10048
rect 1515 -10082 1531 -10048
rect 1455 -10088 1531 -10082
rect 1565 -10120 1599 -9400
rect 1633 -9438 1709 -9432
rect 1633 -9472 1649 -9438
rect 1693 -9472 1709 -9438
rect 1633 -9488 1709 -9472
rect 1633 -10048 1709 -10032
rect 1633 -10082 1649 -10048
rect 1693 -10082 1709 -10048
rect 1633 -10088 1709 -10082
rect 1743 -10120 1777 -9400
rect 1832 -9432 1866 -9426
rect 1811 -9438 1887 -9432
rect 1811 -9472 1827 -9438
rect 1871 -9472 1887 -9438
rect 1811 -9488 1887 -9472
rect 1832 -10032 1866 -9488
rect 1811 -10048 1887 -10032
rect 1811 -10082 1827 -10048
rect 1871 -10082 1887 -10048
rect 1811 -10088 1887 -10082
rect 1921 -10120 1955 -9400
rect 2010 -9432 2044 -9426
rect 1989 -9438 2065 -9432
rect 1989 -9472 2005 -9438
rect 2049 -9472 2065 -9438
rect 1989 -9488 2065 -9472
rect 2010 -10032 2044 -9488
rect 1989 -10048 2065 -10032
rect 1989 -10082 2005 -10048
rect 2049 -10082 2065 -10048
rect 1989 -10088 2065 -10082
rect 2099 -10120 2133 -9400
rect 2188 -9432 2222 -9426
rect 2167 -9438 2243 -9432
rect 2167 -9472 2183 -9438
rect 2227 -9472 2243 -9438
rect 2167 -9488 2243 -9472
rect 2188 -9547 2222 -9488
rect 2168 -9600 2178 -9547
rect 2231 -9600 2241 -9547
rect 2188 -10032 2222 -9600
rect 2167 -10048 2243 -10032
rect 2167 -10082 2183 -10048
rect 2227 -10082 2243 -10048
rect 2167 -10088 2243 -10082
rect 2277 -10120 2311 -9400
rect 2345 -9438 2421 -9432
rect 2345 -9472 2361 -9438
rect 2405 -9472 2421 -9438
rect 2345 -9488 2421 -9472
rect 2366 -9546 2400 -9488
rect 2347 -9599 2357 -9546
rect 2410 -9599 2420 -9546
rect 2346 -9978 2356 -9925
rect 2409 -9978 2419 -9925
rect 2366 -10032 2400 -9978
rect 2345 -10048 2421 -10032
rect 2345 -10082 2361 -10048
rect 2405 -10082 2421 -10048
rect 2345 -10088 2421 -10082
rect 2455 -10120 2489 -9400
rect 2523 -9438 2599 -9432
rect 2523 -9472 2539 -9438
rect 2583 -9472 2599 -9438
rect 2523 -9488 2599 -9472
rect 2544 -9546 2578 -9488
rect 2524 -9599 2534 -9546
rect 2587 -9599 2597 -9546
rect 2524 -9978 2534 -9925
rect 2587 -9978 2597 -9925
rect 2544 -10032 2578 -9978
rect 2523 -10048 2599 -10032
rect 2523 -10082 2539 -10048
rect 2583 -10082 2599 -10048
rect 2523 -10088 2599 -10082
rect 2633 -10120 2667 -9400
rect 2701 -9438 2777 -9432
rect 2701 -9472 2717 -9438
rect 2761 -9472 2777 -9438
rect 2701 -9488 2777 -9472
rect 2722 -9546 2756 -9488
rect 2703 -9599 2713 -9546
rect 2766 -9599 2776 -9546
rect 2702 -9979 2712 -9926
rect 2765 -9979 2775 -9926
rect 2722 -10032 2756 -9979
rect 2701 -10048 2777 -10032
rect 2701 -10082 2717 -10048
rect 2761 -10082 2777 -10048
rect 2701 -10088 2777 -10082
rect 2811 -10120 2845 -9400
rect 2879 -9438 2955 -9432
rect 2879 -9472 2895 -9438
rect 2939 -9472 2955 -9438
rect 2879 -9488 2955 -9472
rect 2881 -9978 2891 -9925
rect 2944 -9978 2954 -9925
rect 2900 -10032 2934 -9978
rect 2879 -10048 2955 -10032
rect 2879 -10082 2895 -10048
rect 2939 -10082 2955 -10048
rect 2879 -10088 2955 -10082
rect 2989 -10120 3023 -9400
rect 3057 -9438 3133 -9432
rect 3057 -9472 3073 -9438
rect 3117 -9472 3133 -9438
rect 3057 -9488 3133 -9472
rect 3059 -9978 3069 -9925
rect 3122 -9978 3132 -9925
rect 3078 -10032 3112 -9978
rect 3057 -10048 3133 -10032
rect 3057 -10082 3073 -10048
rect 3117 -10082 3133 -10048
rect 3057 -10088 3133 -10082
rect 3167 -10120 3201 -9400
rect 3235 -9438 3311 -9432
rect 3235 -9472 3251 -9438
rect 3295 -9472 3311 -9438
rect 3235 -9488 3311 -9472
rect 3256 -9925 3290 -9488
rect 3236 -9978 3246 -9925
rect 3299 -9978 3309 -9925
rect 3256 -10032 3290 -9978
rect 3235 -10048 3311 -10032
rect 3235 -10082 3251 -10048
rect 3295 -10082 3311 -10048
rect 3235 -10088 3311 -10082
rect 3345 -10120 3379 -9400
rect 3413 -9438 3489 -9432
rect 3413 -9472 3429 -9438
rect 3473 -9472 3489 -9438
rect 3413 -9488 3489 -9472
rect 3413 -10048 3489 -10032
rect 3413 -10082 3429 -10048
rect 3473 -10082 3489 -10048
rect 3413 -10088 3489 -10082
rect 3523 -10120 3557 -9400
rect 3591 -9438 3667 -9432
rect 3591 -9472 3607 -9438
rect 3651 -9472 3667 -9438
rect 3591 -9488 3667 -9472
rect 3591 -10048 3667 -10032
rect 3591 -10082 3607 -10048
rect 3651 -10082 3667 -10048
rect 3591 -10088 3667 -10082
rect 3701 -10120 3735 -9400
rect 3769 -9438 3845 -9432
rect 3769 -9472 3785 -9438
rect 3829 -9472 3845 -9438
rect 3769 -9488 3845 -9472
rect 3879 -9439 3913 -9400
rect 3947 -9438 4023 -9432
rect 3947 -9439 3963 -9438
rect 3879 -9472 3963 -9439
rect 4007 -9439 4023 -9438
rect 4056 -9439 4090 -9400
rect 4007 -9472 4090 -9439
rect 3879 -9473 4090 -9472
rect 3769 -10048 3845 -10032
rect 3769 -10082 3785 -10048
rect 3829 -10082 3845 -10048
rect 3769 -10088 3845 -10082
rect 3879 -10047 3913 -9473
rect 3947 -9488 4023 -9473
rect 4208 -9546 4261 -7976
rect 4771 -9262 4823 -7907
rect 4771 -9314 4824 -9262
rect 4761 -9367 4771 -9314
rect 4824 -9367 4834 -9314
rect 4198 -9599 4208 -9546
rect 4261 -9599 4271 -9546
rect 3947 -10047 4023 -10032
rect 3879 -10048 4092 -10047
rect 3879 -10081 3963 -10048
rect 3879 -10120 3913 -10081
rect 3947 -10082 3963 -10081
rect 4007 -10081 4092 -10048
rect 4007 -10082 4023 -10081
rect 3947 -10088 4023 -10082
rect 4058 -10120 4092 -10081
rect -2179 -10132 -2133 -10120
rect -2179 -10388 -2173 -10132
rect -2139 -10388 -2133 -10132
rect -2179 -10400 -2133 -10388
rect -2001 -10132 -1955 -10120
rect -2001 -10388 -1995 -10132
rect -1961 -10388 -1955 -10132
rect -2001 -10400 -1955 -10388
rect -1823 -10132 -1777 -10120
rect -1823 -10388 -1817 -10132
rect -1783 -10388 -1777 -10132
rect -1823 -10400 -1777 -10388
rect -1645 -10132 -1599 -10120
rect -1645 -10388 -1639 -10132
rect -1605 -10388 -1599 -10132
rect -1645 -10400 -1599 -10388
rect -1467 -10132 -1421 -10120
rect -1467 -10388 -1461 -10132
rect -1427 -10388 -1421 -10132
rect -1467 -10400 -1421 -10388
rect -1289 -10132 -1243 -10120
rect -1289 -10388 -1283 -10132
rect -1249 -10388 -1243 -10132
rect -1289 -10400 -1243 -10388
rect -1111 -10132 -1065 -10120
rect -1111 -10388 -1105 -10132
rect -1071 -10388 -1065 -10132
rect -1111 -10400 -1065 -10388
rect -933 -10132 -887 -10120
rect -933 -10388 -927 -10132
rect -893 -10388 -887 -10132
rect -933 -10400 -887 -10388
rect -755 -10132 -709 -10120
rect -755 -10388 -749 -10132
rect -715 -10388 -709 -10132
rect -755 -10400 -709 -10388
rect -577 -10132 -531 -10120
rect -577 -10388 -571 -10132
rect -537 -10388 -531 -10132
rect -577 -10400 -531 -10388
rect -399 -10132 -353 -10120
rect -399 -10388 -393 -10132
rect -359 -10388 -353 -10132
rect -399 -10400 -353 -10388
rect -221 -10132 -175 -10120
rect -221 -10388 -215 -10132
rect -181 -10388 -175 -10132
rect -221 -10400 -175 -10388
rect -43 -10132 3 -10120
rect -43 -10388 -37 -10132
rect -3 -10388 3 -10132
rect -43 -10400 3 -10388
rect 135 -10132 181 -10120
rect 135 -10388 141 -10132
rect 175 -10388 181 -10132
rect 135 -10400 181 -10388
rect 313 -10132 359 -10120
rect 313 -10388 319 -10132
rect 353 -10388 359 -10132
rect 313 -10400 359 -10388
rect 491 -10132 537 -10120
rect 491 -10388 497 -10132
rect 531 -10388 537 -10132
rect 491 -10400 537 -10388
rect 669 -10132 715 -10120
rect 669 -10388 675 -10132
rect 709 -10388 715 -10132
rect 669 -10400 715 -10388
rect 847 -10132 893 -10120
rect 847 -10388 853 -10132
rect 887 -10388 893 -10132
rect 847 -10400 893 -10388
rect 1025 -10132 1071 -10120
rect 1025 -10388 1031 -10132
rect 1065 -10388 1071 -10132
rect 1025 -10400 1071 -10388
rect 1203 -10132 1249 -10120
rect 1203 -10388 1209 -10132
rect 1243 -10388 1249 -10132
rect 1203 -10400 1249 -10388
rect 1381 -10132 1427 -10120
rect 1381 -10388 1387 -10132
rect 1421 -10388 1427 -10132
rect 1381 -10400 1427 -10388
rect 1559 -10132 1605 -10120
rect 1559 -10388 1565 -10132
rect 1599 -10388 1605 -10132
rect 1559 -10400 1605 -10388
rect 1737 -10132 1783 -10120
rect 1737 -10388 1743 -10132
rect 1777 -10388 1783 -10132
rect 1737 -10400 1783 -10388
rect 1915 -10132 1961 -10120
rect 1915 -10388 1921 -10132
rect 1955 -10388 1961 -10132
rect 1915 -10400 1961 -10388
rect 2093 -10132 2139 -10120
rect 2093 -10388 2099 -10132
rect 2133 -10388 2139 -10132
rect 2093 -10400 2139 -10388
rect 2271 -10132 2317 -10120
rect 2271 -10388 2277 -10132
rect 2311 -10388 2317 -10132
rect 2271 -10400 2317 -10388
rect 2449 -10132 2495 -10120
rect 2449 -10388 2455 -10132
rect 2489 -10388 2495 -10132
rect 2449 -10400 2495 -10388
rect 2627 -10132 2673 -10120
rect 2627 -10388 2633 -10132
rect 2667 -10388 2673 -10132
rect 2627 -10400 2673 -10388
rect 2805 -10132 2851 -10120
rect 2805 -10388 2811 -10132
rect 2845 -10388 2851 -10132
rect 2805 -10400 2851 -10388
rect 2983 -10132 3029 -10120
rect 2983 -10388 2989 -10132
rect 3023 -10388 3029 -10132
rect 2983 -10400 3029 -10388
rect 3161 -10132 3207 -10120
rect 3161 -10388 3167 -10132
rect 3201 -10388 3207 -10132
rect 3161 -10400 3207 -10388
rect 3339 -10132 3385 -10120
rect 3339 -10388 3345 -10132
rect 3379 -10388 3385 -10132
rect 3339 -10400 3385 -10388
rect 3517 -10132 3563 -10120
rect 3517 -10388 3523 -10132
rect 3557 -10388 3563 -10132
rect 3517 -10400 3563 -10388
rect 3695 -10132 3741 -10120
rect 3695 -10388 3701 -10132
rect 3735 -10388 3741 -10132
rect 3695 -10400 3741 -10388
rect 3873 -10132 3919 -10120
rect 3873 -10388 3879 -10132
rect 3913 -10388 3919 -10132
rect 3873 -10400 3919 -10388
rect 4051 -10132 4097 -10120
rect 4051 -10388 4057 -10132
rect 4091 -10388 4097 -10132
rect 4051 -10400 4097 -10388
rect -2105 -10438 -2029 -10432
rect -2105 -10472 -2089 -10438
rect -2045 -10472 -2029 -10438
rect -2105 -10488 -2029 -10472
rect -1927 -10438 -1851 -10432
rect -1927 -10472 -1911 -10438
rect -1867 -10472 -1851 -10438
rect -1927 -10488 -1851 -10472
rect -1749 -10438 -1673 -10432
rect -1749 -10472 -1733 -10438
rect -1689 -10472 -1673 -10438
rect -1749 -10488 -1673 -10472
rect -1571 -10438 -1495 -10432
rect -1571 -10472 -1555 -10438
rect -1511 -10472 -1495 -10438
rect -1571 -10488 -1495 -10472
rect -1393 -10438 -1317 -10432
rect -1393 -10472 -1377 -10438
rect -1333 -10472 -1317 -10438
rect -1393 -10488 -1317 -10472
rect -1215 -10438 -1139 -10432
rect -1215 -10472 -1199 -10438
rect -1155 -10472 -1139 -10438
rect -1215 -10488 -1139 -10472
rect -1037 -10438 -961 -10432
rect -1037 -10472 -1021 -10438
rect -977 -10472 -961 -10438
rect -1037 -10488 -961 -10472
rect -859 -10438 -783 -10432
rect -859 -10472 -843 -10438
rect -799 -10472 -783 -10438
rect -859 -10488 -783 -10472
rect -681 -10438 -605 -10432
rect -681 -10472 -665 -10438
rect -621 -10472 -605 -10438
rect -681 -10488 -605 -10472
rect -503 -10438 -427 -10432
rect -503 -10472 -487 -10438
rect -443 -10472 -427 -10438
rect -503 -10488 -427 -10472
rect -325 -10438 -249 -10432
rect -325 -10472 -309 -10438
rect -265 -10472 -249 -10438
rect -325 -10488 -249 -10472
rect -147 -10438 -71 -10432
rect -147 -10472 -131 -10438
rect -87 -10472 -71 -10438
rect -147 -10488 -71 -10472
rect 31 -10438 107 -10432
rect 31 -10472 47 -10438
rect 91 -10472 107 -10438
rect 31 -10488 107 -10472
rect 209 -10438 285 -10432
rect 209 -10472 225 -10438
rect 269 -10472 285 -10438
rect 209 -10488 285 -10472
rect 387 -10438 463 -10432
rect 387 -10472 403 -10438
rect 447 -10472 463 -10438
rect 387 -10488 463 -10472
rect 565 -10438 641 -10432
rect 565 -10472 581 -10438
rect 625 -10472 641 -10438
rect 565 -10488 641 -10472
rect 743 -10438 819 -10432
rect 853 -10438 887 -10400
rect 941 -10432 975 -10431
rect 921 -10438 997 -10432
rect 1031 -10438 1065 -10400
rect 1653 -10432 1687 -10431
rect 1099 -10438 1175 -10432
rect 743 -10472 759 -10438
rect 803 -10472 937 -10438
rect 981 -10472 1115 -10438
rect 1159 -10472 1175 -10438
rect 743 -10488 819 -10472
rect 921 -10488 997 -10472
rect 1099 -10488 1175 -10472
rect 1277 -10438 1353 -10432
rect 1277 -10472 1293 -10438
rect 1337 -10472 1353 -10438
rect 1277 -10488 1353 -10472
rect 1455 -10438 1531 -10432
rect 1455 -10472 1471 -10438
rect 1515 -10472 1531 -10438
rect 1455 -10488 1531 -10472
rect 1633 -10438 1709 -10432
rect 1633 -10472 1649 -10438
rect 1693 -10472 1709 -10438
rect 1633 -10488 1709 -10472
rect 1811 -10438 1887 -10432
rect 1811 -10472 1827 -10438
rect 1871 -10472 1887 -10438
rect 1811 -10488 1887 -10472
rect 1989 -10438 2065 -10432
rect 1989 -10472 2005 -10438
rect 2049 -10472 2065 -10438
rect 1989 -10488 2065 -10472
rect 2167 -10438 2243 -10432
rect 2167 -10472 2183 -10438
rect 2227 -10472 2243 -10438
rect 2167 -10488 2243 -10472
rect 2345 -10438 2421 -10432
rect 2345 -10472 2361 -10438
rect 2405 -10472 2421 -10438
rect 2345 -10488 2421 -10472
rect 2523 -10438 2599 -10432
rect 2523 -10472 2539 -10438
rect 2583 -10472 2599 -10438
rect 2523 -10488 2599 -10472
rect 2701 -10438 2777 -10432
rect 2701 -10472 2717 -10438
rect 2761 -10472 2777 -10438
rect 2701 -10488 2777 -10472
rect 2879 -10438 2955 -10432
rect 2879 -10472 2895 -10438
rect 2939 -10472 2955 -10438
rect 2879 -10488 2955 -10472
rect 3057 -10438 3133 -10432
rect 3057 -10472 3073 -10438
rect 3117 -10472 3133 -10438
rect 3057 -10488 3133 -10472
rect 3235 -10438 3311 -10432
rect 3235 -10472 3251 -10438
rect 3295 -10472 3311 -10438
rect 3235 -10488 3311 -10472
rect 3413 -10438 3489 -10432
rect 3413 -10472 3429 -10438
rect 3473 -10472 3489 -10438
rect 3413 -10488 3489 -10472
rect 3591 -10438 3667 -10432
rect 3591 -10472 3607 -10438
rect 3651 -10472 3667 -10438
rect 3591 -10488 3667 -10472
rect 3769 -10438 3845 -10432
rect 3769 -10472 3785 -10438
rect 3829 -10472 3845 -10438
rect 3769 -10488 3845 -10472
rect 3947 -10438 4023 -10432
rect 3947 -10472 3963 -10438
rect 4007 -10472 4023 -10438
rect 3947 -10488 4023 -10472
rect -1837 -10961 -1827 -10908
rect -1774 -10961 -1764 -10908
rect -1480 -10961 -1470 -10908
rect -1417 -10961 -1407 -10908
rect -2105 -11048 -2029 -11032
rect -2105 -11082 -2089 -11048
rect -2045 -11082 -2029 -11048
rect -2105 -11088 -2029 -11082
rect -1927 -11048 -1851 -11032
rect -1927 -11082 -1911 -11048
rect -1867 -11082 -1851 -11048
rect -1927 -11088 -1851 -11082
rect -1818 -11120 -1784 -10961
rect -1749 -11048 -1673 -11032
rect -1749 -11082 -1733 -11048
rect -1689 -11082 -1673 -11048
rect -1749 -11088 -1673 -11082
rect -1571 -11048 -1495 -11032
rect -1571 -11082 -1555 -11048
rect -1511 -11082 -1495 -11048
rect -1571 -11088 -1495 -11082
rect -1461 -11120 -1427 -10961
rect -1372 -11032 -1338 -10488
rect -1193 -11032 -1159 -10488
rect -1124 -10961 -1114 -10908
rect -1061 -10961 -1051 -10908
rect -1393 -11048 -1317 -11032
rect -1393 -11082 -1377 -11048
rect -1333 -11082 -1317 -11048
rect -1393 -11088 -1317 -11082
rect -1215 -11048 -1139 -11032
rect -1215 -11082 -1199 -11048
rect -1155 -11082 -1139 -11048
rect -1215 -11088 -1139 -11082
rect -1105 -11120 -1071 -10961
rect -1016 -11032 -982 -10488
rect -838 -11032 -804 -10488
rect -768 -10961 -758 -10908
rect -705 -10961 -695 -10908
rect -1037 -11048 -961 -11032
rect -1037 -11082 -1021 -11048
rect -977 -11082 -961 -11048
rect -1037 -11088 -961 -11082
rect -859 -11048 -783 -11032
rect -859 -11082 -843 -11048
rect -799 -11082 -783 -11048
rect -859 -11088 -783 -11082
rect -749 -11120 -715 -10961
rect -659 -11032 -625 -10488
rect -482 -11032 -448 -10488
rect 941 -10908 975 -10488
rect -412 -10961 -402 -10908
rect -349 -10961 -339 -10908
rect -56 -10961 -46 -10908
rect 7 -10961 17 -10908
rect 299 -10961 309 -10908
rect 362 -10961 372 -10908
rect 655 -10961 665 -10908
rect 718 -10961 728 -10908
rect 921 -10961 931 -10908
rect 984 -10961 994 -10908
rect 1189 -10961 1199 -10908
rect 1252 -10961 1262 -10908
rect -681 -11048 -605 -11032
rect -681 -11082 -665 -11048
rect -621 -11082 -605 -11048
rect -681 -11088 -605 -11082
rect -503 -11048 -427 -11032
rect -503 -11082 -487 -11048
rect -443 -11082 -427 -11048
rect -503 -11088 -427 -11082
rect -393 -11120 -359 -10961
rect -325 -11048 -249 -11032
rect -325 -11082 -309 -11048
rect -265 -11082 -249 -11048
rect -325 -11088 -249 -11082
rect -147 -11048 -71 -11032
rect -147 -11082 -131 -11048
rect -87 -11082 -71 -11048
rect -147 -11088 -71 -11082
rect -36 -11120 -2 -10961
rect 31 -11048 107 -11032
rect 31 -11082 47 -11048
rect 91 -11082 107 -11048
rect 31 -11088 107 -11082
rect 209 -11048 285 -11032
rect 209 -11082 225 -11048
rect 269 -11082 285 -11048
rect 209 -11088 285 -11082
rect 319 -11120 353 -10961
rect 387 -11048 463 -11032
rect 387 -11082 403 -11048
rect 447 -11082 463 -11048
rect 387 -11088 463 -11082
rect 565 -11048 641 -11032
rect 565 -11082 581 -11048
rect 625 -11082 641 -11048
rect 565 -11088 641 -11082
rect 675 -11120 709 -10961
rect 941 -11032 975 -10961
rect 743 -11048 819 -11032
rect 743 -11082 759 -11048
rect 803 -11082 819 -11048
rect 743 -11088 819 -11082
rect 921 -11048 997 -11032
rect 921 -11082 937 -11048
rect 981 -11082 997 -11048
rect 921 -11088 997 -11082
rect 1099 -11048 1175 -11032
rect 1099 -11082 1115 -11048
rect 1159 -11082 1175 -11048
rect 1099 -11088 1175 -11082
rect 1209 -11120 1243 -10961
rect 1299 -11032 1333 -10488
rect 1477 -11032 1511 -10488
rect 1546 -10961 1556 -10908
rect 1609 -10961 1619 -10908
rect 1277 -11048 1353 -11032
rect 1277 -11082 1293 -11048
rect 1337 -11082 1353 -11048
rect 1277 -11088 1353 -11082
rect 1455 -11048 1531 -11032
rect 1455 -11082 1471 -11048
rect 1515 -11082 1531 -11048
rect 1455 -11088 1531 -11082
rect 1566 -11120 1600 -10961
rect 1653 -11032 1687 -10488
rect 1832 -11032 1866 -10488
rect 1903 -10961 1913 -10908
rect 1966 -10961 1976 -10908
rect 1633 -11048 1709 -11032
rect 1633 -11082 1649 -11048
rect 1693 -11082 1709 -11048
rect 1633 -11088 1709 -11082
rect 1811 -11048 1887 -11032
rect 1811 -11082 1827 -11048
rect 1871 -11082 1887 -11048
rect 1811 -11088 1887 -11082
rect 1922 -11120 1956 -10961
rect 2010 -11032 2044 -10488
rect 2188 -11032 2222 -10488
rect 2258 -10961 2268 -10908
rect 2321 -10961 2331 -10908
rect 2613 -10961 2623 -10908
rect 2676 -10961 2686 -10908
rect 2970 -10961 2980 -10908
rect 3033 -10961 3043 -10908
rect 3325 -10961 3335 -10908
rect 3388 -10961 3398 -10908
rect 1989 -11048 2065 -11032
rect 1989 -11082 2005 -11048
rect 2049 -11082 2065 -11048
rect 1989 -11088 2065 -11082
rect 2167 -11048 2243 -11032
rect 2167 -11082 2183 -11048
rect 2227 -11082 2243 -11048
rect 2167 -11088 2243 -11082
rect 2277 -11120 2311 -10961
rect 2345 -11048 2421 -11032
rect 2345 -11082 2361 -11048
rect 2405 -11082 2421 -11048
rect 2345 -11088 2421 -11082
rect 2523 -11048 2599 -11032
rect 2523 -11082 2539 -11048
rect 2583 -11082 2599 -11048
rect 2523 -11088 2599 -11082
rect 2633 -11120 2667 -10961
rect 2701 -11048 2777 -11032
rect 2701 -11082 2717 -11048
rect 2761 -11082 2777 -11048
rect 2701 -11088 2777 -11082
rect 2879 -11048 2955 -11032
rect 2879 -11082 2895 -11048
rect 2939 -11082 2955 -11048
rect 2879 -11088 2955 -11082
rect 2989 -11120 3023 -10961
rect 3057 -11048 3133 -11032
rect 3057 -11082 3073 -11048
rect 3117 -11082 3133 -11048
rect 3057 -11088 3133 -11082
rect 3235 -11048 3311 -11032
rect 3235 -11082 3251 -11048
rect 3295 -11082 3311 -11048
rect 3235 -11088 3311 -11082
rect 3345 -11120 3379 -10961
rect 3434 -11032 3468 -10488
rect 3613 -11032 3647 -10488
rect 3682 -10961 3692 -10908
rect 3745 -10961 3755 -10908
rect 3413 -11048 3489 -11032
rect 3413 -11082 3429 -11048
rect 3473 -11082 3489 -11048
rect 3413 -11088 3489 -11082
rect 3591 -11048 3667 -11032
rect 3591 -11082 3607 -11048
rect 3651 -11082 3667 -11048
rect 3591 -11088 3667 -11082
rect 3701 -11120 3735 -10961
rect 3791 -11032 3825 -10488
rect 3769 -11048 3845 -11032
rect 3769 -11082 3785 -11048
rect 3829 -11082 3845 -11048
rect 3769 -11088 3845 -11082
rect 3947 -11048 4023 -11032
rect 3947 -11082 3963 -11048
rect 4007 -11082 4023 -11048
rect 3947 -11088 4023 -11082
rect -2179 -11132 -2133 -11120
rect -2179 -11388 -2173 -11132
rect -2139 -11388 -2133 -11132
rect -2179 -11400 -2133 -11388
rect -2001 -11132 -1955 -11120
rect -2001 -11388 -1995 -11132
rect -1961 -11388 -1955 -11132
rect -2001 -11400 -1955 -11388
rect -1823 -11132 -1777 -11120
rect -1823 -11388 -1817 -11132
rect -1783 -11388 -1777 -11132
rect -1823 -11400 -1777 -11388
rect -1645 -11132 -1599 -11120
rect -1645 -11388 -1639 -11132
rect -1605 -11388 -1599 -11132
rect -1645 -11400 -1599 -11388
rect -1467 -11132 -1421 -11120
rect -1467 -11388 -1461 -11132
rect -1427 -11388 -1421 -11132
rect -1467 -11400 -1421 -11388
rect -1289 -11132 -1243 -11120
rect -1289 -11388 -1283 -11132
rect -1249 -11388 -1243 -11132
rect -1289 -11400 -1243 -11388
rect -1111 -11132 -1065 -11120
rect -1111 -11388 -1105 -11132
rect -1071 -11388 -1065 -11132
rect -1111 -11400 -1065 -11388
rect -933 -11132 -887 -11120
rect -933 -11388 -927 -11132
rect -893 -11388 -887 -11132
rect -933 -11400 -887 -11388
rect -755 -11132 -709 -11120
rect -755 -11388 -749 -11132
rect -715 -11388 -709 -11132
rect -755 -11400 -709 -11388
rect -577 -11132 -531 -11120
rect -577 -11388 -571 -11132
rect -537 -11388 -531 -11132
rect -577 -11400 -531 -11388
rect -399 -11132 -353 -11120
rect -399 -11388 -393 -11132
rect -359 -11388 -353 -11132
rect -399 -11400 -353 -11388
rect -221 -11132 -175 -11120
rect -221 -11388 -215 -11132
rect -181 -11388 -175 -11132
rect -221 -11400 -175 -11388
rect -43 -11132 3 -11120
rect -43 -11388 -37 -11132
rect -3 -11388 3 -11132
rect -43 -11400 3 -11388
rect 135 -11132 181 -11120
rect 135 -11388 141 -11132
rect 175 -11388 181 -11132
rect 135 -11400 181 -11388
rect 313 -11132 359 -11120
rect 313 -11388 319 -11132
rect 353 -11388 359 -11132
rect 313 -11400 359 -11388
rect 491 -11132 537 -11120
rect 491 -11388 497 -11132
rect 531 -11388 537 -11132
rect 491 -11400 537 -11388
rect 669 -11132 715 -11120
rect 669 -11388 675 -11132
rect 709 -11388 715 -11132
rect 669 -11400 715 -11388
rect 847 -11132 893 -11120
rect 847 -11388 853 -11132
rect 887 -11388 893 -11132
rect 847 -11400 893 -11388
rect 1025 -11132 1071 -11120
rect 1025 -11388 1031 -11132
rect 1065 -11388 1071 -11132
rect 1025 -11400 1071 -11388
rect 1203 -11132 1249 -11120
rect 1203 -11388 1209 -11132
rect 1243 -11388 1249 -11132
rect 1203 -11400 1249 -11388
rect 1381 -11132 1427 -11120
rect 1381 -11388 1387 -11132
rect 1421 -11388 1427 -11132
rect 1381 -11400 1427 -11388
rect 1559 -11132 1605 -11120
rect 1559 -11388 1565 -11132
rect 1599 -11388 1605 -11132
rect 1559 -11400 1605 -11388
rect 1737 -11132 1783 -11120
rect 1737 -11388 1743 -11132
rect 1777 -11388 1783 -11132
rect 1737 -11400 1783 -11388
rect 1915 -11132 1961 -11120
rect 1915 -11388 1921 -11132
rect 1955 -11388 1961 -11132
rect 1915 -11400 1961 -11388
rect 2093 -11132 2139 -11120
rect 2093 -11388 2099 -11132
rect 2133 -11388 2139 -11132
rect 2093 -11400 2139 -11388
rect 2271 -11132 2317 -11120
rect 2271 -11388 2277 -11132
rect 2311 -11388 2317 -11132
rect 2271 -11400 2317 -11388
rect 2449 -11132 2495 -11120
rect 2449 -11388 2455 -11132
rect 2489 -11388 2495 -11132
rect 2449 -11400 2495 -11388
rect 2627 -11132 2673 -11120
rect 2627 -11388 2633 -11132
rect 2667 -11388 2673 -11132
rect 2627 -11400 2673 -11388
rect 2805 -11132 2851 -11120
rect 2805 -11388 2811 -11132
rect 2845 -11388 2851 -11132
rect 2805 -11400 2851 -11388
rect 2983 -11132 3029 -11120
rect 2983 -11388 2989 -11132
rect 3023 -11388 3029 -11132
rect 2983 -11400 3029 -11388
rect 3161 -11132 3207 -11120
rect 3161 -11388 3167 -11132
rect 3201 -11388 3207 -11132
rect 3161 -11400 3207 -11388
rect 3339 -11132 3385 -11120
rect 3339 -11388 3345 -11132
rect 3379 -11388 3385 -11132
rect 3339 -11400 3385 -11388
rect 3517 -11132 3563 -11120
rect 3517 -11388 3523 -11132
rect 3557 -11388 3563 -11132
rect 3517 -11400 3563 -11388
rect 3695 -11132 3741 -11120
rect 3695 -11388 3701 -11132
rect 3735 -11388 3741 -11132
rect 3695 -11400 3741 -11388
rect 3873 -11132 3919 -11120
rect 3873 -11388 3879 -11132
rect 3913 -11388 3919 -11132
rect 3873 -11400 3919 -11388
rect 4051 -11132 4097 -11120
rect 4051 -11388 4057 -11132
rect 4091 -11388 4097 -11132
rect 4051 -11400 4097 -11388
rect -2172 -11439 -2138 -11400
rect -2105 -11438 -2029 -11432
rect -2105 -11439 -2089 -11438
rect -2172 -11472 -2089 -11439
rect -2045 -11439 -2029 -11438
rect -1995 -11439 -1961 -11400
rect -2045 -11472 -1961 -11439
rect -2172 -11473 -1961 -11472
rect -2105 -11488 -2029 -11473
rect -1995 -11637 -1961 -11473
rect -1927 -11438 -1851 -11432
rect -1927 -11472 -1911 -11438
rect -1867 -11472 -1851 -11438
rect -1927 -11488 -1851 -11472
rect -2014 -11690 -2004 -11637
rect -1951 -11690 -1941 -11637
rect -2105 -12047 -2029 -12032
rect -1995 -12047 -1961 -11690
rect -1905 -11919 -1871 -11488
rect -1925 -11972 -1915 -11919
rect -1862 -11972 -1852 -11919
rect -1905 -12032 -1871 -11972
rect -2176 -12048 -1961 -12047
rect -2176 -12081 -2089 -12048
rect -2176 -12120 -2142 -12081
rect -2105 -12082 -2089 -12081
rect -2045 -12081 -1961 -12048
rect -2045 -12082 -2029 -12081
rect -2105 -12088 -2029 -12082
rect -1995 -12120 -1961 -12081
rect -1927 -12048 -1851 -12032
rect -1927 -12082 -1911 -12048
rect -1867 -12082 -1851 -12048
rect -1927 -12088 -1851 -12082
rect -1818 -12120 -1784 -11400
rect -1749 -11438 -1673 -11432
rect -1749 -11472 -1733 -11438
rect -1689 -11472 -1673 -11438
rect -1749 -11488 -1673 -11472
rect -1728 -11919 -1694 -11488
rect -1639 -11528 -1605 -11400
rect -1571 -11438 -1495 -11432
rect -1571 -11472 -1555 -11438
rect -1511 -11472 -1495 -11438
rect -1571 -11488 -1495 -11472
rect -1659 -11581 -1649 -11528
rect -1596 -11581 -1586 -11528
rect -1549 -11919 -1515 -11488
rect -1748 -11972 -1738 -11919
rect -1685 -11972 -1675 -11919
rect -1569 -11972 -1559 -11919
rect -1506 -11972 -1496 -11919
rect -1728 -12032 -1694 -11972
rect -1549 -12032 -1515 -11972
rect -1749 -12048 -1673 -12032
rect -1749 -12082 -1733 -12048
rect -1689 -12082 -1673 -12048
rect -1749 -12088 -1673 -12082
rect -1571 -12048 -1495 -12032
rect -1571 -12082 -1555 -12048
rect -1511 -12082 -1495 -12048
rect -1571 -12088 -1495 -12082
rect -1461 -12120 -1427 -11400
rect -1393 -11438 -1317 -11432
rect -1393 -11472 -1377 -11438
rect -1333 -11472 -1317 -11438
rect -1393 -11488 -1317 -11472
rect -1372 -11919 -1338 -11488
rect -1283 -11526 -1249 -11400
rect -1215 -11438 -1139 -11432
rect -1215 -11472 -1199 -11438
rect -1155 -11472 -1139 -11438
rect -1215 -11488 -1139 -11472
rect -1284 -11528 -1249 -11526
rect -1303 -11581 -1293 -11528
rect -1240 -11581 -1230 -11528
rect -1391 -11972 -1381 -11919
rect -1328 -11972 -1318 -11919
rect -1372 -12032 -1338 -11972
rect -1393 -12048 -1317 -12032
rect -1393 -12082 -1377 -12048
rect -1333 -12082 -1317 -12048
rect -1393 -12088 -1317 -12082
rect -1284 -12120 -1250 -11581
rect -1194 -11919 -1160 -11488
rect -1213 -11972 -1203 -11919
rect -1150 -11972 -1140 -11919
rect -1194 -12032 -1160 -11972
rect -1215 -12048 -1139 -12032
rect -1215 -12082 -1199 -12048
rect -1155 -12082 -1139 -12048
rect -1215 -12088 -1139 -12082
rect -1105 -12120 -1071 -11400
rect -1037 -11438 -961 -11432
rect -1037 -11472 -1021 -11438
rect -977 -11472 -961 -11438
rect -1037 -11488 -961 -11472
rect -1016 -11919 -982 -11488
rect -927 -11528 -893 -11400
rect -859 -11438 -783 -11432
rect -859 -11472 -843 -11438
rect -799 -11472 -783 -11438
rect -859 -11488 -783 -11472
rect -947 -11581 -937 -11528
rect -884 -11581 -874 -11528
rect -838 -11919 -804 -11488
rect -1035 -11972 -1025 -11919
rect -972 -11972 -962 -11919
rect -858 -11972 -848 -11919
rect -795 -11972 -785 -11919
rect -1016 -12032 -982 -11972
rect -838 -12032 -804 -11972
rect -1037 -12048 -961 -12032
rect -1037 -12082 -1021 -12048
rect -977 -12082 -961 -12048
rect -1037 -12088 -961 -12082
rect -859 -12048 -783 -12032
rect -859 -12082 -843 -12048
rect -799 -12082 -783 -12048
rect -859 -12088 -783 -12082
rect -749 -12120 -715 -11400
rect -681 -11438 -605 -11432
rect -681 -11472 -665 -11438
rect -621 -11472 -605 -11438
rect -681 -11488 -605 -11472
rect -660 -11919 -626 -11488
rect -571 -11637 -537 -11400
rect -503 -11438 -427 -11432
rect -503 -11472 -487 -11438
rect -443 -11472 -427 -11438
rect -503 -11488 -427 -11472
rect -590 -11690 -580 -11637
rect -527 -11690 -517 -11637
rect -482 -11919 -448 -11488
rect -680 -11972 -670 -11919
rect -617 -11972 -607 -11919
rect -502 -11972 -492 -11919
rect -439 -11972 -429 -11919
rect -660 -12032 -626 -11972
rect -482 -12032 -448 -11972
rect -681 -12048 -605 -12032
rect -681 -12082 -665 -12048
rect -621 -12082 -605 -12048
rect -681 -12088 -605 -12082
rect -503 -12048 -427 -12032
rect -503 -12082 -487 -12048
rect -443 -12082 -427 -12048
rect -503 -12088 -427 -12082
rect -393 -12120 -359 -11400
rect -325 -11438 -249 -11432
rect -325 -11472 -309 -11438
rect -265 -11472 -249 -11438
rect -325 -11488 -249 -11472
rect -304 -11919 -270 -11488
rect -215 -11757 -181 -11400
rect -147 -11438 -71 -11432
rect -147 -11472 -131 -11438
rect -87 -11472 -71 -11438
rect -147 -11488 -71 -11472
rect -234 -11810 -224 -11757
rect -171 -11810 -161 -11757
rect -324 -11972 -314 -11919
rect -261 -11972 -251 -11919
rect -304 -12032 -270 -11972
rect -325 -12048 -249 -12032
rect -325 -12082 -309 -12048
rect -265 -12082 -249 -12048
rect -325 -12088 -249 -12082
rect -215 -12120 -181 -11810
rect -126 -11919 -92 -11488
rect -146 -11972 -136 -11919
rect -83 -11972 -73 -11919
rect -126 -12032 -92 -11972
rect -147 -12048 -71 -12032
rect -147 -12082 -131 -12048
rect -87 -12082 -71 -12048
rect -147 -12088 -71 -12082
rect -36 -12120 -2 -11400
rect 31 -11438 107 -11432
rect 31 -11472 47 -11438
rect 91 -11472 107 -11438
rect 31 -11488 107 -11472
rect 52 -11919 86 -11488
rect 141 -11757 175 -11400
rect 209 -11438 285 -11432
rect 209 -11472 225 -11438
rect 269 -11472 285 -11438
rect 209 -11488 285 -11472
rect 121 -11810 131 -11757
rect 184 -11810 194 -11757
rect 141 -11811 175 -11810
rect 230 -11919 264 -11488
rect 32 -11972 42 -11919
rect 95 -11972 105 -11919
rect 210 -11972 220 -11919
rect 273 -11972 283 -11919
rect 52 -12032 86 -11972
rect 230 -12032 264 -11972
rect 31 -12048 107 -12032
rect 31 -12082 47 -12048
rect 91 -12082 107 -12048
rect 31 -12088 107 -12082
rect 209 -12048 285 -12032
rect 209 -12082 225 -12048
rect 269 -12082 285 -12048
rect 209 -12088 285 -12082
rect 319 -12120 353 -11400
rect 387 -11438 463 -11432
rect 387 -11472 403 -11438
rect 447 -11472 463 -11438
rect 387 -11488 463 -11472
rect 408 -11919 442 -11488
rect 497 -11757 531 -11400
rect 565 -11438 641 -11432
rect 565 -11472 581 -11438
rect 625 -11472 641 -11438
rect 565 -11488 641 -11472
rect 477 -11810 487 -11757
rect 540 -11810 550 -11757
rect 389 -11972 399 -11919
rect 452 -11972 462 -11919
rect 408 -12032 442 -11972
rect 387 -12048 463 -12032
rect 387 -12082 403 -12048
rect 447 -12082 463 -12048
rect 387 -12088 463 -12082
rect 496 -12120 530 -11810
rect 586 -11919 620 -11488
rect 567 -11972 577 -11919
rect 630 -11972 640 -11919
rect 586 -12032 620 -11972
rect 565 -12048 641 -12032
rect 565 -12082 581 -12048
rect 625 -12082 641 -12048
rect 565 -12088 641 -12082
rect 675 -12120 709 -11400
rect 743 -11438 819 -11432
rect 853 -11438 887 -11400
rect 921 -11438 997 -11432
rect 1031 -11438 1065 -11400
rect 1099 -11438 1175 -11432
rect 743 -11472 759 -11438
rect 803 -11472 937 -11438
rect 981 -11472 1115 -11438
rect 1159 -11472 1175 -11438
rect 743 -11488 819 -11472
rect 921 -11488 997 -11472
rect 1099 -11488 1175 -11472
rect 942 -12032 976 -11488
rect 743 -12048 819 -12032
rect 743 -12082 759 -12048
rect 803 -12082 819 -12048
rect 743 -12088 819 -12082
rect 921 -12048 997 -12032
rect 921 -12082 937 -12048
rect 981 -12082 997 -12048
rect 921 -12088 997 -12082
rect 1099 -12048 1175 -12032
rect 1099 -12082 1115 -12048
rect 1159 -12082 1175 -12048
rect 1099 -12088 1175 -12082
rect 1209 -12120 1243 -11400
rect 1277 -11438 1353 -11432
rect 1277 -11472 1293 -11438
rect 1337 -11472 1353 -11438
rect 1277 -11488 1353 -11472
rect 1298 -11919 1332 -11488
rect 1387 -11528 1421 -11400
rect 1455 -11438 1531 -11432
rect 1455 -11472 1471 -11438
rect 1515 -11472 1531 -11438
rect 1455 -11488 1531 -11472
rect 1367 -11581 1377 -11528
rect 1430 -11581 1440 -11528
rect 1477 -11919 1511 -11488
rect 1278 -11972 1288 -11919
rect 1341 -11972 1351 -11919
rect 1458 -11972 1468 -11919
rect 1521 -11972 1531 -11919
rect 1298 -12032 1332 -11972
rect 1477 -12032 1511 -11972
rect 1277 -12048 1353 -12032
rect 1277 -12082 1293 -12048
rect 1337 -12082 1353 -12048
rect 1277 -12088 1353 -12082
rect 1455 -12048 1531 -12032
rect 1455 -12082 1471 -12048
rect 1515 -12082 1531 -12048
rect 1455 -12088 1531 -12082
rect 1566 -12120 1600 -11400
rect 1633 -11438 1709 -11432
rect 1633 -11472 1649 -11438
rect 1693 -11472 1709 -11438
rect 1633 -11488 1709 -11472
rect 1654 -11920 1688 -11488
rect 1743 -11528 1777 -11400
rect 1811 -11438 1887 -11432
rect 1811 -11472 1827 -11438
rect 1871 -11472 1887 -11438
rect 1811 -11488 1887 -11472
rect 1723 -11581 1733 -11528
rect 1786 -11581 1796 -11528
rect 1634 -11973 1644 -11920
rect 1697 -11973 1707 -11920
rect 1654 -12032 1688 -11973
rect 1633 -12048 1709 -12032
rect 1633 -12082 1649 -12048
rect 1693 -12082 1709 -12048
rect 1633 -12088 1709 -12082
rect 1744 -12120 1778 -11581
rect 1832 -11919 1866 -11488
rect 1813 -11972 1823 -11919
rect 1876 -11972 1886 -11919
rect 1832 -12032 1866 -11972
rect 1811 -12048 1887 -12032
rect 1811 -12082 1827 -12048
rect 1871 -12082 1887 -12048
rect 1811 -12088 1887 -12082
rect 1922 -12120 1956 -11400
rect 1989 -11438 2065 -11432
rect 1989 -11472 2005 -11438
rect 2049 -11472 2065 -11438
rect 1989 -11488 2065 -11472
rect 2010 -11919 2044 -11488
rect 2099 -11528 2133 -11400
rect 2167 -11438 2243 -11432
rect 2167 -11472 2183 -11438
rect 2227 -11472 2243 -11438
rect 2167 -11488 2243 -11472
rect 2079 -11581 2089 -11528
rect 2142 -11581 2152 -11528
rect 2188 -11919 2222 -11488
rect 1990 -11972 2000 -11919
rect 2053 -11972 2063 -11919
rect 2168 -11972 2178 -11919
rect 2231 -11972 2241 -11919
rect 2010 -12032 2044 -11972
rect 2188 -12032 2222 -11972
rect 1989 -12048 2065 -12032
rect 1989 -12082 2005 -12048
rect 2049 -12082 2065 -12048
rect 1989 -12088 2065 -12082
rect 2167 -12048 2243 -12032
rect 2167 -12082 2183 -12048
rect 2227 -12082 2243 -12048
rect 2167 -12088 2243 -12082
rect 2277 -12120 2311 -11400
rect 2345 -11438 2421 -11432
rect 2345 -11472 2361 -11438
rect 2405 -11472 2421 -11438
rect 2345 -11488 2421 -11472
rect 2366 -11919 2400 -11488
rect 2456 -11637 2490 -11400
rect 2523 -11438 2599 -11432
rect 2523 -11472 2539 -11438
rect 2583 -11472 2599 -11438
rect 2523 -11488 2599 -11472
rect 2436 -11690 2446 -11637
rect 2499 -11690 2509 -11637
rect 2544 -11919 2578 -11488
rect 2347 -11972 2357 -11919
rect 2410 -11972 2420 -11919
rect 2524 -11972 2534 -11919
rect 2587 -11972 2597 -11919
rect 2366 -12032 2400 -11972
rect 2544 -12032 2578 -11972
rect 2345 -12048 2421 -12032
rect 2345 -12082 2361 -12048
rect 2405 -12082 2421 -12048
rect 2345 -12088 2421 -12082
rect 2523 -12048 2599 -12032
rect 2523 -12082 2539 -12048
rect 2583 -12082 2599 -12048
rect 2523 -12088 2599 -12082
rect 2633 -12120 2667 -11400
rect 2701 -11438 2777 -11432
rect 2701 -11472 2717 -11438
rect 2761 -11472 2777 -11438
rect 2701 -11488 2777 -11472
rect 2722 -11919 2756 -11488
rect 2810 -11757 2844 -11400
rect 2879 -11438 2955 -11432
rect 2879 -11472 2895 -11438
rect 2939 -11472 2955 -11438
rect 2879 -11488 2955 -11472
rect 2790 -11810 2800 -11757
rect 2853 -11810 2863 -11757
rect 2703 -11972 2713 -11919
rect 2766 -11972 2776 -11919
rect 2722 -12032 2756 -11972
rect 2701 -12048 2777 -12032
rect 2701 -12082 2717 -12048
rect 2761 -12082 2777 -12048
rect 2701 -12088 2777 -12082
rect 2811 -12120 2845 -11810
rect 2900 -11919 2934 -11488
rect 2880 -11972 2890 -11919
rect 2943 -11972 2953 -11919
rect 2900 -12032 2934 -11972
rect 2879 -12048 2955 -12032
rect 2879 -12082 2895 -12048
rect 2939 -12082 2955 -12048
rect 2879 -12088 2955 -12082
rect 2989 -12120 3023 -11400
rect 3057 -11438 3133 -11432
rect 3057 -11472 3073 -11438
rect 3117 -11472 3133 -11438
rect 3057 -11488 3133 -11472
rect 3078 -11919 3112 -11488
rect 3166 -11757 3200 -11400
rect 3235 -11438 3311 -11432
rect 3235 -11472 3251 -11438
rect 3295 -11472 3311 -11438
rect 3235 -11488 3311 -11472
rect 3147 -11810 3157 -11757
rect 3210 -11810 3220 -11757
rect 3256 -11919 3290 -11488
rect 3058 -11972 3068 -11919
rect 3121 -11972 3131 -11919
rect 3237 -11972 3247 -11919
rect 3300 -11972 3310 -11919
rect 3078 -12032 3112 -11972
rect 3256 -12032 3290 -11972
rect 3057 -12048 3133 -12032
rect 3057 -12082 3073 -12048
rect 3117 -12082 3133 -12048
rect 3057 -12088 3133 -12082
rect 3235 -12048 3311 -12032
rect 3235 -12082 3251 -12048
rect 3295 -12082 3311 -12048
rect 3235 -12088 3311 -12082
rect 3345 -12120 3379 -11400
rect 3413 -11438 3489 -11432
rect 3413 -11472 3429 -11438
rect 3473 -11472 3489 -11438
rect 3413 -11488 3489 -11472
rect 3434 -11919 3468 -11488
rect 3522 -11757 3556 -11400
rect 3591 -11438 3667 -11432
rect 3591 -11472 3607 -11438
rect 3651 -11472 3667 -11438
rect 3591 -11488 3667 -11472
rect 3503 -11810 3513 -11757
rect 3566 -11810 3576 -11757
rect 3612 -11919 3646 -11488
rect 3415 -11972 3425 -11919
rect 3478 -11972 3488 -11919
rect 3593 -11972 3603 -11919
rect 3656 -11972 3666 -11919
rect 3434 -12032 3468 -11972
rect 3612 -12032 3646 -11972
rect 3413 -12048 3489 -12032
rect 3413 -12082 3429 -12048
rect 3473 -12082 3489 -12048
rect 3413 -12088 3489 -12082
rect 3591 -12048 3667 -12032
rect 3591 -12082 3607 -12048
rect 3651 -12082 3667 -12048
rect 3591 -12088 3667 -12082
rect 3701 -12120 3735 -11400
rect 3769 -11438 3845 -11432
rect 3769 -11472 3785 -11438
rect 3829 -11472 3845 -11438
rect 3769 -11488 3845 -11472
rect 3881 -11437 3915 -11400
rect 3947 -11437 4023 -11432
rect 4056 -11437 4090 -11400
rect 3881 -11438 4090 -11437
rect 3881 -11471 3963 -11438
rect 3790 -11919 3824 -11488
rect 3881 -11638 3915 -11471
rect 3947 -11472 3963 -11471
rect 4007 -11471 4090 -11438
rect 4007 -11472 4023 -11471
rect 3947 -11488 4023 -11472
rect 3861 -11691 3871 -11638
rect 3924 -11691 3934 -11638
rect 3771 -11972 3781 -11919
rect 3834 -11972 3844 -11919
rect 3790 -12032 3824 -11972
rect 3769 -12048 3845 -12032
rect 3769 -12082 3785 -12048
rect 3829 -12082 3845 -12048
rect 3769 -12088 3845 -12082
rect 3881 -12120 3915 -11691
rect 3947 -12048 4023 -12032
rect 3947 -12082 3963 -12048
rect 4007 -12082 4023 -12048
rect 3947 -12088 4023 -12082
rect -2179 -12132 -2133 -12120
rect -2179 -12388 -2173 -12132
rect -2139 -12388 -2133 -12132
rect -2179 -12400 -2133 -12388
rect -2001 -12132 -1955 -12120
rect -2001 -12388 -1995 -12132
rect -1961 -12388 -1955 -12132
rect -2001 -12400 -1955 -12388
rect -1823 -12132 -1777 -12120
rect -1823 -12388 -1817 -12132
rect -1783 -12388 -1777 -12132
rect -1823 -12400 -1777 -12388
rect -1645 -12132 -1599 -12120
rect -1645 -12388 -1639 -12132
rect -1605 -12388 -1599 -12132
rect -1645 -12400 -1599 -12388
rect -1467 -12132 -1421 -12120
rect -1467 -12388 -1461 -12132
rect -1427 -12388 -1421 -12132
rect -1467 -12400 -1421 -12388
rect -1289 -12132 -1243 -12120
rect -1289 -12388 -1283 -12132
rect -1249 -12388 -1243 -12132
rect -1289 -12400 -1243 -12388
rect -1111 -12132 -1065 -12120
rect -1111 -12388 -1105 -12132
rect -1071 -12388 -1065 -12132
rect -1111 -12400 -1065 -12388
rect -933 -12132 -887 -12120
rect -933 -12388 -927 -12132
rect -893 -12388 -887 -12132
rect -933 -12400 -887 -12388
rect -755 -12132 -709 -12120
rect -755 -12388 -749 -12132
rect -715 -12388 -709 -12132
rect -755 -12400 -709 -12388
rect -577 -12132 -531 -12120
rect -577 -12388 -571 -12132
rect -537 -12388 -531 -12132
rect -577 -12400 -531 -12388
rect -399 -12132 -353 -12120
rect -399 -12388 -393 -12132
rect -359 -12388 -353 -12132
rect -399 -12400 -353 -12388
rect -221 -12132 -175 -12120
rect -221 -12388 -215 -12132
rect -181 -12388 -175 -12132
rect -221 -12400 -175 -12388
rect -43 -12132 3 -12120
rect -43 -12388 -37 -12132
rect -3 -12388 3 -12132
rect -43 -12400 3 -12388
rect 135 -12132 181 -12120
rect 135 -12388 141 -12132
rect 175 -12388 181 -12132
rect 135 -12400 181 -12388
rect 313 -12132 359 -12120
rect 313 -12388 319 -12132
rect 353 -12388 359 -12132
rect 313 -12400 359 -12388
rect 491 -12132 537 -12120
rect 491 -12388 497 -12132
rect 531 -12388 537 -12132
rect 491 -12400 537 -12388
rect 669 -12132 715 -12120
rect 669 -12388 675 -12132
rect 709 -12388 715 -12132
rect 669 -12400 715 -12388
rect 847 -12132 893 -12120
rect 847 -12388 853 -12132
rect 887 -12388 893 -12132
rect 847 -12400 893 -12388
rect 1025 -12132 1071 -12120
rect 1025 -12388 1031 -12132
rect 1065 -12388 1071 -12132
rect 1025 -12400 1071 -12388
rect 1203 -12132 1249 -12120
rect 1203 -12388 1209 -12132
rect 1243 -12388 1249 -12132
rect 1203 -12400 1249 -12388
rect 1381 -12132 1427 -12120
rect 1381 -12388 1387 -12132
rect 1421 -12388 1427 -12132
rect 1381 -12400 1427 -12388
rect 1559 -12132 1605 -12120
rect 1559 -12388 1565 -12132
rect 1599 -12388 1605 -12132
rect 1559 -12400 1605 -12388
rect 1737 -12132 1783 -12120
rect 1737 -12388 1743 -12132
rect 1777 -12388 1783 -12132
rect 1737 -12400 1783 -12388
rect 1915 -12132 1961 -12120
rect 1915 -12388 1921 -12132
rect 1955 -12388 1961 -12132
rect 1915 -12400 1961 -12388
rect 2093 -12132 2139 -12120
rect 2093 -12388 2099 -12132
rect 2133 -12388 2139 -12132
rect 2093 -12400 2139 -12388
rect 2271 -12132 2317 -12120
rect 2271 -12388 2277 -12132
rect 2311 -12388 2317 -12132
rect 2271 -12400 2317 -12388
rect 2449 -12132 2495 -12120
rect 2449 -12388 2455 -12132
rect 2489 -12388 2495 -12132
rect 2449 -12400 2495 -12388
rect 2627 -12132 2673 -12120
rect 2627 -12388 2633 -12132
rect 2667 -12388 2673 -12132
rect 2627 -12400 2673 -12388
rect 2805 -12132 2851 -12120
rect 2805 -12388 2811 -12132
rect 2845 -12388 2851 -12132
rect 2805 -12400 2851 -12388
rect 2983 -12132 3029 -12120
rect 2983 -12388 2989 -12132
rect 3023 -12388 3029 -12132
rect 2983 -12400 3029 -12388
rect 3161 -12132 3207 -12120
rect 3161 -12388 3167 -12132
rect 3201 -12388 3207 -12132
rect 3161 -12400 3207 -12388
rect 3339 -12132 3385 -12120
rect 3339 -12388 3345 -12132
rect 3379 -12388 3385 -12132
rect 3339 -12400 3385 -12388
rect 3517 -12132 3563 -12120
rect 3517 -12388 3523 -12132
rect 3557 -12388 3563 -12132
rect 3517 -12400 3563 -12388
rect 3695 -12132 3741 -12120
rect 3695 -12388 3701 -12132
rect 3735 -12388 3741 -12132
rect 3695 -12400 3741 -12388
rect 3873 -12132 3919 -12120
rect 3873 -12388 3879 -12132
rect 3913 -12388 3919 -12132
rect 3873 -12400 3919 -12388
rect 4051 -12132 4097 -12120
rect 4051 -12388 4057 -12132
rect 4091 -12388 4097 -12132
rect 4051 -12400 4097 -12388
rect -2105 -12438 -2029 -12432
rect -2105 -12472 -2089 -12438
rect -2045 -12472 -2029 -12438
rect -2105 -12488 -2029 -12472
rect -1995 -12542 -1961 -12400
rect -1927 -12438 -1851 -12432
rect -1927 -12472 -1911 -12438
rect -1867 -12472 -1851 -12438
rect -1927 -12488 -1851 -12472
rect -2015 -12595 -2005 -12542
rect -1952 -12595 -1942 -12542
rect -2105 -13046 -2029 -13032
rect -1995 -13046 -1961 -12595
rect -1906 -13032 -1872 -12488
rect -2174 -13048 -1961 -13046
rect -2174 -13080 -2089 -13048
rect -2174 -13120 -2140 -13080
rect -2105 -13082 -2089 -13080
rect -2045 -13080 -1961 -13048
rect -2045 -13082 -2029 -13080
rect -2105 -13088 -2029 -13082
rect -1995 -13120 -1961 -13080
rect -1927 -13048 -1851 -13032
rect -1927 -13082 -1911 -13048
rect -1867 -13082 -1851 -13048
rect -1927 -13088 -1851 -13082
rect -1818 -13120 -1784 -12400
rect -1749 -12438 -1673 -12432
rect -1749 -12472 -1733 -12438
rect -1689 -12472 -1673 -12438
rect -1749 -12488 -1673 -12472
rect -1728 -13032 -1694 -12488
rect -1639 -12542 -1605 -12400
rect -1571 -12438 -1495 -12432
rect -1571 -12472 -1555 -12438
rect -1511 -12472 -1495 -12438
rect -1571 -12488 -1495 -12472
rect -1659 -12595 -1649 -12542
rect -1596 -12595 -1586 -12542
rect -1549 -13032 -1515 -12488
rect -1749 -13048 -1673 -13032
rect -1749 -13082 -1733 -13048
rect -1689 -13082 -1673 -13048
rect -1749 -13088 -1673 -13082
rect -1571 -13048 -1495 -13032
rect -1571 -13082 -1555 -13048
rect -1511 -13082 -1495 -13048
rect -1571 -13088 -1495 -13082
rect -1461 -13120 -1427 -12400
rect -1393 -12438 -1317 -12432
rect -1393 -12472 -1377 -12438
rect -1333 -12472 -1317 -12438
rect -1393 -12488 -1317 -12472
rect -1372 -13032 -1338 -12488
rect -1284 -12654 -1250 -12400
rect -1215 -12438 -1139 -12432
rect -1215 -12472 -1199 -12438
rect -1155 -12472 -1139 -12438
rect -1215 -12488 -1139 -12472
rect -1304 -12707 -1294 -12654
rect -1241 -12707 -1231 -12654
rect -1194 -13032 -1160 -12488
rect -1393 -13048 -1317 -13032
rect -1393 -13082 -1377 -13048
rect -1333 -13082 -1317 -13048
rect -1393 -13088 -1317 -13082
rect -1215 -13048 -1139 -13032
rect -1215 -13082 -1199 -13048
rect -1155 -13082 -1139 -13048
rect -1215 -13088 -1139 -13082
rect -1105 -13120 -1071 -12400
rect -1037 -12438 -961 -12432
rect -1037 -12472 -1021 -12438
rect -977 -12472 -961 -12438
rect -1037 -12488 -961 -12472
rect -1016 -13032 -982 -12488
rect -927 -12783 -893 -12400
rect -859 -12438 -783 -12432
rect -859 -12472 -843 -12438
rect -799 -12472 -783 -12438
rect -859 -12488 -783 -12472
rect -947 -12836 -937 -12783
rect -884 -12836 -874 -12783
rect -1037 -13048 -961 -13032
rect -1037 -13082 -1021 -13048
rect -977 -13082 -961 -13048
rect -1037 -13088 -961 -13082
rect -927 -13120 -893 -12836
rect -838 -13032 -804 -12488
rect -859 -13048 -783 -13032
rect -859 -13082 -843 -13048
rect -799 -13082 -783 -13048
rect -859 -13088 -783 -13082
rect -749 -13120 -715 -12400
rect -681 -12438 -605 -12432
rect -681 -12472 -665 -12438
rect -621 -12472 -605 -12438
rect -681 -12488 -605 -12472
rect -660 -13032 -626 -12488
rect -571 -12653 -537 -12400
rect -503 -12438 -427 -12432
rect -503 -12472 -487 -12438
rect -443 -12472 -427 -12438
rect -503 -12488 -427 -12472
rect -592 -12706 -582 -12653
rect -529 -12706 -519 -12653
rect -482 -13032 -448 -12488
rect -681 -13048 -605 -13032
rect -681 -13082 -665 -13048
rect -621 -13082 -605 -13048
rect -681 -13088 -605 -13082
rect -503 -13048 -427 -13032
rect -503 -13082 -487 -13048
rect -443 -13082 -427 -13048
rect -503 -13088 -427 -13082
rect -393 -13120 -359 -12400
rect -325 -12438 -249 -12432
rect -325 -12472 -309 -12438
rect -265 -12472 -249 -12438
rect -325 -12488 -249 -12472
rect -304 -13032 -270 -12488
rect -215 -12783 -181 -12400
rect -147 -12438 -71 -12432
rect -147 -12472 -131 -12438
rect -87 -12472 -71 -12438
rect -147 -12488 -71 -12472
rect -234 -12836 -224 -12783
rect -171 -12836 -161 -12783
rect -126 -13032 -92 -12488
rect -325 -13048 -249 -13032
rect -325 -13082 -309 -13048
rect -265 -13082 -249 -13048
rect -325 -13088 -249 -13082
rect -147 -13048 -71 -13032
rect -147 -13082 -131 -13048
rect -87 -13082 -71 -13048
rect -147 -13088 -71 -13082
rect -36 -13120 -2 -12400
rect 31 -12438 107 -12432
rect 31 -12472 47 -12438
rect 91 -12472 107 -12438
rect 31 -12488 107 -12472
rect 52 -13032 86 -12488
rect 141 -12653 175 -12400
rect 209 -12438 285 -12432
rect 209 -12472 225 -12438
rect 269 -12472 285 -12438
rect 209 -12488 285 -12472
rect 120 -12706 130 -12653
rect 183 -12706 193 -12653
rect 31 -13048 107 -13032
rect 31 -13082 47 -13048
rect 91 -13082 107 -13048
rect 31 -13088 107 -13082
rect 141 -13120 175 -12706
rect 230 -13032 264 -12488
rect 209 -13048 285 -13032
rect 209 -13082 225 -13048
rect 269 -13082 285 -13048
rect 209 -13088 285 -13082
rect 319 -13120 353 -12400
rect 387 -12438 463 -12432
rect 387 -12472 403 -12438
rect 447 -12472 463 -12438
rect 387 -12488 463 -12472
rect 408 -13032 442 -12488
rect 496 -12784 530 -12400
rect 565 -12438 641 -12432
rect 565 -12472 581 -12438
rect 625 -12472 641 -12438
rect 565 -12488 641 -12472
rect 476 -12837 486 -12784
rect 539 -12837 549 -12784
rect 587 -13032 621 -12488
rect 387 -13048 463 -13032
rect 387 -13082 403 -13048
rect 447 -13082 463 -13048
rect 387 -13088 463 -13082
rect 565 -13048 641 -13032
rect 565 -13082 581 -13048
rect 625 -13082 641 -13048
rect 565 -13088 641 -13082
rect 675 -13120 709 -12400
rect 743 -12438 819 -12432
rect 852 -12438 886 -12400
rect 921 -12438 997 -12432
rect 1031 -12438 1065 -12400
rect 1099 -12438 1175 -12432
rect 743 -12472 759 -12438
rect 803 -12472 937 -12438
rect 981 -12472 1115 -12438
rect 1159 -12472 1175 -12438
rect 743 -12488 819 -12472
rect 921 -12488 997 -12472
rect 1099 -12488 1175 -12472
rect 942 -13032 976 -12488
rect 743 -13048 819 -13032
rect 921 -13048 997 -13032
rect 1099 -13048 1175 -13032
rect 743 -13082 759 -13048
rect 803 -13082 937 -13048
rect 981 -13082 1115 -13048
rect 1159 -13082 1175 -13048
rect 743 -13088 819 -13082
rect 852 -13120 886 -13082
rect 921 -13088 997 -13082
rect 1032 -13120 1066 -13082
rect 1099 -13088 1175 -13082
rect 1209 -13120 1243 -12400
rect 1277 -12438 1353 -12432
rect 1277 -12472 1293 -12438
rect 1337 -12472 1353 -12438
rect 1277 -12488 1353 -12472
rect 1299 -13032 1333 -12488
rect 1388 -12783 1422 -12400
rect 1455 -12438 1531 -12432
rect 1455 -12472 1471 -12438
rect 1515 -12472 1531 -12438
rect 1455 -12488 1531 -12472
rect 1368 -12836 1378 -12783
rect 1431 -12836 1441 -12783
rect 1277 -13048 1353 -13032
rect 1277 -13082 1293 -13048
rect 1337 -13082 1353 -13048
rect 1277 -13088 1353 -13082
rect 1388 -13120 1422 -12836
rect 1476 -13032 1510 -12488
rect 1455 -13048 1531 -13032
rect 1455 -13082 1471 -13048
rect 1515 -13082 1531 -13048
rect 1455 -13088 1531 -13082
rect 1566 -13120 1600 -12400
rect 1633 -12438 1709 -12432
rect 1633 -12472 1649 -12438
rect 1693 -12472 1709 -12438
rect 1633 -12488 1709 -12472
rect 1655 -13032 1689 -12488
rect 1744 -12654 1778 -12400
rect 1811 -12438 1887 -12432
rect 1811 -12472 1827 -12438
rect 1871 -12472 1887 -12438
rect 1811 -12488 1887 -12472
rect 1725 -12707 1735 -12654
rect 1788 -12707 1798 -12654
rect 1833 -13032 1867 -12488
rect 1633 -13048 1709 -13032
rect 1633 -13082 1649 -13048
rect 1693 -13082 1709 -13048
rect 1633 -13088 1709 -13082
rect 1811 -13048 1887 -13032
rect 1811 -13082 1827 -13048
rect 1871 -13082 1887 -13048
rect 1811 -13088 1887 -13082
rect 1922 -13120 1956 -12400
rect 1989 -12438 2065 -12432
rect 1989 -12472 2005 -12438
rect 2049 -12472 2065 -12438
rect 1989 -12488 2065 -12472
rect 2009 -13032 2043 -12488
rect 2098 -12782 2132 -12400
rect 2167 -12438 2243 -12432
rect 2167 -12472 2183 -12438
rect 2227 -12472 2243 -12438
rect 2167 -12488 2243 -12472
rect 2078 -12835 2088 -12782
rect 2141 -12835 2151 -12782
rect 1989 -13048 2065 -13032
rect 1989 -13082 2005 -13048
rect 2049 -13082 2065 -13048
rect 1989 -13088 2065 -13082
rect 2098 -13120 2132 -12835
rect 2188 -13032 2222 -12488
rect 2167 -13048 2243 -13032
rect 2167 -13082 2183 -13048
rect 2227 -13082 2243 -13048
rect 2167 -13088 2243 -13082
rect 2277 -13120 2311 -12400
rect 2345 -12438 2421 -12432
rect 2345 -12472 2361 -12438
rect 2405 -12472 2421 -12438
rect 2345 -12488 2421 -12472
rect 2366 -13032 2400 -12488
rect 2455 -12653 2489 -12400
rect 2523 -12438 2599 -12432
rect 2523 -12472 2539 -12438
rect 2583 -12472 2599 -12438
rect 2523 -12488 2599 -12472
rect 2435 -12706 2445 -12653
rect 2498 -12706 2508 -12653
rect 2544 -13032 2578 -12488
rect 2345 -13048 2421 -13032
rect 2345 -13082 2361 -13048
rect 2405 -13082 2421 -13048
rect 2345 -13088 2421 -13082
rect 2523 -13048 2599 -13032
rect 2523 -13082 2539 -13048
rect 2583 -13082 2599 -13048
rect 2523 -13088 2599 -13082
rect 2633 -13120 2667 -12400
rect 2701 -12438 2777 -12432
rect 2701 -12472 2717 -12438
rect 2761 -12472 2777 -12438
rect 2701 -12488 2777 -12472
rect 2722 -13032 2756 -12488
rect 2811 -12782 2845 -12400
rect 2879 -12438 2955 -12432
rect 2879 -12472 2895 -12438
rect 2939 -12472 2955 -12438
rect 2879 -12488 2955 -12472
rect 2791 -12835 2801 -12782
rect 2854 -12835 2864 -12782
rect 2900 -13032 2934 -12488
rect 2701 -13048 2777 -13032
rect 2701 -13082 2717 -13048
rect 2761 -13082 2777 -13048
rect 2701 -13088 2777 -13082
rect 2879 -13048 2955 -13032
rect 2879 -13082 2895 -13048
rect 2939 -13082 2955 -13048
rect 2879 -13088 2955 -13082
rect 2989 -13120 3023 -12400
rect 3057 -12438 3133 -12432
rect 3057 -12472 3073 -12438
rect 3117 -12472 3133 -12438
rect 3057 -12488 3133 -12472
rect 3078 -13032 3112 -12488
rect 3167 -12650 3201 -12400
rect 3235 -12438 3311 -12432
rect 3235 -12472 3251 -12438
rect 3295 -12472 3311 -12438
rect 3235 -12488 3311 -12472
rect 3166 -12652 3201 -12650
rect 3148 -12705 3158 -12652
rect 3211 -12705 3221 -12652
rect 3057 -13048 3133 -13032
rect 3057 -13082 3073 -13048
rect 3117 -13082 3133 -13048
rect 3057 -13088 3133 -13082
rect 3166 -13120 3200 -12705
rect 3256 -13032 3290 -12488
rect 3235 -13048 3311 -13032
rect 3235 -13082 3251 -13048
rect 3295 -13082 3311 -13048
rect 3235 -13088 3311 -13082
rect 3345 -13120 3379 -12400
rect 3413 -12438 3489 -12432
rect 3413 -12472 3429 -12438
rect 3473 -12472 3489 -12438
rect 3413 -12488 3489 -12472
rect 3434 -13032 3468 -12488
rect 3524 -12542 3558 -12400
rect 3591 -12438 3667 -12432
rect 3591 -12472 3607 -12438
rect 3651 -12472 3667 -12438
rect 3591 -12488 3667 -12472
rect 3504 -12595 3514 -12542
rect 3567 -12595 3577 -12542
rect 3613 -13032 3647 -12488
rect 3413 -13048 3489 -13032
rect 3413 -13082 3429 -13048
rect 3473 -13082 3489 -13048
rect 3413 -13088 3489 -13082
rect 3591 -13048 3667 -13032
rect 3591 -13082 3607 -13048
rect 3651 -13082 3667 -13048
rect 3591 -13088 3667 -13082
rect 3701 -13120 3735 -12400
rect 3769 -12438 3845 -12432
rect 3769 -12472 3785 -12438
rect 3829 -12472 3845 -12438
rect 3769 -12488 3845 -12472
rect 3881 -12436 3915 -12400
rect 3947 -12436 4023 -12432
rect 4058 -12436 4092 -12400
rect 3881 -12438 4092 -12436
rect 3881 -12470 3963 -12438
rect 3790 -13032 3824 -12488
rect 3881 -12542 3915 -12470
rect 3947 -12472 3963 -12470
rect 4007 -12470 4092 -12438
rect 4007 -12472 4023 -12470
rect 3947 -12488 4023 -12472
rect 3861 -12595 3871 -12542
rect 3924 -12595 3934 -12542
rect 3769 -13048 3845 -13032
rect 3769 -13082 3785 -13048
rect 3829 -13082 3845 -13048
rect 3769 -13088 3845 -13082
rect 3881 -13047 3915 -12595
rect 3947 -13047 4023 -13032
rect 3881 -13048 4090 -13047
rect 3881 -13081 3963 -13048
rect 3881 -13120 3915 -13081
rect 3947 -13082 3963 -13081
rect 4007 -13081 4090 -13048
rect 4007 -13082 4023 -13081
rect 3947 -13088 4023 -13082
rect 4056 -13120 4090 -13081
rect -2179 -13132 -2133 -13120
rect -2179 -13388 -2173 -13132
rect -2139 -13388 -2133 -13132
rect -2179 -13400 -2133 -13388
rect -2001 -13132 -1955 -13120
rect -2001 -13388 -1995 -13132
rect -1961 -13388 -1955 -13132
rect -2001 -13400 -1955 -13388
rect -1823 -13132 -1777 -13120
rect -1823 -13388 -1817 -13132
rect -1783 -13388 -1777 -13132
rect -1823 -13400 -1777 -13388
rect -1645 -13132 -1599 -13120
rect -1645 -13388 -1639 -13132
rect -1605 -13388 -1599 -13132
rect -1645 -13400 -1599 -13388
rect -1467 -13132 -1421 -13120
rect -1467 -13388 -1461 -13132
rect -1427 -13388 -1421 -13132
rect -1467 -13400 -1421 -13388
rect -1289 -13132 -1243 -13120
rect -1289 -13388 -1283 -13132
rect -1249 -13388 -1243 -13132
rect -1289 -13400 -1243 -13388
rect -1111 -13132 -1065 -13120
rect -1111 -13388 -1105 -13132
rect -1071 -13388 -1065 -13132
rect -1111 -13400 -1065 -13388
rect -933 -13132 -887 -13120
rect -933 -13388 -927 -13132
rect -893 -13388 -887 -13132
rect -933 -13400 -887 -13388
rect -755 -13132 -709 -13120
rect -755 -13388 -749 -13132
rect -715 -13388 -709 -13132
rect -755 -13400 -709 -13388
rect -577 -13132 -531 -13120
rect -577 -13388 -571 -13132
rect -537 -13388 -531 -13132
rect -577 -13400 -531 -13388
rect -399 -13132 -353 -13120
rect -399 -13388 -393 -13132
rect -359 -13388 -353 -13132
rect -399 -13400 -353 -13388
rect -221 -13132 -175 -13120
rect -221 -13388 -215 -13132
rect -181 -13388 -175 -13132
rect -221 -13400 -175 -13388
rect -43 -13132 3 -13120
rect -43 -13388 -37 -13132
rect -3 -13388 3 -13132
rect -43 -13400 3 -13388
rect 135 -13132 181 -13120
rect 135 -13388 141 -13132
rect 175 -13388 181 -13132
rect 135 -13400 181 -13388
rect 313 -13132 359 -13120
rect 313 -13388 319 -13132
rect 353 -13388 359 -13132
rect 313 -13400 359 -13388
rect 491 -13132 537 -13120
rect 491 -13388 497 -13132
rect 531 -13388 537 -13132
rect 491 -13400 537 -13388
rect 669 -13132 715 -13120
rect 669 -13388 675 -13132
rect 709 -13388 715 -13132
rect 669 -13400 715 -13388
rect 847 -13132 893 -13120
rect 847 -13388 853 -13132
rect 887 -13388 893 -13132
rect 847 -13400 893 -13388
rect 1025 -13132 1071 -13120
rect 1025 -13388 1031 -13132
rect 1065 -13388 1071 -13132
rect 1025 -13400 1071 -13388
rect 1203 -13132 1249 -13120
rect 1203 -13388 1209 -13132
rect 1243 -13388 1249 -13132
rect 1203 -13400 1249 -13388
rect 1381 -13132 1427 -13120
rect 1381 -13388 1387 -13132
rect 1421 -13388 1427 -13132
rect 1381 -13400 1427 -13388
rect 1559 -13132 1605 -13120
rect 1559 -13388 1565 -13132
rect 1599 -13388 1605 -13132
rect 1559 -13400 1605 -13388
rect 1737 -13132 1783 -13120
rect 1737 -13388 1743 -13132
rect 1777 -13388 1783 -13132
rect 1737 -13400 1783 -13388
rect 1915 -13132 1961 -13120
rect 1915 -13388 1921 -13132
rect 1955 -13388 1961 -13132
rect 1915 -13400 1961 -13388
rect 2093 -13132 2139 -13120
rect 2093 -13388 2099 -13132
rect 2133 -13388 2139 -13132
rect 2093 -13400 2139 -13388
rect 2271 -13132 2317 -13120
rect 2271 -13388 2277 -13132
rect 2311 -13388 2317 -13132
rect 2271 -13400 2317 -13388
rect 2449 -13132 2495 -13120
rect 2449 -13388 2455 -13132
rect 2489 -13388 2495 -13132
rect 2449 -13400 2495 -13388
rect 2627 -13132 2673 -13120
rect 2627 -13388 2633 -13132
rect 2667 -13388 2673 -13132
rect 2627 -13400 2673 -13388
rect 2805 -13132 2851 -13120
rect 2805 -13388 2811 -13132
rect 2845 -13388 2851 -13132
rect 2805 -13400 2851 -13388
rect 2983 -13132 3029 -13120
rect 2983 -13388 2989 -13132
rect 3023 -13388 3029 -13132
rect 2983 -13400 3029 -13388
rect 3161 -13132 3207 -13120
rect 3161 -13388 3167 -13132
rect 3201 -13388 3207 -13132
rect 3161 -13400 3207 -13388
rect 3339 -13132 3385 -13120
rect 3339 -13388 3345 -13132
rect 3379 -13388 3385 -13132
rect 3339 -13400 3385 -13388
rect 3517 -13132 3563 -13120
rect 3517 -13388 3523 -13132
rect 3557 -13388 3563 -13132
rect 3517 -13400 3563 -13388
rect 3695 -13132 3741 -13120
rect 3695 -13388 3701 -13132
rect 3735 -13388 3741 -13132
rect 3695 -13400 3741 -13388
rect 3873 -13132 3919 -13120
rect 3873 -13388 3879 -13132
rect 3913 -13388 3919 -13132
rect 3873 -13400 3919 -13388
rect 4051 -13132 4097 -13120
rect 4051 -13388 4057 -13132
rect 4091 -13388 4097 -13132
rect 4051 -13400 4097 -13388
rect -2105 -13438 -2029 -13432
rect -2105 -13472 -2089 -13438
rect -2045 -13472 -2029 -13438
rect -2105 -13488 -2029 -13472
rect -1995 -13545 -1961 -13400
rect -1927 -13438 -1851 -13432
rect -1927 -13472 -1911 -13438
rect -1867 -13472 -1851 -13438
rect -1927 -13488 -1851 -13472
rect -1749 -13438 -1673 -13432
rect -1749 -13472 -1733 -13438
rect -1689 -13472 -1673 -13438
rect -1749 -13488 -1673 -13472
rect -2014 -13598 -2004 -13545
rect -1951 -13598 -1941 -13545
rect -1905 -14032 -1871 -13488
rect -1728 -14032 -1694 -13488
rect -1638 -13672 -1604 -13400
rect -1571 -13438 -1495 -13432
rect -1571 -13472 -1555 -13438
rect -1511 -13472 -1495 -13438
rect -1571 -13488 -1495 -13472
rect -1393 -13438 -1317 -13432
rect -1393 -13472 -1377 -13438
rect -1333 -13472 -1317 -13438
rect -1393 -13488 -1317 -13472
rect -1658 -13725 -1648 -13672
rect -1595 -13725 -1585 -13672
rect -1550 -14032 -1516 -13488
rect -1282 -13672 -1248 -13400
rect -1215 -13438 -1139 -13432
rect -1215 -13472 -1199 -13438
rect -1155 -13472 -1139 -13438
rect -1215 -13488 -1139 -13472
rect -1037 -13438 -961 -13432
rect -1037 -13472 -1021 -13438
rect -977 -13472 -961 -13438
rect -1037 -13488 -961 -13472
rect -927 -13672 -893 -13400
rect -859 -13438 -783 -13432
rect -859 -13472 -843 -13438
rect -799 -13472 -783 -13438
rect -859 -13488 -783 -13472
rect -681 -13438 -605 -13432
rect -681 -13472 -665 -13438
rect -621 -13472 -605 -13438
rect -681 -13488 -605 -13472
rect -571 -13545 -537 -13400
rect -503 -13438 -427 -13432
rect -503 -13472 -487 -13438
rect -443 -13472 -427 -13438
rect -503 -13488 -427 -13472
rect -325 -13438 -249 -13432
rect -325 -13472 -309 -13438
rect -265 -13472 -249 -13438
rect -325 -13488 -249 -13472
rect -591 -13598 -581 -13545
rect -528 -13598 -518 -13545
rect -1301 -13725 -1291 -13672
rect -1238 -13725 -1228 -13672
rect -947 -13725 -937 -13672
rect -884 -13725 -874 -13672
rect -927 -13726 -893 -13725
rect -304 -14032 -270 -13488
rect -216 -13794 -182 -13400
rect -147 -13438 -71 -13432
rect -147 -13472 -131 -13438
rect -87 -13472 -71 -13438
rect -147 -13488 -71 -13472
rect 31 -13438 107 -13432
rect 31 -13472 47 -13438
rect 91 -13472 107 -13438
rect 31 -13488 107 -13472
rect -235 -13847 -225 -13794
rect -172 -13847 -162 -13794
rect -125 -14032 -91 -13488
rect 52 -14032 86 -13488
rect 141 -13794 175 -13400
rect 209 -13438 285 -13432
rect 209 -13472 225 -13438
rect 269 -13472 285 -13438
rect 209 -13488 285 -13472
rect 387 -13438 463 -13432
rect 387 -13472 403 -13438
rect 447 -13472 463 -13438
rect 387 -13488 463 -13472
rect 123 -13847 133 -13794
rect 186 -13847 196 -13794
rect 230 -14032 264 -13488
rect 408 -14032 442 -13488
rect 496 -13795 530 -13400
rect 942 -13432 976 -13430
rect 565 -13438 641 -13432
rect 565 -13472 581 -13438
rect 625 -13472 641 -13438
rect 565 -13488 641 -13472
rect 743 -13438 819 -13432
rect 743 -13472 759 -13438
rect 803 -13472 819 -13438
rect 743 -13488 819 -13472
rect 921 -13438 997 -13432
rect 921 -13472 937 -13438
rect 981 -13472 997 -13438
rect 921 -13488 997 -13472
rect 1099 -13438 1175 -13432
rect 1099 -13472 1115 -13438
rect 1159 -13472 1175 -13438
rect 1099 -13488 1175 -13472
rect 1277 -13438 1353 -13432
rect 1277 -13472 1293 -13438
rect 1337 -13472 1353 -13438
rect 1277 -13488 1353 -13472
rect 477 -13848 487 -13795
rect 540 -13848 550 -13795
rect 587 -14032 621 -13488
rect 942 -14032 976 -13488
rect 1388 -13672 1422 -13400
rect 1455 -13438 1531 -13432
rect 1455 -13472 1471 -13438
rect 1515 -13472 1531 -13438
rect 1455 -13488 1531 -13472
rect 1633 -13438 1709 -13432
rect 1633 -13472 1649 -13438
rect 1693 -13472 1709 -13438
rect 1633 -13488 1709 -13472
rect 1743 -13672 1777 -13400
rect 1811 -13438 1887 -13432
rect 1811 -13472 1827 -13438
rect 1871 -13472 1887 -13438
rect 1811 -13488 1887 -13472
rect 1989 -13438 2065 -13432
rect 1989 -13472 2005 -13438
rect 2049 -13472 2065 -13438
rect 1989 -13488 2065 -13472
rect 2100 -13672 2134 -13400
rect 2167 -13438 2243 -13432
rect 2167 -13472 2183 -13438
rect 2227 -13472 2243 -13438
rect 2167 -13488 2243 -13472
rect 2345 -13438 2421 -13432
rect 2345 -13472 2361 -13438
rect 2405 -13472 2421 -13438
rect 2345 -13488 2421 -13472
rect 1369 -13725 1379 -13672
rect 1432 -13725 1442 -13672
rect 1722 -13725 1732 -13672
rect 1785 -13725 1795 -13672
rect 2081 -13725 2091 -13672
rect 2144 -13725 2154 -13672
rect 2366 -14032 2400 -13488
rect 2455 -13545 2489 -13400
rect 2523 -13438 2599 -13432
rect 2523 -13472 2539 -13438
rect 2583 -13472 2599 -13438
rect 2523 -13488 2599 -13472
rect 2701 -13438 2777 -13432
rect 2701 -13472 2717 -13438
rect 2761 -13472 2777 -13438
rect 2701 -13488 2777 -13472
rect 2436 -13598 2446 -13545
rect 2499 -13598 2509 -13545
rect 2544 -14032 2578 -13488
rect 2723 -14032 2757 -13488
rect 2812 -13794 2846 -13400
rect 2879 -13438 2955 -13432
rect 2879 -13472 2895 -13438
rect 2939 -13472 2955 -13438
rect 2879 -13488 2955 -13472
rect 3057 -13438 3133 -13432
rect 3057 -13472 3073 -13438
rect 3117 -13472 3133 -13438
rect 3057 -13488 3133 -13472
rect 2792 -13847 2802 -13794
rect 2855 -13847 2865 -13794
rect 2901 -14032 2935 -13488
rect 3078 -14032 3112 -13488
rect 3166 -13795 3200 -13400
rect 3257 -13432 3291 -13431
rect 3235 -13438 3311 -13432
rect 3235 -13472 3251 -13438
rect 3295 -13472 3311 -13438
rect 3235 -13488 3311 -13472
rect 3413 -13438 3489 -13432
rect 3413 -13472 3429 -13438
rect 3473 -13472 3489 -13438
rect 3413 -13488 3489 -13472
rect 3147 -13848 3157 -13795
rect 3210 -13848 3220 -13795
rect 3257 -14032 3291 -13488
rect 3523 -13794 3557 -13400
rect 3591 -13438 3667 -13432
rect 3591 -13472 3607 -13438
rect 3651 -13472 3667 -13438
rect 3591 -13488 3667 -13472
rect 3769 -13438 3845 -13432
rect 3769 -13472 3785 -13438
rect 3829 -13472 3845 -13438
rect 3769 -13488 3845 -13472
rect 3879 -13545 3913 -13400
rect 3947 -13438 4023 -13432
rect 3947 -13472 3963 -13438
rect 4007 -13472 4023 -13438
rect 3947 -13488 4023 -13472
rect 3860 -13598 3870 -13545
rect 3923 -13598 3933 -13545
rect 3502 -13847 3512 -13794
rect 3565 -13847 3575 -13794
rect 3523 -13848 3557 -13847
rect -2105 -14048 -2029 -14032
rect -2105 -14082 -2089 -14048
rect -2045 -14082 -2029 -14048
rect -2105 -14088 -2029 -14082
rect -1927 -14048 -1851 -14032
rect -1927 -14082 -1911 -14048
rect -1867 -14082 -1851 -14048
rect -1927 -14088 -1851 -14082
rect -1749 -14048 -1673 -14032
rect -1749 -14082 -1733 -14048
rect -1689 -14082 -1673 -14048
rect -1749 -14088 -1673 -14082
rect -1571 -14048 -1495 -14032
rect -1571 -14082 -1555 -14048
rect -1511 -14082 -1495 -14048
rect -1571 -14088 -1495 -14082
rect -1393 -14048 -1317 -14032
rect -1393 -14082 -1377 -14048
rect -1333 -14082 -1317 -14048
rect -1393 -14088 -1317 -14082
rect -1215 -14048 -1139 -14032
rect -1215 -14082 -1199 -14048
rect -1155 -14082 -1139 -14048
rect -1215 -14088 -1139 -14082
rect -1037 -14048 -961 -14032
rect -1037 -14082 -1021 -14048
rect -977 -14082 -961 -14048
rect -1037 -14088 -961 -14082
rect -859 -14048 -783 -14032
rect -859 -14082 -843 -14048
rect -799 -14082 -783 -14048
rect -859 -14088 -783 -14082
rect -681 -14048 -605 -14032
rect -681 -14082 -665 -14048
rect -621 -14082 -605 -14048
rect -681 -14088 -605 -14082
rect -503 -14048 -427 -14032
rect -503 -14082 -487 -14048
rect -443 -14082 -427 -14048
rect -503 -14088 -427 -14082
rect -325 -14048 -249 -14032
rect -325 -14082 -309 -14048
rect -265 -14082 -249 -14048
rect -325 -14088 -249 -14082
rect -147 -14048 -71 -14032
rect -147 -14082 -131 -14048
rect -87 -14082 -71 -14048
rect -147 -14088 -71 -14082
rect 31 -14048 107 -14032
rect 31 -14082 47 -14048
rect 91 -14082 107 -14048
rect 31 -14088 107 -14082
rect 209 -14048 285 -14032
rect 209 -14082 225 -14048
rect 269 -14082 285 -14048
rect 209 -14088 285 -14082
rect 387 -14048 463 -14032
rect 387 -14082 403 -14048
rect 447 -14082 463 -14048
rect 387 -14088 463 -14082
rect 565 -14048 641 -14032
rect 565 -14082 581 -14048
rect 625 -14082 641 -14048
rect 565 -14088 641 -14082
rect 743 -14048 819 -14032
rect 921 -14048 997 -14032
rect 1099 -14048 1175 -14032
rect 743 -14082 759 -14048
rect 803 -14082 937 -14048
rect 981 -14082 1115 -14048
rect 1159 -14082 1175 -14048
rect 743 -14088 819 -14082
rect 853 -14120 887 -14082
rect 921 -14088 997 -14082
rect 1032 -14120 1066 -14082
rect 1099 -14088 1175 -14082
rect 1277 -14048 1353 -14032
rect 1277 -14082 1293 -14048
rect 1337 -14082 1353 -14048
rect 1277 -14088 1353 -14082
rect 1455 -14048 1531 -14032
rect 1455 -14082 1471 -14048
rect 1515 -14082 1531 -14048
rect 1455 -14088 1531 -14082
rect 1633 -14048 1709 -14032
rect 1633 -14082 1649 -14048
rect 1693 -14082 1709 -14048
rect 1633 -14088 1709 -14082
rect 1811 -14048 1887 -14032
rect 1811 -14082 1827 -14048
rect 1871 -14082 1887 -14048
rect 1811 -14088 1887 -14082
rect 1989 -14048 2065 -14032
rect 1989 -14082 2005 -14048
rect 2049 -14082 2065 -14048
rect 1989 -14088 2065 -14082
rect 2167 -14048 2243 -14032
rect 2167 -14082 2183 -14048
rect 2227 -14082 2243 -14048
rect 2167 -14088 2243 -14082
rect 2345 -14048 2421 -14032
rect 2345 -14082 2361 -14048
rect 2405 -14082 2421 -14048
rect 2345 -14088 2421 -14082
rect 2523 -14048 2599 -14032
rect 2523 -14082 2539 -14048
rect 2583 -14082 2599 -14048
rect 2523 -14088 2599 -14082
rect 2701 -14048 2777 -14032
rect 2701 -14082 2717 -14048
rect 2761 -14082 2777 -14048
rect 2701 -14088 2777 -14082
rect 2879 -14048 2955 -14032
rect 2879 -14082 2895 -14048
rect 2939 -14082 2955 -14048
rect 2879 -14088 2955 -14082
rect 3057 -14048 3133 -14032
rect 3057 -14082 3073 -14048
rect 3117 -14082 3133 -14048
rect 3057 -14088 3133 -14082
rect 3235 -14048 3311 -14032
rect 3235 -14082 3251 -14048
rect 3295 -14082 3311 -14048
rect 3235 -14088 3311 -14082
rect 3413 -14048 3489 -14032
rect 3413 -14082 3429 -14048
rect 3473 -14082 3489 -14048
rect 3413 -14088 3489 -14082
rect 3591 -14048 3667 -14032
rect 3591 -14082 3607 -14048
rect 3651 -14082 3667 -14048
rect 3591 -14088 3667 -14082
rect 3769 -14048 3845 -14032
rect 3769 -14082 3785 -14048
rect 3829 -14082 3845 -14048
rect 3769 -14088 3845 -14082
rect 3947 -14048 4023 -14032
rect 3947 -14082 3963 -14048
rect 4007 -14082 4023 -14048
rect 3947 -14088 4023 -14082
rect -2179 -14132 -2133 -14120
rect -2179 -14388 -2173 -14132
rect -2139 -14388 -2133 -14132
rect -2179 -14400 -2133 -14388
rect -2001 -14132 -1955 -14120
rect -2001 -14388 -1995 -14132
rect -1961 -14388 -1955 -14132
rect -2001 -14400 -1955 -14388
rect -1823 -14132 -1777 -14120
rect -1823 -14388 -1817 -14132
rect -1783 -14388 -1777 -14132
rect -1823 -14400 -1777 -14388
rect -1645 -14132 -1599 -14120
rect -1645 -14388 -1639 -14132
rect -1605 -14388 -1599 -14132
rect -1645 -14400 -1599 -14388
rect -1467 -14132 -1421 -14120
rect -1467 -14388 -1461 -14132
rect -1427 -14388 -1421 -14132
rect -1467 -14400 -1421 -14388
rect -1289 -14132 -1243 -14120
rect -1289 -14388 -1283 -14132
rect -1249 -14388 -1243 -14132
rect -1289 -14400 -1243 -14388
rect -1111 -14132 -1065 -14120
rect -1111 -14388 -1105 -14132
rect -1071 -14388 -1065 -14132
rect -1111 -14400 -1065 -14388
rect -933 -14132 -887 -14120
rect -933 -14388 -927 -14132
rect -893 -14388 -887 -14132
rect -933 -14400 -887 -14388
rect -755 -14132 -709 -14120
rect -755 -14388 -749 -14132
rect -715 -14388 -709 -14132
rect -755 -14400 -709 -14388
rect -577 -14132 -531 -14120
rect -577 -14388 -571 -14132
rect -537 -14388 -531 -14132
rect -577 -14400 -531 -14388
rect -399 -14132 -353 -14120
rect -399 -14388 -393 -14132
rect -359 -14388 -353 -14132
rect -399 -14400 -353 -14388
rect -221 -14132 -175 -14120
rect -221 -14388 -215 -14132
rect -181 -14388 -175 -14132
rect -221 -14400 -175 -14388
rect -43 -14132 3 -14120
rect -43 -14388 -37 -14132
rect -3 -14388 3 -14132
rect -43 -14400 3 -14388
rect 135 -14132 181 -14120
rect 135 -14388 141 -14132
rect 175 -14388 181 -14132
rect 135 -14400 181 -14388
rect 313 -14132 359 -14120
rect 313 -14388 319 -14132
rect 353 -14388 359 -14132
rect 313 -14400 359 -14388
rect 491 -14132 537 -14120
rect 491 -14388 497 -14132
rect 531 -14388 537 -14132
rect 491 -14400 537 -14388
rect 669 -14132 715 -14120
rect 669 -14388 675 -14132
rect 709 -14388 715 -14132
rect 669 -14400 715 -14388
rect 847 -14132 893 -14120
rect 847 -14388 853 -14132
rect 887 -14388 893 -14132
rect 847 -14400 893 -14388
rect 1025 -14132 1071 -14120
rect 1025 -14388 1031 -14132
rect 1065 -14388 1071 -14132
rect 1025 -14400 1071 -14388
rect 1203 -14132 1249 -14120
rect 1203 -14388 1209 -14132
rect 1243 -14388 1249 -14132
rect 1203 -14400 1249 -14388
rect 1381 -14132 1427 -14120
rect 1381 -14388 1387 -14132
rect 1421 -14388 1427 -14132
rect 1381 -14400 1427 -14388
rect 1559 -14132 1605 -14120
rect 1559 -14388 1565 -14132
rect 1599 -14388 1605 -14132
rect 1559 -14400 1605 -14388
rect 1737 -14132 1783 -14120
rect 1737 -14388 1743 -14132
rect 1777 -14388 1783 -14132
rect 1737 -14400 1783 -14388
rect 1915 -14132 1961 -14120
rect 1915 -14388 1921 -14132
rect 1955 -14388 1961 -14132
rect 1915 -14400 1961 -14388
rect 2093 -14132 2139 -14120
rect 2093 -14388 2099 -14132
rect 2133 -14388 2139 -14132
rect 2093 -14400 2139 -14388
rect 2271 -14132 2317 -14120
rect 2271 -14388 2277 -14132
rect 2311 -14388 2317 -14132
rect 2271 -14400 2317 -14388
rect 2449 -14132 2495 -14120
rect 2449 -14388 2455 -14132
rect 2489 -14388 2495 -14132
rect 2449 -14400 2495 -14388
rect 2627 -14132 2673 -14120
rect 2627 -14388 2633 -14132
rect 2667 -14388 2673 -14132
rect 2627 -14400 2673 -14388
rect 2805 -14132 2851 -14120
rect 2805 -14388 2811 -14132
rect 2845 -14388 2851 -14132
rect 2805 -14400 2851 -14388
rect 2983 -14132 3029 -14120
rect 2983 -14388 2989 -14132
rect 3023 -14388 3029 -14132
rect 2983 -14400 3029 -14388
rect 3161 -14132 3207 -14120
rect 3161 -14388 3167 -14132
rect 3201 -14388 3207 -14132
rect 3161 -14400 3207 -14388
rect 3339 -14132 3385 -14120
rect 3339 -14388 3345 -14132
rect 3379 -14388 3385 -14132
rect 3339 -14400 3385 -14388
rect 3517 -14132 3563 -14120
rect 3517 -14388 3523 -14132
rect 3557 -14388 3563 -14132
rect 3517 -14400 3563 -14388
rect 3695 -14132 3741 -14120
rect 3695 -14388 3701 -14132
rect 3735 -14388 3741 -14132
rect 3695 -14400 3741 -14388
rect 3873 -14132 3919 -14120
rect 3873 -14388 3879 -14132
rect 3913 -14388 3919 -14132
rect 3873 -14400 3919 -14388
rect 4051 -14132 4097 -14120
rect 4051 -14388 4057 -14132
rect 4091 -14388 4097 -14132
rect 4051 -14400 4097 -14388
rect -2173 -14441 -2139 -14400
rect -2105 -14438 -2029 -14432
rect -2105 -14441 -2089 -14438
rect -2173 -14472 -2089 -14441
rect -2045 -14441 -2029 -14438
rect -1995 -14441 -1961 -14400
rect -2045 -14472 -1961 -14441
rect -2173 -14475 -1961 -14472
rect -2105 -14488 -2029 -14475
rect -2325 -14596 -2315 -14543
rect -2262 -14596 -2252 -14543
rect -2105 -15045 -2029 -15032
rect -1995 -15045 -1961 -14475
rect -1927 -14438 -1851 -14432
rect -1927 -14472 -1911 -14438
rect -1867 -14472 -1851 -14438
rect -1927 -14488 -1851 -14472
rect -2176 -15048 -1961 -15045
rect -2176 -15079 -2089 -15048
rect -2176 -15120 -2142 -15079
rect -2105 -15082 -2089 -15079
rect -2045 -15079 -1961 -15048
rect -2045 -15082 -2029 -15079
rect -2105 -15088 -2029 -15082
rect -1995 -15120 -1961 -15079
rect -1927 -15048 -1851 -15032
rect -1927 -15082 -1911 -15048
rect -1867 -15082 -1851 -15048
rect -1927 -15088 -1851 -15082
rect -1817 -15120 -1783 -14400
rect -1749 -14438 -1673 -14432
rect -1749 -14472 -1733 -14438
rect -1689 -14472 -1673 -14438
rect -1749 -14488 -1673 -14472
rect -1749 -15048 -1673 -15032
rect -1749 -15082 -1733 -15048
rect -1689 -15082 -1673 -15048
rect -1749 -15088 -1673 -15082
rect -1639 -15120 -1605 -14400
rect -1571 -14438 -1495 -14432
rect -1571 -14472 -1555 -14438
rect -1511 -14472 -1495 -14438
rect -1571 -14488 -1495 -14472
rect -1571 -15048 -1495 -15032
rect -1571 -15082 -1555 -15048
rect -1511 -15082 -1495 -15048
rect -1571 -15088 -1495 -15082
rect -1461 -15120 -1427 -14400
rect -1393 -14438 -1317 -14432
rect -1393 -14472 -1377 -14438
rect -1333 -14472 -1317 -14438
rect -1393 -14488 -1317 -14472
rect -1371 -14543 -1337 -14488
rect -1391 -14596 -1381 -14543
rect -1328 -14596 -1318 -14543
rect -1371 -15032 -1337 -14596
rect -1393 -15048 -1317 -15032
rect -1393 -15082 -1377 -15048
rect -1333 -15082 -1317 -15048
rect -1393 -15088 -1317 -15082
rect -1283 -15120 -1249 -14400
rect -1215 -14438 -1139 -14432
rect -1215 -14472 -1199 -14438
rect -1155 -14472 -1139 -14438
rect -1215 -14488 -1139 -14472
rect -1194 -14543 -1160 -14488
rect -1214 -14596 -1204 -14543
rect -1151 -14596 -1141 -14543
rect -1215 -15048 -1139 -15032
rect -1215 -15082 -1199 -15048
rect -1155 -15082 -1139 -15048
rect -1215 -15088 -1139 -15082
rect -1104 -15120 -1070 -14400
rect -1037 -14438 -961 -14432
rect -1037 -14472 -1021 -14438
rect -977 -14472 -961 -14438
rect -1037 -14488 -961 -14472
rect -1016 -14543 -982 -14488
rect -1036 -14596 -1026 -14543
rect -973 -14596 -963 -14543
rect -1037 -15048 -961 -15032
rect -1037 -15082 -1021 -15048
rect -977 -15082 -961 -15048
rect -1037 -15088 -961 -15082
rect -927 -15120 -893 -14400
rect -859 -14438 -783 -14432
rect -859 -14472 -843 -14438
rect -799 -14472 -783 -14438
rect -859 -14488 -783 -14472
rect -838 -14543 -804 -14488
rect -858 -14596 -848 -14543
rect -795 -14596 -785 -14543
rect -857 -14979 -847 -14926
rect -794 -14979 -784 -14926
rect -838 -15032 -804 -14979
rect -859 -15048 -783 -15032
rect -859 -15082 -843 -15048
rect -799 -15082 -783 -15048
rect -859 -15088 -783 -15082
rect -749 -15120 -715 -14400
rect -681 -14438 -605 -14432
rect -681 -14472 -665 -14438
rect -621 -14472 -605 -14438
rect -681 -14488 -605 -14472
rect -659 -14543 -625 -14488
rect -679 -14596 -669 -14543
rect -616 -14596 -606 -14543
rect -679 -14979 -669 -14926
rect -616 -14979 -606 -14926
rect -660 -15032 -626 -14979
rect -681 -15048 -605 -15032
rect -681 -15082 -665 -15048
rect -621 -15082 -605 -15048
rect -681 -15088 -605 -15082
rect -571 -15120 -537 -14400
rect -503 -14438 -427 -14432
rect -503 -14472 -487 -14438
rect -443 -14472 -427 -14438
rect -503 -14488 -427 -14472
rect -482 -14543 -448 -14488
rect -501 -14596 -491 -14543
rect -438 -14596 -428 -14543
rect -501 -14979 -491 -14926
rect -438 -14979 -428 -14926
rect -481 -15032 -447 -14979
rect -503 -15048 -427 -15032
rect -503 -15082 -487 -15048
rect -443 -15082 -427 -15048
rect -503 -15088 -427 -15082
rect -393 -15120 -359 -14400
rect -325 -14438 -249 -14432
rect -325 -14472 -309 -14438
rect -265 -14472 -249 -14438
rect -325 -14488 -249 -14472
rect -304 -14927 -270 -14488
rect -324 -14980 -314 -14927
rect -261 -14980 -251 -14927
rect -304 -15032 -270 -14980
rect -325 -15048 -249 -15032
rect -325 -15082 -309 -15048
rect -265 -15082 -249 -15048
rect -325 -15088 -249 -15082
rect -215 -15120 -181 -14400
rect -147 -14438 -71 -14432
rect -147 -14472 -131 -14438
rect -87 -14472 -71 -14438
rect -147 -14488 -71 -14472
rect -126 -14926 -92 -14488
rect -147 -14979 -137 -14926
rect -84 -14979 -74 -14926
rect -126 -15032 -92 -14979
rect -147 -15048 -71 -15032
rect -147 -15082 -131 -15048
rect -87 -15082 -71 -15048
rect -147 -15088 -71 -15082
rect -37 -15120 -3 -14400
rect 31 -14438 107 -14432
rect 31 -14472 47 -14438
rect 91 -14472 107 -14438
rect 31 -14488 107 -14472
rect 52 -14926 86 -14488
rect 33 -14979 43 -14926
rect 96 -14979 106 -14926
rect 52 -15032 86 -14979
rect 31 -15048 107 -15032
rect 31 -15082 47 -15048
rect 91 -15082 107 -15048
rect 31 -15088 107 -15082
rect 141 -15120 175 -14400
rect 209 -14438 285 -14432
rect 209 -14472 225 -14438
rect 269 -14472 285 -14438
rect 209 -14488 285 -14472
rect 209 -15048 285 -15032
rect 209 -15082 225 -15048
rect 269 -15082 285 -15048
rect 209 -15088 285 -15082
rect 319 -15120 353 -14400
rect 387 -14438 463 -14432
rect 387 -14472 403 -14438
rect 447 -14472 463 -14438
rect 387 -14488 463 -14472
rect 387 -15048 463 -15032
rect 387 -15082 403 -15048
rect 447 -15082 463 -15048
rect 387 -15088 463 -15082
rect 497 -15120 531 -14400
rect 565 -14438 641 -14432
rect 565 -14472 581 -14438
rect 625 -14472 641 -14438
rect 565 -14488 641 -14472
rect 565 -15048 641 -15032
rect 565 -15082 581 -15048
rect 625 -15082 641 -15048
rect 565 -15088 641 -15082
rect 675 -15120 709 -14400
rect 743 -14438 819 -14432
rect 743 -14472 759 -14438
rect 803 -14472 819 -14438
rect 743 -14488 819 -14472
rect 921 -14438 997 -14432
rect 921 -14472 937 -14438
rect 981 -14472 997 -14438
rect 921 -14488 997 -14472
rect 743 -15048 819 -15032
rect 743 -15082 759 -15048
rect 803 -15082 819 -15048
rect 743 -15088 819 -15082
rect 921 -15048 997 -15032
rect 921 -15082 937 -15048
rect 981 -15082 997 -15048
rect 921 -15088 997 -15082
rect 1031 -15120 1065 -14400
rect 1099 -14438 1175 -14432
rect 1099 -14472 1115 -14438
rect 1159 -14472 1175 -14438
rect 1099 -14488 1175 -14472
rect 1099 -15048 1175 -15032
rect 1099 -15082 1115 -15048
rect 1159 -15082 1175 -15048
rect 1099 -15088 1175 -15082
rect 1209 -15120 1243 -14400
rect 1277 -14438 1353 -14432
rect 1277 -14472 1293 -14438
rect 1337 -14472 1353 -14438
rect 1277 -14488 1353 -14472
rect 1298 -14543 1332 -14488
rect 1278 -14596 1288 -14543
rect 1341 -14596 1351 -14543
rect 1279 -14980 1289 -14927
rect 1342 -14980 1352 -14927
rect 1298 -15032 1332 -14980
rect 1277 -15048 1353 -15032
rect 1277 -15082 1293 -15048
rect 1337 -15082 1353 -15048
rect 1277 -15088 1353 -15082
rect 1387 -15120 1421 -14400
rect 1455 -14438 1531 -14432
rect 1455 -14472 1471 -14438
rect 1515 -14472 1531 -14438
rect 1455 -14488 1531 -14472
rect 1477 -14543 1511 -14488
rect 1456 -14596 1466 -14543
rect 1519 -14596 1529 -14543
rect 1457 -14979 1467 -14926
rect 1520 -14979 1530 -14926
rect 1476 -15032 1510 -14979
rect 1455 -15048 1531 -15032
rect 1455 -15082 1471 -15048
rect 1515 -15082 1531 -15048
rect 1455 -15088 1531 -15082
rect 1565 -15120 1599 -14400
rect 1633 -14438 1709 -14432
rect 1633 -14472 1649 -14438
rect 1693 -14472 1709 -14438
rect 1633 -14488 1709 -14472
rect 1654 -14543 1688 -14488
rect 1634 -14596 1644 -14543
rect 1697 -14596 1707 -14543
rect 1634 -14979 1644 -14926
rect 1697 -14979 1707 -14926
rect 1654 -15032 1688 -14979
rect 1633 -15048 1709 -15032
rect 1633 -15082 1649 -15048
rect 1693 -15082 1709 -15048
rect 1633 -15088 1709 -15082
rect 1744 -15120 1778 -14400
rect 1811 -14438 1887 -14432
rect 1811 -14472 1827 -14438
rect 1871 -14472 1887 -14438
rect 1811 -14488 1887 -14472
rect 1832 -14542 1866 -14488
rect 1813 -14595 1823 -14542
rect 1876 -14595 1886 -14542
rect 1812 -14979 1822 -14926
rect 1875 -14979 1885 -14926
rect 1833 -15032 1867 -14979
rect 1811 -15048 1887 -15032
rect 1811 -15082 1827 -15048
rect 1871 -15082 1887 -15048
rect 1811 -15088 1887 -15082
rect 1921 -15120 1955 -14400
rect 1989 -14438 2065 -14432
rect 1989 -14472 2005 -14438
rect 2049 -14472 2065 -14438
rect 1989 -14488 2065 -14472
rect 2010 -14543 2044 -14488
rect 1990 -14596 2000 -14543
rect 2053 -14596 2063 -14543
rect 1989 -14979 1999 -14926
rect 2052 -14979 2062 -14926
rect 2010 -15032 2044 -14979
rect 1989 -15048 2065 -15032
rect 1989 -15082 2005 -15048
rect 2049 -15082 2065 -15048
rect 1989 -15088 2065 -15082
rect 2100 -15120 2134 -14400
rect 2167 -14438 2243 -14432
rect 2167 -14472 2183 -14438
rect 2227 -14472 2243 -14438
rect 2167 -14488 2243 -14472
rect 2188 -14543 2222 -14488
rect 2168 -14596 2178 -14543
rect 2231 -14596 2241 -14543
rect 2170 -14979 2180 -14926
rect 2233 -14979 2243 -14926
rect 2189 -15032 2223 -14979
rect 2167 -15048 2243 -15032
rect 2167 -15082 2183 -15048
rect 2227 -15082 2243 -15048
rect 2167 -15088 2243 -15082
rect 2277 -15120 2311 -14400
rect 2345 -14438 2421 -14432
rect 2345 -14472 2361 -14438
rect 2405 -14472 2421 -14438
rect 2345 -14488 2421 -14472
rect 2345 -15048 2421 -15032
rect 2345 -15082 2361 -15048
rect 2405 -15082 2421 -15048
rect 2345 -15088 2421 -15082
rect 2455 -15120 2489 -14400
rect 2523 -14438 2599 -14432
rect 2523 -14472 2539 -14438
rect 2583 -14472 2599 -14438
rect 2523 -14488 2599 -14472
rect 2523 -15048 2599 -15032
rect 2523 -15082 2539 -15048
rect 2583 -15082 2599 -15048
rect 2523 -15088 2599 -15082
rect 2633 -15120 2667 -14400
rect 2701 -14438 2777 -14432
rect 2701 -14472 2717 -14438
rect 2761 -14472 2777 -14438
rect 2701 -14488 2777 -14472
rect 2701 -15048 2777 -15032
rect 2701 -15082 2717 -15048
rect 2761 -15082 2777 -15048
rect 2701 -15088 2777 -15082
rect 2811 -15120 2845 -14400
rect 2879 -14438 2955 -14432
rect 2879 -14472 2895 -14438
rect 2939 -14472 2955 -14438
rect 2879 -14488 2955 -14472
rect 2879 -15048 2955 -15032
rect 2879 -15082 2895 -15048
rect 2939 -15082 2955 -15048
rect 2879 -15088 2955 -15082
rect 2989 -15120 3023 -14400
rect 3057 -14438 3133 -14432
rect 3057 -14472 3073 -14438
rect 3117 -14472 3133 -14438
rect 3057 -14488 3133 -14472
rect 3057 -15048 3133 -15032
rect 3057 -15082 3073 -15048
rect 3117 -15082 3133 -15048
rect 3057 -15088 3133 -15082
rect 3167 -15120 3201 -14400
rect 3235 -14438 3311 -14432
rect 3235 -14472 3251 -14438
rect 3295 -14472 3311 -14438
rect 3235 -14488 3311 -14472
rect 3236 -14597 3246 -14544
rect 3299 -14597 3309 -14544
rect 3256 -15032 3290 -14597
rect 3235 -15048 3311 -15032
rect 3235 -15082 3251 -15048
rect 3295 -15082 3311 -15048
rect 3235 -15088 3311 -15082
rect 3345 -15120 3379 -14400
rect 3413 -14438 3489 -14432
rect 3413 -14472 3429 -14438
rect 3473 -14472 3489 -14438
rect 3413 -14488 3489 -14472
rect 3434 -14543 3468 -14488
rect 3414 -14596 3424 -14543
rect 3477 -14596 3487 -14543
rect 3415 -14979 3425 -14926
rect 3478 -14979 3488 -14926
rect 3434 -15032 3468 -14979
rect 3413 -15048 3489 -15032
rect 3413 -15082 3429 -15048
rect 3473 -15082 3489 -15048
rect 3413 -15088 3489 -15082
rect 3524 -15120 3558 -14400
rect 3591 -14438 3667 -14432
rect 3591 -14472 3607 -14438
rect 3651 -14472 3667 -14438
rect 3591 -14488 3667 -14472
rect 3612 -14543 3646 -14488
rect 3592 -14596 3602 -14543
rect 3655 -14596 3665 -14543
rect 3593 -14979 3603 -14926
rect 3656 -14979 3666 -14926
rect 3612 -15032 3646 -14979
rect 3591 -15048 3667 -15032
rect 3591 -15082 3607 -15048
rect 3651 -15082 3667 -15048
rect 3591 -15088 3667 -15082
rect 3701 -15120 3735 -14400
rect 3769 -14438 3845 -14432
rect 3769 -14472 3785 -14438
rect 3829 -14472 3845 -14438
rect 3769 -14488 3845 -14472
rect 3879 -14439 3913 -14400
rect 3947 -14438 4023 -14432
rect 3947 -14439 3963 -14438
rect 3879 -14472 3963 -14439
rect 4007 -14439 4023 -14438
rect 4057 -14439 4091 -14400
rect 4007 -14472 4091 -14439
rect 3879 -14473 4091 -14472
rect 3791 -14543 3825 -14488
rect 3771 -14596 3781 -14543
rect 3834 -14596 3844 -14543
rect 3770 -14979 3780 -14926
rect 3833 -14979 3843 -14926
rect 3790 -15032 3824 -14979
rect 3769 -15048 3845 -15032
rect 3769 -15082 3785 -15048
rect 3829 -15082 3845 -15048
rect 3769 -15088 3845 -15082
rect 3879 -15047 3913 -14473
rect 3947 -14488 4023 -14473
rect 4905 -14545 4958 -7905
rect 5037 -13296 5090 -7903
rect 5174 -7908 5184 -7855
rect 5237 -7908 5247 -7855
rect 5327 -7903 5337 -7850
rect 5390 -7903 5400 -7850
rect 5185 -8635 5237 -7908
rect 5175 -8687 5185 -8635
rect 5237 -8687 5247 -8635
rect 5337 -9925 5390 -7903
rect 11647 -8716 11681 -8715
rect 6690 -8760 6815 -8726
rect 6580 -8810 6656 -8794
rect 6580 -8844 6596 -8810
rect 6640 -8844 6656 -8810
rect 6580 -8850 6656 -8844
rect 6690 -8882 6724 -8760
rect 6781 -8794 6815 -8760
rect 11044 -8769 11054 -8716
rect 11107 -8769 11117 -8716
rect 11335 -8769 11345 -8716
rect 11398 -8769 11408 -8716
rect 11628 -8769 11638 -8716
rect 11691 -8769 11701 -8716
rect 11922 -8769 11932 -8716
rect 11985 -8769 11995 -8716
rect 12212 -8769 12222 -8716
rect 12275 -8769 12285 -8716
rect 6758 -8810 6834 -8794
rect 6758 -8844 6774 -8810
rect 6818 -8844 6834 -8810
rect 6758 -8850 6834 -8844
rect 6936 -8810 7012 -8794
rect 6936 -8844 6952 -8810
rect 6996 -8844 7012 -8810
rect 6936 -8850 7012 -8844
rect 7114 -8810 7190 -8794
rect 7114 -8844 7130 -8810
rect 7174 -8844 7190 -8810
rect 7114 -8850 7190 -8844
rect 7292 -8810 7368 -8794
rect 7292 -8844 7308 -8810
rect 7352 -8844 7368 -8810
rect 7292 -8850 7368 -8844
rect 7470 -8810 7546 -8794
rect 7470 -8844 7486 -8810
rect 7530 -8844 7546 -8810
rect 7470 -8850 7546 -8844
rect 7648 -8810 7724 -8794
rect 7648 -8844 7664 -8810
rect 7708 -8844 7724 -8810
rect 7648 -8850 7724 -8844
rect 7826 -8810 7902 -8794
rect 7826 -8844 7842 -8810
rect 7886 -8844 7902 -8810
rect 7826 -8850 7902 -8844
rect 8004 -8810 8080 -8794
rect 8004 -8844 8020 -8810
rect 8064 -8844 8080 -8810
rect 8004 -8850 8080 -8844
rect 8182 -8810 8258 -8794
rect 8182 -8844 8198 -8810
rect 8242 -8844 8258 -8810
rect 8182 -8850 8258 -8844
rect 8360 -8810 8436 -8794
rect 8360 -8844 8376 -8810
rect 8420 -8844 8436 -8810
rect 8360 -8850 8436 -8844
rect 8538 -8810 8614 -8794
rect 8538 -8844 8554 -8810
rect 8598 -8844 8614 -8810
rect 8538 -8850 8614 -8844
rect 8716 -8810 8792 -8794
rect 8716 -8844 8732 -8810
rect 8776 -8844 8792 -8810
rect 8716 -8850 8792 -8844
rect 8894 -8810 8970 -8794
rect 9072 -8808 9148 -8794
rect 9250 -8808 9326 -8794
rect 8894 -8844 8910 -8810
rect 8954 -8844 8970 -8810
rect 8894 -8850 8970 -8844
rect 9004 -8810 9395 -8808
rect 9004 -8842 9088 -8810
rect 9004 -8882 9038 -8842
rect 9072 -8844 9088 -8842
rect 9132 -8842 9266 -8810
rect 9132 -8844 9148 -8842
rect 9072 -8850 9148 -8844
rect 9183 -8882 9217 -8842
rect 9250 -8844 9266 -8842
rect 9310 -8842 9395 -8810
rect 9310 -8844 9326 -8842
rect 9250 -8850 9326 -8844
rect 9361 -8882 9395 -8842
rect 10840 -8840 10916 -8824
rect 10840 -8874 10856 -8840
rect 10900 -8874 10916 -8840
rect 10840 -8880 10916 -8874
rect 6506 -8894 6552 -8882
rect 6506 -9150 6512 -8894
rect 6546 -9150 6552 -8894
rect 6506 -9162 6552 -9150
rect 6684 -8894 6730 -8882
rect 6684 -9150 6690 -8894
rect 6724 -9150 6730 -8894
rect 6684 -9162 6730 -9150
rect 6862 -8894 6908 -8882
rect 6862 -9150 6868 -8894
rect 6902 -9150 6908 -8894
rect 6862 -9162 6908 -9150
rect 7040 -8894 7086 -8882
rect 7040 -9150 7046 -8894
rect 7080 -9150 7086 -8894
rect 7040 -9162 7086 -9150
rect 7218 -8894 7264 -8882
rect 7218 -9150 7224 -8894
rect 7258 -9150 7264 -8894
rect 7218 -9162 7264 -9150
rect 7396 -8894 7442 -8882
rect 7396 -9150 7402 -8894
rect 7436 -9150 7442 -8894
rect 7396 -9162 7442 -9150
rect 7574 -8894 7620 -8882
rect 7574 -9150 7580 -8894
rect 7614 -9150 7620 -8894
rect 7574 -9162 7620 -9150
rect 7752 -8894 7798 -8882
rect 7752 -9150 7758 -8894
rect 7792 -9150 7798 -8894
rect 7752 -9162 7798 -9150
rect 7930 -8894 7976 -8882
rect 7930 -9150 7936 -8894
rect 7970 -9150 7976 -8894
rect 7930 -9162 7976 -9150
rect 8108 -8894 8154 -8882
rect 8108 -9150 8114 -8894
rect 8148 -9150 8154 -8894
rect 8108 -9162 8154 -9150
rect 8286 -8894 8332 -8882
rect 8286 -9150 8292 -8894
rect 8326 -9150 8332 -8894
rect 8286 -9162 8332 -9150
rect 8464 -8894 8510 -8882
rect 8464 -9150 8470 -8894
rect 8504 -9150 8510 -8894
rect 8464 -9162 8510 -9150
rect 8642 -8894 8688 -8882
rect 8642 -9150 8648 -8894
rect 8682 -9150 8688 -8894
rect 8642 -9162 8688 -9150
rect 8820 -8894 8866 -8882
rect 8820 -9150 8826 -8894
rect 8860 -9150 8866 -8894
rect 8820 -9162 8866 -9150
rect 8998 -8894 9044 -8882
rect 8998 -9150 9004 -8894
rect 9038 -9150 9044 -8894
rect 8998 -9162 9044 -9150
rect 9176 -8894 9222 -8882
rect 9176 -9150 9182 -8894
rect 9216 -9150 9222 -8894
rect 9176 -9162 9222 -9150
rect 9354 -8894 9400 -8882
rect 9354 -9150 9360 -8894
rect 9394 -9150 9400 -8894
rect 11063 -8912 11097 -8769
rect 11132 -8840 11208 -8824
rect 11132 -8874 11148 -8840
rect 11192 -8874 11208 -8840
rect 11132 -8880 11208 -8874
rect 11354 -8912 11388 -8769
rect 11424 -8840 11500 -8824
rect 11424 -8874 11440 -8840
rect 11484 -8874 11500 -8840
rect 11424 -8880 11500 -8874
rect 11647 -8912 11681 -8769
rect 11716 -8840 11792 -8824
rect 11716 -8874 11732 -8840
rect 11776 -8874 11792 -8840
rect 11716 -8880 11792 -8874
rect 11941 -8912 11975 -8769
rect 12008 -8840 12084 -8824
rect 12008 -8874 12024 -8840
rect 12068 -8874 12084 -8840
rect 12008 -8880 12084 -8874
rect 12231 -8840 12265 -8769
rect 12300 -8840 12376 -8824
rect 12592 -8840 12668 -8824
rect 12231 -8874 12316 -8840
rect 12360 -8874 12608 -8840
rect 12652 -8874 12738 -8840
rect 12231 -8912 12265 -8874
rect 12300 -8880 12376 -8874
rect 12522 -8912 12556 -8874
rect 12592 -8880 12668 -8874
rect 12704 -8912 12738 -8874
rect 9354 -9162 9400 -9150
rect 10766 -8924 10812 -8912
rect 6513 -9201 6547 -9162
rect 6580 -9200 6656 -9194
rect 6580 -9201 6596 -9200
rect 6513 -9234 6596 -9201
rect 6640 -9201 6656 -9200
rect 6689 -9201 6723 -9162
rect 6640 -9234 6723 -9201
rect 6513 -9235 6723 -9234
rect 6758 -9200 6834 -9194
rect 6758 -9234 6774 -9200
rect 6818 -9234 6834 -9200
rect 6580 -9250 6656 -9235
rect 6758 -9250 6834 -9234
rect 6779 -9314 6813 -9250
rect 6759 -9367 6769 -9314
rect 6822 -9367 6832 -9314
rect 6669 -9598 6679 -9545
rect 6732 -9598 6742 -9545
rect 6580 -9710 6656 -9694
rect 6580 -9744 6596 -9710
rect 6640 -9744 6656 -9710
rect 6580 -9750 6656 -9744
rect 6690 -9782 6724 -9598
rect 6779 -9694 6813 -9367
rect 6758 -9710 6834 -9694
rect 6758 -9744 6774 -9710
rect 6818 -9744 6834 -9710
rect 6758 -9750 6834 -9744
rect 6868 -9782 6902 -9162
rect 6936 -9200 7012 -9194
rect 6936 -9234 6952 -9200
rect 6996 -9234 7012 -9200
rect 6936 -9250 7012 -9234
rect 6957 -9315 6991 -9250
rect 6937 -9368 6947 -9315
rect 7000 -9368 7010 -9315
rect 6957 -9621 6991 -9368
rect 7046 -9621 7080 -9162
rect 7114 -9200 7190 -9194
rect 7114 -9234 7130 -9200
rect 7174 -9234 7190 -9200
rect 7114 -9250 7190 -9234
rect 7135 -9315 7169 -9250
rect 7116 -9368 7126 -9315
rect 7179 -9368 7189 -9315
rect 6957 -9655 7080 -9621
rect 6957 -9694 6991 -9655
rect 6936 -9710 7012 -9694
rect 6936 -9744 6952 -9710
rect 6996 -9744 7012 -9710
rect 6936 -9750 7012 -9744
rect 7046 -9782 7080 -9655
rect 7135 -9694 7169 -9368
rect 7114 -9710 7190 -9694
rect 7114 -9744 7130 -9710
rect 7174 -9744 7190 -9710
rect 7114 -9750 7190 -9744
rect 7224 -9782 7258 -9162
rect 7292 -9200 7368 -9194
rect 7292 -9234 7308 -9200
rect 7352 -9234 7368 -9200
rect 7292 -9250 7368 -9234
rect 7313 -9313 7347 -9250
rect 7293 -9366 7303 -9313
rect 7356 -9366 7366 -9313
rect 7313 -9694 7347 -9366
rect 7292 -9710 7368 -9694
rect 7292 -9744 7308 -9710
rect 7352 -9744 7368 -9710
rect 7292 -9750 7368 -9744
rect 7402 -9782 7436 -9162
rect 7470 -9200 7546 -9194
rect 7470 -9234 7486 -9200
rect 7530 -9234 7546 -9200
rect 7470 -9250 7546 -9234
rect 7491 -9313 7525 -9250
rect 7472 -9366 7482 -9313
rect 7535 -9366 7545 -9313
rect 7491 -9694 7525 -9366
rect 7470 -9710 7546 -9694
rect 7470 -9744 7486 -9710
rect 7530 -9744 7546 -9710
rect 7470 -9750 7546 -9744
rect 7580 -9782 7614 -9162
rect 7648 -9200 7724 -9194
rect 7648 -9234 7664 -9200
rect 7708 -9234 7724 -9200
rect 7648 -9250 7724 -9234
rect 7669 -9315 7703 -9250
rect 7649 -9368 7659 -9315
rect 7712 -9368 7722 -9315
rect 7669 -9694 7703 -9368
rect 7648 -9710 7724 -9694
rect 7648 -9744 7664 -9710
rect 7708 -9744 7724 -9710
rect 7648 -9750 7724 -9744
rect 7758 -9782 7792 -9162
rect 7826 -9200 7902 -9194
rect 7826 -9234 7842 -9200
rect 7886 -9234 7902 -9200
rect 7826 -9250 7902 -9234
rect 7847 -9314 7881 -9250
rect 7827 -9367 7837 -9314
rect 7890 -9367 7900 -9314
rect 7847 -9694 7881 -9367
rect 7826 -9710 7902 -9694
rect 7826 -9744 7842 -9710
rect 7886 -9744 7902 -9710
rect 7826 -9750 7902 -9744
rect 7936 -9782 7970 -9162
rect 8004 -9200 8080 -9194
rect 8004 -9234 8020 -9200
rect 8064 -9234 8080 -9200
rect 8004 -9250 8080 -9234
rect 8025 -9315 8059 -9250
rect 8005 -9368 8015 -9315
rect 8068 -9368 8078 -9315
rect 8025 -9694 8059 -9368
rect 8004 -9710 8080 -9694
rect 8004 -9744 8020 -9710
rect 8064 -9744 8080 -9710
rect 8004 -9750 8080 -9744
rect 8113 -9782 8147 -9162
rect 8182 -9200 8258 -9194
rect 8182 -9234 8198 -9200
rect 8242 -9234 8258 -9200
rect 8182 -9250 8258 -9234
rect 8203 -9314 8237 -9250
rect 8184 -9367 8194 -9314
rect 8247 -9367 8257 -9314
rect 8203 -9694 8237 -9367
rect 8182 -9710 8258 -9694
rect 8182 -9744 8198 -9710
rect 8242 -9744 8258 -9710
rect 8182 -9750 8258 -9744
rect 8292 -9782 8326 -9162
rect 8360 -9200 8436 -9194
rect 8360 -9234 8376 -9200
rect 8420 -9234 8436 -9200
rect 8360 -9250 8436 -9234
rect 8381 -9314 8415 -9250
rect 8361 -9367 8371 -9314
rect 8424 -9367 8434 -9314
rect 8381 -9694 8415 -9367
rect 8360 -9710 8436 -9694
rect 8360 -9744 8376 -9710
rect 8420 -9744 8436 -9710
rect 8360 -9750 8436 -9744
rect 8470 -9782 8504 -9162
rect 8538 -9200 8614 -9194
rect 8538 -9234 8554 -9200
rect 8598 -9234 8614 -9200
rect 8538 -9250 8614 -9234
rect 8559 -9314 8593 -9250
rect 8539 -9367 8549 -9314
rect 8602 -9367 8612 -9314
rect 8559 -9694 8593 -9367
rect 8538 -9710 8614 -9694
rect 8538 -9744 8554 -9710
rect 8598 -9744 8614 -9710
rect 8538 -9750 8614 -9744
rect 8648 -9782 8682 -9162
rect 8716 -9200 8792 -9194
rect 8716 -9234 8732 -9200
rect 8776 -9234 8792 -9200
rect 8716 -9250 8792 -9234
rect 8737 -9315 8771 -9250
rect 8717 -9368 8727 -9315
rect 8780 -9368 8790 -9315
rect 8737 -9694 8771 -9368
rect 8716 -9710 8792 -9694
rect 8716 -9744 8732 -9710
rect 8776 -9744 8792 -9710
rect 8716 -9750 8792 -9744
rect 8826 -9782 8860 -9162
rect 8894 -9200 8970 -9194
rect 8894 -9234 8910 -9200
rect 8954 -9234 8970 -9200
rect 8894 -9250 8970 -9234
rect 8915 -9314 8949 -9250
rect 8896 -9367 8906 -9314
rect 8959 -9367 8969 -9314
rect 8915 -9694 8949 -9367
rect 8894 -9710 8970 -9694
rect 8894 -9744 8910 -9710
rect 8954 -9744 8970 -9710
rect 8894 -9750 8970 -9744
rect 9004 -9709 9038 -9162
rect 10766 -9180 10772 -8924
rect 10806 -9180 10812 -8924
rect 9970 -9191 10172 -9185
rect 9072 -9200 9148 -9194
rect 9072 -9234 9088 -9200
rect 9132 -9234 9148 -9200
rect 9072 -9250 9148 -9234
rect 9250 -9200 9326 -9194
rect 9250 -9234 9266 -9200
rect 9310 -9234 9326 -9200
rect 9250 -9250 9326 -9234
rect 9970 -9369 9982 -9191
rect 10160 -9369 10172 -9191
rect 10766 -9192 10812 -9180
rect 10944 -8924 10990 -8912
rect 10944 -9180 10950 -8924
rect 10984 -9145 10990 -8924
rect 11058 -8924 11104 -8912
rect 11058 -9145 11064 -8924
rect 10984 -9179 11064 -9145
rect 10984 -9180 10990 -9179
rect 10944 -9192 10990 -9180
rect 11058 -9180 11064 -9179
rect 11098 -9180 11104 -8924
rect 11058 -9192 11104 -9180
rect 11236 -8924 11282 -8912
rect 11236 -9180 11242 -8924
rect 11276 -9180 11282 -8924
rect 11236 -9192 11282 -9180
rect 11350 -8924 11396 -8912
rect 11350 -9180 11356 -8924
rect 11390 -9180 11396 -8924
rect 11350 -9192 11396 -9180
rect 11528 -8924 11574 -8912
rect 11528 -9180 11534 -8924
rect 11568 -9180 11574 -8924
rect 11528 -9192 11574 -9180
rect 11642 -8924 11688 -8912
rect 11642 -9180 11648 -8924
rect 11682 -9180 11688 -8924
rect 11642 -9192 11688 -9180
rect 11820 -8924 11866 -8912
rect 11820 -9180 11826 -8924
rect 11860 -9180 11866 -8924
rect 11820 -9192 11866 -9180
rect 11934 -8924 11980 -8912
rect 11934 -9180 11940 -8924
rect 11974 -9180 11980 -8924
rect 11934 -9192 11980 -9180
rect 12112 -8924 12158 -8912
rect 12112 -9180 12118 -8924
rect 12152 -9180 12158 -8924
rect 12112 -9192 12158 -9180
rect 12226 -8924 12272 -8912
rect 12226 -9180 12232 -8924
rect 12266 -9180 12272 -8924
rect 12226 -9192 12272 -9180
rect 12404 -8924 12450 -8912
rect 12404 -9180 12410 -8924
rect 12444 -9180 12450 -8924
rect 12404 -9192 12450 -9180
rect 12518 -8924 12564 -8912
rect 12518 -9180 12524 -8924
rect 12558 -9180 12564 -8924
rect 12518 -9192 12564 -9180
rect 12696 -8924 12742 -8912
rect 12696 -9180 12702 -8924
rect 12736 -9180 12742 -8924
rect 12696 -9192 12742 -9180
rect 10772 -9230 10806 -9192
rect 10840 -9230 10916 -9224
rect 10950 -9230 10984 -9192
rect 10772 -9264 10856 -9230
rect 10900 -9264 10984 -9230
rect 10840 -9280 10916 -9264
rect 9970 -9375 10172 -9369
rect 10861 -9594 10895 -9280
rect 11063 -9387 11097 -9192
rect 11132 -9230 11208 -9224
rect 11132 -9264 11148 -9230
rect 11192 -9264 11208 -9230
rect 11132 -9280 11208 -9264
rect 11154 -9374 11188 -9280
rect 11134 -9387 11144 -9374
rect 11063 -9421 11144 -9387
rect 11134 -9427 11144 -9421
rect 11197 -9427 11207 -9374
rect 11154 -9594 11188 -9427
rect 10840 -9610 10916 -9594
rect 10840 -9644 10856 -9610
rect 10900 -9644 10916 -9610
rect 10840 -9650 10916 -9644
rect 11132 -9610 11208 -9594
rect 11132 -9644 11148 -9610
rect 11192 -9644 11208 -9610
rect 11132 -9650 11208 -9644
rect 11242 -9682 11276 -9192
rect 11424 -9230 11500 -9224
rect 11424 -9264 11440 -9230
rect 11484 -9264 11500 -9230
rect 11424 -9280 11500 -9264
rect 11445 -9375 11479 -9280
rect 11426 -9428 11436 -9375
rect 11489 -9428 11499 -9375
rect 11445 -9594 11479 -9428
rect 11424 -9610 11500 -9594
rect 11424 -9644 11440 -9610
rect 11484 -9644 11500 -9610
rect 11424 -9650 11500 -9644
rect 11534 -9682 11568 -9192
rect 11716 -9230 11792 -9224
rect 11716 -9264 11732 -9230
rect 11776 -9264 11792 -9230
rect 11716 -9280 11792 -9264
rect 11738 -9375 11772 -9280
rect 11718 -9428 11728 -9375
rect 11781 -9428 11791 -9375
rect 11738 -9594 11772 -9428
rect 11716 -9610 11792 -9594
rect 11716 -9644 11732 -9610
rect 11776 -9644 11792 -9610
rect 11716 -9650 11792 -9644
rect 11825 -9682 11859 -9192
rect 12008 -9230 12084 -9224
rect 12008 -9264 12024 -9230
rect 12068 -9264 12084 -9230
rect 12008 -9280 12084 -9264
rect 12030 -9376 12064 -9280
rect 12010 -9429 12020 -9376
rect 12073 -9429 12083 -9376
rect 12030 -9594 12064 -9429
rect 12008 -9610 12084 -9594
rect 12008 -9644 12024 -9610
rect 12068 -9644 12084 -9610
rect 12008 -9650 12084 -9644
rect 12118 -9682 12152 -9192
rect 12300 -9230 12376 -9224
rect 12300 -9264 12316 -9230
rect 12360 -9264 12376 -9230
rect 12300 -9280 12376 -9264
rect 12321 -9375 12355 -9280
rect 12302 -9428 12312 -9375
rect 12365 -9428 12375 -9375
rect 12321 -9594 12355 -9428
rect 12300 -9610 12376 -9594
rect 12300 -9644 12316 -9610
rect 12360 -9644 12376 -9610
rect 12300 -9650 12376 -9644
rect 12410 -9682 12444 -9192
rect 12592 -9230 12668 -9224
rect 12592 -9264 12608 -9230
rect 12652 -9264 12668 -9230
rect 12592 -9280 12668 -9264
rect 12613 -9594 12647 -9280
rect 12592 -9610 12668 -9594
rect 12525 -9644 12608 -9610
rect 12652 -9644 12736 -9610
rect 12525 -9682 12559 -9644
rect 12592 -9650 12668 -9644
rect 12702 -9682 12736 -9644
rect 10766 -9694 10812 -9682
rect 9072 -9709 9148 -9694
rect 9250 -9709 9326 -9694
rect 9004 -9710 9394 -9709
rect 9004 -9743 9088 -9710
rect 9004 -9782 9038 -9743
rect 9072 -9744 9088 -9743
rect 9132 -9743 9266 -9710
rect 9132 -9744 9148 -9743
rect 9072 -9750 9148 -9744
rect 9182 -9782 9216 -9743
rect 9250 -9744 9266 -9743
rect 9310 -9743 9394 -9710
rect 9310 -9744 9326 -9743
rect 9250 -9750 9326 -9744
rect 9360 -9782 9394 -9743
rect 6506 -9794 6552 -9782
rect 5327 -9978 5337 -9925
rect 5390 -9978 5400 -9925
rect 6506 -10050 6512 -9794
rect 6546 -10050 6552 -9794
rect 6506 -10062 6552 -10050
rect 6684 -9794 6730 -9782
rect 6684 -10050 6690 -9794
rect 6724 -10050 6730 -9794
rect 6684 -10062 6730 -10050
rect 6862 -9794 6908 -9782
rect 6862 -10050 6868 -9794
rect 6902 -10050 6908 -9794
rect 6862 -10062 6908 -10050
rect 7040 -9794 7086 -9782
rect 7040 -10050 7046 -9794
rect 7080 -10050 7086 -9794
rect 7040 -10062 7086 -10050
rect 7218 -9794 7264 -9782
rect 7218 -10050 7224 -9794
rect 7258 -10050 7264 -9794
rect 7218 -10062 7264 -10050
rect 7396 -9794 7442 -9782
rect 7396 -10050 7402 -9794
rect 7436 -10050 7442 -9794
rect 7396 -10062 7442 -10050
rect 7574 -9794 7620 -9782
rect 7574 -10050 7580 -9794
rect 7614 -10050 7620 -9794
rect 7574 -10062 7620 -10050
rect 7752 -9794 7798 -9782
rect 7752 -10050 7758 -9794
rect 7792 -10050 7798 -9794
rect 7752 -10062 7798 -10050
rect 7930 -9794 7976 -9782
rect 7930 -10050 7936 -9794
rect 7970 -10050 7976 -9794
rect 7930 -10062 7976 -10050
rect 8108 -9794 8154 -9782
rect 8108 -10050 8114 -9794
rect 8148 -10050 8154 -9794
rect 8108 -10062 8154 -10050
rect 8286 -9794 8332 -9782
rect 8286 -10050 8292 -9794
rect 8326 -10050 8332 -9794
rect 8286 -10062 8332 -10050
rect 8464 -9794 8510 -9782
rect 8464 -10050 8470 -9794
rect 8504 -10050 8510 -9794
rect 8464 -10062 8510 -10050
rect 8642 -9794 8688 -9782
rect 8642 -10050 8648 -9794
rect 8682 -10050 8688 -9794
rect 8642 -10062 8688 -10050
rect 8820 -9794 8866 -9782
rect 8820 -10050 8826 -9794
rect 8860 -10050 8866 -9794
rect 8820 -10062 8866 -10050
rect 8998 -9794 9044 -9782
rect 8998 -10050 9004 -9794
rect 9038 -10050 9044 -9794
rect 8998 -10062 9044 -10050
rect 9176 -9794 9222 -9782
rect 9176 -10050 9182 -9794
rect 9216 -10050 9222 -9794
rect 9176 -10062 9222 -10050
rect 9354 -9794 9400 -9782
rect 9354 -10050 9360 -9794
rect 9394 -10050 9400 -9794
rect 10766 -9950 10772 -9694
rect 10806 -9950 10812 -9694
rect 10766 -9962 10812 -9950
rect 10944 -9694 10990 -9682
rect 10944 -9950 10950 -9694
rect 10984 -9950 10990 -9694
rect 10944 -9962 10990 -9950
rect 11058 -9694 11104 -9682
rect 11058 -9950 11064 -9694
rect 11098 -9950 11104 -9694
rect 11058 -9962 11104 -9950
rect 11236 -9694 11282 -9682
rect 11236 -9950 11242 -9694
rect 11276 -9950 11282 -9694
rect 11236 -9962 11282 -9950
rect 11350 -9694 11396 -9682
rect 11350 -9950 11356 -9694
rect 11390 -9950 11396 -9694
rect 11350 -9962 11396 -9950
rect 11528 -9694 11574 -9682
rect 11528 -9950 11534 -9694
rect 11568 -9950 11574 -9694
rect 11528 -9962 11574 -9950
rect 11642 -9694 11688 -9682
rect 11642 -9950 11648 -9694
rect 11682 -9950 11688 -9694
rect 11642 -9962 11688 -9950
rect 11820 -9694 11866 -9682
rect 11820 -9950 11826 -9694
rect 11860 -9950 11866 -9694
rect 11820 -9962 11866 -9950
rect 11934 -9694 11980 -9682
rect 11934 -9950 11940 -9694
rect 11974 -9950 11980 -9694
rect 11934 -9962 11980 -9950
rect 12112 -9694 12158 -9682
rect 12112 -9950 12118 -9694
rect 12152 -9950 12158 -9694
rect 12112 -9962 12158 -9950
rect 12226 -9694 12272 -9682
rect 12226 -9950 12232 -9694
rect 12266 -9950 12272 -9694
rect 12226 -9962 12272 -9950
rect 12404 -9694 12450 -9682
rect 12404 -9950 12410 -9694
rect 12444 -9950 12450 -9694
rect 12404 -9962 12450 -9950
rect 12518 -9694 12564 -9682
rect 12518 -9950 12524 -9694
rect 12558 -9950 12564 -9694
rect 12518 -9962 12564 -9950
rect 12696 -9694 12742 -9682
rect 12696 -9950 12702 -9694
rect 12736 -9950 12742 -9694
rect 12696 -9962 12742 -9950
rect 10773 -10001 10807 -9962
rect 10840 -10000 10916 -9994
rect 10840 -10001 10856 -10000
rect 10773 -10034 10856 -10001
rect 10900 -10001 10916 -10000
rect 10951 -10001 10985 -9962
rect 10900 -10034 10985 -10001
rect 10773 -10035 10985 -10034
rect 10840 -10050 10916 -10035
rect 9354 -10062 9400 -10050
rect 6513 -10099 6547 -10062
rect 6580 -10099 6656 -10094
rect 6690 -10099 6724 -10062
rect 6513 -10100 6724 -10099
rect 6513 -10133 6596 -10100
rect 6580 -10134 6596 -10133
rect 6640 -10133 6724 -10100
rect 6640 -10134 6656 -10133
rect 6580 -10150 6656 -10134
rect 6690 -10313 6724 -10133
rect 6758 -10100 6834 -10094
rect 6758 -10134 6774 -10100
rect 6818 -10134 6834 -10100
rect 6758 -10150 6834 -10134
rect 6670 -10366 6680 -10313
rect 6733 -10366 6743 -10313
rect 6868 -10467 6902 -10062
rect 6936 -10100 7012 -10094
rect 6936 -10134 6952 -10100
rect 6996 -10134 7012 -10100
rect 6936 -10150 7012 -10134
rect 6848 -10520 6858 -10467
rect 6911 -10520 6921 -10467
rect 6580 -10610 6656 -10594
rect 6580 -10644 6596 -10610
rect 6640 -10644 6656 -10610
rect 6580 -10650 6656 -10644
rect 6758 -10610 6834 -10594
rect 6758 -10644 6774 -10610
rect 6818 -10644 6834 -10610
rect 6758 -10650 6834 -10644
rect 6868 -10682 6902 -10520
rect 6958 -10594 6992 -10150
rect 6936 -10610 7012 -10594
rect 6936 -10644 6952 -10610
rect 6996 -10644 7012 -10610
rect 6936 -10650 7012 -10644
rect 7046 -10682 7080 -10062
rect 7114 -10100 7190 -10094
rect 7114 -10134 7130 -10100
rect 7174 -10134 7190 -10100
rect 7114 -10150 7190 -10134
rect 7136 -10594 7170 -10150
rect 7224 -10466 7258 -10062
rect 7292 -10100 7368 -10094
rect 7292 -10134 7308 -10100
rect 7352 -10134 7368 -10100
rect 7292 -10150 7368 -10134
rect 7204 -10519 7214 -10466
rect 7267 -10519 7277 -10466
rect 7114 -10610 7190 -10594
rect 7114 -10644 7130 -10610
rect 7174 -10644 7190 -10610
rect 7114 -10650 7190 -10644
rect 7224 -10682 7258 -10519
rect 7313 -10594 7347 -10150
rect 7292 -10610 7368 -10594
rect 7292 -10644 7308 -10610
rect 7352 -10644 7368 -10610
rect 7292 -10650 7368 -10644
rect 7402 -10682 7436 -10062
rect 7470 -10100 7546 -10094
rect 7470 -10134 7486 -10100
rect 7530 -10134 7546 -10100
rect 7470 -10150 7546 -10134
rect 7492 -10594 7526 -10150
rect 7580 -10466 7614 -10062
rect 7648 -10100 7724 -10094
rect 7648 -10134 7664 -10100
rect 7708 -10134 7724 -10100
rect 7648 -10150 7724 -10134
rect 7561 -10519 7571 -10466
rect 7624 -10519 7634 -10466
rect 7470 -10610 7546 -10594
rect 7470 -10644 7486 -10610
rect 7530 -10644 7546 -10610
rect 7470 -10650 7546 -10644
rect 7580 -10682 7614 -10519
rect 7669 -10594 7703 -10150
rect 7648 -10610 7724 -10594
rect 7648 -10644 7664 -10610
rect 7708 -10644 7724 -10610
rect 7648 -10650 7724 -10644
rect 7758 -10682 7792 -10062
rect 7826 -10100 7902 -10094
rect 7826 -10134 7842 -10100
rect 7886 -10134 7902 -10100
rect 7826 -10150 7902 -10134
rect 7847 -10594 7881 -10150
rect 7936 -10466 7970 -10062
rect 8004 -10100 8080 -10094
rect 8004 -10134 8020 -10100
rect 8064 -10134 8080 -10100
rect 8004 -10150 8080 -10134
rect 7917 -10519 7927 -10466
rect 7980 -10519 7990 -10466
rect 7826 -10610 7902 -10594
rect 7826 -10644 7842 -10610
rect 7886 -10644 7902 -10610
rect 7826 -10650 7902 -10644
rect 7936 -10682 7970 -10519
rect 8025 -10594 8059 -10150
rect 8004 -10610 8080 -10594
rect 8004 -10644 8020 -10610
rect 8064 -10644 8080 -10610
rect 8004 -10650 8080 -10644
rect 8113 -10682 8147 -10062
rect 8182 -10100 8258 -10094
rect 8182 -10134 8198 -10100
rect 8242 -10134 8258 -10100
rect 8182 -10150 8258 -10134
rect 8203 -10594 8237 -10150
rect 8292 -10467 8326 -10062
rect 8360 -10100 8436 -10094
rect 8360 -10134 8376 -10100
rect 8420 -10134 8436 -10100
rect 8360 -10150 8436 -10134
rect 8273 -10520 8283 -10467
rect 8336 -10520 8346 -10467
rect 8182 -10610 8258 -10594
rect 8182 -10644 8198 -10610
rect 8242 -10644 8258 -10610
rect 8182 -10650 8258 -10644
rect 8292 -10682 8326 -10520
rect 8382 -10594 8416 -10150
rect 8360 -10610 8436 -10594
rect 8360 -10644 8376 -10610
rect 8420 -10644 8436 -10610
rect 8360 -10650 8436 -10644
rect 8470 -10682 8504 -10062
rect 8538 -10100 8614 -10094
rect 8538 -10134 8554 -10100
rect 8598 -10134 8614 -10100
rect 8538 -10150 8614 -10134
rect 8559 -10594 8593 -10150
rect 8648 -10466 8682 -10062
rect 8716 -10100 8792 -10094
rect 8716 -10134 8732 -10100
rect 8776 -10134 8792 -10100
rect 8716 -10150 8792 -10134
rect 8628 -10519 8638 -10466
rect 8691 -10519 8701 -10466
rect 8538 -10610 8614 -10594
rect 8538 -10644 8554 -10610
rect 8598 -10644 8614 -10610
rect 8538 -10650 8614 -10644
rect 8648 -10682 8682 -10519
rect 8737 -10594 8771 -10150
rect 8716 -10610 8792 -10594
rect 8716 -10644 8732 -10610
rect 8776 -10644 8792 -10610
rect 8716 -10650 8792 -10644
rect 8826 -10682 8860 -10062
rect 8894 -10100 8970 -10094
rect 8894 -10134 8910 -10100
rect 8954 -10134 8970 -10100
rect 8894 -10150 8970 -10134
rect 8915 -10594 8949 -10150
rect 9004 -10467 9038 -10062
rect 9072 -10100 9148 -10094
rect 9072 -10134 9088 -10100
rect 9132 -10134 9148 -10100
rect 9072 -10150 9148 -10134
rect 9250 -10100 9326 -10094
rect 9250 -10134 9266 -10100
rect 9310 -10134 9326 -10100
rect 9250 -10150 9326 -10134
rect 9161 -10367 9171 -10314
rect 9224 -10367 9234 -10314
rect 10862 -10364 10896 -10050
rect 8985 -10520 8995 -10467
rect 9048 -10520 9058 -10467
rect 8894 -10610 8970 -10594
rect 8894 -10644 8910 -10610
rect 8954 -10644 8970 -10610
rect 8894 -10650 8970 -10644
rect 9004 -10682 9038 -10520
rect 9072 -10610 9148 -10594
rect 9072 -10644 9088 -10610
rect 9132 -10644 9148 -10610
rect 9072 -10650 9148 -10644
rect 9181 -10614 9215 -10367
rect 10840 -10380 10916 -10364
rect 10772 -10414 10856 -10380
rect 10900 -10414 10986 -10380
rect 10772 -10452 10806 -10414
rect 10840 -10420 10916 -10414
rect 10952 -10452 10986 -10414
rect 11063 -10452 11097 -9962
rect 11132 -10000 11208 -9994
rect 11132 -10034 11148 -10000
rect 11192 -10034 11208 -10000
rect 11132 -10050 11208 -10034
rect 11153 -10364 11187 -10050
rect 11132 -10380 11208 -10364
rect 11132 -10414 11148 -10380
rect 11192 -10414 11208 -10380
rect 11132 -10420 11208 -10414
rect 11356 -10452 11390 -9962
rect 11424 -10000 11500 -9994
rect 11424 -10034 11440 -10000
rect 11484 -10034 11500 -10000
rect 11424 -10050 11500 -10034
rect 11446 -10364 11480 -10050
rect 11424 -10380 11500 -10364
rect 11424 -10414 11440 -10380
rect 11484 -10414 11500 -10380
rect 11424 -10420 11500 -10414
rect 11648 -10452 11682 -9962
rect 11716 -10000 11792 -9994
rect 11716 -10034 11732 -10000
rect 11776 -10034 11792 -10000
rect 11716 -10050 11792 -10034
rect 11737 -10364 11771 -10050
rect 11716 -10380 11792 -10364
rect 11716 -10414 11732 -10380
rect 11776 -10414 11792 -10380
rect 11716 -10420 11792 -10414
rect 11940 -10452 11974 -9962
rect 12008 -10000 12084 -9994
rect 12008 -10034 12024 -10000
rect 12068 -10034 12084 -10000
rect 12008 -10050 12084 -10034
rect 12028 -10364 12062 -10050
rect 12008 -10380 12084 -10364
rect 12008 -10414 12024 -10380
rect 12068 -10414 12084 -10380
rect 12008 -10420 12084 -10414
rect 12232 -10452 12266 -9962
rect 12300 -10000 12376 -9994
rect 12300 -10034 12316 -10000
rect 12360 -10034 12376 -10000
rect 12300 -10050 12376 -10034
rect 12592 -10000 12668 -9994
rect 12592 -10034 12608 -10000
rect 12652 -10034 12668 -10000
rect 12592 -10050 12668 -10034
rect 12320 -10364 12354 -10050
rect 12613 -10364 12647 -10050
rect 12300 -10380 12376 -10364
rect 12300 -10414 12316 -10380
rect 12360 -10414 12376 -10380
rect 12300 -10420 12376 -10414
rect 12592 -10380 12668 -10364
rect 12592 -10414 12608 -10380
rect 12652 -10414 12668 -10380
rect 12592 -10420 12668 -10414
rect 10766 -10464 10812 -10452
rect 9250 -10610 9326 -10594
rect 9250 -10614 9266 -10610
rect 9181 -10644 9266 -10614
rect 9310 -10614 9326 -10610
rect 9310 -10644 9393 -10614
rect 9181 -10648 9393 -10644
rect 9181 -10682 9215 -10648
rect 9250 -10650 9326 -10648
rect 9359 -10682 9393 -10648
rect 6506 -10694 6552 -10682
rect 6506 -10950 6512 -10694
rect 6546 -10950 6552 -10694
rect 6506 -10962 6552 -10950
rect 6684 -10694 6730 -10682
rect 6684 -10950 6690 -10694
rect 6724 -10950 6730 -10694
rect 6684 -10962 6730 -10950
rect 6862 -10694 6908 -10682
rect 6862 -10950 6868 -10694
rect 6902 -10950 6908 -10694
rect 6862 -10962 6908 -10950
rect 7040 -10694 7086 -10682
rect 7040 -10950 7046 -10694
rect 7080 -10950 7086 -10694
rect 7040 -10962 7086 -10950
rect 7218 -10694 7264 -10682
rect 7218 -10950 7224 -10694
rect 7258 -10950 7264 -10694
rect 7218 -10962 7264 -10950
rect 7396 -10694 7442 -10682
rect 7396 -10950 7402 -10694
rect 7436 -10950 7442 -10694
rect 7396 -10962 7442 -10950
rect 7574 -10694 7620 -10682
rect 7574 -10950 7580 -10694
rect 7614 -10950 7620 -10694
rect 7574 -10962 7620 -10950
rect 7752 -10694 7798 -10682
rect 7752 -10950 7758 -10694
rect 7792 -10950 7798 -10694
rect 7752 -10962 7798 -10950
rect 7930 -10694 7976 -10682
rect 7930 -10950 7936 -10694
rect 7970 -10950 7976 -10694
rect 7930 -10962 7976 -10950
rect 8108 -10694 8154 -10682
rect 8108 -10950 8114 -10694
rect 8148 -10950 8154 -10694
rect 8108 -10962 8154 -10950
rect 8286 -10694 8332 -10682
rect 8286 -10950 8292 -10694
rect 8326 -10950 8332 -10694
rect 8286 -10962 8332 -10950
rect 8464 -10694 8510 -10682
rect 8464 -10950 8470 -10694
rect 8504 -10950 8510 -10694
rect 8464 -10962 8510 -10950
rect 8642 -10694 8688 -10682
rect 8642 -10950 8648 -10694
rect 8682 -10950 8688 -10694
rect 8642 -10962 8688 -10950
rect 8820 -10694 8866 -10682
rect 8820 -10950 8826 -10694
rect 8860 -10950 8866 -10694
rect 8820 -10962 8866 -10950
rect 8998 -10694 9044 -10682
rect 8998 -10950 9004 -10694
rect 9038 -10950 9044 -10694
rect 8998 -10962 9044 -10950
rect 9176 -10694 9222 -10682
rect 9176 -10950 9182 -10694
rect 9216 -10950 9222 -10694
rect 9176 -10962 9222 -10950
rect 9354 -10694 9400 -10682
rect 9354 -10950 9360 -10694
rect 9394 -10950 9400 -10694
rect 10766 -10720 10772 -10464
rect 10806 -10720 10812 -10464
rect 10766 -10732 10812 -10720
rect 10944 -10464 10990 -10452
rect 10944 -10720 10950 -10464
rect 10984 -10720 10990 -10464
rect 10944 -10732 10990 -10720
rect 11058 -10464 11104 -10452
rect 11058 -10720 11064 -10464
rect 11098 -10720 11104 -10464
rect 11058 -10732 11104 -10720
rect 11236 -10464 11282 -10452
rect 11236 -10720 11242 -10464
rect 11276 -10720 11282 -10464
rect 11236 -10732 11282 -10720
rect 11350 -10464 11396 -10452
rect 11350 -10720 11356 -10464
rect 11390 -10720 11396 -10464
rect 11350 -10732 11396 -10720
rect 11528 -10464 11574 -10452
rect 11528 -10720 11534 -10464
rect 11568 -10720 11574 -10464
rect 11528 -10732 11574 -10720
rect 11642 -10464 11688 -10452
rect 11642 -10720 11648 -10464
rect 11682 -10720 11688 -10464
rect 11642 -10732 11688 -10720
rect 11820 -10464 11866 -10452
rect 11820 -10720 11826 -10464
rect 11860 -10720 11866 -10464
rect 11820 -10732 11866 -10720
rect 11934 -10464 11980 -10452
rect 11934 -10720 11940 -10464
rect 11974 -10720 11980 -10464
rect 11934 -10732 11980 -10720
rect 12112 -10464 12158 -10452
rect 12112 -10720 12118 -10464
rect 12152 -10720 12158 -10464
rect 12112 -10732 12158 -10720
rect 12226 -10464 12272 -10452
rect 12226 -10720 12232 -10464
rect 12266 -10720 12272 -10464
rect 12226 -10732 12272 -10720
rect 12404 -10464 12450 -10452
rect 12404 -10720 12410 -10464
rect 12444 -10720 12450 -10464
rect 12404 -10732 12450 -10720
rect 12518 -10464 12564 -10452
rect 12518 -10720 12524 -10464
rect 12558 -10720 12564 -10464
rect 12518 -10732 12564 -10720
rect 12696 -10464 12742 -10452
rect 12696 -10720 12702 -10464
rect 12736 -10720 12742 -10464
rect 12696 -10732 12742 -10720
rect 10840 -10770 10916 -10764
rect 10840 -10804 10856 -10770
rect 10900 -10804 10916 -10770
rect 10840 -10820 10916 -10804
rect 11132 -10770 11208 -10764
rect 11132 -10804 11148 -10770
rect 11192 -10804 11208 -10770
rect 11132 -10820 11208 -10804
rect 9354 -10962 9400 -10950
rect 6510 -11003 6544 -10962
rect 6580 -11000 6656 -10994
rect 6580 -11003 6596 -11000
rect 6510 -11034 6596 -11003
rect 6640 -11003 6656 -11000
rect 6688 -11003 6722 -10962
rect 6758 -11000 6834 -10994
rect 6758 -11003 6774 -11000
rect 6640 -11034 6774 -11003
rect 6818 -11003 6834 -11000
rect 6868 -11003 6902 -10962
rect 6818 -11034 6902 -11003
rect 6510 -11037 6902 -11034
rect 6580 -11050 6656 -11037
rect 6758 -11050 6834 -11037
rect 5674 -11151 5876 -11145
rect 5674 -11329 5686 -11151
rect 5864 -11329 5876 -11151
rect 5674 -11335 5876 -11329
rect 6580 -11510 6656 -11494
rect 6580 -11544 6596 -11510
rect 6640 -11544 6656 -11510
rect 6580 -11550 6656 -11544
rect 6758 -11510 6834 -11494
rect 6758 -11544 6774 -11510
rect 6818 -11544 6834 -11510
rect 6758 -11550 6834 -11544
rect 6868 -11582 6902 -11037
rect 6936 -11000 7012 -10994
rect 6936 -11034 6952 -11000
rect 6996 -11034 7012 -11000
rect 6936 -11050 7012 -11034
rect 6958 -11494 6992 -11050
rect 7046 -11366 7080 -10962
rect 7114 -11000 7190 -10994
rect 7114 -11034 7130 -11000
rect 7174 -11034 7190 -11000
rect 7114 -11050 7190 -11034
rect 7027 -11419 7037 -11366
rect 7090 -11419 7100 -11366
rect 6936 -11510 7012 -11494
rect 6936 -11544 6952 -11510
rect 6996 -11544 7012 -11510
rect 6936 -11550 7012 -11544
rect 7046 -11582 7080 -11419
rect 7135 -11494 7169 -11050
rect 7114 -11510 7190 -11494
rect 7114 -11544 7130 -11510
rect 7174 -11544 7190 -11510
rect 7114 -11550 7190 -11544
rect 7224 -11582 7258 -10962
rect 7313 -10994 7347 -10993
rect 7292 -11000 7368 -10994
rect 7292 -11034 7308 -11000
rect 7352 -11034 7368 -11000
rect 7292 -11050 7368 -11034
rect 7313 -11494 7347 -11050
rect 7402 -11366 7436 -10962
rect 7491 -10994 7525 -10993
rect 7470 -11000 7546 -10994
rect 7470 -11034 7486 -11000
rect 7530 -11034 7546 -11000
rect 7470 -11050 7546 -11034
rect 7383 -11419 7393 -11366
rect 7446 -11419 7456 -11366
rect 7292 -11510 7368 -11494
rect 7292 -11544 7308 -11510
rect 7352 -11544 7368 -11510
rect 7292 -11550 7368 -11544
rect 7402 -11582 7436 -11419
rect 7491 -11494 7525 -11050
rect 7470 -11510 7546 -11494
rect 7470 -11544 7486 -11510
rect 7530 -11544 7546 -11510
rect 7470 -11550 7546 -11544
rect 7580 -11582 7614 -10962
rect 7669 -10994 7703 -10993
rect 7648 -11000 7724 -10994
rect 7648 -11034 7664 -11000
rect 7708 -11034 7724 -11000
rect 7648 -11050 7724 -11034
rect 7669 -11494 7703 -11050
rect 7758 -11367 7792 -10962
rect 7848 -10994 7882 -10993
rect 7826 -11000 7902 -10994
rect 7826 -11034 7842 -11000
rect 7886 -11034 7902 -11000
rect 7826 -11050 7902 -11034
rect 7738 -11420 7748 -11367
rect 7801 -11420 7811 -11367
rect 7648 -11510 7724 -11494
rect 7648 -11544 7664 -11510
rect 7708 -11544 7724 -11510
rect 7648 -11550 7724 -11544
rect 7758 -11582 7792 -11420
rect 7848 -11494 7882 -11050
rect 7826 -11510 7902 -11494
rect 7826 -11544 7842 -11510
rect 7886 -11544 7902 -11510
rect 7826 -11550 7902 -11544
rect 7936 -11582 7970 -10962
rect 8004 -11000 8080 -10994
rect 8004 -11034 8020 -11000
rect 8064 -11034 8080 -11000
rect 8004 -11050 8080 -11034
rect 8024 -11494 8058 -11050
rect 8113 -11366 8147 -10962
rect 8182 -11000 8258 -10994
rect 8182 -11034 8198 -11000
rect 8242 -11034 8258 -11000
rect 8182 -11050 8258 -11034
rect 8093 -11419 8103 -11366
rect 8156 -11419 8166 -11366
rect 8004 -11510 8080 -11494
rect 8004 -11544 8020 -11510
rect 8064 -11544 8080 -11510
rect 8004 -11550 8080 -11544
rect 8113 -11582 8147 -11419
rect 8203 -11494 8237 -11050
rect 8182 -11510 8258 -11494
rect 8182 -11544 8198 -11510
rect 8242 -11544 8258 -11510
rect 8182 -11550 8258 -11544
rect 8292 -11582 8326 -10962
rect 8360 -11000 8436 -10994
rect 8360 -11034 8376 -11000
rect 8420 -11034 8436 -11000
rect 8360 -11050 8436 -11034
rect 8381 -11494 8415 -11050
rect 8470 -11366 8504 -10962
rect 8538 -11000 8614 -10994
rect 8538 -11034 8554 -11000
rect 8598 -11034 8614 -11000
rect 8538 -11050 8614 -11034
rect 8451 -11419 8461 -11366
rect 8514 -11419 8524 -11366
rect 8360 -11510 8436 -11494
rect 8360 -11544 8376 -11510
rect 8420 -11544 8436 -11510
rect 8360 -11550 8436 -11544
rect 8470 -11582 8504 -11419
rect 8559 -11494 8593 -11050
rect 8538 -11510 8614 -11494
rect 8538 -11544 8554 -11510
rect 8598 -11544 8614 -11510
rect 8538 -11550 8614 -11544
rect 8648 -11582 8682 -10962
rect 8716 -11000 8792 -10994
rect 8716 -11034 8732 -11000
rect 8776 -11034 8792 -11000
rect 8716 -11050 8792 -11034
rect 8737 -11494 8771 -11050
rect 8826 -11366 8860 -10962
rect 8894 -11000 8970 -10994
rect 8894 -11034 8910 -11000
rect 8954 -11034 8970 -11000
rect 8894 -11050 8970 -11034
rect 8807 -11419 8817 -11366
rect 8870 -11419 8880 -11366
rect 8716 -11510 8792 -11494
rect 8716 -11544 8732 -11510
rect 8776 -11544 8792 -11510
rect 8716 -11550 8792 -11544
rect 8826 -11582 8860 -11419
rect 8915 -11494 8949 -11050
rect 8894 -11510 8970 -11494
rect 8894 -11544 8910 -11510
rect 8954 -11544 8970 -11510
rect 8894 -11550 8970 -11544
rect 9004 -11582 9038 -10962
rect 9072 -11000 9148 -10994
rect 9072 -11034 9088 -11000
rect 9132 -11034 9148 -11000
rect 9072 -11050 9148 -11034
rect 9250 -11000 9326 -10994
rect 9250 -11034 9266 -11000
rect 9310 -11034 9326 -11000
rect 9250 -11050 9326 -11034
rect 9093 -11494 9127 -11050
rect 10860 -11134 10894 -10820
rect 11152 -11134 11186 -10820
rect 10772 -11149 10806 -11148
rect 10840 -11149 10916 -11134
rect 10772 -11150 10986 -11149
rect 10772 -11183 10856 -11150
rect 9970 -11191 10172 -11185
rect 9970 -11369 9982 -11191
rect 10160 -11369 10172 -11191
rect 10772 -11222 10806 -11183
rect 10840 -11184 10856 -11183
rect 10900 -11183 10986 -11150
rect 10900 -11184 10916 -11183
rect 10840 -11190 10916 -11184
rect 10952 -11222 10986 -11183
rect 11132 -11150 11208 -11134
rect 11132 -11184 11148 -11150
rect 11192 -11184 11208 -11150
rect 11132 -11190 11208 -11184
rect 11244 -11222 11278 -10732
rect 11424 -10770 11500 -10764
rect 11424 -10804 11440 -10770
rect 11484 -10804 11500 -10770
rect 11424 -10820 11500 -10804
rect 11446 -11134 11480 -10820
rect 11424 -11150 11500 -11134
rect 11424 -11184 11440 -11150
rect 11484 -11184 11500 -11150
rect 11424 -11190 11500 -11184
rect 11534 -11222 11568 -10732
rect 11716 -10770 11792 -10764
rect 11716 -10804 11732 -10770
rect 11776 -10804 11792 -10770
rect 11716 -10820 11792 -10804
rect 11737 -11134 11771 -10820
rect 11716 -11150 11792 -11134
rect 11716 -11184 11732 -11150
rect 11776 -11184 11792 -11150
rect 11716 -11190 11792 -11184
rect 11826 -11222 11860 -10732
rect 12008 -10770 12084 -10764
rect 12008 -10804 12024 -10770
rect 12068 -10804 12084 -10770
rect 12008 -10820 12084 -10804
rect 12029 -11134 12063 -10820
rect 12008 -11150 12084 -11134
rect 12008 -11184 12024 -11150
rect 12068 -11184 12084 -11150
rect 12008 -11190 12084 -11184
rect 12118 -11222 12152 -10732
rect 12300 -10770 12376 -10764
rect 12300 -10804 12316 -10770
rect 12360 -10804 12376 -10770
rect 12300 -10820 12376 -10804
rect 12322 -11134 12356 -10820
rect 12300 -11150 12376 -11134
rect 12300 -11184 12316 -11150
rect 12360 -11184 12376 -11150
rect 12300 -11190 12376 -11184
rect 12410 -11222 12444 -10732
rect 12525 -10772 12559 -10732
rect 12592 -10770 12668 -10764
rect 12592 -10772 12608 -10770
rect 12525 -10804 12608 -10772
rect 12652 -10772 12668 -10770
rect 12700 -10772 12734 -10732
rect 12652 -10804 12734 -10772
rect 12525 -10806 12734 -10804
rect 12592 -10820 12668 -10806
rect 12613 -11134 12647 -10820
rect 12592 -11150 12668 -11134
rect 12592 -11184 12608 -11150
rect 12652 -11184 12668 -11150
rect 12592 -11190 12668 -11184
rect 9970 -11375 10172 -11369
rect 10766 -11234 10812 -11222
rect 10766 -11490 10772 -11234
rect 10806 -11490 10812 -11234
rect 9072 -11510 9148 -11494
rect 9250 -11510 9326 -11494
rect 10766 -11502 10812 -11490
rect 10944 -11234 10990 -11222
rect 10944 -11490 10950 -11234
rect 10984 -11490 10990 -11234
rect 10944 -11502 10990 -11490
rect 11058 -11234 11104 -11222
rect 11058 -11490 11064 -11234
rect 11098 -11490 11104 -11234
rect 11058 -11502 11104 -11490
rect 11236 -11234 11282 -11222
rect 11236 -11490 11242 -11234
rect 11276 -11490 11282 -11234
rect 11236 -11502 11282 -11490
rect 11350 -11234 11396 -11222
rect 11350 -11490 11356 -11234
rect 11390 -11490 11396 -11234
rect 11350 -11502 11396 -11490
rect 11528 -11234 11574 -11222
rect 11528 -11490 11534 -11234
rect 11568 -11490 11574 -11234
rect 11528 -11502 11574 -11490
rect 11642 -11234 11688 -11222
rect 11642 -11490 11648 -11234
rect 11682 -11490 11688 -11234
rect 11642 -11502 11688 -11490
rect 11820 -11234 11866 -11222
rect 11820 -11490 11826 -11234
rect 11860 -11490 11866 -11234
rect 11820 -11502 11866 -11490
rect 11934 -11234 11980 -11222
rect 11934 -11490 11940 -11234
rect 11974 -11490 11980 -11234
rect 11934 -11502 11980 -11490
rect 12112 -11234 12158 -11222
rect 12112 -11490 12118 -11234
rect 12152 -11490 12158 -11234
rect 12112 -11502 12158 -11490
rect 12226 -11234 12272 -11222
rect 12226 -11490 12232 -11234
rect 12266 -11490 12272 -11234
rect 12226 -11502 12272 -11490
rect 12404 -11234 12450 -11222
rect 12404 -11490 12410 -11234
rect 12444 -11490 12450 -11234
rect 12404 -11502 12450 -11490
rect 12518 -11234 12564 -11222
rect 12518 -11490 12524 -11234
rect 12558 -11490 12564 -11234
rect 12518 -11502 12564 -11490
rect 12696 -11234 12742 -11222
rect 12696 -11490 12702 -11234
rect 12736 -11490 12742 -11234
rect 12696 -11502 12742 -11490
rect 9072 -11544 9088 -11510
rect 9132 -11544 9148 -11510
rect 9072 -11550 9148 -11544
rect 9182 -11544 9266 -11510
rect 9310 -11544 9394 -11510
rect 9182 -11582 9216 -11544
rect 9250 -11550 9326 -11544
rect 9360 -11582 9394 -11544
rect 10840 -11540 10916 -11534
rect 10840 -11574 10856 -11540
rect 10900 -11574 10916 -11540
rect 6506 -11594 6552 -11582
rect 6506 -11850 6512 -11594
rect 6546 -11850 6552 -11594
rect 6506 -11862 6552 -11850
rect 6684 -11594 6730 -11582
rect 6684 -11850 6690 -11594
rect 6724 -11850 6730 -11594
rect 6684 -11862 6730 -11850
rect 6862 -11594 6908 -11582
rect 6862 -11850 6868 -11594
rect 6902 -11850 6908 -11594
rect 6862 -11862 6908 -11850
rect 7040 -11594 7086 -11582
rect 7040 -11850 7046 -11594
rect 7080 -11850 7086 -11594
rect 7040 -11862 7086 -11850
rect 7218 -11594 7264 -11582
rect 7218 -11850 7224 -11594
rect 7258 -11850 7264 -11594
rect 7218 -11862 7264 -11850
rect 7396 -11594 7442 -11582
rect 7396 -11850 7402 -11594
rect 7436 -11850 7442 -11594
rect 7396 -11862 7442 -11850
rect 7574 -11594 7620 -11582
rect 7574 -11850 7580 -11594
rect 7614 -11850 7620 -11594
rect 7574 -11862 7620 -11850
rect 7752 -11594 7798 -11582
rect 7752 -11850 7758 -11594
rect 7792 -11850 7798 -11594
rect 7752 -11862 7798 -11850
rect 7930 -11594 7976 -11582
rect 7930 -11850 7936 -11594
rect 7970 -11850 7976 -11594
rect 7930 -11862 7976 -11850
rect 8108 -11594 8154 -11582
rect 8108 -11850 8114 -11594
rect 8148 -11850 8154 -11594
rect 8108 -11862 8154 -11850
rect 8286 -11594 8332 -11582
rect 8286 -11850 8292 -11594
rect 8326 -11850 8332 -11594
rect 8286 -11862 8332 -11850
rect 8464 -11594 8510 -11582
rect 8464 -11850 8470 -11594
rect 8504 -11850 8510 -11594
rect 8464 -11862 8510 -11850
rect 8642 -11594 8688 -11582
rect 8642 -11850 8648 -11594
rect 8682 -11850 8688 -11594
rect 8642 -11862 8688 -11850
rect 8820 -11594 8866 -11582
rect 8820 -11850 8826 -11594
rect 8860 -11850 8866 -11594
rect 8820 -11862 8866 -11850
rect 8998 -11594 9044 -11582
rect 8998 -11850 9004 -11594
rect 9038 -11850 9044 -11594
rect 8998 -11862 9044 -11850
rect 9176 -11594 9222 -11582
rect 9176 -11850 9182 -11594
rect 9216 -11850 9222 -11594
rect 9176 -11862 9222 -11850
rect 9354 -11594 9400 -11582
rect 10840 -11590 10916 -11574
rect 9354 -11850 9360 -11594
rect 9394 -11850 9400 -11594
rect 11063 -11674 11097 -11502
rect 11132 -11540 11208 -11534
rect 11132 -11574 11148 -11540
rect 11192 -11574 11208 -11540
rect 11132 -11590 11208 -11574
rect 11043 -11727 11053 -11674
rect 11106 -11727 11116 -11674
rect 11356 -11675 11390 -11502
rect 11424 -11540 11500 -11534
rect 11424 -11574 11440 -11540
rect 11484 -11574 11500 -11540
rect 11424 -11590 11500 -11574
rect 11648 -11674 11682 -11502
rect 11716 -11540 11792 -11534
rect 11716 -11574 11732 -11540
rect 11776 -11574 11792 -11540
rect 11716 -11590 11792 -11574
rect 11940 -11674 11974 -11502
rect 12008 -11540 12084 -11534
rect 12008 -11574 12024 -11540
rect 12068 -11574 12084 -11540
rect 12008 -11590 12084 -11574
rect 12233 -11674 12267 -11502
rect 12300 -11540 12376 -11534
rect 12300 -11574 12316 -11540
rect 12360 -11574 12376 -11540
rect 12300 -11590 12376 -11574
rect 12525 -11541 12559 -11502
rect 12592 -11540 12668 -11534
rect 12592 -11541 12608 -11540
rect 12525 -11574 12608 -11541
rect 12652 -11541 12668 -11540
rect 12701 -11541 12735 -11502
rect 12652 -11574 12735 -11541
rect 12525 -11575 12735 -11574
rect 12592 -11590 12668 -11575
rect 11337 -11728 11347 -11675
rect 11400 -11728 11410 -11675
rect 11628 -11727 11638 -11674
rect 11691 -11727 11701 -11674
rect 11921 -11727 11931 -11674
rect 11984 -11727 11994 -11674
rect 12213 -11727 12223 -11674
rect 12276 -11727 12286 -11674
rect 13012 -11726 13022 -11673
rect 13075 -11726 13085 -11673
rect 9354 -11862 9400 -11850
rect 6511 -11900 6545 -11862
rect 6580 -11900 6656 -11894
rect 6688 -11900 6722 -11862
rect 6758 -11900 6834 -11894
rect 6868 -11900 6902 -11862
rect 6511 -11934 6596 -11900
rect 6640 -11934 6774 -11900
rect 6818 -11934 6902 -11900
rect 6580 -11950 6656 -11934
rect 6758 -11950 6834 -11934
rect 6868 -12040 6902 -11934
rect 6936 -11900 7012 -11894
rect 6936 -11934 6952 -11900
rect 6996 -11934 7012 -11900
rect 6936 -11950 7012 -11934
rect 7114 -11900 7190 -11894
rect 7114 -11934 7130 -11900
rect 7174 -11934 7190 -11900
rect 7114 -11950 7190 -11934
rect 7224 -12040 7258 -11862
rect 7292 -11900 7368 -11894
rect 7292 -11934 7308 -11900
rect 7352 -11934 7368 -11900
rect 7292 -11950 7368 -11934
rect 7470 -11900 7546 -11894
rect 7470 -11934 7486 -11900
rect 7530 -11934 7546 -11900
rect 7470 -11950 7546 -11934
rect 7580 -12040 7614 -11862
rect 7648 -11900 7724 -11894
rect 7648 -11934 7664 -11900
rect 7708 -11934 7724 -11900
rect 7648 -11950 7724 -11934
rect 7826 -11900 7902 -11894
rect 7826 -11934 7842 -11900
rect 7886 -11934 7902 -11900
rect 7826 -11950 7902 -11934
rect 7936 -12040 7970 -11862
rect 8004 -11900 8080 -11894
rect 8004 -11934 8020 -11900
rect 8064 -11934 8080 -11900
rect 8004 -11950 8080 -11934
rect 8182 -11900 8258 -11894
rect 8182 -11934 8198 -11900
rect 8242 -11934 8258 -11900
rect 8182 -11950 8258 -11934
rect 8292 -12040 8326 -11862
rect 8360 -11900 8436 -11894
rect 8360 -11934 8376 -11900
rect 8420 -11934 8436 -11900
rect 8360 -11950 8436 -11934
rect 8538 -11900 8614 -11894
rect 8538 -11934 8554 -11900
rect 8598 -11934 8614 -11900
rect 8538 -11950 8614 -11934
rect 8648 -12040 8682 -11862
rect 8716 -11900 8792 -11894
rect 8716 -11934 8732 -11900
rect 8776 -11934 8792 -11900
rect 8716 -11950 8792 -11934
rect 8894 -11900 8970 -11894
rect 8894 -11934 8910 -11900
rect 8954 -11934 8970 -11900
rect 8894 -11950 8970 -11934
rect 9072 -11900 9148 -11894
rect 9072 -11934 9088 -11900
rect 9132 -11934 9148 -11900
rect 9072 -11950 9148 -11934
rect 8912 -11985 8946 -11950
rect 9095 -11985 9129 -11950
rect 9182 -11985 9216 -11862
rect 9250 -11900 9326 -11894
rect 9250 -11934 9266 -11900
rect 9310 -11934 9326 -11900
rect 9250 -11950 9326 -11934
rect 8912 -12019 9216 -11985
rect 6868 -12074 8682 -12040
rect 5027 -13349 5037 -13296
rect 5090 -13349 5100 -13296
rect 5524 -13349 5534 -13296
rect 5587 -13349 5597 -13296
rect 5021 -13486 5031 -13433
rect 5084 -13486 5094 -13433
rect 4895 -14598 4905 -14545
rect 4958 -14598 4968 -14545
rect 4531 -14869 4733 -14863
rect 4229 -14979 4239 -14926
rect 4292 -14979 4302 -14926
rect 3947 -15047 4023 -15032
rect 3879 -15048 4091 -15047
rect 3879 -15081 3963 -15048
rect 3879 -15120 3913 -15081
rect 3947 -15082 3963 -15081
rect 4007 -15081 4091 -15048
rect 4007 -15082 4023 -15081
rect 3947 -15088 4023 -15082
rect 4057 -15120 4091 -15081
rect -2179 -15132 -2133 -15120
rect -2179 -15388 -2173 -15132
rect -2139 -15388 -2133 -15132
rect -2179 -15400 -2133 -15388
rect -2001 -15132 -1955 -15120
rect -2001 -15388 -1995 -15132
rect -1961 -15388 -1955 -15132
rect -2001 -15400 -1955 -15388
rect -1823 -15132 -1777 -15120
rect -1823 -15388 -1817 -15132
rect -1783 -15388 -1777 -15132
rect -1823 -15400 -1777 -15388
rect -1645 -15132 -1599 -15120
rect -1645 -15388 -1639 -15132
rect -1605 -15388 -1599 -15132
rect -1645 -15400 -1599 -15388
rect -1467 -15132 -1421 -15120
rect -1467 -15388 -1461 -15132
rect -1427 -15388 -1421 -15132
rect -1467 -15400 -1421 -15388
rect -1289 -15132 -1243 -15120
rect -1289 -15388 -1283 -15132
rect -1249 -15388 -1243 -15132
rect -1289 -15400 -1243 -15388
rect -1111 -15132 -1065 -15120
rect -1111 -15388 -1105 -15132
rect -1071 -15388 -1065 -15132
rect -1111 -15400 -1065 -15388
rect -933 -15132 -887 -15120
rect -933 -15388 -927 -15132
rect -893 -15388 -887 -15132
rect -933 -15400 -887 -15388
rect -755 -15132 -709 -15120
rect -755 -15388 -749 -15132
rect -715 -15388 -709 -15132
rect -755 -15400 -709 -15388
rect -577 -15132 -531 -15120
rect -577 -15388 -571 -15132
rect -537 -15388 -531 -15132
rect -577 -15400 -531 -15388
rect -399 -15132 -353 -15120
rect -399 -15388 -393 -15132
rect -359 -15388 -353 -15132
rect -399 -15400 -353 -15388
rect -221 -15132 -175 -15120
rect -221 -15388 -215 -15132
rect -181 -15388 -175 -15132
rect -221 -15400 -175 -15388
rect -43 -15132 3 -15120
rect -43 -15388 -37 -15132
rect -3 -15388 3 -15132
rect -43 -15400 3 -15388
rect 135 -15132 181 -15120
rect 135 -15388 141 -15132
rect 175 -15388 181 -15132
rect 135 -15400 181 -15388
rect 313 -15132 359 -15120
rect 313 -15388 319 -15132
rect 353 -15388 359 -15132
rect 313 -15400 359 -15388
rect 491 -15132 537 -15120
rect 491 -15388 497 -15132
rect 531 -15388 537 -15132
rect 491 -15400 537 -15388
rect 669 -15132 715 -15120
rect 669 -15388 675 -15132
rect 709 -15388 715 -15132
rect 669 -15400 715 -15388
rect 847 -15132 893 -15120
rect 847 -15388 853 -15132
rect 887 -15388 893 -15132
rect 847 -15400 893 -15388
rect 1025 -15132 1071 -15120
rect 1025 -15388 1031 -15132
rect 1065 -15388 1071 -15132
rect 1025 -15400 1071 -15388
rect 1203 -15132 1249 -15120
rect 1203 -15388 1209 -15132
rect 1243 -15388 1249 -15132
rect 1203 -15400 1249 -15388
rect 1381 -15132 1427 -15120
rect 1381 -15388 1387 -15132
rect 1421 -15388 1427 -15132
rect 1381 -15400 1427 -15388
rect 1559 -15132 1605 -15120
rect 1559 -15388 1565 -15132
rect 1599 -15388 1605 -15132
rect 1559 -15400 1605 -15388
rect 1737 -15132 1783 -15120
rect 1737 -15388 1743 -15132
rect 1777 -15388 1783 -15132
rect 1737 -15400 1783 -15388
rect 1915 -15132 1961 -15120
rect 1915 -15388 1921 -15132
rect 1955 -15388 1961 -15132
rect 1915 -15400 1961 -15388
rect 2093 -15132 2139 -15120
rect 2093 -15388 2099 -15132
rect 2133 -15388 2139 -15132
rect 2093 -15400 2139 -15388
rect 2271 -15132 2317 -15120
rect 2271 -15388 2277 -15132
rect 2311 -15388 2317 -15132
rect 2271 -15400 2317 -15388
rect 2449 -15132 2495 -15120
rect 2449 -15388 2455 -15132
rect 2489 -15388 2495 -15132
rect 2449 -15400 2495 -15388
rect 2627 -15132 2673 -15120
rect 2627 -15388 2633 -15132
rect 2667 -15388 2673 -15132
rect 2627 -15400 2673 -15388
rect 2805 -15132 2851 -15120
rect 2805 -15388 2811 -15132
rect 2845 -15388 2851 -15132
rect 2805 -15400 2851 -15388
rect 2983 -15132 3029 -15120
rect 2983 -15388 2989 -15132
rect 3023 -15388 3029 -15132
rect 2983 -15400 3029 -15388
rect 3161 -15132 3207 -15120
rect 3161 -15388 3167 -15132
rect 3201 -15388 3207 -15132
rect 3161 -15400 3207 -15388
rect 3339 -15132 3385 -15120
rect 3339 -15388 3345 -15132
rect 3379 -15388 3385 -15132
rect 3339 -15400 3385 -15388
rect 3517 -15132 3563 -15120
rect 3517 -15388 3523 -15132
rect 3557 -15388 3563 -15132
rect 3517 -15400 3563 -15388
rect 3695 -15132 3741 -15120
rect 3695 -15388 3701 -15132
rect 3735 -15388 3741 -15132
rect 3695 -15400 3741 -15388
rect 3873 -15132 3919 -15120
rect 3873 -15388 3879 -15132
rect 3913 -15388 3919 -15132
rect 3873 -15400 3919 -15388
rect 4051 -15132 4097 -15120
rect 4051 -15388 4057 -15132
rect 4091 -15388 4097 -15132
rect 4051 -15400 4097 -15388
rect -2105 -15438 -2029 -15432
rect -2105 -15472 -2089 -15438
rect -2045 -15472 -2029 -15438
rect -2105 -15488 -2029 -15472
rect -2457 -15874 -2447 -15821
rect -2394 -15874 -2384 -15821
rect -1995 -15822 -1961 -15400
rect -1927 -15438 -1851 -15432
rect -1927 -15472 -1911 -15438
rect -1867 -15472 -1851 -15438
rect -1927 -15488 -1851 -15472
rect -2015 -15875 -2005 -15822
rect -1952 -15875 -1942 -15822
rect -2105 -16048 -2029 -16032
rect -2105 -16050 -2089 -16048
rect -2173 -16082 -2089 -16050
rect -2045 -16050 -2029 -16048
rect -1995 -16050 -1961 -15875
rect -1906 -15933 -1872 -15488
rect -1925 -15986 -1915 -15933
rect -1862 -15986 -1852 -15933
rect -2045 -16082 -1961 -16050
rect -2173 -16084 -1961 -16082
rect -2173 -16120 -2139 -16084
rect -2105 -16088 -2029 -16084
rect -1995 -16120 -1961 -16084
rect -1927 -16048 -1851 -16032
rect -1927 -16082 -1911 -16048
rect -1867 -16082 -1851 -16048
rect -1927 -16088 -1851 -16082
rect -1817 -16120 -1783 -15400
rect -1749 -15438 -1673 -15432
rect -1749 -15472 -1733 -15438
rect -1689 -15472 -1673 -15438
rect -1749 -15488 -1673 -15472
rect -1728 -15933 -1694 -15488
rect -1639 -15822 -1605 -15400
rect -1571 -15438 -1495 -15432
rect -1571 -15472 -1555 -15438
rect -1511 -15472 -1495 -15438
rect -1571 -15488 -1495 -15472
rect -1659 -15875 -1649 -15822
rect -1596 -15875 -1586 -15822
rect -1748 -15986 -1738 -15933
rect -1685 -15986 -1675 -15933
rect -1749 -16048 -1673 -16032
rect -1749 -16082 -1733 -16048
rect -1689 -16082 -1673 -16048
rect -1749 -16088 -1673 -16082
rect -1639 -16120 -1605 -15875
rect -1550 -15933 -1516 -15488
rect -1570 -15986 -1560 -15933
rect -1507 -15986 -1497 -15933
rect -1571 -16048 -1495 -16032
rect -1571 -16082 -1555 -16048
rect -1511 -16082 -1495 -16048
rect -1571 -16088 -1495 -16082
rect -1461 -16120 -1427 -15400
rect -1393 -15438 -1317 -15432
rect -1393 -15472 -1377 -15438
rect -1333 -15472 -1317 -15438
rect -1393 -15488 -1317 -15472
rect -1372 -15933 -1338 -15488
rect -1283 -15822 -1249 -15400
rect -1215 -15438 -1139 -15432
rect -1215 -15472 -1199 -15438
rect -1155 -15472 -1139 -15438
rect -1215 -15488 -1139 -15472
rect -1303 -15875 -1293 -15822
rect -1240 -15875 -1230 -15822
rect -1392 -15986 -1382 -15933
rect -1329 -15986 -1319 -15933
rect -1393 -16048 -1317 -16032
rect -1393 -16082 -1377 -16048
rect -1333 -16082 -1317 -16048
rect -1393 -16088 -1317 -16082
rect -1283 -16120 -1249 -15875
rect -1194 -15933 -1160 -15488
rect -1214 -15986 -1204 -15933
rect -1151 -15986 -1141 -15933
rect -1215 -16048 -1139 -16032
rect -1215 -16082 -1199 -16048
rect -1155 -16082 -1139 -16048
rect -1215 -16088 -1139 -16082
rect -1104 -16120 -1070 -15400
rect -1037 -15438 -961 -15432
rect -1037 -15472 -1021 -15438
rect -977 -15472 -961 -15438
rect -1037 -15488 -961 -15472
rect -1015 -15933 -981 -15488
rect -927 -15822 -893 -15400
rect -859 -15438 -783 -15432
rect -859 -15472 -843 -15438
rect -799 -15472 -783 -15438
rect -859 -15488 -783 -15472
rect -947 -15875 -937 -15822
rect -884 -15875 -874 -15822
rect -1035 -15986 -1025 -15933
rect -972 -15986 -962 -15933
rect -1037 -16048 -961 -16032
rect -1037 -16082 -1021 -16048
rect -977 -16082 -961 -16048
rect -1037 -16088 -961 -16082
rect -927 -16120 -893 -15875
rect -857 -15986 -847 -15933
rect -794 -15986 -784 -15933
rect -838 -16032 -804 -15986
rect -859 -16048 -783 -16032
rect -859 -16082 -843 -16048
rect -799 -16082 -783 -16048
rect -859 -16088 -783 -16082
rect -749 -16120 -715 -15400
rect -681 -15438 -605 -15432
rect -681 -15472 -665 -15438
rect -621 -15472 -605 -15438
rect -681 -15488 -605 -15472
rect -571 -15822 -537 -15400
rect -503 -15438 -427 -15432
rect -503 -15472 -487 -15438
rect -443 -15472 -427 -15438
rect -503 -15488 -427 -15472
rect -591 -15875 -581 -15822
rect -528 -15875 -518 -15822
rect -680 -15986 -670 -15933
rect -617 -15986 -607 -15933
rect -660 -16032 -626 -15986
rect -681 -16048 -605 -16032
rect -681 -16082 -665 -16048
rect -621 -16082 -605 -16048
rect -681 -16088 -605 -16082
rect -571 -16120 -537 -15875
rect -501 -15986 -491 -15933
rect -438 -15986 -428 -15933
rect -482 -16032 -448 -15986
rect -503 -16048 -427 -16032
rect -503 -16082 -487 -16048
rect -443 -16082 -427 -16048
rect -503 -16088 -427 -16082
rect -393 -16120 -359 -15400
rect -325 -15438 -249 -15432
rect -325 -15472 -309 -15438
rect -265 -15472 -249 -15438
rect -325 -15488 -249 -15472
rect -215 -15822 -181 -15400
rect -147 -15438 -71 -15432
rect -147 -15472 -131 -15438
rect -87 -15472 -71 -15438
rect -147 -15488 -71 -15472
rect -235 -15875 -225 -15822
rect -172 -15875 -162 -15822
rect -323 -15986 -313 -15933
rect -260 -15986 -250 -15933
rect -304 -16032 -270 -15986
rect -325 -16048 -249 -16032
rect -325 -16082 -309 -16048
rect -265 -16082 -249 -16048
rect -325 -16088 -249 -16082
rect -215 -16120 -181 -15875
rect -146 -15986 -136 -15933
rect -83 -15986 -73 -15933
rect -126 -16032 -92 -15986
rect -147 -16048 -71 -16032
rect -147 -16082 -131 -16048
rect -87 -16082 -71 -16048
rect -147 -16088 -71 -16082
rect -37 -16120 -3 -15400
rect 31 -15438 107 -15432
rect 31 -15472 47 -15438
rect 91 -15472 107 -15438
rect 31 -15488 107 -15472
rect 141 -15821 175 -15400
rect 209 -15438 285 -15432
rect 209 -15472 225 -15438
rect 269 -15472 285 -15438
rect 209 -15488 285 -15472
rect 122 -15874 132 -15821
rect 185 -15874 195 -15821
rect 33 -15986 43 -15933
rect 96 -15986 106 -15933
rect 52 -16032 86 -15986
rect 31 -16048 107 -16032
rect 31 -16082 47 -16048
rect 91 -16082 107 -16048
rect 31 -16088 107 -16082
rect 141 -16120 175 -15874
rect 230 -15933 264 -15488
rect 211 -15986 221 -15933
rect 274 -15986 284 -15933
rect 209 -16048 285 -16032
rect 209 -16082 225 -16048
rect 269 -16082 285 -16048
rect 209 -16088 285 -16082
rect 319 -16120 353 -15400
rect 387 -15438 463 -15432
rect 387 -15472 403 -15438
rect 447 -15472 463 -15438
rect 387 -15488 463 -15472
rect 408 -15933 442 -15488
rect 497 -15822 531 -15400
rect 565 -15438 641 -15432
rect 565 -15472 581 -15438
rect 625 -15472 641 -15438
rect 565 -15488 641 -15472
rect 477 -15875 487 -15822
rect 540 -15875 550 -15822
rect 388 -15986 398 -15933
rect 451 -15986 461 -15933
rect 387 -16048 463 -16032
rect 387 -16082 403 -16048
rect 447 -16082 463 -16048
rect 387 -16088 463 -16082
rect 497 -16120 531 -15875
rect 585 -15933 619 -15488
rect 565 -15986 575 -15933
rect 628 -15986 638 -15933
rect 565 -16048 641 -16032
rect 565 -16082 581 -16048
rect 625 -16082 641 -16048
rect 565 -16088 641 -16082
rect 675 -16120 709 -15400
rect 743 -15438 819 -15432
rect 743 -15472 759 -15438
rect 803 -15472 819 -15438
rect 743 -15488 819 -15472
rect 764 -15933 798 -15488
rect 853 -15822 887 -15400
rect 921 -15438 997 -15432
rect 921 -15472 937 -15438
rect 981 -15472 997 -15438
rect 921 -15488 997 -15472
rect 833 -15875 843 -15822
rect 896 -15875 906 -15822
rect 745 -15986 755 -15933
rect 808 -15986 818 -15933
rect 743 -16048 819 -16032
rect 743 -16082 759 -16048
rect 803 -16082 819 -16048
rect 743 -16088 819 -16082
rect 853 -16120 887 -15875
rect 941 -15933 975 -15488
rect 921 -15986 931 -15933
rect 984 -15986 994 -15933
rect 921 -16048 997 -16032
rect 921 -16082 937 -16048
rect 981 -16082 997 -16048
rect 921 -16088 997 -16082
rect 1031 -16120 1065 -15400
rect 1099 -15438 1175 -15432
rect 1099 -15472 1115 -15438
rect 1159 -15472 1175 -15438
rect 1099 -15488 1175 -15472
rect 1120 -15933 1154 -15488
rect 1209 -15822 1243 -15400
rect 1277 -15438 1353 -15432
rect 1277 -15472 1293 -15438
rect 1337 -15472 1353 -15438
rect 1277 -15488 1353 -15472
rect 1191 -15875 1201 -15822
rect 1254 -15875 1264 -15822
rect 1100 -15986 1110 -15933
rect 1163 -15986 1173 -15933
rect 1099 -16048 1175 -16032
rect 1099 -16082 1115 -16048
rect 1159 -16082 1175 -16048
rect 1099 -16088 1175 -16082
rect 1209 -16120 1243 -15875
rect 1279 -15986 1289 -15933
rect 1342 -15986 1352 -15933
rect 1298 -16032 1332 -15986
rect 1277 -16048 1353 -16032
rect 1277 -16082 1293 -16048
rect 1337 -16082 1353 -16048
rect 1277 -16088 1353 -16082
rect 1387 -16120 1421 -15400
rect 1455 -15438 1531 -15432
rect 1455 -15472 1471 -15438
rect 1515 -15472 1531 -15438
rect 1455 -15488 1531 -15472
rect 1565 -15822 1599 -15400
rect 1633 -15438 1709 -15432
rect 1633 -15472 1649 -15438
rect 1693 -15472 1709 -15438
rect 1633 -15488 1709 -15472
rect 1545 -15875 1555 -15822
rect 1608 -15875 1618 -15822
rect 1456 -15986 1466 -15933
rect 1519 -15986 1529 -15933
rect 1476 -16032 1510 -15986
rect 1455 -16048 1531 -16032
rect 1455 -16082 1471 -16048
rect 1515 -16082 1531 -16048
rect 1455 -16088 1531 -16082
rect 1565 -16120 1599 -15875
rect 1633 -15986 1643 -15933
rect 1696 -15986 1706 -15933
rect 1653 -16032 1687 -15986
rect 1633 -16048 1709 -16032
rect 1633 -16082 1649 -16048
rect 1693 -16082 1709 -16048
rect 1633 -16088 1709 -16082
rect 1744 -16120 1778 -15400
rect 1811 -15438 1887 -15432
rect 1811 -15472 1827 -15438
rect 1871 -15472 1887 -15438
rect 1811 -15488 1887 -15472
rect 1921 -15822 1955 -15400
rect 1989 -15438 2065 -15432
rect 1989 -15472 2005 -15438
rect 2049 -15472 2065 -15438
rect 1989 -15488 2065 -15472
rect 1900 -15875 1910 -15822
rect 1963 -15875 1973 -15822
rect 1812 -15986 1822 -15933
rect 1875 -15986 1885 -15933
rect 1832 -16032 1866 -15986
rect 1811 -16048 1887 -16032
rect 1811 -16082 1827 -16048
rect 1871 -16082 1887 -16048
rect 1811 -16088 1887 -16082
rect 1921 -16120 1955 -15875
rect 1990 -15986 2000 -15933
rect 2053 -15986 2063 -15933
rect 2010 -16032 2044 -15986
rect 1989 -16048 2065 -16032
rect 1989 -16082 2005 -16048
rect 2049 -16082 2065 -16048
rect 1989 -16088 2065 -16082
rect 2100 -16120 2134 -15400
rect 2167 -15438 2243 -15432
rect 2167 -15472 2183 -15438
rect 2227 -15472 2243 -15438
rect 2167 -15488 2243 -15472
rect 2277 -15822 2311 -15400
rect 2345 -15438 2421 -15432
rect 2345 -15472 2361 -15438
rect 2405 -15472 2421 -15438
rect 2345 -15488 2421 -15472
rect 2257 -15875 2267 -15822
rect 2320 -15875 2330 -15822
rect 2169 -15986 2179 -15933
rect 2232 -15986 2242 -15933
rect 2189 -16032 2223 -15986
rect 2167 -16048 2243 -16032
rect 2167 -16082 2183 -16048
rect 2227 -16082 2243 -16048
rect 2167 -16088 2243 -16082
rect 2277 -16120 2311 -15875
rect 2366 -15933 2400 -15488
rect 2346 -15986 2356 -15933
rect 2409 -15986 2419 -15933
rect 2345 -16048 2421 -16032
rect 2345 -16082 2361 -16048
rect 2405 -16082 2421 -16048
rect 2345 -16088 2421 -16082
rect 2455 -16120 2489 -15400
rect 2523 -15438 2599 -15432
rect 2523 -15472 2539 -15438
rect 2583 -15472 2599 -15438
rect 2523 -15488 2599 -15472
rect 2544 -15933 2578 -15488
rect 2633 -15822 2667 -15400
rect 2701 -15438 2777 -15432
rect 2701 -15472 2717 -15438
rect 2761 -15472 2777 -15438
rect 2701 -15488 2777 -15472
rect 2614 -15875 2624 -15822
rect 2677 -15875 2687 -15822
rect 2524 -15986 2534 -15933
rect 2587 -15986 2597 -15933
rect 2523 -16048 2599 -16032
rect 2523 -16082 2539 -16048
rect 2583 -16082 2599 -16048
rect 2523 -16088 2599 -16082
rect 2633 -16120 2667 -15875
rect 2722 -15933 2756 -15488
rect 2702 -15986 2712 -15933
rect 2765 -15986 2775 -15933
rect 2701 -16048 2777 -16032
rect 2701 -16082 2717 -16048
rect 2761 -16082 2777 -16048
rect 2701 -16088 2777 -16082
rect 2811 -16120 2845 -15400
rect 2879 -15438 2955 -15432
rect 2879 -15472 2895 -15438
rect 2939 -15472 2955 -15438
rect 2879 -15488 2955 -15472
rect 2900 -15933 2934 -15488
rect 2989 -15822 3023 -15400
rect 3057 -15438 3133 -15432
rect 3057 -15472 3073 -15438
rect 3117 -15472 3133 -15438
rect 3057 -15488 3133 -15472
rect 2969 -15875 2979 -15822
rect 3032 -15875 3042 -15822
rect 2881 -15986 2891 -15933
rect 2944 -15986 2954 -15933
rect 2879 -16048 2955 -16032
rect 2879 -16082 2895 -16048
rect 2939 -16082 2955 -16048
rect 2879 -16088 2955 -16082
rect 2989 -16120 3023 -15875
rect 3078 -15933 3112 -15488
rect 3058 -15986 3068 -15933
rect 3121 -15986 3131 -15933
rect 3057 -16048 3133 -16032
rect 3057 -16082 3073 -16048
rect 3117 -16082 3133 -16048
rect 3057 -16088 3133 -16082
rect 3167 -16120 3201 -15400
rect 3235 -15438 3311 -15432
rect 3235 -15472 3251 -15438
rect 3295 -15472 3311 -15438
rect 3235 -15488 3311 -15472
rect 3256 -15933 3290 -15488
rect 3345 -15822 3379 -15400
rect 3413 -15438 3489 -15432
rect 3413 -15472 3429 -15438
rect 3473 -15472 3489 -15438
rect 3413 -15488 3489 -15472
rect 3325 -15875 3335 -15822
rect 3388 -15875 3398 -15822
rect 3237 -15986 3247 -15933
rect 3300 -15986 3310 -15933
rect 3235 -16048 3311 -16032
rect 3235 -16082 3251 -16048
rect 3295 -16082 3311 -16048
rect 3235 -16088 3311 -16082
rect 3345 -16120 3379 -15875
rect 3414 -15986 3424 -15933
rect 3477 -15986 3487 -15933
rect 3434 -16032 3468 -15986
rect 3413 -16048 3489 -16032
rect 3413 -16082 3429 -16048
rect 3473 -16082 3489 -16048
rect 3413 -16088 3489 -16082
rect 3524 -16120 3558 -15400
rect 3591 -15438 3667 -15432
rect 3591 -15472 3607 -15438
rect 3651 -15472 3667 -15438
rect 3591 -15488 3667 -15472
rect 3701 -15822 3735 -15400
rect 3769 -15438 3845 -15432
rect 3769 -15472 3785 -15438
rect 3829 -15472 3845 -15438
rect 3769 -15488 3845 -15472
rect 3682 -15875 3692 -15822
rect 3745 -15875 3755 -15822
rect 3593 -15986 3603 -15933
rect 3656 -15986 3666 -15933
rect 3612 -16032 3646 -15986
rect 3591 -16048 3667 -16032
rect 3591 -16082 3607 -16048
rect 3651 -16082 3667 -16048
rect 3591 -16088 3667 -16082
rect 3701 -16120 3735 -15875
rect 3770 -15986 3780 -15933
rect 3833 -15986 3843 -15933
rect 3790 -16032 3824 -15986
rect 3769 -16048 3845 -16032
rect 3769 -16082 3785 -16048
rect 3829 -16082 3845 -16048
rect 3769 -16088 3845 -16082
rect 3879 -16047 3913 -15400
rect 3947 -15438 4023 -15432
rect 3947 -15472 3963 -15438
rect 4007 -15472 4023 -15438
rect 3947 -15488 4023 -15472
rect 4238 -15539 4291 -14979
rect 4531 -15047 4543 -14869
rect 4721 -15047 4733 -14869
rect 4531 -15053 4733 -15047
rect 4228 -15592 4238 -15539
rect 4291 -15592 4301 -15539
rect 5031 -15540 5084 -13486
rect 5390 -13598 5400 -13545
rect 5453 -13598 5463 -13545
rect 5132 -13847 5142 -13794
rect 5195 -13847 5205 -13794
rect 5142 -14658 5195 -13847
rect 5133 -14711 5143 -14658
rect 5196 -14711 5206 -14658
rect 3947 -16047 4023 -16032
rect 3879 -16048 4090 -16047
rect 3879 -16081 3963 -16048
rect 3879 -16120 3913 -16081
rect 3947 -16082 3963 -16081
rect 4007 -16081 4090 -16048
rect 4007 -16082 4023 -16081
rect 3947 -16088 4023 -16082
rect 4056 -16120 4090 -16081
rect -2179 -16132 -2133 -16120
rect -3945 -16347 -3935 -16295
rect -3883 -16347 -3873 -16295
rect -4180 -16410 -4104 -16394
rect -4180 -16444 -4164 -16410
rect -4120 -16444 -4104 -16410
rect -4180 -16450 -4104 -16444
rect -6034 -16494 -5988 -16482
rect -6034 -16750 -6028 -16494
rect -5994 -16750 -5988 -16494
rect -6034 -16762 -5988 -16750
rect -5856 -16494 -5810 -16482
rect -5856 -16750 -5850 -16494
rect -5816 -16750 -5810 -16494
rect -5856 -16762 -5810 -16750
rect -5678 -16494 -5632 -16482
rect -5678 -16750 -5672 -16494
rect -5638 -16750 -5632 -16494
rect -5678 -16762 -5632 -16750
rect -5500 -16494 -5454 -16482
rect -5500 -16750 -5494 -16494
rect -5460 -16750 -5454 -16494
rect -5500 -16762 -5454 -16750
rect -5322 -16494 -5276 -16482
rect -5322 -16750 -5316 -16494
rect -5282 -16750 -5276 -16494
rect -5322 -16762 -5276 -16750
rect -5144 -16494 -5098 -16482
rect -5144 -16750 -5138 -16494
rect -5104 -16750 -5098 -16494
rect -5144 -16762 -5098 -16750
rect -4966 -16494 -4920 -16482
rect -4966 -16750 -4960 -16494
rect -4926 -16750 -4920 -16494
rect -4966 -16762 -4920 -16750
rect -4788 -16494 -4742 -16482
rect -4788 -16750 -4782 -16494
rect -4748 -16750 -4742 -16494
rect -4788 -16762 -4742 -16750
rect -4610 -16494 -4564 -16482
rect -4610 -16750 -4604 -16494
rect -4570 -16750 -4564 -16494
rect -4610 -16762 -4564 -16750
rect -4432 -16494 -4386 -16482
rect -4432 -16750 -4426 -16494
rect -4392 -16750 -4386 -16494
rect -4432 -16762 -4386 -16750
rect -4254 -16494 -4208 -16482
rect -4254 -16750 -4248 -16494
rect -4214 -16750 -4208 -16494
rect -4254 -16762 -4208 -16750
rect -4076 -16494 -4030 -16482
rect -4076 -16750 -4070 -16494
rect -4036 -16750 -4030 -16494
rect -4076 -16762 -4030 -16750
rect -6028 -16886 -5994 -16762
rect -5960 -16800 -5884 -16794
rect -5960 -16834 -5944 -16800
rect -5900 -16834 -5884 -16800
rect -5960 -16850 -5884 -16834
rect -5939 -16886 -5905 -16850
rect -5850 -16886 -5816 -16762
rect -5782 -16800 -5706 -16794
rect -5782 -16834 -5766 -16800
rect -5722 -16834 -5706 -16800
rect -5782 -16850 -5706 -16834
rect -5672 -16886 -5638 -16762
rect -5604 -16800 -5528 -16794
rect -5604 -16834 -5588 -16800
rect -5544 -16834 -5528 -16800
rect -5604 -16850 -5528 -16834
rect -6028 -16920 -5816 -16886
rect -5850 -17007 -5816 -16920
rect -5692 -16939 -5682 -16886
rect -5629 -16939 -5619 -16886
rect -6169 -17060 -6159 -17007
rect -6106 -17060 -6096 -17007
rect -5869 -17060 -5859 -17007
rect -5806 -17060 -5796 -17007
rect -5494 -17118 -5460 -16762
rect -5426 -16800 -5350 -16794
rect -5426 -16834 -5410 -16800
rect -5366 -16834 -5350 -16800
rect -5426 -16850 -5350 -16834
rect -5316 -16886 -5282 -16762
rect -5248 -16800 -5172 -16794
rect -5248 -16834 -5232 -16800
rect -5188 -16834 -5172 -16800
rect -5248 -16850 -5172 -16834
rect -5336 -16939 -5326 -16886
rect -5273 -16939 -5263 -16886
rect -5138 -17007 -5104 -16762
rect -5070 -16800 -4994 -16794
rect -5070 -16834 -5054 -16800
rect -5010 -16834 -4994 -16800
rect -5070 -16850 -4994 -16834
rect -4960 -16886 -4926 -16762
rect -4892 -16800 -4816 -16794
rect -4892 -16834 -4876 -16800
rect -4832 -16834 -4816 -16800
rect -4892 -16850 -4816 -16834
rect -4980 -16939 -4970 -16886
rect -4917 -16939 -4907 -16886
rect -5158 -17060 -5148 -17007
rect -5095 -17060 -5085 -17007
rect -5514 -17171 -5504 -17118
rect -5451 -17171 -5441 -17118
rect -7605 -17251 -7329 -17250
rect -4970 -17251 -4917 -16939
rect -4782 -17118 -4748 -16762
rect -4714 -16800 -4638 -16794
rect -4714 -16834 -4698 -16800
rect -4654 -16834 -4638 -16800
rect -4714 -16850 -4638 -16834
rect -4604 -16886 -4570 -16762
rect -4536 -16800 -4460 -16794
rect -4536 -16834 -4520 -16800
rect -4476 -16834 -4460 -16800
rect -4536 -16850 -4460 -16834
rect -4624 -16939 -4614 -16886
rect -4561 -16939 -4551 -16886
rect -4426 -17007 -4392 -16762
rect -4358 -16800 -4282 -16794
rect -4358 -16834 -4342 -16800
rect -4298 -16834 -4282 -16800
rect -4358 -16850 -4282 -16834
rect -4248 -16886 -4214 -16762
rect -4180 -16800 -4104 -16794
rect -4180 -16834 -4164 -16800
rect -4120 -16834 -4104 -16800
rect -4180 -16850 -4104 -16834
rect -4159 -16886 -4125 -16850
rect -4070 -16886 -4036 -16762
rect -4268 -16939 -4258 -16886
rect -4205 -16939 -4036 -16886
rect -4447 -17060 -4437 -17007
rect -4384 -17060 -4374 -17007
rect -3935 -17118 -3883 -16347
rect -2179 -16388 -2173 -16132
rect -2139 -16388 -2133 -16132
rect -2179 -16400 -2133 -16388
rect -2001 -16132 -1955 -16120
rect -2001 -16388 -1995 -16132
rect -1961 -16388 -1955 -16132
rect -2001 -16400 -1955 -16388
rect -1823 -16132 -1777 -16120
rect -1823 -16388 -1817 -16132
rect -1783 -16388 -1777 -16132
rect -1823 -16400 -1777 -16388
rect -1645 -16132 -1599 -16120
rect -1645 -16388 -1639 -16132
rect -1605 -16388 -1599 -16132
rect -1645 -16400 -1599 -16388
rect -1467 -16132 -1421 -16120
rect -1467 -16388 -1461 -16132
rect -1427 -16388 -1421 -16132
rect -1467 -16400 -1421 -16388
rect -1289 -16132 -1243 -16120
rect -1289 -16388 -1283 -16132
rect -1249 -16388 -1243 -16132
rect -1289 -16400 -1243 -16388
rect -1111 -16132 -1065 -16120
rect -1111 -16388 -1105 -16132
rect -1071 -16388 -1065 -16132
rect -1111 -16400 -1065 -16388
rect -933 -16132 -887 -16120
rect -933 -16388 -927 -16132
rect -893 -16388 -887 -16132
rect -933 -16400 -887 -16388
rect -755 -16132 -709 -16120
rect -755 -16388 -749 -16132
rect -715 -16388 -709 -16132
rect -755 -16400 -709 -16388
rect -577 -16132 -531 -16120
rect -577 -16388 -571 -16132
rect -537 -16388 -531 -16132
rect -577 -16400 -531 -16388
rect -399 -16132 -353 -16120
rect -399 -16388 -393 -16132
rect -359 -16388 -353 -16132
rect -399 -16400 -353 -16388
rect -221 -16132 -175 -16120
rect -221 -16388 -215 -16132
rect -181 -16388 -175 -16132
rect -221 -16400 -175 -16388
rect -43 -16132 3 -16120
rect -43 -16388 -37 -16132
rect -3 -16388 3 -16132
rect -43 -16400 3 -16388
rect 135 -16132 181 -16120
rect 135 -16388 141 -16132
rect 175 -16388 181 -16132
rect 135 -16400 181 -16388
rect 313 -16132 359 -16120
rect 313 -16388 319 -16132
rect 353 -16388 359 -16132
rect 313 -16400 359 -16388
rect 491 -16132 537 -16120
rect 491 -16388 497 -16132
rect 531 -16388 537 -16132
rect 491 -16400 537 -16388
rect 669 -16132 715 -16120
rect 669 -16388 675 -16132
rect 709 -16388 715 -16132
rect 669 -16400 715 -16388
rect 847 -16132 893 -16120
rect 847 -16388 853 -16132
rect 887 -16388 893 -16132
rect 847 -16400 893 -16388
rect 1025 -16132 1071 -16120
rect 1025 -16388 1031 -16132
rect 1065 -16388 1071 -16132
rect 1025 -16400 1071 -16388
rect 1203 -16132 1249 -16120
rect 1203 -16388 1209 -16132
rect 1243 -16388 1249 -16132
rect 1203 -16400 1249 -16388
rect 1381 -16132 1427 -16120
rect 1381 -16388 1387 -16132
rect 1421 -16388 1427 -16132
rect 1381 -16400 1427 -16388
rect 1559 -16132 1605 -16120
rect 1559 -16388 1565 -16132
rect 1599 -16388 1605 -16132
rect 1559 -16400 1605 -16388
rect 1737 -16132 1783 -16120
rect 1737 -16388 1743 -16132
rect 1777 -16388 1783 -16132
rect 1737 -16400 1783 -16388
rect 1915 -16132 1961 -16120
rect 1915 -16388 1921 -16132
rect 1955 -16388 1961 -16132
rect 1915 -16400 1961 -16388
rect 2093 -16132 2139 -16120
rect 2093 -16388 2099 -16132
rect 2133 -16388 2139 -16132
rect 2093 -16400 2139 -16388
rect 2271 -16132 2317 -16120
rect 2271 -16388 2277 -16132
rect 2311 -16388 2317 -16132
rect 2271 -16400 2317 -16388
rect 2449 -16132 2495 -16120
rect 2449 -16388 2455 -16132
rect 2489 -16388 2495 -16132
rect 2449 -16400 2495 -16388
rect 2627 -16132 2673 -16120
rect 2627 -16388 2633 -16132
rect 2667 -16388 2673 -16132
rect 2627 -16400 2673 -16388
rect 2805 -16132 2851 -16120
rect 2805 -16388 2811 -16132
rect 2845 -16388 2851 -16132
rect 2805 -16400 2851 -16388
rect 2983 -16132 3029 -16120
rect 2983 -16388 2989 -16132
rect 3023 -16388 3029 -16132
rect 2983 -16400 3029 -16388
rect 3161 -16132 3207 -16120
rect 3161 -16388 3167 -16132
rect 3201 -16388 3207 -16132
rect 3161 -16400 3207 -16388
rect 3339 -16132 3385 -16120
rect 3339 -16388 3345 -16132
rect 3379 -16388 3385 -16132
rect 3339 -16400 3385 -16388
rect 3517 -16132 3563 -16120
rect 3517 -16388 3523 -16132
rect 3557 -16388 3563 -16132
rect 3517 -16400 3563 -16388
rect 3695 -16132 3741 -16120
rect 3695 -16388 3701 -16132
rect 3735 -16388 3741 -16132
rect 3695 -16400 3741 -16388
rect 3873 -16132 3919 -16120
rect 3873 -16388 3879 -16132
rect 3913 -16388 3919 -16132
rect 3873 -16400 3919 -16388
rect 4051 -16132 4097 -16120
rect 4051 -16388 4057 -16132
rect 4091 -16388 4097 -16132
rect 4051 -16400 4097 -16388
rect -2105 -16438 -2029 -16432
rect -2105 -16472 -2089 -16438
rect -2045 -16472 -2029 -16438
rect -2105 -16488 -2029 -16472
rect -1927 -16438 -1851 -16432
rect -1927 -16472 -1911 -16438
rect -1867 -16472 -1851 -16438
rect -1927 -16488 -1851 -16472
rect -1906 -16542 -1872 -16488
rect -1927 -16595 -1917 -16542
rect -1864 -16595 -1854 -16542
rect -1817 -16665 -1783 -16400
rect -1749 -16438 -1673 -16432
rect -1749 -16472 -1733 -16438
rect -1689 -16472 -1673 -16438
rect -1749 -16488 -1673 -16472
rect -1571 -16438 -1495 -16432
rect -1571 -16472 -1555 -16438
rect -1511 -16472 -1495 -16438
rect -1571 -16488 -1495 -16472
rect -1728 -16542 -1694 -16488
rect -1550 -16541 -1516 -16488
rect -1748 -16595 -1738 -16542
rect -1685 -16595 -1675 -16542
rect -1571 -16594 -1561 -16541
rect -1508 -16594 -1498 -16541
rect -1837 -16718 -1827 -16665
rect -1774 -16718 -1764 -16665
rect -1461 -16666 -1427 -16400
rect -1393 -16438 -1317 -16432
rect -1393 -16472 -1377 -16438
rect -1333 -16472 -1317 -16438
rect -1393 -16488 -1317 -16472
rect -1215 -16438 -1139 -16432
rect -1215 -16472 -1199 -16438
rect -1155 -16472 -1139 -16438
rect -1215 -16488 -1139 -16472
rect -1372 -16543 -1338 -16488
rect -1194 -16542 -1160 -16488
rect -1391 -16596 -1381 -16543
rect -1328 -16596 -1318 -16543
rect -1214 -16595 -1204 -16542
rect -1151 -16595 -1141 -16542
rect -1104 -16665 -1070 -16400
rect -1037 -16438 -961 -16432
rect -1037 -16472 -1021 -16438
rect -977 -16472 -961 -16438
rect -1037 -16488 -961 -16472
rect -859 -16438 -783 -16432
rect -859 -16472 -843 -16438
rect -799 -16472 -783 -16438
rect -859 -16488 -783 -16472
rect -1016 -16542 -982 -16488
rect -1036 -16595 -1026 -16542
rect -973 -16595 -963 -16542
rect -749 -16664 -715 -16400
rect -681 -16438 -605 -16432
rect -681 -16472 -665 -16438
rect -621 -16472 -605 -16438
rect -681 -16488 -605 -16472
rect -503 -16438 -427 -16432
rect -503 -16472 -487 -16438
rect -443 -16472 -427 -16438
rect -503 -16488 -427 -16472
rect -1481 -16719 -1471 -16666
rect -1418 -16719 -1408 -16666
rect -1124 -16718 -1114 -16665
rect -1061 -16718 -1051 -16665
rect -769 -16717 -759 -16664
rect -706 -16717 -696 -16664
rect -393 -16665 -359 -16400
rect -325 -16438 -249 -16432
rect -325 -16472 -309 -16438
rect -265 -16472 -249 -16438
rect -325 -16488 -249 -16472
rect -147 -16438 -71 -16432
rect -147 -16472 -131 -16438
rect -87 -16472 -71 -16438
rect -147 -16488 -71 -16472
rect -37 -16665 -3 -16400
rect 31 -16438 107 -16432
rect 31 -16472 47 -16438
rect 91 -16472 107 -16438
rect 31 -16488 107 -16472
rect 209 -16438 285 -16432
rect 209 -16472 225 -16438
rect 269 -16472 285 -16438
rect 209 -16488 285 -16472
rect 230 -16542 264 -16488
rect 210 -16595 220 -16542
rect 273 -16595 283 -16542
rect -413 -16718 -403 -16665
rect -350 -16718 -340 -16665
rect -57 -16718 -47 -16665
rect 6 -16718 16 -16665
rect 319 -16666 353 -16400
rect 387 -16438 463 -16432
rect 387 -16472 403 -16438
rect 447 -16472 463 -16438
rect 387 -16488 463 -16472
rect 565 -16438 641 -16432
rect 565 -16472 581 -16438
rect 625 -16472 641 -16438
rect 565 -16488 641 -16472
rect 408 -16542 442 -16488
rect 586 -16542 620 -16488
rect 387 -16595 397 -16542
rect 450 -16595 460 -16542
rect 566 -16595 576 -16542
rect 629 -16595 639 -16542
rect 675 -16665 709 -16400
rect 743 -16438 819 -16432
rect 743 -16472 759 -16438
rect 803 -16472 819 -16438
rect 743 -16488 819 -16472
rect 921 -16438 997 -16432
rect 921 -16472 937 -16438
rect 981 -16472 997 -16438
rect 921 -16488 997 -16472
rect 765 -16542 799 -16488
rect 943 -16542 977 -16488
rect 745 -16595 755 -16542
rect 808 -16595 818 -16542
rect 923 -16595 933 -16542
rect 986 -16595 996 -16542
rect 1031 -16665 1065 -16400
rect 1099 -16438 1175 -16432
rect 1099 -16472 1115 -16438
rect 1159 -16472 1175 -16438
rect 1099 -16488 1175 -16472
rect 1277 -16438 1353 -16432
rect 1277 -16472 1293 -16438
rect 1337 -16472 1353 -16438
rect 1277 -16488 1353 -16472
rect 1120 -16542 1154 -16488
rect 1101 -16595 1111 -16542
rect 1164 -16595 1174 -16542
rect 1387 -16665 1421 -16400
rect 1455 -16438 1531 -16432
rect 1455 -16472 1471 -16438
rect 1515 -16472 1531 -16438
rect 1455 -16488 1531 -16472
rect 1633 -16438 1709 -16432
rect 1633 -16472 1649 -16438
rect 1693 -16472 1709 -16438
rect 1633 -16488 1709 -16472
rect 1744 -16665 1778 -16400
rect 1811 -16438 1887 -16432
rect 1811 -16472 1827 -16438
rect 1871 -16472 1887 -16438
rect 1811 -16488 1887 -16472
rect 1989 -16438 2065 -16432
rect 1989 -16472 2005 -16438
rect 2049 -16472 2065 -16438
rect 1989 -16488 2065 -16472
rect 2100 -16664 2134 -16400
rect 2167 -16438 2243 -16432
rect 2167 -16472 2183 -16438
rect 2227 -16472 2243 -16438
rect 2167 -16488 2243 -16472
rect 2345 -16438 2421 -16432
rect 2345 -16472 2361 -16438
rect 2405 -16472 2421 -16438
rect 2345 -16488 2421 -16472
rect 2366 -16542 2400 -16488
rect 2346 -16595 2356 -16542
rect 2409 -16595 2419 -16542
rect 299 -16719 309 -16666
rect 362 -16719 372 -16666
rect 655 -16718 665 -16665
rect 718 -16718 728 -16665
rect 835 -16718 845 -16665
rect 898 -16718 908 -16665
rect 1011 -16718 1021 -16665
rect 1074 -16718 1084 -16665
rect 1367 -16718 1377 -16665
rect 1430 -16718 1440 -16665
rect 1725 -16718 1735 -16665
rect 1788 -16718 1798 -16665
rect 2080 -16717 2090 -16664
rect 2143 -16717 2153 -16664
rect 2455 -16665 2489 -16400
rect 2523 -16438 2599 -16432
rect 2523 -16472 2539 -16438
rect 2583 -16472 2599 -16438
rect 2523 -16488 2599 -16472
rect 2701 -16438 2777 -16432
rect 2701 -16472 2717 -16438
rect 2761 -16472 2777 -16438
rect 2701 -16488 2777 -16472
rect 2544 -16542 2578 -16488
rect 2722 -16541 2756 -16488
rect 2524 -16595 2534 -16542
rect 2587 -16595 2597 -16542
rect 2703 -16594 2713 -16541
rect 2766 -16594 2776 -16541
rect 2811 -16665 2845 -16400
rect 2879 -16438 2955 -16432
rect 2879 -16472 2895 -16438
rect 2939 -16472 2955 -16438
rect 2879 -16488 2955 -16472
rect 3057 -16438 3133 -16432
rect 3057 -16472 3073 -16438
rect 3117 -16472 3133 -16438
rect 3057 -16488 3133 -16472
rect 2901 -16542 2935 -16488
rect 3079 -16542 3113 -16488
rect 2881 -16595 2891 -16542
rect 2944 -16595 2954 -16542
rect 3060 -16595 3070 -16542
rect 3123 -16595 3133 -16542
rect 3167 -16664 3201 -16400
rect 3235 -16438 3311 -16432
rect 3235 -16472 3251 -16438
rect 3295 -16472 3311 -16438
rect 3235 -16488 3311 -16472
rect 3413 -16438 3489 -16432
rect 3413 -16472 3429 -16438
rect 3473 -16472 3489 -16438
rect 3413 -16488 3489 -16472
rect 3257 -16542 3291 -16488
rect 3239 -16595 3249 -16542
rect 3302 -16595 3312 -16542
rect 2435 -16718 2445 -16665
rect 2498 -16718 2508 -16665
rect 2791 -16718 2801 -16665
rect 2854 -16718 2864 -16665
rect 3147 -16717 3157 -16664
rect 3210 -16717 3220 -16664
rect 3524 -16666 3558 -16400
rect 3591 -16438 3667 -16432
rect 3591 -16472 3607 -16438
rect 3651 -16472 3667 -16438
rect 3591 -16488 3667 -16472
rect 3769 -16438 3845 -16432
rect 3769 -16472 3785 -16438
rect 3829 -16472 3845 -16438
rect 3769 -16488 3845 -16472
rect 3879 -16665 3913 -16400
rect 3947 -16438 4023 -16432
rect 3947 -16472 3963 -16438
rect 4007 -16472 4023 -16438
rect 3947 -16488 4023 -16472
rect 4238 -16542 4291 -15592
rect 5021 -15593 5031 -15540
rect 5084 -15593 5094 -15540
rect 4228 -16595 4238 -16542
rect 4291 -16595 4301 -16542
rect -4802 -17171 -4792 -17118
rect -4739 -17171 -4729 -17118
rect -3945 -17170 -3935 -17118
rect -3883 -17170 -3873 -17118
rect 846 -17251 899 -16718
rect 3504 -16719 3514 -16666
rect 3567 -16719 3577 -16666
rect 3858 -16718 3868 -16665
rect 3921 -16718 3931 -16665
rect 5031 -16782 5084 -15593
rect 5400 -15653 5453 -13598
rect 5534 -13672 5587 -13349
rect 5524 -13725 5534 -13672
rect 5587 -13725 5597 -13672
rect 6912 -13922 6946 -12074
rect 8425 -12554 8627 -12548
rect 8425 -12732 8437 -12554
rect 8615 -12732 8627 -12554
rect 8425 -12738 8627 -12732
rect 11425 -12554 11627 -12548
rect 11425 -12732 11437 -12554
rect 11615 -12732 11627 -12554
rect 11425 -12738 11627 -12732
rect 8940 -13486 8950 -13433
rect 9003 -13486 9013 -13433
rect 9295 -13486 9305 -13433
rect 9358 -13486 9368 -13433
rect 8762 -13609 8772 -13556
rect 8825 -13609 8835 -13556
rect 7516 -13725 7526 -13672
rect 7579 -13725 7589 -13672
rect 7338 -13849 7348 -13796
rect 7401 -13849 7411 -13796
rect 5823 -13975 5833 -13922
rect 5886 -13975 5896 -13922
rect 6003 -13975 6013 -13922
rect 6066 -13975 6076 -13922
rect 5843 -14032 5877 -13975
rect 6022 -14032 6056 -13975
rect 6180 -13976 6190 -13923
rect 6243 -13976 6253 -13923
rect 6359 -13975 6369 -13922
rect 6422 -13975 6432 -13922
rect 6200 -14032 6234 -13976
rect 6378 -14032 6412 -13975
rect 6537 -13976 6547 -13923
rect 6600 -13976 6610 -13923
rect 6715 -13975 6725 -13922
rect 6778 -13975 6788 -13922
rect 6892 -13975 6902 -13922
rect 6955 -13975 6965 -13922
rect 6556 -14032 6590 -13976
rect 6734 -14032 6768 -13975
rect 6912 -14032 6946 -13975
rect 5645 -14048 5721 -14032
rect 5823 -14048 5899 -14032
rect 5577 -14082 5661 -14048
rect 5705 -14082 5790 -14048
rect 5577 -14120 5611 -14082
rect 5645 -14088 5721 -14082
rect 5756 -14120 5790 -14082
rect 5823 -14082 5839 -14048
rect 5883 -14082 5899 -14048
rect 5823 -14088 5899 -14082
rect 6001 -14048 6077 -14032
rect 6001 -14082 6017 -14048
rect 6061 -14082 6077 -14048
rect 6001 -14088 6077 -14082
rect 6179 -14048 6255 -14032
rect 6179 -14082 6195 -14048
rect 6239 -14082 6255 -14048
rect 6179 -14088 6255 -14082
rect 6357 -14048 6433 -14032
rect 6357 -14082 6373 -14048
rect 6417 -14082 6433 -14048
rect 6357 -14088 6433 -14082
rect 6535 -14048 6611 -14032
rect 6535 -14082 6551 -14048
rect 6595 -14082 6611 -14048
rect 6535 -14088 6611 -14082
rect 6713 -14048 6789 -14032
rect 6713 -14082 6729 -14048
rect 6773 -14082 6789 -14048
rect 6713 -14088 6789 -14082
rect 6891 -14048 6967 -14032
rect 6891 -14082 6907 -14048
rect 6951 -14082 6967 -14048
rect 6891 -14088 6967 -14082
rect 7069 -14048 7145 -14032
rect 7247 -14048 7323 -14032
rect 7069 -14082 7085 -14048
rect 7129 -14082 7263 -14048
rect 7307 -14082 7323 -14048
rect 7069 -14088 7145 -14082
rect 7179 -14120 7213 -14082
rect 7247 -14088 7323 -14082
rect 7357 -14120 7391 -13849
rect 7427 -13975 7437 -13922
rect 7490 -13975 7500 -13922
rect 7446 -14032 7480 -13975
rect 7425 -14048 7501 -14032
rect 7425 -14082 7441 -14048
rect 7485 -14082 7501 -14048
rect 7425 -14088 7501 -14082
rect 7535 -14120 7569 -13725
rect 7872 -13726 7882 -13673
rect 7935 -13726 7945 -13673
rect 8228 -13724 8238 -13671
rect 8291 -13724 8301 -13671
rect 7694 -13848 7704 -13795
rect 7757 -13848 7767 -13795
rect 7605 -13975 7615 -13922
rect 7668 -13975 7678 -13922
rect 7624 -14032 7658 -13975
rect 7603 -14048 7679 -14032
rect 7603 -14082 7619 -14048
rect 7663 -14082 7679 -14048
rect 7603 -14088 7679 -14082
rect 7713 -14120 7747 -13848
rect 7783 -13976 7793 -13923
rect 7846 -13976 7856 -13923
rect 7802 -14032 7836 -13976
rect 7781 -14048 7857 -14032
rect 7781 -14082 7797 -14048
rect 7841 -14082 7857 -14048
rect 7781 -14088 7857 -14082
rect 7892 -14120 7926 -13726
rect 8051 -13849 8061 -13796
rect 8114 -13849 8124 -13796
rect 7960 -13975 7970 -13922
rect 8023 -13975 8033 -13922
rect 7980 -14032 8014 -13975
rect 7959 -14048 8035 -14032
rect 7959 -14082 7975 -14048
rect 8019 -14082 8035 -14048
rect 7959 -14088 8035 -14082
rect 8069 -14120 8103 -13849
rect 8138 -13975 8148 -13922
rect 8201 -13975 8211 -13922
rect 8158 -14032 8192 -13975
rect 8137 -14048 8213 -14032
rect 8137 -14082 8153 -14048
rect 8197 -14082 8213 -14048
rect 8137 -14088 8213 -14082
rect 8248 -14120 8282 -13724
rect 8405 -13849 8415 -13796
rect 8468 -13849 8478 -13796
rect 8316 -13975 8326 -13922
rect 8379 -13975 8389 -13922
rect 8336 -14032 8370 -13975
rect 8315 -14048 8391 -14032
rect 8315 -14082 8331 -14048
rect 8375 -14082 8391 -14048
rect 8315 -14088 8391 -14082
rect 8425 -14120 8459 -13849
rect 8493 -14048 8569 -14032
rect 8671 -14048 8747 -14032
rect 8493 -14082 8509 -14048
rect 8553 -14082 8687 -14048
rect 8731 -14082 8747 -14048
rect 8493 -14088 8569 -14082
rect 8603 -14120 8637 -14082
rect 8671 -14088 8747 -14082
rect 8781 -14120 8815 -13609
rect 8851 -13975 8861 -13922
rect 8914 -13975 8924 -13922
rect 8871 -14032 8905 -13975
rect 8849 -14048 8925 -14032
rect 8849 -14082 8865 -14048
rect 8909 -14082 8925 -14048
rect 8849 -14088 8925 -14082
rect 8960 -14120 8994 -13486
rect 9117 -13609 9127 -13556
rect 9180 -13609 9190 -13556
rect 9028 -13975 9038 -13922
rect 9091 -13975 9101 -13922
rect 9048 -14032 9082 -13975
rect 9027 -14048 9103 -14032
rect 9027 -14082 9043 -14048
rect 9087 -14082 9103 -14048
rect 9027 -14088 9103 -14082
rect 9137 -14120 9171 -13609
rect 9207 -13975 9217 -13922
rect 9270 -13975 9280 -13922
rect 9227 -14032 9261 -13975
rect 9205 -14048 9281 -14032
rect 9205 -14082 9221 -14048
rect 9265 -14082 9281 -14048
rect 9205 -14088 9281 -14082
rect 9315 -14120 9349 -13486
rect 9473 -13609 9483 -13556
rect 9536 -13609 9546 -13556
rect 9384 -13975 9394 -13922
rect 9447 -13975 9457 -13922
rect 9404 -14032 9438 -13975
rect 9383 -14048 9459 -14032
rect 9383 -14082 9399 -14048
rect 9443 -14082 9459 -14048
rect 9383 -14088 9459 -14082
rect 9493 -14120 9527 -13609
rect 11432 -13725 11442 -13672
rect 11495 -13725 11505 -13672
rect 11788 -13725 11798 -13672
rect 11851 -13725 11861 -13672
rect 11254 -13849 11264 -13796
rect 11317 -13849 11327 -13796
rect 9919 -13976 9929 -13923
rect 9982 -13976 9992 -13923
rect 10098 -13975 10108 -13922
rect 10161 -13975 10171 -13922
rect 9938 -14032 9972 -13976
rect 10117 -14032 10151 -13975
rect 10274 -13976 10284 -13923
rect 10337 -13976 10347 -13923
rect 10452 -13976 10462 -13923
rect 10515 -13976 10525 -13923
rect 10630 -13975 10640 -13922
rect 10693 -13975 10703 -13922
rect 10294 -14032 10328 -13976
rect 10472 -14032 10506 -13976
rect 10650 -14032 10684 -13975
rect 10809 -13976 10819 -13923
rect 10872 -13976 10882 -13923
rect 10828 -14032 10862 -13976
rect 9561 -14048 9637 -14032
rect 9739 -14048 9815 -14032
rect 9561 -14082 9577 -14048
rect 9621 -14082 9755 -14048
rect 9799 -14082 9815 -14048
rect 9561 -14088 9637 -14082
rect 9671 -14120 9705 -14082
rect 9739 -14088 9815 -14082
rect 9917 -14048 9993 -14032
rect 9917 -14082 9933 -14048
rect 9977 -14082 9993 -14048
rect 9917 -14088 9993 -14082
rect 10095 -14048 10171 -14032
rect 10095 -14082 10111 -14048
rect 10155 -14082 10171 -14048
rect 10095 -14088 10171 -14082
rect 10273 -14048 10349 -14032
rect 10273 -14082 10289 -14048
rect 10333 -14082 10349 -14048
rect 10273 -14088 10349 -14082
rect 10451 -14048 10527 -14032
rect 10451 -14082 10467 -14048
rect 10511 -14082 10527 -14048
rect 10451 -14088 10527 -14082
rect 10629 -14048 10705 -14032
rect 10629 -14082 10645 -14048
rect 10689 -14082 10705 -14048
rect 10629 -14088 10705 -14082
rect 10807 -14048 10883 -14032
rect 10807 -14082 10823 -14048
rect 10867 -14082 10883 -14048
rect 10807 -14088 10883 -14082
rect 10985 -14048 11061 -14032
rect 11163 -14048 11239 -14032
rect 10985 -14082 11001 -14048
rect 11045 -14082 11179 -14048
rect 11223 -14082 11239 -14048
rect 10985 -14088 11061 -14082
rect 11095 -14120 11129 -14082
rect 11163 -14088 11239 -14082
rect 11273 -14120 11307 -13849
rect 11343 -13975 11353 -13922
rect 11406 -13975 11416 -13922
rect 11362 -14032 11396 -13975
rect 11341 -14048 11417 -14032
rect 11341 -14082 11357 -14048
rect 11401 -14082 11417 -14048
rect 11341 -14088 11417 -14082
rect 11452 -14120 11486 -13725
rect 11610 -13850 11620 -13797
rect 11673 -13850 11683 -13797
rect 11520 -13975 11530 -13922
rect 11583 -13975 11593 -13922
rect 11540 -14032 11574 -13975
rect 11519 -14048 11595 -14032
rect 11519 -14082 11535 -14048
rect 11579 -14082 11595 -14048
rect 11519 -14088 11595 -14082
rect 11630 -14120 11664 -13850
rect 11699 -13975 11709 -13922
rect 11762 -13975 11772 -13922
rect 11719 -14032 11753 -13975
rect 11697 -14048 11773 -14032
rect 11697 -14082 11713 -14048
rect 11757 -14082 11773 -14048
rect 11697 -14088 11773 -14082
rect 11807 -14120 11841 -13725
rect 12142 -13726 12152 -13673
rect 12205 -13726 12215 -13673
rect 12499 -13725 12509 -13672
rect 12562 -13725 12572 -13672
rect 11967 -13849 11977 -13796
rect 12030 -13849 12040 -13796
rect 11876 -13976 11886 -13923
rect 11939 -13976 11949 -13923
rect 11895 -14032 11929 -13976
rect 11875 -14048 11951 -14032
rect 11875 -14082 11891 -14048
rect 11935 -14082 11951 -14048
rect 11875 -14088 11951 -14082
rect 11986 -14120 12020 -13849
rect 12054 -13975 12064 -13922
rect 12117 -13975 12127 -13922
rect 12073 -14032 12107 -13975
rect 12053 -14048 12129 -14032
rect 12053 -14082 12069 -14048
rect 12113 -14082 12129 -14048
rect 12053 -14088 12129 -14082
rect 12162 -14120 12196 -13726
rect 12324 -13849 12334 -13796
rect 12387 -13849 12397 -13796
rect 12232 -13976 12242 -13923
rect 12295 -13976 12305 -13923
rect 12252 -14032 12286 -13976
rect 12231 -14048 12307 -14032
rect 12231 -14082 12247 -14048
rect 12291 -14082 12307 -14048
rect 12231 -14088 12307 -14082
rect 12342 -14120 12376 -13849
rect 12410 -13975 12420 -13922
rect 12473 -13975 12483 -13922
rect 12430 -14032 12464 -13975
rect 12409 -14048 12485 -14032
rect 12409 -14082 12425 -14048
rect 12469 -14082 12485 -14048
rect 12409 -14088 12485 -14082
rect 12519 -14048 12553 -13725
rect 12587 -14048 12663 -14032
rect 12519 -14082 12603 -14048
rect 12647 -14082 12731 -14048
rect 12519 -14120 12553 -14082
rect 12587 -14088 12663 -14082
rect 12697 -14120 12731 -14082
rect 5571 -14132 5617 -14120
rect 5571 -14388 5577 -14132
rect 5611 -14388 5617 -14132
rect 5571 -14400 5617 -14388
rect 5749 -14132 5795 -14120
rect 5749 -14388 5755 -14132
rect 5789 -14388 5795 -14132
rect 5749 -14400 5795 -14388
rect 5927 -14132 5973 -14120
rect 5927 -14388 5933 -14132
rect 5967 -14388 5973 -14132
rect 5927 -14400 5973 -14388
rect 6105 -14132 6151 -14120
rect 6105 -14388 6111 -14132
rect 6145 -14388 6151 -14132
rect 6105 -14400 6151 -14388
rect 6283 -14132 6329 -14120
rect 6283 -14388 6289 -14132
rect 6323 -14388 6329 -14132
rect 6283 -14400 6329 -14388
rect 6461 -14132 6507 -14120
rect 6461 -14388 6467 -14132
rect 6501 -14388 6507 -14132
rect 6461 -14400 6507 -14388
rect 6639 -14132 6685 -14120
rect 6639 -14388 6645 -14132
rect 6679 -14388 6685 -14132
rect 6639 -14400 6685 -14388
rect 6817 -14132 6863 -14120
rect 6817 -14388 6823 -14132
rect 6857 -14388 6863 -14132
rect 6817 -14400 6863 -14388
rect 6995 -14132 7041 -14120
rect 6995 -14388 7001 -14132
rect 7035 -14388 7041 -14132
rect 6995 -14400 7041 -14388
rect 7173 -14132 7219 -14120
rect 7173 -14388 7179 -14132
rect 7213 -14388 7219 -14132
rect 7173 -14400 7219 -14388
rect 7351 -14132 7397 -14120
rect 7351 -14388 7357 -14132
rect 7391 -14388 7397 -14132
rect 7351 -14400 7397 -14388
rect 7529 -14132 7575 -14120
rect 7529 -14388 7535 -14132
rect 7569 -14388 7575 -14132
rect 7529 -14400 7575 -14388
rect 7707 -14132 7753 -14120
rect 7707 -14388 7713 -14132
rect 7747 -14388 7753 -14132
rect 7707 -14400 7753 -14388
rect 7885 -14132 7931 -14120
rect 7885 -14388 7891 -14132
rect 7925 -14388 7931 -14132
rect 7885 -14400 7931 -14388
rect 8063 -14132 8109 -14120
rect 8063 -14388 8069 -14132
rect 8103 -14388 8109 -14132
rect 8063 -14400 8109 -14388
rect 8241 -14132 8287 -14120
rect 8241 -14388 8247 -14132
rect 8281 -14388 8287 -14132
rect 8241 -14400 8287 -14388
rect 8419 -14132 8465 -14120
rect 8419 -14388 8425 -14132
rect 8459 -14388 8465 -14132
rect 8419 -14400 8465 -14388
rect 8597 -14132 8643 -14120
rect 8597 -14388 8603 -14132
rect 8637 -14388 8643 -14132
rect 8597 -14400 8643 -14388
rect 8775 -14132 8821 -14120
rect 8775 -14388 8781 -14132
rect 8815 -14388 8821 -14132
rect 8775 -14400 8821 -14388
rect 8953 -14132 8999 -14120
rect 8953 -14388 8959 -14132
rect 8993 -14388 8999 -14132
rect 8953 -14400 8999 -14388
rect 9131 -14132 9177 -14120
rect 9131 -14388 9137 -14132
rect 9171 -14388 9177 -14132
rect 9131 -14400 9177 -14388
rect 9309 -14132 9355 -14120
rect 9309 -14388 9315 -14132
rect 9349 -14388 9355 -14132
rect 9309 -14400 9355 -14388
rect 9487 -14132 9533 -14120
rect 9487 -14388 9493 -14132
rect 9527 -14388 9533 -14132
rect 9487 -14400 9533 -14388
rect 9665 -14132 9711 -14120
rect 9665 -14388 9671 -14132
rect 9705 -14388 9711 -14132
rect 9665 -14400 9711 -14388
rect 9843 -14132 9889 -14120
rect 9843 -14388 9849 -14132
rect 9883 -14388 9889 -14132
rect 9843 -14400 9889 -14388
rect 10021 -14132 10067 -14120
rect 10021 -14388 10027 -14132
rect 10061 -14388 10067 -14132
rect 10021 -14400 10067 -14388
rect 10199 -14132 10245 -14120
rect 10199 -14388 10205 -14132
rect 10239 -14388 10245 -14132
rect 10199 -14400 10245 -14388
rect 10377 -14132 10423 -14120
rect 10377 -14388 10383 -14132
rect 10417 -14388 10423 -14132
rect 10377 -14400 10423 -14388
rect 10555 -14132 10601 -14120
rect 10555 -14388 10561 -14132
rect 10595 -14388 10601 -14132
rect 10555 -14400 10601 -14388
rect 10733 -14132 10779 -14120
rect 10733 -14388 10739 -14132
rect 10773 -14388 10779 -14132
rect 10733 -14400 10779 -14388
rect 10911 -14132 10957 -14120
rect 10911 -14388 10917 -14132
rect 10951 -14388 10957 -14132
rect 10911 -14400 10957 -14388
rect 11089 -14132 11135 -14120
rect 11089 -14388 11095 -14132
rect 11129 -14388 11135 -14132
rect 11089 -14400 11135 -14388
rect 11267 -14132 11313 -14120
rect 11267 -14388 11273 -14132
rect 11307 -14388 11313 -14132
rect 11267 -14400 11313 -14388
rect 11445 -14132 11491 -14120
rect 11445 -14388 11451 -14132
rect 11485 -14388 11491 -14132
rect 11445 -14400 11491 -14388
rect 11623 -14132 11669 -14120
rect 11623 -14388 11629 -14132
rect 11663 -14388 11669 -14132
rect 11623 -14400 11669 -14388
rect 11801 -14132 11847 -14120
rect 11801 -14388 11807 -14132
rect 11841 -14388 11847 -14132
rect 11801 -14400 11847 -14388
rect 11979 -14132 12025 -14120
rect 11979 -14388 11985 -14132
rect 12019 -14388 12025 -14132
rect 11979 -14400 12025 -14388
rect 12157 -14132 12203 -14120
rect 12157 -14388 12163 -14132
rect 12197 -14388 12203 -14132
rect 12157 -14400 12203 -14388
rect 12335 -14132 12381 -14120
rect 12335 -14388 12341 -14132
rect 12375 -14388 12381 -14132
rect 12335 -14400 12381 -14388
rect 12513 -14132 12559 -14120
rect 12513 -14388 12519 -14132
rect 12553 -14388 12559 -14132
rect 12513 -14400 12559 -14388
rect 12691 -14132 12737 -14120
rect 12691 -14388 12697 -14132
rect 12731 -14388 12737 -14132
rect 12691 -14400 12737 -14388
rect 5645 -14438 5721 -14432
rect 5645 -14472 5661 -14438
rect 5705 -14472 5721 -14438
rect 5645 -14488 5721 -14472
rect 5756 -14545 5790 -14400
rect 5823 -14438 5899 -14432
rect 5823 -14472 5839 -14438
rect 5883 -14472 5899 -14438
rect 5823 -14488 5899 -14472
rect 5736 -14598 5746 -14545
rect 5799 -14598 5809 -14545
rect 5843 -15032 5877 -14488
rect 5933 -14658 5967 -14400
rect 6001 -14438 6077 -14432
rect 6001 -14472 6017 -14438
rect 6061 -14472 6077 -14438
rect 6001 -14488 6077 -14472
rect 5914 -14711 5924 -14658
rect 5977 -14711 5987 -14658
rect 6022 -15032 6056 -14488
rect 6111 -14545 6145 -14400
rect 6179 -14438 6255 -14432
rect 6179 -14472 6195 -14438
rect 6239 -14472 6255 -14438
rect 6179 -14488 6255 -14472
rect 6091 -14598 6101 -14545
rect 6154 -14598 6164 -14545
rect 6200 -15032 6234 -14488
rect 6289 -14658 6323 -14400
rect 6357 -14438 6433 -14432
rect 6357 -14472 6373 -14438
rect 6417 -14472 6433 -14438
rect 6357 -14488 6433 -14472
rect 6269 -14711 6279 -14658
rect 6332 -14711 6342 -14658
rect 6378 -15032 6412 -14488
rect 6468 -14545 6502 -14400
rect 6535 -14438 6611 -14432
rect 6535 -14472 6551 -14438
rect 6595 -14472 6611 -14438
rect 6535 -14488 6611 -14472
rect 6449 -14598 6459 -14545
rect 6512 -14598 6522 -14545
rect 6557 -15032 6591 -14488
rect 6645 -14658 6679 -14400
rect 6713 -14438 6789 -14432
rect 6713 -14472 6729 -14438
rect 6773 -14472 6789 -14438
rect 6713 -14488 6789 -14472
rect 6823 -14545 6857 -14400
rect 6891 -14438 6967 -14432
rect 6891 -14472 6907 -14438
rect 6951 -14472 6967 -14438
rect 6891 -14488 6967 -14472
rect 6803 -14598 6813 -14545
rect 6866 -14598 6876 -14545
rect 7000 -14658 7034 -14400
rect 7069 -14438 7145 -14432
rect 7069 -14472 7085 -14438
rect 7129 -14472 7145 -14438
rect 7069 -14488 7145 -14472
rect 6626 -14711 6636 -14658
rect 6689 -14711 6699 -14658
rect 6981 -14711 6991 -14658
rect 7044 -14711 7054 -14658
rect 7179 -14749 7213 -14400
rect 7247 -14438 7323 -14432
rect 7247 -14472 7263 -14438
rect 7307 -14472 7323 -14438
rect 7247 -14488 7323 -14472
rect 6822 -14783 7213 -14749
rect 5645 -15047 5721 -15032
rect 5575 -15048 5789 -15047
rect 5575 -15081 5661 -15048
rect 5575 -15120 5609 -15081
rect 5645 -15082 5661 -15081
rect 5705 -15081 5789 -15048
rect 5705 -15082 5721 -15081
rect 5645 -15088 5721 -15082
rect 5755 -15120 5789 -15081
rect 5823 -15048 5899 -15032
rect 5823 -15082 5839 -15048
rect 5883 -15082 5899 -15048
rect 5823 -15088 5899 -15082
rect 6001 -15048 6077 -15032
rect 6001 -15082 6017 -15048
rect 6061 -15082 6077 -15048
rect 6001 -15088 6077 -15082
rect 6179 -15048 6255 -15032
rect 6179 -15082 6195 -15048
rect 6239 -15082 6255 -15048
rect 6179 -15088 6255 -15082
rect 6357 -15048 6433 -15032
rect 6357 -15082 6373 -15048
rect 6417 -15082 6433 -15048
rect 6357 -15088 6433 -15082
rect 6535 -15048 6611 -15032
rect 6535 -15082 6551 -15048
rect 6595 -15082 6611 -15048
rect 6535 -15088 6611 -15082
rect 6713 -15048 6789 -15032
rect 6713 -15082 6729 -15048
rect 6773 -15082 6789 -15048
rect 6713 -15088 6789 -15082
rect 6822 -15120 6856 -14783
rect 7357 -14824 7391 -14400
rect 7425 -14438 7501 -14432
rect 7425 -14472 7441 -14438
rect 7485 -14472 7501 -14438
rect 7425 -14488 7501 -14472
rect 6983 -14877 6993 -14824
rect 7046 -14877 7056 -14824
rect 7337 -14877 7347 -14824
rect 7400 -14877 7410 -14824
rect 6891 -15048 6967 -15032
rect 6891 -15082 6907 -15048
rect 6951 -15082 6967 -15048
rect 6891 -15088 6967 -15082
rect 7002 -15120 7036 -14877
rect 7070 -14976 7080 -14923
rect 7133 -14976 7143 -14923
rect 7090 -15032 7124 -14976
rect 7250 -14977 7260 -14924
rect 7313 -14977 7323 -14924
rect 7269 -15032 7303 -14977
rect 7069 -15048 7145 -15032
rect 7069 -15082 7085 -15048
rect 7129 -15082 7145 -15048
rect 7069 -15088 7145 -15082
rect 7247 -15048 7323 -15032
rect 7247 -15082 7263 -15048
rect 7307 -15082 7323 -15048
rect 7247 -15088 7323 -15082
rect 7357 -15120 7391 -14877
rect 7447 -14923 7481 -14488
rect 7429 -14976 7439 -14923
rect 7492 -14976 7502 -14923
rect 7447 -15032 7481 -14976
rect 7425 -15048 7501 -15032
rect 7425 -15082 7441 -15048
rect 7485 -15082 7501 -15048
rect 7425 -15088 7501 -15082
rect 7535 -15120 7569 -14400
rect 7603 -14438 7679 -14432
rect 7603 -14472 7619 -14438
rect 7663 -14472 7679 -14438
rect 7603 -14488 7679 -14472
rect 7781 -14438 7857 -14432
rect 7781 -14472 7797 -14438
rect 7841 -14472 7857 -14438
rect 7781 -14488 7857 -14472
rect 7959 -14438 8035 -14432
rect 7959 -14472 7975 -14438
rect 8019 -14472 8035 -14438
rect 7959 -14488 8035 -14472
rect 8137 -14438 8213 -14432
rect 8137 -14472 8153 -14438
rect 8197 -14472 8213 -14438
rect 8137 -14488 8213 -14472
rect 8315 -14438 8391 -14432
rect 8315 -14472 8331 -14438
rect 8375 -14472 8391 -14438
rect 8315 -14488 8391 -14472
rect 8493 -14438 8569 -14432
rect 8493 -14472 8509 -14438
rect 8553 -14472 8569 -14438
rect 8493 -14488 8569 -14472
rect 8671 -14438 8747 -14432
rect 8671 -14472 8687 -14438
rect 8731 -14472 8747 -14438
rect 8671 -14488 8747 -14472
rect 8849 -14438 8925 -14432
rect 8849 -14472 8865 -14438
rect 8909 -14472 8925 -14438
rect 8849 -14488 8925 -14472
rect 9027 -14438 9103 -14432
rect 9027 -14472 9043 -14438
rect 9087 -14472 9103 -14438
rect 9027 -14488 9103 -14472
rect 9205 -14438 9281 -14432
rect 9205 -14472 9221 -14438
rect 9265 -14472 9281 -14438
rect 9205 -14488 9281 -14472
rect 9383 -14438 9459 -14432
rect 9383 -14472 9399 -14438
rect 9443 -14472 9459 -14438
rect 9383 -14488 9459 -14472
rect 9561 -14438 9637 -14432
rect 9561 -14472 9577 -14438
rect 9621 -14472 9637 -14438
rect 9561 -14488 9637 -14472
rect 9739 -14438 9815 -14432
rect 9739 -14472 9755 -14438
rect 9799 -14472 9815 -14438
rect 9739 -14488 9815 -14472
rect 7625 -15032 7659 -14488
rect 7694 -14878 7704 -14825
rect 7757 -14878 7767 -14825
rect 7603 -15048 7679 -15032
rect 7603 -15082 7619 -15048
rect 7663 -15082 7679 -15048
rect 7603 -15088 7679 -15082
rect 7714 -15120 7748 -14878
rect 7802 -15032 7836 -14488
rect 8226 -14598 8236 -14545
rect 8289 -14598 8299 -14545
rect 8050 -14874 8060 -14821
rect 8113 -14874 8123 -14821
rect 7781 -15048 7857 -15032
rect 7781 -15082 7797 -15048
rect 7841 -15082 7857 -15048
rect 7781 -15088 7857 -15082
rect 7959 -15048 8035 -15032
rect 7959 -15082 7975 -15048
rect 8019 -15082 8035 -15048
rect 7959 -15088 8035 -15082
rect 8069 -15120 8103 -14874
rect 8137 -15048 8213 -15032
rect 8137 -15082 8153 -15048
rect 8197 -15082 8213 -15048
rect 8137 -15088 8213 -15082
rect 8247 -15120 8281 -14598
rect 8336 -14923 8370 -14488
rect 8407 -14710 8417 -14657
rect 8470 -14710 8480 -14657
rect 8317 -14976 8327 -14923
rect 8380 -14976 8390 -14923
rect 8336 -15032 8370 -14976
rect 8315 -15048 8391 -15032
rect 8315 -15082 8331 -15048
rect 8375 -15082 8391 -15048
rect 8315 -15088 8391 -15082
rect 8426 -15120 8460 -14710
rect 8514 -14806 8548 -14488
rect 8585 -14598 8595 -14545
rect 8648 -14598 8658 -14545
rect 8494 -14859 8504 -14806
rect 8557 -14859 8567 -14806
rect 8514 -14871 8548 -14859
rect 8495 -14977 8505 -14924
rect 8558 -14977 8568 -14924
rect 8514 -15032 8548 -14977
rect 8493 -15048 8569 -15032
rect 8493 -15082 8509 -15048
rect 8553 -15082 8569 -15048
rect 8493 -15088 8569 -15082
rect 8604 -15120 8638 -14598
rect 8762 -14711 8772 -14658
rect 8825 -14711 8835 -14658
rect 8692 -14924 8726 -14923
rect 8673 -14977 8683 -14924
rect 8736 -14977 8746 -14924
rect 8692 -15032 8726 -14977
rect 8671 -15048 8747 -15032
rect 8671 -15082 8687 -15048
rect 8731 -15082 8747 -15048
rect 8671 -15088 8747 -15082
rect 8781 -15120 8815 -14711
rect 8870 -15032 8904 -14488
rect 8940 -14599 8950 -14546
rect 9003 -14599 9013 -14546
rect 8849 -15048 8925 -15032
rect 8849 -15082 8865 -15048
rect 8909 -15082 8925 -15048
rect 8849 -15088 8925 -15082
rect 8960 -15120 8994 -14599
rect 9048 -15032 9082 -14488
rect 9117 -14712 9127 -14659
rect 9180 -14712 9190 -14659
rect 9027 -15048 9103 -15032
rect 9027 -15082 9043 -15048
rect 9087 -15082 9103 -15048
rect 9027 -15088 9103 -15082
rect 9137 -15120 9171 -14712
rect 9226 -15032 9260 -14488
rect 9294 -14598 9304 -14545
rect 9357 -14598 9367 -14545
rect 9205 -15048 9281 -15032
rect 9205 -15082 9221 -15048
rect 9265 -15082 9281 -15048
rect 9205 -15088 9281 -15082
rect 9314 -15120 9348 -14598
rect 9404 -15032 9438 -14488
rect 9651 -14598 9661 -14545
rect 9714 -14598 9724 -14545
rect 9473 -14711 9483 -14658
rect 9536 -14711 9546 -14658
rect 9383 -15048 9459 -15032
rect 9383 -15082 9399 -15048
rect 9443 -15082 9459 -15048
rect 9383 -15088 9459 -15082
rect 9493 -15120 9527 -14711
rect 9562 -14976 9572 -14923
rect 9625 -14976 9635 -14923
rect 9582 -15032 9616 -14976
rect 9561 -15048 9637 -15032
rect 9561 -15082 9577 -15048
rect 9621 -15082 9637 -15048
rect 9561 -15088 9637 -15082
rect 9671 -15120 9705 -14598
rect 9763 -14806 9797 -14488
rect 9848 -14659 9882 -14400
rect 9917 -14438 9993 -14432
rect 9917 -14472 9933 -14438
rect 9977 -14472 9993 -14438
rect 9917 -14488 9993 -14472
rect 9827 -14712 9837 -14659
rect 9890 -14712 9900 -14659
rect 9743 -14859 9753 -14806
rect 9806 -14859 9816 -14806
rect 9763 -14871 9797 -14859
rect 9740 -14976 9750 -14923
rect 9803 -14976 9813 -14923
rect 9760 -15032 9794 -14976
rect 9739 -15048 9815 -15032
rect 9739 -15082 9755 -15048
rect 9799 -15082 9815 -15048
rect 9739 -15088 9815 -15082
rect 9848 -15120 9882 -14712
rect 9939 -14923 9973 -14488
rect 10026 -14545 10060 -14400
rect 10095 -14438 10171 -14432
rect 10095 -14472 10111 -14438
rect 10155 -14472 10171 -14438
rect 10095 -14488 10171 -14472
rect 10006 -14598 10016 -14545
rect 10069 -14598 10079 -14545
rect 9919 -14976 9929 -14923
rect 9982 -14976 9992 -14923
rect 9939 -15032 9973 -14976
rect 9917 -15048 9993 -15032
rect 9917 -15082 9933 -15048
rect 9977 -15082 9993 -15048
rect 9917 -15088 9993 -15082
rect 10026 -15120 10060 -14598
rect 10205 -14658 10239 -14400
rect 10273 -14438 10349 -14432
rect 10273 -14472 10289 -14438
rect 10333 -14472 10349 -14438
rect 10273 -14488 10349 -14472
rect 10383 -14546 10417 -14400
rect 10451 -14438 10527 -14432
rect 10451 -14472 10467 -14438
rect 10511 -14472 10527 -14438
rect 10451 -14488 10527 -14472
rect 10363 -14599 10373 -14546
rect 10426 -14599 10436 -14546
rect 10186 -14711 10196 -14658
rect 10249 -14711 10259 -14658
rect 10185 -14875 10195 -14822
rect 10248 -14875 10258 -14822
rect 10095 -15048 10171 -15032
rect 10095 -15082 10111 -15048
rect 10155 -15082 10171 -15048
rect 10095 -15088 10171 -15082
rect 10205 -15120 10239 -14875
rect 10472 -15032 10506 -14488
rect 10560 -14658 10594 -14400
rect 10629 -14438 10705 -14432
rect 10629 -14472 10645 -14438
rect 10689 -14472 10705 -14438
rect 10629 -14488 10705 -14472
rect 10540 -14711 10550 -14658
rect 10603 -14711 10613 -14658
rect 10542 -14868 10552 -14815
rect 10605 -14868 10615 -14815
rect 10273 -15048 10349 -15032
rect 10273 -15082 10289 -15048
rect 10333 -15082 10349 -15048
rect 10273 -15088 10349 -15082
rect 10451 -15048 10527 -15032
rect 10451 -15082 10467 -15048
rect 10511 -15082 10527 -15048
rect 10451 -15088 10527 -15082
rect 10561 -15120 10595 -14868
rect 10650 -15032 10684 -14488
rect 10738 -14545 10772 -14400
rect 10807 -14438 10883 -14432
rect 10807 -14472 10823 -14438
rect 10867 -14472 10883 -14438
rect 10807 -14488 10883 -14472
rect 10719 -14598 10729 -14545
rect 10782 -14598 10792 -14545
rect 10828 -14923 10862 -14488
rect 10917 -14658 10951 -14400
rect 10985 -14438 11061 -14432
rect 10985 -14472 11001 -14438
rect 11045 -14472 11061 -14438
rect 10985 -14488 11061 -14472
rect 11096 -14658 11130 -14400
rect 11163 -14438 11239 -14432
rect 11163 -14472 11179 -14438
rect 11223 -14472 11239 -14438
rect 11163 -14488 11239 -14472
rect 10898 -14711 10908 -14658
rect 10961 -14711 10971 -14658
rect 11077 -14711 11087 -14658
rect 11140 -14711 11150 -14658
rect 10898 -14866 10908 -14813
rect 10961 -14866 10971 -14813
rect 11273 -14815 11307 -14400
rect 11341 -14438 11417 -14432
rect 11341 -14472 11357 -14438
rect 11401 -14472 11417 -14438
rect 11341 -14488 11417 -14472
rect 11519 -14438 11595 -14432
rect 11519 -14472 11535 -14438
rect 11579 -14472 11595 -14438
rect 11519 -14488 11595 -14472
rect 11697 -14438 11773 -14432
rect 11697 -14472 11713 -14438
rect 11757 -14472 11773 -14438
rect 11697 -14488 11773 -14472
rect 11875 -14438 11951 -14432
rect 11875 -14472 11891 -14438
rect 11935 -14472 11951 -14438
rect 11875 -14488 11951 -14472
rect 12053 -14438 12129 -14432
rect 12053 -14472 12069 -14438
rect 12113 -14472 12129 -14438
rect 12053 -14488 12129 -14472
rect 12231 -14438 12307 -14432
rect 12231 -14472 12247 -14438
rect 12291 -14472 12307 -14438
rect 12231 -14488 12307 -14472
rect 12409 -14438 12485 -14432
rect 12409 -14472 12425 -14438
rect 12469 -14472 12485 -14438
rect 12409 -14488 12485 -14472
rect 12587 -14438 12663 -14432
rect 12587 -14472 12603 -14438
rect 12647 -14472 12663 -14438
rect 12587 -14488 12663 -14472
rect 11430 -14709 11440 -14656
rect 11493 -14709 11503 -14656
rect 10809 -14976 10819 -14923
rect 10872 -14976 10882 -14923
rect 10828 -15032 10862 -14976
rect 10629 -15048 10705 -15032
rect 10629 -15082 10645 -15048
rect 10689 -15082 10705 -15048
rect 10629 -15088 10705 -15082
rect 10807 -15048 10883 -15032
rect 10807 -15082 10823 -15048
rect 10867 -15082 10883 -15048
rect 10807 -15088 10883 -15082
rect 10916 -15120 10950 -14866
rect 11254 -14868 11264 -14815
rect 11317 -14868 11327 -14815
rect 10986 -14976 10996 -14923
rect 11049 -14976 11059 -14923
rect 11165 -14976 11175 -14923
rect 11228 -14976 11238 -14923
rect 11006 -15032 11040 -14976
rect 11184 -15032 11218 -14976
rect 10985 -15048 11061 -15032
rect 10985 -15082 11001 -15048
rect 11045 -15082 11061 -15048
rect 10985 -15088 11061 -15082
rect 11163 -15048 11239 -15032
rect 11163 -15082 11179 -15048
rect 11223 -15082 11239 -15048
rect 11163 -15088 11239 -15082
rect 11273 -15120 11307 -14868
rect 11341 -15048 11417 -15032
rect 11341 -15082 11357 -15048
rect 11401 -15082 11417 -15048
rect 11341 -15088 11417 -15082
rect 11451 -15120 11485 -14709
rect 11717 -15032 11751 -14488
rect 11897 -15032 11931 -14488
rect 12075 -15032 12109 -14488
rect 12253 -15032 12287 -14488
rect 12430 -15032 12464 -14488
rect 11519 -15048 11595 -15032
rect 11519 -15082 11535 -15048
rect 11579 -15082 11595 -15048
rect 11519 -15088 11595 -15082
rect 11697 -15048 11773 -15032
rect 11697 -15082 11713 -15048
rect 11757 -15082 11773 -15048
rect 11697 -15088 11773 -15082
rect 11875 -15048 11951 -15032
rect 11875 -15082 11891 -15048
rect 11935 -15082 11951 -15048
rect 11875 -15088 11951 -15082
rect 12053 -15048 12129 -15032
rect 12053 -15082 12069 -15048
rect 12113 -15082 12129 -15048
rect 12053 -15088 12129 -15082
rect 12231 -15048 12307 -15032
rect 12231 -15082 12247 -15048
rect 12291 -15082 12307 -15048
rect 12231 -15088 12307 -15082
rect 12409 -15048 12485 -15032
rect 12409 -15082 12425 -15048
rect 12469 -15082 12485 -15048
rect 12587 -15048 12663 -15032
rect 12587 -15049 12603 -15048
rect 12409 -15088 12485 -15082
rect 12520 -15082 12603 -15049
rect 12647 -15049 12663 -15048
rect 12647 -15082 12730 -15049
rect 12520 -15083 12730 -15082
rect 12520 -15120 12554 -15083
rect 12587 -15088 12663 -15083
rect 12696 -15120 12730 -15083
rect 5571 -15132 5617 -15120
rect 5571 -15388 5577 -15132
rect 5611 -15388 5617 -15132
rect 5571 -15400 5617 -15388
rect 5749 -15132 5795 -15120
rect 5749 -15388 5755 -15132
rect 5789 -15388 5795 -15132
rect 5749 -15400 5795 -15388
rect 5927 -15132 5973 -15120
rect 5927 -15388 5933 -15132
rect 5967 -15388 5973 -15132
rect 5927 -15400 5973 -15388
rect 6105 -15132 6151 -15120
rect 6105 -15388 6111 -15132
rect 6145 -15388 6151 -15132
rect 6105 -15400 6151 -15388
rect 6283 -15132 6329 -15120
rect 6283 -15388 6289 -15132
rect 6323 -15388 6329 -15132
rect 6283 -15400 6329 -15388
rect 6461 -15132 6507 -15120
rect 6461 -15388 6467 -15132
rect 6501 -15388 6507 -15132
rect 6461 -15400 6507 -15388
rect 6639 -15132 6685 -15120
rect 6639 -15388 6645 -15132
rect 6679 -15388 6685 -15132
rect 6639 -15400 6685 -15388
rect 6817 -15132 6863 -15120
rect 6817 -15388 6823 -15132
rect 6857 -15388 6863 -15132
rect 6817 -15400 6863 -15388
rect 6995 -15132 7041 -15120
rect 6995 -15388 7001 -15132
rect 7035 -15388 7041 -15132
rect 6995 -15400 7041 -15388
rect 7173 -15132 7219 -15120
rect 7173 -15388 7179 -15132
rect 7213 -15388 7219 -15132
rect 7173 -15400 7219 -15388
rect 7351 -15132 7397 -15120
rect 7351 -15388 7357 -15132
rect 7391 -15388 7397 -15132
rect 7351 -15400 7397 -15388
rect 7529 -15132 7575 -15120
rect 7529 -15388 7535 -15132
rect 7569 -15388 7575 -15132
rect 7529 -15400 7575 -15388
rect 7707 -15132 7753 -15120
rect 7707 -15388 7713 -15132
rect 7747 -15388 7753 -15132
rect 7707 -15400 7753 -15388
rect 7885 -15132 7931 -15120
rect 7885 -15388 7891 -15132
rect 7925 -15388 7931 -15132
rect 7885 -15400 7931 -15388
rect 8063 -15132 8109 -15120
rect 8063 -15388 8069 -15132
rect 8103 -15388 8109 -15132
rect 8063 -15400 8109 -15388
rect 8241 -15132 8287 -15120
rect 8241 -15388 8247 -15132
rect 8281 -15388 8287 -15132
rect 8241 -15400 8287 -15388
rect 8419 -15132 8465 -15120
rect 8419 -15388 8425 -15132
rect 8459 -15388 8465 -15132
rect 8419 -15400 8465 -15388
rect 8597 -15132 8643 -15120
rect 8597 -15388 8603 -15132
rect 8637 -15388 8643 -15132
rect 8597 -15400 8643 -15388
rect 8775 -15132 8821 -15120
rect 8775 -15388 8781 -15132
rect 8815 -15388 8821 -15132
rect 8775 -15400 8821 -15388
rect 8953 -15132 8999 -15120
rect 8953 -15388 8959 -15132
rect 8993 -15388 8999 -15132
rect 8953 -15400 8999 -15388
rect 9131 -15132 9177 -15120
rect 9131 -15388 9137 -15132
rect 9171 -15388 9177 -15132
rect 9131 -15400 9177 -15388
rect 9309 -15132 9355 -15120
rect 9309 -15388 9315 -15132
rect 9349 -15388 9355 -15132
rect 9309 -15400 9355 -15388
rect 9487 -15132 9533 -15120
rect 9487 -15388 9493 -15132
rect 9527 -15388 9533 -15132
rect 9487 -15400 9533 -15388
rect 9665 -15132 9711 -15120
rect 9665 -15388 9671 -15132
rect 9705 -15388 9711 -15132
rect 9665 -15400 9711 -15388
rect 9843 -15132 9889 -15120
rect 9843 -15388 9849 -15132
rect 9883 -15388 9889 -15132
rect 9843 -15400 9889 -15388
rect 10021 -15132 10067 -15120
rect 10021 -15388 10027 -15132
rect 10061 -15388 10067 -15132
rect 10021 -15400 10067 -15388
rect 10199 -15132 10245 -15120
rect 10199 -15388 10205 -15132
rect 10239 -15388 10245 -15132
rect 10199 -15400 10245 -15388
rect 10377 -15132 10423 -15120
rect 10377 -15388 10383 -15132
rect 10417 -15388 10423 -15132
rect 10377 -15400 10423 -15388
rect 10555 -15132 10601 -15120
rect 10555 -15388 10561 -15132
rect 10595 -15388 10601 -15132
rect 10555 -15400 10601 -15388
rect 10733 -15132 10779 -15120
rect 10733 -15388 10739 -15132
rect 10773 -15388 10779 -15132
rect 10733 -15400 10779 -15388
rect 10911 -15132 10957 -15120
rect 10911 -15388 10917 -15132
rect 10951 -15388 10957 -15132
rect 10911 -15400 10957 -15388
rect 11089 -15132 11135 -15120
rect 11089 -15388 11095 -15132
rect 11129 -15388 11135 -15132
rect 11089 -15400 11135 -15388
rect 11267 -15132 11313 -15120
rect 11267 -15388 11273 -15132
rect 11307 -15388 11313 -15132
rect 11267 -15400 11313 -15388
rect 11445 -15132 11491 -15120
rect 11445 -15388 11451 -15132
rect 11485 -15388 11491 -15132
rect 11445 -15400 11491 -15388
rect 11623 -15132 11669 -15120
rect 11623 -15388 11629 -15132
rect 11663 -15388 11669 -15132
rect 11623 -15400 11669 -15388
rect 11801 -15132 11847 -15120
rect 11801 -15388 11807 -15132
rect 11841 -15388 11847 -15132
rect 11801 -15400 11847 -15388
rect 11979 -15132 12025 -15120
rect 11979 -15388 11985 -15132
rect 12019 -15388 12025 -15132
rect 11979 -15400 12025 -15388
rect 12157 -15132 12203 -15120
rect 12157 -15388 12163 -15132
rect 12197 -15388 12203 -15132
rect 12157 -15400 12203 -15388
rect 12335 -15132 12381 -15120
rect 12335 -15388 12341 -15132
rect 12375 -15388 12381 -15132
rect 12335 -15400 12381 -15388
rect 12513 -15132 12559 -15120
rect 12513 -15388 12519 -15132
rect 12553 -15388 12559 -15132
rect 12513 -15400 12559 -15388
rect 12691 -15132 12737 -15120
rect 12691 -15388 12697 -15132
rect 12731 -15388 12737 -15132
rect 12691 -15400 12737 -15388
rect 5645 -15438 5721 -15432
rect 5645 -15472 5661 -15438
rect 5705 -15472 5721 -15438
rect 5645 -15488 5721 -15472
rect 5755 -15539 5789 -15400
rect 5823 -15438 5899 -15432
rect 5823 -15472 5839 -15438
rect 5883 -15472 5899 -15438
rect 5823 -15488 5899 -15472
rect 5735 -15592 5745 -15539
rect 5798 -15592 5808 -15539
rect 5390 -15706 5400 -15653
rect 5453 -15706 5463 -15653
rect 5400 -16667 5453 -15706
rect 5737 -15803 5747 -15750
rect 5800 -15803 5810 -15750
rect 5645 -16048 5721 -16032
rect 5645 -16082 5661 -16048
rect 5705 -16082 5721 -16048
rect 5645 -16088 5721 -16082
rect 5756 -16120 5790 -15803
rect 5844 -16032 5878 -15488
rect 5933 -15652 5967 -15400
rect 6001 -15438 6077 -15432
rect 6001 -15472 6017 -15438
rect 6061 -15472 6077 -15438
rect 6001 -15488 6077 -15472
rect 5913 -15705 5923 -15652
rect 5976 -15705 5986 -15652
rect 5911 -16001 5921 -15948
rect 5974 -16001 5984 -15948
rect 5823 -16048 5899 -16032
rect 5823 -16082 5839 -16048
rect 5883 -16082 5899 -16048
rect 5823 -16088 5899 -16082
rect 5931 -16120 5965 -16001
rect 6022 -16032 6056 -15488
rect 6111 -15539 6145 -15400
rect 6179 -15438 6255 -15432
rect 6179 -15472 6195 -15438
rect 6239 -15472 6255 -15438
rect 6179 -15488 6255 -15472
rect 6091 -15592 6101 -15539
rect 6154 -15592 6164 -15539
rect 6091 -15802 6101 -15749
rect 6154 -15802 6164 -15749
rect 6001 -16048 6077 -16032
rect 6001 -16082 6017 -16048
rect 6061 -16082 6077 -16048
rect 6001 -16088 6077 -16082
rect 6112 -16120 6146 -15802
rect 6201 -16032 6235 -15488
rect 6289 -15652 6323 -15400
rect 6357 -15438 6433 -15432
rect 6357 -15472 6373 -15438
rect 6417 -15472 6433 -15438
rect 6357 -15488 6433 -15472
rect 6269 -15705 6279 -15652
rect 6332 -15705 6342 -15652
rect 6269 -16001 6279 -15948
rect 6332 -16001 6342 -15948
rect 6179 -16048 6255 -16032
rect 6179 -16082 6195 -16048
rect 6239 -16082 6255 -16048
rect 6179 -16088 6255 -16082
rect 6288 -16120 6322 -16001
rect 6379 -16032 6413 -15488
rect 6468 -15539 6502 -15400
rect 6535 -15438 6611 -15432
rect 6535 -15472 6551 -15438
rect 6595 -15472 6611 -15438
rect 6535 -15488 6611 -15472
rect 6448 -15592 6458 -15539
rect 6511 -15592 6521 -15539
rect 6446 -15803 6456 -15750
rect 6509 -15803 6519 -15750
rect 6357 -16048 6433 -16032
rect 6357 -16082 6373 -16048
rect 6417 -16082 6433 -16048
rect 6357 -16088 6433 -16082
rect 6467 -16120 6501 -15803
rect 6556 -16032 6590 -15488
rect 6645 -15652 6679 -15400
rect 6713 -15438 6789 -15432
rect 6822 -15438 6857 -15400
rect 6891 -15438 6967 -15432
rect 6713 -15472 6729 -15438
rect 6773 -15472 6907 -15438
rect 6951 -15472 6967 -15438
rect 6713 -15488 6789 -15472
rect 6625 -15705 6635 -15652
rect 6688 -15705 6698 -15652
rect 6703 -15804 6713 -15751
rect 6766 -15804 6776 -15751
rect 6624 -16001 6634 -15948
rect 6687 -16001 6697 -15948
rect 6734 -15956 6768 -15804
rect 6822 -15851 6856 -15472
rect 6891 -15488 6967 -15472
rect 6803 -15904 6813 -15851
rect 6866 -15904 6876 -15851
rect 7002 -15951 7036 -15400
rect 7069 -15438 7145 -15432
rect 7069 -15472 7085 -15438
rect 7129 -15472 7145 -15438
rect 7069 -15488 7145 -15472
rect 7179 -15750 7213 -15400
rect 7247 -15438 7323 -15432
rect 7247 -15472 7263 -15438
rect 7307 -15472 7323 -15438
rect 7247 -15488 7323 -15472
rect 7425 -15438 7501 -15432
rect 7425 -15472 7441 -15438
rect 7485 -15472 7501 -15438
rect 7425 -15488 7501 -15472
rect 7159 -15803 7169 -15750
rect 7222 -15803 7232 -15750
rect 7159 -15905 7169 -15852
rect 7222 -15905 7232 -15852
rect 6734 -15990 6858 -15956
rect 6535 -16048 6611 -16032
rect 6535 -16082 6551 -16048
rect 6595 -16082 6611 -16048
rect 6535 -16088 6611 -16082
rect 6644 -16120 6678 -16001
rect 6713 -16048 6789 -16032
rect 6713 -16082 6729 -16048
rect 6773 -16082 6789 -16048
rect 6713 -16088 6789 -16082
rect 6824 -16120 6858 -15990
rect 6984 -16004 6994 -15951
rect 7047 -16004 7057 -15951
rect 6891 -16048 6967 -16032
rect 6891 -16082 6907 -16048
rect 6951 -16082 6967 -16048
rect 6891 -16088 6967 -16082
rect 7002 -16120 7036 -16004
rect 7069 -16048 7145 -16032
rect 7069 -16082 7085 -16048
rect 7129 -16082 7145 -16048
rect 7069 -16088 7145 -16082
rect 7178 -16120 7212 -15905
rect 7447 -16032 7481 -15488
rect 7536 -15749 7570 -15400
rect 7603 -15438 7679 -15432
rect 7603 -15472 7619 -15438
rect 7663 -15472 7679 -15438
rect 7603 -15488 7679 -15472
rect 7781 -15438 7857 -15432
rect 7781 -15472 7797 -15438
rect 7841 -15472 7857 -15438
rect 7781 -15488 7857 -15472
rect 7516 -15802 7526 -15749
rect 7579 -15802 7589 -15749
rect 7516 -16006 7526 -15953
rect 7579 -16006 7589 -15953
rect 7247 -16048 7323 -16032
rect 7247 -16082 7263 -16048
rect 7307 -16082 7323 -16048
rect 7247 -16088 7323 -16082
rect 7425 -16048 7501 -16032
rect 7425 -16082 7441 -16048
rect 7485 -16082 7501 -16048
rect 7425 -16088 7501 -16082
rect 7535 -16120 7569 -16006
rect 7624 -16032 7658 -15488
rect 7803 -16032 7837 -15488
rect 7891 -15749 7925 -15400
rect 7959 -15438 8035 -15432
rect 8069 -15438 8103 -15400
rect 8137 -15438 8213 -15432
rect 7959 -15472 7975 -15438
rect 8019 -15472 8153 -15438
rect 8197 -15472 8213 -15438
rect 7959 -15488 8035 -15472
rect 7872 -15802 7882 -15749
rect 7935 -15802 7945 -15749
rect 8069 -15851 8103 -15472
rect 8137 -15488 8213 -15472
rect 8050 -15904 8060 -15851
rect 8113 -15904 8123 -15851
rect 8247 -15952 8281 -15400
rect 8315 -15438 8391 -15432
rect 8315 -15472 8331 -15438
rect 8375 -15472 8391 -15438
rect 8315 -15488 8391 -15472
rect 7871 -16005 7881 -15952
rect 7934 -16005 7944 -15952
rect 8227 -16005 8237 -15952
rect 8290 -16005 8300 -15952
rect 7603 -16048 7679 -16032
rect 7603 -16082 7619 -16048
rect 7663 -16082 7679 -16048
rect 7603 -16088 7679 -16082
rect 7781 -16048 7857 -16032
rect 7781 -16082 7797 -16048
rect 7841 -16082 7857 -16048
rect 7781 -16088 7857 -16082
rect 7891 -16120 7925 -16005
rect 7959 -16048 8035 -16032
rect 7959 -16082 7975 -16048
rect 8019 -16082 8035 -16048
rect 7959 -16088 8035 -16082
rect 8137 -16048 8213 -16032
rect 8137 -16082 8153 -16048
rect 8197 -16082 8213 -16048
rect 8137 -16088 8213 -16082
rect 8247 -16120 8281 -16005
rect 8336 -16032 8370 -15488
rect 8315 -16048 8391 -16032
rect 8315 -16082 8331 -16048
rect 8375 -16082 8391 -16048
rect 8315 -16088 8391 -16082
rect 8426 -16120 8460 -15400
rect 8493 -15438 8569 -15432
rect 8493 -15472 8509 -15438
rect 8553 -15472 8569 -15438
rect 8493 -15488 8569 -15472
rect 8671 -15438 8747 -15432
rect 8671 -15472 8687 -15438
rect 8731 -15472 8747 -15438
rect 8671 -15488 8747 -15472
rect 8849 -15438 8925 -15432
rect 8849 -15472 8865 -15438
rect 8909 -15472 8925 -15438
rect 8849 -15488 8925 -15472
rect 9027 -15438 9103 -15432
rect 9027 -15472 9043 -15438
rect 9087 -15472 9103 -15438
rect 9027 -15488 9103 -15472
rect 9205 -15438 9281 -15432
rect 9205 -15472 9221 -15438
rect 9265 -15472 9281 -15438
rect 9205 -15488 9281 -15472
rect 9383 -15438 9459 -15432
rect 9383 -15472 9399 -15438
rect 9443 -15472 9459 -15438
rect 9383 -15488 9459 -15472
rect 9561 -15438 9637 -15432
rect 9561 -15472 9577 -15438
rect 9621 -15472 9637 -15438
rect 9561 -15488 9637 -15472
rect 9739 -15438 9815 -15432
rect 9739 -15472 9755 -15438
rect 9799 -15472 9815 -15438
rect 9739 -15488 9815 -15472
rect 9917 -15438 9993 -15432
rect 9917 -15472 9933 -15438
rect 9977 -15472 9993 -15438
rect 9917 -15488 9993 -15472
rect 10095 -15438 10171 -15432
rect 10205 -15438 10239 -15400
rect 10273 -15438 10349 -15432
rect 10095 -15472 10111 -15438
rect 10155 -15472 10289 -15438
rect 10333 -15472 10349 -15438
rect 10095 -15488 10171 -15472
rect 8583 -15905 8593 -15852
rect 8646 -15905 8656 -15852
rect 8493 -16048 8569 -16032
rect 8493 -16082 8509 -16048
rect 8553 -16082 8569 -16048
rect 8493 -16088 8569 -16082
rect 8603 -16120 8637 -15905
rect 8870 -16032 8904 -15488
rect 9049 -16032 9083 -15488
rect 9226 -16032 9260 -15488
rect 9404 -16032 9438 -15488
rect 9653 -15905 9663 -15852
rect 9716 -15905 9726 -15852
rect 8671 -16048 8747 -16032
rect 8671 -16082 8687 -16048
rect 8731 -16082 8747 -16048
rect 8671 -16088 8747 -16082
rect 8849 -16048 8925 -16032
rect 8849 -16082 8865 -16048
rect 8909 -16082 8925 -16048
rect 8849 -16088 8925 -16082
rect 9027 -16048 9103 -16032
rect 9027 -16082 9043 -16048
rect 9087 -16082 9103 -16048
rect 9027 -16088 9103 -16082
rect 9205 -16048 9281 -16032
rect 9205 -16082 9221 -16048
rect 9265 -16082 9281 -16048
rect 9205 -16088 9281 -16082
rect 9383 -16048 9459 -16032
rect 9383 -16082 9399 -16048
rect 9443 -16082 9459 -16048
rect 9383 -16088 9459 -16082
rect 9561 -16048 9637 -16032
rect 9561 -16082 9577 -16048
rect 9621 -16082 9637 -16048
rect 9561 -16088 9637 -16082
rect 9672 -16120 9706 -15905
rect 9939 -16032 9973 -15488
rect 10205 -15852 10239 -15472
rect 10273 -15488 10349 -15472
rect 10383 -15751 10417 -15400
rect 10451 -15438 10527 -15432
rect 10451 -15472 10467 -15438
rect 10511 -15472 10527 -15438
rect 10451 -15488 10527 -15472
rect 10629 -15438 10705 -15432
rect 10629 -15472 10645 -15438
rect 10689 -15472 10705 -15438
rect 10629 -15488 10705 -15472
rect 10363 -15804 10373 -15751
rect 10426 -15804 10436 -15751
rect 10184 -15905 10194 -15852
rect 10247 -15905 10257 -15852
rect 10472 -16032 10506 -15488
rect 10650 -16032 10684 -15488
rect 10739 -15750 10773 -15400
rect 10807 -15438 10883 -15432
rect 10807 -15472 10823 -15438
rect 10867 -15472 10883 -15438
rect 10807 -15488 10883 -15472
rect 10720 -15803 10730 -15750
rect 10783 -15803 10793 -15750
rect 9739 -16048 9815 -16032
rect 9739 -16082 9755 -16048
rect 9799 -16082 9815 -16048
rect 9739 -16088 9815 -16082
rect 9917 -16048 9993 -16032
rect 9917 -16082 9933 -16048
rect 9977 -16082 9993 -16048
rect 9917 -16088 9993 -16082
rect 10095 -16048 10171 -16032
rect 10095 -16082 10111 -16048
rect 10155 -16082 10171 -16048
rect 10095 -16088 10171 -16082
rect 10273 -16048 10349 -16032
rect 10273 -16082 10289 -16048
rect 10333 -16082 10349 -16048
rect 10273 -16088 10349 -16082
rect 10451 -16048 10527 -16032
rect 10451 -16082 10467 -16048
rect 10511 -16082 10527 -16048
rect 10451 -16088 10527 -16082
rect 10629 -16048 10705 -16032
rect 10629 -16082 10645 -16048
rect 10689 -16082 10705 -16048
rect 10629 -16088 10705 -16082
rect 10739 -16120 10773 -15803
rect 10828 -16032 10862 -15488
rect 10807 -16048 10883 -16032
rect 10807 -16082 10823 -16048
rect 10867 -16082 10883 -16048
rect 10807 -16088 10883 -16082
rect 10916 -16120 10950 -15400
rect 10985 -15438 11061 -15432
rect 10985 -15472 11001 -15438
rect 11045 -15472 11061 -15438
rect 10985 -15488 11061 -15472
rect 11095 -15750 11129 -15400
rect 11163 -15438 11239 -15432
rect 11163 -15472 11179 -15438
rect 11223 -15472 11239 -15438
rect 11163 -15488 11239 -15472
rect 11341 -15438 11417 -15432
rect 11451 -15438 11485 -15400
rect 11519 -15438 11595 -15432
rect 11341 -15472 11357 -15438
rect 11401 -15472 11535 -15438
rect 11579 -15472 11595 -15438
rect 11341 -15488 11417 -15472
rect 11076 -15803 11086 -15750
rect 11139 -15803 11149 -15750
rect 11451 -15841 11485 -15472
rect 11519 -15488 11595 -15472
rect 11629 -15652 11663 -15400
rect 11697 -15438 11773 -15432
rect 11697 -15472 11713 -15438
rect 11757 -15472 11773 -15438
rect 11697 -15488 11773 -15472
rect 11609 -15705 11619 -15652
rect 11672 -15705 11682 -15652
rect 11629 -15706 11663 -15705
rect 11074 -15905 11084 -15852
rect 11137 -15905 11147 -15852
rect 11430 -15894 11440 -15841
rect 11493 -15894 11503 -15841
rect 11451 -15902 11485 -15894
rect 10985 -16048 11061 -16032
rect 10985 -16082 11001 -16048
rect 11045 -16082 11061 -16048
rect 10985 -16088 11061 -16082
rect 11094 -16120 11128 -15905
rect 11431 -16005 11441 -15952
rect 11494 -16005 11504 -15952
rect 11163 -16048 11239 -16032
rect 11163 -16082 11179 -16048
rect 11223 -16082 11239 -16048
rect 11163 -16088 11239 -16082
rect 11341 -16048 11417 -16032
rect 11341 -16082 11357 -16048
rect 11401 -16082 11417 -16048
rect 11341 -16088 11417 -16082
rect 11451 -16120 11485 -16005
rect 11718 -16032 11752 -15488
rect 11808 -15540 11842 -15400
rect 11875 -15438 11951 -15432
rect 11875 -15472 11891 -15438
rect 11935 -15472 11951 -15438
rect 11875 -15488 11951 -15472
rect 11788 -15593 11798 -15540
rect 11851 -15593 11861 -15540
rect 11787 -16005 11797 -15952
rect 11850 -16005 11860 -15952
rect 11519 -16048 11595 -16032
rect 11519 -16082 11535 -16048
rect 11579 -16082 11595 -16048
rect 11519 -16088 11595 -16082
rect 11697 -16048 11773 -16032
rect 11697 -16082 11713 -16048
rect 11757 -16082 11773 -16048
rect 11697 -16088 11773 -16082
rect 11806 -16120 11840 -16005
rect 11897 -16032 11931 -15488
rect 11985 -15652 12019 -15400
rect 12053 -15438 12129 -15432
rect 12053 -15472 12069 -15438
rect 12113 -15472 12129 -15438
rect 12053 -15488 12129 -15472
rect 11965 -15705 11975 -15652
rect 12028 -15705 12038 -15652
rect 12074 -16032 12108 -15488
rect 12165 -15539 12199 -15400
rect 12231 -15438 12307 -15432
rect 12231 -15472 12247 -15438
rect 12291 -15472 12307 -15438
rect 12231 -15488 12307 -15472
rect 12145 -15592 12155 -15539
rect 12208 -15592 12218 -15539
rect 12144 -16005 12154 -15952
rect 12207 -16005 12217 -15952
rect 11875 -16048 11951 -16032
rect 11875 -16082 11891 -16048
rect 11935 -16082 11951 -16048
rect 11875 -16088 11951 -16082
rect 12053 -16048 12129 -16032
rect 12053 -16082 12069 -16048
rect 12113 -16082 12129 -16048
rect 12053 -16088 12129 -16082
rect 12163 -16120 12197 -16005
rect 12252 -16032 12286 -15488
rect 12342 -15652 12376 -15400
rect 12409 -15438 12485 -15432
rect 12409 -15472 12425 -15438
rect 12469 -15472 12485 -15438
rect 12409 -15488 12485 -15472
rect 12322 -15705 12332 -15652
rect 12385 -15705 12395 -15652
rect 12431 -16032 12465 -15488
rect 12520 -15539 12554 -15400
rect 12587 -15438 12663 -15432
rect 12587 -15472 12603 -15438
rect 12647 -15472 12663 -15438
rect 12587 -15488 12663 -15472
rect 12501 -15592 12511 -15539
rect 12564 -15592 12574 -15539
rect 12501 -16005 12511 -15952
rect 12564 -16005 12574 -15952
rect 12231 -16048 12307 -16032
rect 12231 -16082 12247 -16048
rect 12291 -16082 12307 -16048
rect 12231 -16088 12307 -16082
rect 12409 -16048 12485 -16032
rect 12409 -16082 12425 -16048
rect 12469 -16082 12485 -16048
rect 12409 -16088 12485 -16082
rect 12520 -16120 12554 -16005
rect 12587 -16048 12663 -16032
rect 12587 -16082 12603 -16048
rect 12647 -16082 12663 -16048
rect 12587 -16088 12663 -16082
rect 5571 -16132 5617 -16120
rect 5571 -16388 5577 -16132
rect 5611 -16388 5617 -16132
rect 5571 -16400 5617 -16388
rect 5749 -16132 5795 -16120
rect 5749 -16388 5755 -16132
rect 5789 -16388 5795 -16132
rect 5749 -16400 5795 -16388
rect 5927 -16132 5973 -16120
rect 5927 -16388 5933 -16132
rect 5967 -16388 5973 -16132
rect 5927 -16400 5973 -16388
rect 6105 -16132 6151 -16120
rect 6105 -16388 6111 -16132
rect 6145 -16388 6151 -16132
rect 6105 -16400 6151 -16388
rect 6283 -16132 6329 -16120
rect 6283 -16388 6289 -16132
rect 6323 -16388 6329 -16132
rect 6283 -16400 6329 -16388
rect 6461 -16132 6507 -16120
rect 6461 -16388 6467 -16132
rect 6501 -16388 6507 -16132
rect 6461 -16400 6507 -16388
rect 6639 -16132 6685 -16120
rect 6639 -16388 6645 -16132
rect 6679 -16388 6685 -16132
rect 6639 -16400 6685 -16388
rect 6817 -16132 6863 -16120
rect 6817 -16388 6823 -16132
rect 6857 -16388 6863 -16132
rect 6817 -16400 6863 -16388
rect 6995 -16132 7041 -16120
rect 6995 -16388 7001 -16132
rect 7035 -16388 7041 -16132
rect 6995 -16400 7041 -16388
rect 7173 -16132 7219 -16120
rect 7173 -16388 7179 -16132
rect 7213 -16388 7219 -16132
rect 7173 -16400 7219 -16388
rect 7351 -16132 7397 -16120
rect 7351 -16388 7357 -16132
rect 7391 -16388 7397 -16132
rect 7351 -16400 7397 -16388
rect 7529 -16132 7575 -16120
rect 7529 -16388 7535 -16132
rect 7569 -16388 7575 -16132
rect 7529 -16400 7575 -16388
rect 7707 -16132 7753 -16120
rect 7707 -16388 7713 -16132
rect 7747 -16388 7753 -16132
rect 7707 -16400 7753 -16388
rect 7885 -16132 7931 -16120
rect 7885 -16388 7891 -16132
rect 7925 -16388 7931 -16132
rect 7885 -16400 7931 -16388
rect 8063 -16132 8109 -16120
rect 8063 -16388 8069 -16132
rect 8103 -16388 8109 -16132
rect 8063 -16400 8109 -16388
rect 8241 -16132 8287 -16120
rect 8241 -16388 8247 -16132
rect 8281 -16388 8287 -16132
rect 8241 -16400 8287 -16388
rect 8419 -16132 8465 -16120
rect 8419 -16388 8425 -16132
rect 8459 -16388 8465 -16132
rect 8419 -16400 8465 -16388
rect 8597 -16132 8643 -16120
rect 8597 -16388 8603 -16132
rect 8637 -16388 8643 -16132
rect 8597 -16400 8643 -16388
rect 8775 -16132 8821 -16120
rect 8775 -16388 8781 -16132
rect 8815 -16388 8821 -16132
rect 8775 -16400 8821 -16388
rect 8953 -16132 8999 -16120
rect 8953 -16388 8959 -16132
rect 8993 -16388 8999 -16132
rect 8953 -16400 8999 -16388
rect 9131 -16132 9177 -16120
rect 9131 -16388 9137 -16132
rect 9171 -16388 9177 -16132
rect 9131 -16400 9177 -16388
rect 9309 -16132 9355 -16120
rect 9309 -16388 9315 -16132
rect 9349 -16388 9355 -16132
rect 9309 -16400 9355 -16388
rect 9487 -16132 9533 -16120
rect 9487 -16388 9493 -16132
rect 9527 -16388 9533 -16132
rect 9487 -16400 9533 -16388
rect 9665 -16132 9711 -16120
rect 9665 -16388 9671 -16132
rect 9705 -16388 9711 -16132
rect 9665 -16400 9711 -16388
rect 9843 -16132 9889 -16120
rect 9843 -16388 9849 -16132
rect 9883 -16388 9889 -16132
rect 9843 -16400 9889 -16388
rect 10021 -16132 10067 -16120
rect 10021 -16388 10027 -16132
rect 10061 -16388 10067 -16132
rect 10021 -16400 10067 -16388
rect 10199 -16132 10245 -16120
rect 10199 -16388 10205 -16132
rect 10239 -16388 10245 -16132
rect 10199 -16400 10245 -16388
rect 10377 -16132 10423 -16120
rect 10377 -16388 10383 -16132
rect 10417 -16388 10423 -16132
rect 10377 -16400 10423 -16388
rect 10555 -16132 10601 -16120
rect 10555 -16388 10561 -16132
rect 10595 -16388 10601 -16132
rect 10555 -16400 10601 -16388
rect 10733 -16132 10779 -16120
rect 10733 -16388 10739 -16132
rect 10773 -16388 10779 -16132
rect 10733 -16400 10779 -16388
rect 10911 -16132 10957 -16120
rect 10911 -16388 10917 -16132
rect 10951 -16388 10957 -16132
rect 10911 -16400 10957 -16388
rect 11089 -16132 11135 -16120
rect 11089 -16388 11095 -16132
rect 11129 -16388 11135 -16132
rect 11089 -16400 11135 -16388
rect 11267 -16132 11313 -16120
rect 11267 -16388 11273 -16132
rect 11307 -16388 11313 -16132
rect 11267 -16400 11313 -16388
rect 11445 -16132 11491 -16120
rect 11445 -16388 11451 -16132
rect 11485 -16388 11491 -16132
rect 11445 -16400 11491 -16388
rect 11623 -16132 11669 -16120
rect 11623 -16388 11629 -16132
rect 11663 -16388 11669 -16132
rect 11623 -16400 11669 -16388
rect 11801 -16132 11847 -16120
rect 11801 -16388 11807 -16132
rect 11841 -16388 11847 -16132
rect 11801 -16400 11847 -16388
rect 11979 -16132 12025 -16120
rect 11979 -16388 11985 -16132
rect 12019 -16388 12025 -16132
rect 11979 -16400 12025 -16388
rect 12157 -16132 12203 -16120
rect 12157 -16388 12163 -16132
rect 12197 -16388 12203 -16132
rect 12157 -16400 12203 -16388
rect 12335 -16132 12381 -16120
rect 12335 -16388 12341 -16132
rect 12375 -16388 12381 -16132
rect 12335 -16400 12381 -16388
rect 12513 -16132 12559 -16120
rect 12513 -16388 12519 -16132
rect 12553 -16388 12559 -16132
rect 12513 -16400 12559 -16388
rect 12691 -16132 12737 -16120
rect 12691 -16388 12697 -16132
rect 12731 -16388 12737 -16132
rect 12691 -16400 12737 -16388
rect 5576 -16438 5610 -16400
rect 5645 -16438 5721 -16432
rect 5756 -16438 5790 -16400
rect 5576 -16472 5661 -16438
rect 5705 -16472 5790 -16438
rect 5823 -16438 5899 -16432
rect 5823 -16472 5839 -16438
rect 5883 -16472 5899 -16438
rect 5645 -16488 5721 -16472
rect 5823 -16488 5899 -16472
rect 6001 -16438 6077 -16432
rect 6001 -16472 6017 -16438
rect 6061 -16472 6077 -16438
rect 6001 -16488 6077 -16472
rect 6179 -16438 6255 -16432
rect 6179 -16472 6195 -16438
rect 6239 -16472 6255 -16438
rect 6179 -16488 6255 -16472
rect 6357 -16438 6433 -16432
rect 6357 -16472 6373 -16438
rect 6417 -16472 6433 -16438
rect 6357 -16488 6433 -16472
rect 6535 -16438 6611 -16432
rect 6535 -16472 6551 -16438
rect 6595 -16472 6611 -16438
rect 6535 -16488 6611 -16472
rect 6713 -16438 6789 -16432
rect 6713 -16472 6729 -16438
rect 6773 -16472 6789 -16438
rect 6713 -16488 6789 -16472
rect 6891 -16438 6967 -16432
rect 6891 -16472 6907 -16438
rect 6951 -16472 6967 -16438
rect 6891 -16488 6967 -16472
rect 7069 -16438 7145 -16432
rect 7178 -16438 7212 -16400
rect 7247 -16438 7323 -16432
rect 7069 -16472 7085 -16438
rect 7129 -16472 7263 -16438
rect 7307 -16472 7323 -16438
rect 7069 -16488 7145 -16472
rect 7247 -16488 7323 -16472
rect 6557 -16544 6591 -16488
rect 6735 -16544 6769 -16488
rect 6538 -16597 6548 -16544
rect 6601 -16597 6611 -16544
rect 6716 -16597 6726 -16544
rect 6779 -16597 6789 -16544
rect 6912 -16545 6946 -16488
rect 6893 -16598 6903 -16545
rect 6956 -16598 6966 -16545
rect 5389 -16720 5399 -16667
rect 5452 -16720 5462 -16667
rect 5021 -16835 5031 -16782
rect 5084 -16835 5094 -16782
rect 7357 -16890 7391 -16400
rect 7425 -16438 7501 -16432
rect 7425 -16472 7441 -16438
rect 7485 -16472 7501 -16438
rect 7425 -16488 7501 -16472
rect 7603 -16438 7679 -16432
rect 7603 -16472 7619 -16438
rect 7663 -16472 7679 -16438
rect 7603 -16488 7679 -16472
rect 7713 -16890 7747 -16400
rect 7781 -16438 7857 -16432
rect 7781 -16472 7797 -16438
rect 7841 -16472 7857 -16438
rect 7781 -16488 7857 -16472
rect 7959 -16438 8035 -16432
rect 7959 -16472 7975 -16438
rect 8019 -16472 8035 -16438
rect 7959 -16488 8035 -16472
rect 7980 -16545 8014 -16488
rect 7960 -16598 7970 -16545
rect 8023 -16598 8033 -16545
rect 8069 -16890 8103 -16400
rect 8137 -16438 8213 -16432
rect 8137 -16472 8153 -16438
rect 8197 -16472 8213 -16438
rect 8137 -16488 8213 -16472
rect 8315 -16438 8391 -16432
rect 8315 -16472 8331 -16438
rect 8375 -16472 8391 -16438
rect 8315 -16488 8391 -16472
rect 8158 -16544 8192 -16488
rect 8139 -16597 8149 -16544
rect 8202 -16597 8212 -16544
rect 8426 -16890 8460 -16400
rect 8493 -16438 8569 -16432
rect 8603 -16438 8637 -16400
rect 8671 -16438 8747 -16432
rect 8493 -16472 8509 -16438
rect 8553 -16472 8687 -16438
rect 8731 -16472 8747 -16438
rect 8493 -16488 8569 -16472
rect 8671 -16488 8747 -16472
rect 8781 -16666 8815 -16400
rect 8849 -16438 8925 -16432
rect 8849 -16472 8865 -16438
rect 8909 -16472 8925 -16438
rect 8849 -16488 8925 -16472
rect 8761 -16719 8771 -16666
rect 8824 -16719 8834 -16666
rect 8960 -16782 8994 -16400
rect 9027 -16438 9103 -16432
rect 9027 -16472 9043 -16438
rect 9087 -16472 9103 -16438
rect 9027 -16488 9103 -16472
rect 9138 -16666 9172 -16400
rect 9205 -16438 9281 -16432
rect 9205 -16472 9221 -16438
rect 9265 -16472 9281 -16438
rect 9205 -16488 9281 -16472
rect 9118 -16719 9128 -16666
rect 9181 -16719 9191 -16666
rect 9315 -16782 9349 -16400
rect 9383 -16438 9459 -16432
rect 9383 -16472 9399 -16438
rect 9443 -16472 9459 -16438
rect 9383 -16488 9459 -16472
rect 9493 -16666 9527 -16400
rect 9561 -16438 9637 -16432
rect 9672 -16438 9706 -16400
rect 9739 -16438 9815 -16432
rect 9561 -16472 9577 -16438
rect 9621 -16472 9755 -16438
rect 9799 -16472 9815 -16438
rect 9561 -16488 9637 -16472
rect 9474 -16719 9484 -16666
rect 9537 -16719 9547 -16666
rect 8940 -16835 8950 -16782
rect 9003 -16835 9013 -16782
rect 9295 -16835 9305 -16782
rect 9358 -16835 9368 -16782
rect 7337 -16943 7347 -16890
rect 7400 -16943 7410 -16890
rect 7694 -16943 7704 -16890
rect 7757 -16943 7767 -16890
rect 8050 -16943 8060 -16890
rect 8113 -16943 8123 -16890
rect 8406 -16943 8416 -16890
rect 8469 -16943 8479 -16890
rect 9672 -17251 9706 -16472
rect 9739 -16488 9815 -16472
rect 9848 -16666 9882 -16400
rect 9917 -16438 9993 -16432
rect 9917 -16472 9933 -16438
rect 9977 -16472 9993 -16438
rect 9917 -16488 9993 -16472
rect 9938 -16544 9972 -16488
rect 9919 -16597 9929 -16544
rect 9982 -16597 9992 -16544
rect 9828 -16719 9838 -16666
rect 9891 -16719 9901 -16666
rect 10028 -16781 10062 -16400
rect 10095 -16438 10171 -16432
rect 10095 -16472 10111 -16438
rect 10155 -16472 10171 -16438
rect 10095 -16488 10171 -16472
rect 10117 -16545 10151 -16488
rect 10097 -16598 10107 -16545
rect 10160 -16598 10170 -16545
rect 10205 -16665 10239 -16400
rect 10273 -16438 10349 -16432
rect 10273 -16472 10289 -16438
rect 10333 -16472 10349 -16438
rect 10273 -16488 10349 -16472
rect 10296 -16545 10330 -16488
rect 10277 -16598 10287 -16545
rect 10340 -16598 10350 -16545
rect 10185 -16718 10195 -16665
rect 10248 -16718 10258 -16665
rect 10383 -16781 10417 -16400
rect 10451 -16438 10527 -16432
rect 10451 -16472 10467 -16438
rect 10511 -16472 10527 -16438
rect 10451 -16488 10527 -16472
rect 10561 -16665 10595 -16400
rect 10629 -16438 10705 -16432
rect 10629 -16472 10645 -16438
rect 10689 -16472 10705 -16438
rect 10629 -16488 10705 -16472
rect 10540 -16718 10550 -16665
rect 10603 -16718 10613 -16665
rect 10739 -16779 10773 -16400
rect 10807 -16438 10883 -16432
rect 10807 -16472 10823 -16438
rect 10867 -16472 10883 -16438
rect 10807 -16488 10883 -16472
rect 10917 -16665 10951 -16400
rect 10985 -16437 11061 -16432
rect 11094 -16437 11128 -16400
rect 11163 -16437 11239 -16432
rect 10985 -16438 11239 -16437
rect 10985 -16472 11001 -16438
rect 11045 -16471 11179 -16438
rect 11045 -16472 11061 -16471
rect 10985 -16488 11061 -16472
rect 11163 -16472 11179 -16471
rect 11223 -16472 11239 -16438
rect 11163 -16488 11239 -16472
rect 10897 -16718 10907 -16665
rect 10960 -16718 10970 -16665
rect 10007 -16834 10017 -16781
rect 10070 -16834 10080 -16781
rect 10364 -16834 10374 -16781
rect 10427 -16834 10437 -16781
rect 10721 -16832 10731 -16779
rect 10784 -16832 10794 -16779
rect 11273 -16890 11307 -16400
rect 11341 -16438 11417 -16432
rect 11341 -16472 11357 -16438
rect 11401 -16472 11417 -16438
rect 11341 -16488 11417 -16472
rect 11519 -16438 11595 -16432
rect 11519 -16472 11535 -16438
rect 11579 -16472 11595 -16438
rect 11519 -16488 11595 -16472
rect 11362 -16545 11396 -16488
rect 11342 -16598 11352 -16545
rect 11405 -16598 11415 -16545
rect 11540 -16546 11574 -16488
rect 11520 -16599 11530 -16546
rect 11583 -16599 11593 -16546
rect 11630 -16890 11664 -16400
rect 11697 -16438 11773 -16432
rect 11697 -16472 11713 -16438
rect 11757 -16472 11773 -16438
rect 11697 -16488 11773 -16472
rect 11875 -16438 11951 -16432
rect 11875 -16472 11891 -16438
rect 11935 -16472 11951 -16438
rect 11875 -16488 11951 -16472
rect 11718 -16545 11752 -16488
rect 11699 -16598 11709 -16545
rect 11762 -16598 11772 -16545
rect 11985 -16889 12019 -16400
rect 12053 -16438 12129 -16432
rect 12053 -16472 12069 -16438
rect 12113 -16472 12129 -16438
rect 12053 -16488 12129 -16472
rect 12231 -16438 12307 -16432
rect 12231 -16472 12247 -16438
rect 12291 -16472 12307 -16438
rect 12231 -16488 12307 -16472
rect 12340 -16889 12374 -16400
rect 12409 -16438 12485 -16432
rect 12409 -16472 12425 -16438
rect 12469 -16472 12485 -16438
rect 12409 -16488 12485 -16472
rect 12520 -16440 12554 -16400
rect 12587 -16438 12663 -16432
rect 12587 -16440 12603 -16438
rect 12520 -16472 12603 -16440
rect 12647 -16440 12663 -16438
rect 12698 -16440 12732 -16400
rect 12647 -16472 12732 -16440
rect 12520 -16474 12732 -16472
rect 12587 -16488 12663 -16474
rect 11253 -16943 11263 -16890
rect 11316 -16943 11326 -16890
rect 11610 -16943 11620 -16890
rect 11673 -16943 11683 -16890
rect 11965 -16942 11975 -16889
rect 12028 -16942 12038 -16889
rect 12321 -16942 12331 -16889
rect 12384 -16942 12394 -16889
rect 13022 -17251 13075 -11726
rect 18337 -13421 18412 -6822
rect 18327 -13496 18337 -13421
rect 18412 -13496 18422 -13421
rect 18337 -13506 18412 -13496
rect -7605 -17459 13720 -17251
rect -7605 -17559 -7323 -17459
rect 13384 -17527 13720 -17459
rect 13384 -17559 13719 -17527
rect -7605 -17587 13719 -17559
<< via1 >>
rect 7145 2707 7197 2717
rect 7145 2673 7154 2707
rect 7154 2673 7188 2707
rect 7188 2673 7197 2707
rect 7145 2665 7197 2673
rect 7337 2707 7389 2717
rect 7337 2673 7346 2707
rect 7346 2673 7380 2707
rect 7380 2673 7389 2707
rect 7337 2665 7389 2673
rect 7529 2707 7581 2717
rect 7529 2673 7538 2707
rect 7538 2673 7572 2707
rect 7572 2673 7581 2707
rect 7529 2665 7581 2673
rect 7721 2707 7773 2717
rect 7721 2673 7730 2707
rect 7730 2673 7764 2707
rect 7764 2673 7773 2707
rect 7721 2665 7773 2673
rect 7912 2707 7964 2717
rect 7912 2673 7922 2707
rect 7922 2673 7956 2707
rect 7956 2673 7964 2707
rect 7912 2665 7964 2673
rect 8105 2707 8157 2717
rect 8105 2673 8114 2707
rect 8114 2673 8148 2707
rect 8148 2673 8157 2707
rect 8105 2665 8157 2673
rect -5867 -1963 -5814 -1910
rect -5689 -1963 -5636 -1910
rect -5510 -1963 -5457 -1910
rect -5333 -1963 -5280 -1910
rect -5155 -1963 -5102 -1910
rect -4976 -1963 -4923 -1910
rect -4799 -1963 -4746 -1910
rect -4621 -1963 -4568 -1910
rect -4443 -1963 -4390 -1910
rect -4265 -1963 -4212 -1910
rect -4086 -1963 -4033 -1910
rect -3909 -1963 -3856 -1910
rect -1109 -1963 -1056 -1910
rect -6498 -2582 -6445 -2529
rect -6625 -3454 -6572 -3401
rect -6044 -2833 -5991 -2780
rect -5777 -2583 -5724 -2530
rect -5866 -2833 -5813 -2780
rect -5421 -2721 -5368 -2668
rect -5066 -2583 -5013 -2530
rect -4710 -2721 -4657 -2668
rect -4354 -2583 -4301 -2530
rect -3998 -2721 -3945 -2668
rect -3908 -2833 -3855 -2780
rect -1109 -2478 -1056 -2425
rect -752 -2478 -699 -2425
rect -2624 -2611 -2571 -2558
rect -1285 -2611 -1232 -2558
rect -3298 -2721 -3245 -2668
rect -3731 -2833 -3678 -2780
rect -6134 -3454 -6081 -3401
rect -6498 -3693 -6445 -3640
rect -5777 -3569 -5724 -3516
rect -5422 -3693 -5369 -3640
rect -5066 -3454 -5013 -3401
rect -4710 -3454 -4657 -3401
rect -4353 -3693 -4300 -3640
rect -3998 -3569 -3945 -3516
rect -3642 -3454 -3589 -3401
rect -3131 -3454 -3078 -3401
rect -3298 -3569 -3245 -3516
rect -6498 -4324 -6445 -4271
rect -6134 -4443 -6081 -4390
rect -5778 -4324 -5725 -4271
rect -5422 -4559 -5369 -4506
rect -5066 -4443 -5013 -4390
rect -4709 -4443 -4656 -4390
rect -4353 -4559 -4300 -4506
rect -3998 -4324 -3945 -4271
rect -3642 -4443 -3589 -4390
rect -3298 -4559 -3245 -4506
rect -6498 -5194 -6445 -5141
rect -6625 -5375 -6572 -5322
rect -6134 -5285 -6081 -5232
rect -5777 -5468 -5724 -5415
rect -5422 -5194 -5369 -5141
rect -5066 -5286 -5013 -5233
rect -4710 -5375 -4657 -5322
rect -4353 -5194 -4300 -5141
rect -3997 -5468 -3944 -5415
rect -3642 -5372 -3589 -5319
rect -3130 -5286 -3077 -5233
rect -1197 -2718 -1144 -2665
rect -930 -2611 -877 -2558
rect -1019 -2718 -966 -2665
rect -841 -2718 -788 -2665
rect -129 -2718 -76 -2665
rect 50 -2718 103 -2665
rect 227 -2718 280 -2665
rect 5337 -2258 5390 -2205
rect 1919 -2479 1972 -2426
rect 2275 -2479 2328 -2426
rect 940 -2718 993 -2665
rect 1117 -2718 1170 -2665
rect 1295 -2718 1348 -2665
rect 2097 -2607 2150 -2554
rect 2007 -2718 2060 -2665
rect 2186 -2718 2239 -2665
rect 3193 -2480 3246 -2427
rect 2453 -2607 2506 -2554
rect 2363 -2718 2416 -2665
rect -1645 -3510 -1584 -3449
rect -2004 -4465 -1951 -4412
rect -2624 -5377 -2571 -5324
rect -3298 -5469 -3245 -5416
rect -5956 -6069 -5903 -6016
rect -5601 -6069 -5548 -6016
rect -5778 -6184 -5725 -6131
rect -5244 -6069 -5191 -6016
rect -5065 -6184 -5012 -6131
rect -6498 -6301 -6445 -6248
rect -5421 -6301 -5368 -6248
rect -4888 -6069 -4835 -6016
rect -4710 -6301 -4657 -6248
rect -4532 -6069 -4479 -6016
rect -4175 -6069 -4122 -6016
rect -4354 -6184 -4301 -6131
rect -3820 -6069 -3767 -6016
rect -2624 -6060 -2571 -6007
rect -3298 -6184 -3245 -6131
rect -3998 -6300 -3945 -6247
rect -4786 -6431 -4733 -6378
rect -1876 -5285 -1823 -5232
rect -1286 -3624 -1233 -3571
rect -1108 -3509 -1055 -3456
rect -929 -3624 -876 -3571
rect -484 -3354 -431 -3301
rect -750 -3509 -697 -3456
rect -396 -3509 -343 -3456
rect -573 -3624 -520 -3571
rect -217 -3624 -164 -3571
rect 583 -3354 636 -3301
rect -39 -3509 14 -3456
rect 317 -3509 370 -3456
rect 850 -3509 903 -3456
rect 1206 -3509 1259 -3456
rect 1654 -3354 1707 -3301
rect 1562 -3509 1615 -3456
rect 1919 -3509 1972 -3456
rect 1384 -3617 1437 -3564
rect 1741 -3617 1794 -3564
rect 2097 -3617 2150 -3564
rect 2275 -3509 2328 -3456
rect 2451 -3617 2504 -3564
rect -841 -4245 -788 -4192
rect -662 -4245 -609 -4192
rect -483 -4245 -430 -4192
rect -306 -4245 -253 -4192
rect 407 -4245 460 -4192
rect 317 -4357 370 -4304
rect 583 -4245 636 -4192
rect 495 -4465 548 -4412
rect 761 -4245 814 -4192
rect 673 -4357 726 -4304
rect 850 -4465 903 -4412
rect 1474 -4245 1527 -4192
rect 1652 -4245 1705 -4192
rect 1830 -4245 1883 -4192
rect 2008 -4245 2061 -4192
rect 2538 -4327 2599 -4266
rect 2746 -4507 2807 -4446
rect -1287 -5150 -1234 -5097
rect -1646 -5339 -1585 -5278
rect -1105 -5266 -1052 -5213
rect -929 -5150 -876 -5097
rect -572 -5150 -519 -5097
rect -218 -5150 -165 -5097
rect -751 -5266 -698 -5213
rect -396 -5266 -343 -5213
rect -41 -5266 12 -5213
rect 316 -5266 369 -5213
rect -128 -5433 -75 -5380
rect 50 -5433 103 -5380
rect 228 -5433 281 -5380
rect 850 -5266 903 -5213
rect 1207 -5266 1260 -5213
rect 940 -5434 993 -5381
rect 1119 -5433 1172 -5380
rect 1385 -5146 1438 -5093
rect 1296 -5433 1349 -5380
rect 1740 -5146 1793 -5093
rect 1563 -5266 1616 -5213
rect 1917 -5266 1970 -5213
rect 2096 -5146 2149 -5093
rect 2274 -5266 2327 -5213
rect 2453 -5146 2506 -5093
rect -1876 -6417 -1823 -6364
rect -1282 -6417 -1229 -6364
rect -928 -6417 -876 -6365
rect -1110 -6532 -1057 -6479
rect -752 -6532 -699 -6479
rect 227 -6303 280 -6250
rect 942 -6303 995 -6250
rect 2096 -6060 2149 -6007
rect 2452 -6060 2505 -6007
rect 1918 -6177 1971 -6124
rect 2275 -6177 2328 -6124
rect 3194 -4857 3246 -4805
rect 4771 -4857 4823 -4805
rect 2879 -6417 2931 -6365
rect 5037 -5059 5090 -5006
rect 4905 -5265 4958 -5212
rect -753 -6651 -700 -6598
rect 4772 -6650 4825 -6597
rect -2003 -6767 -1950 -6714
rect 8080 2162 8144 2226
rect 8382 2665 8434 2717
rect 16145 2707 16197 2717
rect 16145 2673 16154 2707
rect 16154 2673 16188 2707
rect 16188 2673 16197 2707
rect 16145 2665 16197 2673
rect 16337 2707 16389 2717
rect 16337 2673 16346 2707
rect 16346 2673 16380 2707
rect 16380 2673 16389 2707
rect 16337 2665 16389 2673
rect 16529 2707 16581 2717
rect 16529 2673 16538 2707
rect 16538 2673 16572 2707
rect 16572 2673 16581 2707
rect 16529 2665 16581 2673
rect 16721 2707 16773 2717
rect 16721 2673 16730 2707
rect 16730 2673 16764 2707
rect 16764 2673 16773 2707
rect 16721 2665 16773 2673
rect 16912 2707 16964 2717
rect 16912 2673 16922 2707
rect 16922 2673 16956 2707
rect 16956 2673 16964 2707
rect 16912 2665 16964 2673
rect 17105 2707 17157 2717
rect 17105 2673 17114 2707
rect 17114 2673 17148 2707
rect 17148 2673 17157 2707
rect 17105 2665 17157 2673
rect 7145 1899 7197 1909
rect 7145 1865 7154 1899
rect 7154 1865 7188 1899
rect 7188 1865 7197 1899
rect 7145 1857 7197 1865
rect 7337 1899 7389 1909
rect 7337 1865 7346 1899
rect 7346 1865 7380 1899
rect 7380 1865 7389 1899
rect 7337 1857 7389 1865
rect 7530 1899 7582 1910
rect 7530 1865 7538 1899
rect 7538 1865 7572 1899
rect 7572 1865 7582 1899
rect 7530 1858 7582 1865
rect 7722 1899 7774 1910
rect 7722 1865 7730 1899
rect 7730 1865 7764 1899
rect 7764 1865 7774 1899
rect 7722 1858 7774 1865
rect 7914 1899 7966 1910
rect 7914 1865 7922 1899
rect 7922 1865 7956 1899
rect 7956 1865 7966 1899
rect 7914 1858 7966 1865
rect 8105 1899 8157 1910
rect 8105 1865 8114 1899
rect 8114 1865 8148 1899
rect 8148 1865 8157 1899
rect 8105 1858 8157 1865
rect 15793 2164 15857 2228
rect 8382 1858 8434 1910
rect 7145 907 7197 917
rect 7145 873 7154 907
rect 7154 873 7188 907
rect 7188 873 7197 907
rect 7145 865 7197 873
rect 7337 907 7389 917
rect 7337 873 7346 907
rect 7346 873 7380 907
rect 7380 873 7389 907
rect 7337 865 7389 873
rect 7529 907 7581 917
rect 7529 873 7538 907
rect 7538 873 7572 907
rect 7572 873 7581 907
rect 7529 865 7581 873
rect 7721 907 7773 917
rect 7721 873 7730 907
rect 7730 873 7764 907
rect 7764 873 7773 907
rect 7721 865 7773 873
rect 7912 907 7964 917
rect 7912 873 7922 907
rect 7922 873 7956 907
rect 7956 873 7964 907
rect 7912 865 7964 873
rect 8105 907 8157 917
rect 8105 873 8114 907
rect 8114 873 8148 907
rect 8148 873 8157 907
rect 8105 865 8157 873
rect 8074 362 8138 426
rect 10730 943 10794 1007
rect 8382 865 8434 917
rect 7145 99 7197 109
rect 7145 65 7154 99
rect 7154 65 7188 99
rect 7188 65 7197 99
rect 7145 57 7197 65
rect 7337 99 7389 109
rect 7337 65 7346 99
rect 7346 65 7380 99
rect 7380 65 7389 99
rect 7337 57 7389 65
rect 7530 99 7582 110
rect 7530 65 7538 99
rect 7538 65 7572 99
rect 7572 65 7582 99
rect 7530 58 7582 65
rect 7722 99 7774 110
rect 7722 65 7730 99
rect 7730 65 7764 99
rect 7764 65 7774 99
rect 7722 58 7774 65
rect 7914 99 7966 110
rect 7914 65 7922 99
rect 7922 65 7956 99
rect 7956 65 7966 99
rect 7914 58 7966 65
rect 8105 99 8157 110
rect 8105 65 8114 99
rect 8114 65 8148 99
rect 8148 65 8157 99
rect 8105 58 8157 65
rect 8625 360 8689 424
rect 8382 58 8434 110
rect 7145 -893 7197 -883
rect 7145 -927 7154 -893
rect 7154 -927 7188 -893
rect 7188 -927 7197 -893
rect 7145 -935 7197 -927
rect 7337 -893 7389 -883
rect 7337 -927 7346 -893
rect 7346 -927 7380 -893
rect 7380 -927 7389 -893
rect 7337 -935 7389 -927
rect 7529 -893 7581 -883
rect 7529 -927 7538 -893
rect 7538 -927 7572 -893
rect 7572 -927 7581 -893
rect 7529 -935 7581 -927
rect 7721 -893 7773 -883
rect 7721 -927 7730 -893
rect 7730 -927 7764 -893
rect 7764 -927 7773 -893
rect 7721 -935 7773 -927
rect 7912 -893 7964 -883
rect 7912 -927 7922 -893
rect 7922 -927 7956 -893
rect 7956 -927 7964 -893
rect 7912 -935 7964 -927
rect 8105 -893 8157 -883
rect 8105 -927 8114 -893
rect 8114 -927 8148 -893
rect 8148 -927 8157 -893
rect 8105 -935 8157 -927
rect 8078 -1438 8142 -1374
rect 8382 -935 8434 -883
rect 7145 -1701 7197 -1691
rect 7145 -1735 7154 -1701
rect 7154 -1735 7188 -1701
rect 7188 -1735 7197 -1701
rect 7145 -1743 7197 -1735
rect 7337 -1701 7389 -1691
rect 7337 -1735 7346 -1701
rect 7346 -1735 7380 -1701
rect 7380 -1735 7389 -1701
rect 7337 -1743 7389 -1735
rect 7530 -1701 7582 -1690
rect 7530 -1735 7538 -1701
rect 7538 -1735 7572 -1701
rect 7572 -1735 7582 -1701
rect 7530 -1742 7582 -1735
rect 7722 -1701 7774 -1690
rect 7722 -1735 7730 -1701
rect 7730 -1735 7764 -1701
rect 7764 -1735 7774 -1701
rect 7722 -1742 7774 -1735
rect 7914 -1701 7966 -1690
rect 7914 -1735 7922 -1701
rect 7922 -1735 7956 -1701
rect 7956 -1735 7966 -1701
rect 7914 -1742 7966 -1735
rect 8105 -1701 8157 -1690
rect 8105 -1735 8114 -1701
rect 8114 -1735 8148 -1701
rect 8148 -1735 8157 -1701
rect 8105 -1742 8157 -1735
rect 8668 -1439 8732 -1375
rect 17382 2665 17434 2717
rect 16145 1899 16197 1909
rect 16145 1865 16154 1899
rect 16154 1865 16188 1899
rect 16188 1865 16197 1899
rect 16145 1857 16197 1865
rect 16337 1899 16389 1909
rect 16337 1865 16346 1899
rect 16346 1865 16380 1899
rect 16380 1865 16389 1899
rect 16337 1857 16389 1865
rect 16530 1899 16582 1910
rect 16530 1865 16538 1899
rect 16538 1865 16572 1899
rect 16572 1865 16582 1899
rect 16530 1858 16582 1865
rect 16722 1899 16774 1910
rect 16722 1865 16730 1899
rect 16730 1865 16764 1899
rect 16764 1865 16774 1899
rect 16722 1858 16774 1865
rect 16914 1899 16966 1910
rect 16914 1865 16922 1899
rect 16922 1865 16956 1899
rect 16956 1865 16966 1899
rect 16914 1858 16966 1865
rect 17105 1899 17157 1910
rect 17105 1865 17114 1899
rect 17114 1865 17148 1899
rect 17148 1865 17157 1899
rect 17105 1858 17157 1865
rect 17382 1858 17434 1910
rect 16145 907 16197 917
rect 16145 873 16154 907
rect 16154 873 16188 907
rect 16188 873 16197 907
rect 16145 865 16197 873
rect 16337 907 16389 917
rect 16337 873 16346 907
rect 16346 873 16380 907
rect 16380 873 16389 907
rect 16337 865 16389 873
rect 16529 907 16581 917
rect 16529 873 16538 907
rect 16538 873 16572 907
rect 16572 873 16581 907
rect 16529 865 16581 873
rect 16721 907 16773 917
rect 16721 873 16730 907
rect 16730 873 16764 907
rect 16764 873 16773 907
rect 16721 865 16773 873
rect 16912 907 16964 917
rect 16912 873 16922 907
rect 16922 873 16956 907
rect 16956 873 16964 907
rect 16912 865 16964 873
rect 17105 907 17157 917
rect 17105 873 17114 907
rect 17114 873 17148 907
rect 17148 873 17157 907
rect 17105 865 17157 873
rect 15806 362 15870 426
rect 12259 25 12323 89
rect 17382 865 17434 917
rect 16145 99 16197 109
rect 16145 65 16154 99
rect 16154 65 16188 99
rect 16188 65 16197 99
rect 16145 57 16197 65
rect 16337 99 16389 109
rect 16337 65 16346 99
rect 16346 65 16380 99
rect 16380 65 16389 99
rect 16337 57 16389 65
rect 16530 99 16582 110
rect 16530 65 16538 99
rect 16538 65 16572 99
rect 16572 65 16582 99
rect 16530 58 16582 65
rect 16722 99 16774 110
rect 16722 65 16730 99
rect 16730 65 16764 99
rect 16764 65 16774 99
rect 16722 58 16774 65
rect 16914 99 16966 110
rect 16914 65 16922 99
rect 16922 65 16956 99
rect 16956 65 16966 99
rect 16914 58 16966 65
rect 17105 99 17157 110
rect 17105 65 17114 99
rect 17114 65 17148 99
rect 17148 65 17157 99
rect 17105 58 17157 65
rect 17382 58 17434 110
rect 12259 -449 12323 -385
rect 12870 -605 12934 -541
rect 15268 -601 15332 -537
rect 12208 -970 12272 -906
rect 14309 -1143 14373 -1079
rect 12410 -1321 12474 -1257
rect 8382 -1742 8434 -1690
rect 9435 -2050 9499 -1986
rect 10733 -2050 10797 -1986
rect 6680 -2263 6744 -2199
rect 9435 -2379 9499 -2315
rect 7145 -2693 7197 -2683
rect 7145 -2727 7154 -2693
rect 7154 -2727 7188 -2693
rect 7188 -2727 7197 -2693
rect 7145 -2735 7197 -2727
rect 7337 -2693 7389 -2683
rect 7337 -2727 7346 -2693
rect 7346 -2727 7380 -2693
rect 7380 -2727 7389 -2693
rect 7337 -2735 7389 -2727
rect 7529 -2693 7581 -2683
rect 7529 -2727 7538 -2693
rect 7538 -2727 7572 -2693
rect 7572 -2727 7581 -2693
rect 7529 -2735 7581 -2727
rect 7721 -2693 7773 -2683
rect 7721 -2727 7730 -2693
rect 7730 -2727 7764 -2693
rect 7764 -2727 7773 -2693
rect 7721 -2735 7773 -2727
rect 7912 -2693 7964 -2683
rect 7912 -2727 7922 -2693
rect 7922 -2727 7956 -2693
rect 7956 -2727 7964 -2693
rect 7912 -2735 7964 -2727
rect 8105 -2693 8157 -2683
rect 8105 -2727 8114 -2693
rect 8114 -2727 8148 -2693
rect 8148 -2727 8157 -2693
rect 8105 -2735 8157 -2727
rect 6222 -3515 6286 -3451
rect 8075 -3238 8139 -3174
rect 8382 -2735 8434 -2683
rect 7145 -3501 7197 -3491
rect 7145 -3535 7154 -3501
rect 7154 -3535 7188 -3501
rect 7188 -3535 7197 -3501
rect 7145 -3543 7197 -3535
rect 7337 -3501 7389 -3491
rect 7337 -3535 7346 -3501
rect 7346 -3535 7380 -3501
rect 7380 -3535 7389 -3501
rect 7337 -3543 7389 -3535
rect 7530 -3501 7582 -3490
rect 7530 -3535 7538 -3501
rect 7538 -3535 7572 -3501
rect 7572 -3535 7582 -3501
rect 7530 -3542 7582 -3535
rect 7722 -3501 7774 -3490
rect 7722 -3535 7730 -3501
rect 7730 -3535 7764 -3501
rect 7764 -3535 7774 -3501
rect 7722 -3542 7774 -3535
rect 7914 -3501 7966 -3490
rect 7914 -3535 7922 -3501
rect 7922 -3535 7956 -3501
rect 7956 -3535 7966 -3501
rect 7914 -3542 7966 -3535
rect 8105 -3501 8157 -3490
rect 8105 -3535 8114 -3501
rect 8114 -3535 8148 -3501
rect 8148 -3535 8157 -3501
rect 8105 -3542 8157 -3535
rect 8668 -3242 8732 -3178
rect 16145 -893 16197 -883
rect 16145 -927 16154 -893
rect 16154 -927 16188 -893
rect 16188 -927 16197 -893
rect 16145 -935 16197 -927
rect 16337 -893 16389 -883
rect 16337 -927 16346 -893
rect 16346 -927 16380 -893
rect 16380 -927 16389 -893
rect 16337 -935 16389 -927
rect 16529 -893 16581 -883
rect 16529 -927 16538 -893
rect 16538 -927 16572 -893
rect 16572 -927 16581 -893
rect 16529 -935 16581 -927
rect 16721 -893 16773 -883
rect 16721 -927 16730 -893
rect 16730 -927 16764 -893
rect 16764 -927 16773 -893
rect 16721 -935 16773 -927
rect 16912 -893 16964 -883
rect 16912 -927 16922 -893
rect 16922 -927 16956 -893
rect 16956 -927 16964 -893
rect 16912 -935 16964 -927
rect 17105 -893 17157 -883
rect 17105 -927 17114 -893
rect 17114 -927 17148 -893
rect 17148 -927 17157 -893
rect 17105 -935 17157 -927
rect 15861 -1438 15925 -1374
rect 17382 -935 17434 -883
rect 13976 -1891 14040 -1827
rect 16145 -1701 16197 -1691
rect 16145 -1735 16154 -1701
rect 16154 -1735 16188 -1701
rect 16188 -1735 16197 -1701
rect 16145 -1743 16197 -1735
rect 16337 -1701 16389 -1691
rect 16337 -1735 16346 -1701
rect 16346 -1735 16380 -1701
rect 16380 -1735 16389 -1701
rect 16337 -1743 16389 -1735
rect 16530 -1701 16582 -1690
rect 16530 -1735 16538 -1701
rect 16538 -1735 16572 -1701
rect 16572 -1735 16582 -1701
rect 16530 -1742 16582 -1735
rect 16722 -1701 16774 -1690
rect 16722 -1735 16730 -1701
rect 16730 -1735 16764 -1701
rect 16764 -1735 16774 -1701
rect 16722 -1742 16774 -1735
rect 16914 -1701 16966 -1690
rect 16914 -1735 16922 -1701
rect 16922 -1735 16956 -1701
rect 16956 -1735 16966 -1701
rect 16914 -1742 16966 -1735
rect 17105 -1701 17157 -1690
rect 17105 -1735 17114 -1701
rect 17114 -1735 17148 -1701
rect 17148 -1735 17157 -1701
rect 17105 -1742 17157 -1735
rect 17382 -1742 17434 -1690
rect 16145 -2693 16197 -2683
rect 16145 -2727 16154 -2693
rect 16154 -2727 16188 -2693
rect 16188 -2727 16197 -2693
rect 16145 -2735 16197 -2727
rect 16337 -2693 16389 -2683
rect 16337 -2727 16346 -2693
rect 16346 -2727 16380 -2693
rect 16380 -2727 16389 -2693
rect 16337 -2735 16389 -2727
rect 16529 -2693 16581 -2683
rect 16529 -2727 16538 -2693
rect 16538 -2727 16572 -2693
rect 16572 -2727 16581 -2693
rect 16529 -2735 16581 -2727
rect 16721 -2693 16773 -2683
rect 16721 -2727 16730 -2693
rect 16730 -2727 16764 -2693
rect 16764 -2727 16773 -2693
rect 16721 -2735 16773 -2727
rect 16912 -2693 16964 -2683
rect 16912 -2727 16922 -2693
rect 16922 -2727 16956 -2693
rect 16956 -2727 16964 -2693
rect 16912 -2735 16964 -2727
rect 17105 -2693 17157 -2683
rect 17105 -2727 17114 -2693
rect 17114 -2727 17148 -2693
rect 17148 -2727 17157 -2693
rect 17105 -2735 17157 -2727
rect 15866 -3236 15930 -3172
rect 12410 -3310 12474 -3246
rect 8382 -3542 8434 -3490
rect 17382 -2735 17434 -2683
rect 16145 -3501 16197 -3491
rect 16145 -3535 16154 -3501
rect 16154 -3535 16188 -3501
rect 16188 -3535 16197 -3501
rect 16145 -3543 16197 -3535
rect 16337 -3501 16389 -3491
rect 16337 -3535 16346 -3501
rect 16346 -3535 16380 -3501
rect 16380 -3535 16389 -3501
rect 16337 -3543 16389 -3535
rect 16530 -3501 16582 -3490
rect 16530 -3535 16538 -3501
rect 16538 -3535 16572 -3501
rect 16572 -3535 16582 -3501
rect 16530 -3542 16582 -3535
rect 16722 -3501 16774 -3490
rect 16722 -3535 16730 -3501
rect 16730 -3535 16764 -3501
rect 16764 -3535 16774 -3501
rect 16722 -3542 16774 -3535
rect 16914 -3501 16966 -3490
rect 16914 -3535 16922 -3501
rect 16922 -3535 16956 -3501
rect 16956 -3535 16966 -3501
rect 16914 -3542 16966 -3535
rect 17105 -3501 17157 -3490
rect 17105 -3535 17114 -3501
rect 17114 -3535 17148 -3501
rect 17148 -3535 17157 -3501
rect 17105 -3542 17157 -3535
rect 17382 -3542 17434 -3490
rect 11432 -3893 11496 -3829
rect 7145 -4493 7197 -4483
rect 7145 -4527 7154 -4493
rect 7154 -4527 7188 -4493
rect 7188 -4527 7197 -4493
rect 7145 -4535 7197 -4527
rect 7337 -4493 7389 -4483
rect 7337 -4527 7346 -4493
rect 7346 -4527 7380 -4493
rect 7380 -4527 7389 -4493
rect 7337 -4535 7389 -4527
rect 7529 -4493 7581 -4483
rect 7529 -4527 7538 -4493
rect 7538 -4527 7572 -4493
rect 7572 -4527 7581 -4493
rect 7529 -4535 7581 -4527
rect 7721 -4493 7773 -4483
rect 7721 -4527 7730 -4493
rect 7730 -4527 7764 -4493
rect 7764 -4527 7773 -4493
rect 7721 -4535 7773 -4527
rect 7912 -4493 7964 -4483
rect 7912 -4527 7922 -4493
rect 7922 -4527 7956 -4493
rect 7956 -4527 7964 -4493
rect 7912 -4535 7964 -4527
rect 8105 -4493 8157 -4483
rect 8105 -4527 8114 -4493
rect 8114 -4527 8148 -4493
rect 8148 -4527 8157 -4493
rect 8105 -4535 8157 -4527
rect 5614 -5271 5678 -5207
rect 5337 -5580 5390 -5527
rect 8082 -5036 8146 -4972
rect 8382 -4535 8434 -4483
rect 12704 -4007 12768 -3943
rect 15254 -4007 15318 -3943
rect 9272 -4192 9336 -4128
rect 13428 -4192 13492 -4128
rect 16145 -4493 16197 -4483
rect 16145 -4527 16154 -4493
rect 16154 -4527 16188 -4493
rect 16188 -4527 16197 -4493
rect 16145 -4535 16197 -4527
rect 16337 -4493 16389 -4483
rect 16337 -4527 16346 -4493
rect 16346 -4527 16380 -4493
rect 16380 -4527 16389 -4493
rect 16337 -4535 16389 -4527
rect 16529 -4493 16581 -4483
rect 16529 -4527 16538 -4493
rect 16538 -4527 16572 -4493
rect 16572 -4527 16581 -4493
rect 16529 -4535 16581 -4527
rect 16721 -4493 16773 -4483
rect 16721 -4527 16730 -4493
rect 16730 -4527 16764 -4493
rect 16764 -4527 16773 -4493
rect 16721 -4535 16773 -4527
rect 16912 -4493 16964 -4483
rect 16912 -4527 16922 -4493
rect 16922 -4527 16956 -4493
rect 16956 -4527 16964 -4493
rect 16912 -4535 16964 -4527
rect 17105 -4493 17157 -4483
rect 17105 -4527 17114 -4493
rect 17114 -4527 17148 -4493
rect 17148 -4527 17157 -4493
rect 17105 -4535 17157 -4527
rect 7145 -5301 7197 -5291
rect 7145 -5335 7154 -5301
rect 7154 -5335 7188 -5301
rect 7188 -5335 7197 -5301
rect 7145 -5343 7197 -5335
rect 7337 -5301 7389 -5291
rect 7337 -5335 7346 -5301
rect 7346 -5335 7380 -5301
rect 7380 -5335 7389 -5301
rect 7337 -5343 7389 -5335
rect 7530 -5301 7582 -5290
rect 7530 -5335 7538 -5301
rect 7538 -5335 7572 -5301
rect 7572 -5335 7582 -5301
rect 7530 -5342 7582 -5335
rect 7722 -5301 7774 -5290
rect 7722 -5335 7730 -5301
rect 7730 -5335 7764 -5301
rect 7764 -5335 7774 -5301
rect 7722 -5342 7774 -5335
rect 7914 -5301 7966 -5290
rect 7914 -5335 7922 -5301
rect 7922 -5335 7956 -5301
rect 7956 -5335 7966 -5301
rect 7914 -5342 7966 -5335
rect 8105 -5301 8157 -5290
rect 8105 -5335 8114 -5301
rect 8114 -5335 8148 -5301
rect 8148 -5335 8157 -5301
rect 8105 -5342 8157 -5335
rect 15802 -5040 15866 -4976
rect 8382 -5342 8434 -5290
rect 17382 -4535 17434 -4483
rect 16145 -5301 16197 -5291
rect 16145 -5335 16154 -5301
rect 16154 -5335 16188 -5301
rect 16188 -5335 16197 -5301
rect 16145 -5343 16197 -5335
rect 16337 -5301 16389 -5291
rect 16337 -5335 16346 -5301
rect 16346 -5335 16380 -5301
rect 16380 -5335 16389 -5301
rect 16337 -5343 16389 -5335
rect 16530 -5301 16582 -5290
rect 16530 -5335 16538 -5301
rect 16538 -5335 16572 -5301
rect 16572 -5335 16582 -5301
rect 16530 -5342 16582 -5335
rect 16722 -5301 16774 -5290
rect 16722 -5335 16730 -5301
rect 16730 -5335 16764 -5301
rect 16764 -5335 16774 -5301
rect 16722 -5342 16774 -5335
rect 16914 -5301 16966 -5290
rect 16914 -5335 16922 -5301
rect 16922 -5335 16956 -5301
rect 16956 -5335 16966 -5301
rect 16914 -5342 16966 -5335
rect 17105 -5301 17157 -5290
rect 17105 -5335 17114 -5301
rect 17114 -5335 17148 -5301
rect 17148 -5335 17157 -5301
rect 17105 -5342 17157 -5335
rect 17382 -5342 17434 -5290
rect 7145 -6293 7197 -6283
rect 7145 -6327 7154 -6293
rect 7154 -6327 7188 -6293
rect 7188 -6327 7197 -6293
rect 7145 -6335 7197 -6327
rect 7337 -6293 7389 -6283
rect 7337 -6327 7346 -6293
rect 7346 -6327 7380 -6293
rect 7380 -6327 7389 -6293
rect 7337 -6335 7389 -6327
rect 7529 -6293 7581 -6283
rect 7529 -6327 7538 -6293
rect 7538 -6327 7572 -6293
rect 7572 -6327 7581 -6293
rect 7529 -6335 7581 -6327
rect 7721 -6293 7773 -6283
rect 7721 -6327 7730 -6293
rect 7730 -6327 7764 -6293
rect 7764 -6327 7773 -6293
rect 7721 -6335 7773 -6327
rect 7912 -6293 7964 -6283
rect 7912 -6327 7922 -6293
rect 7922 -6327 7956 -6293
rect 7956 -6327 7964 -6293
rect 7912 -6335 7964 -6327
rect 8105 -6293 8157 -6283
rect 8105 -6327 8114 -6293
rect 8114 -6327 8148 -6293
rect 8148 -6327 8157 -6293
rect 8105 -6335 8157 -6327
rect 4770 -6944 4823 -6891
rect 4906 -6942 4959 -6889
rect 5038 -6940 5091 -6887
rect 8083 -6837 8147 -6773
rect 8382 -6335 8434 -6283
rect 16145 -6293 16197 -6283
rect 16145 -6327 16154 -6293
rect 16154 -6327 16188 -6293
rect 16188 -6327 16197 -6293
rect 16145 -6335 16197 -6327
rect 16337 -6293 16389 -6283
rect 16337 -6327 16346 -6293
rect 16346 -6327 16380 -6293
rect 16380 -6327 16389 -6293
rect 16337 -6335 16389 -6327
rect 16529 -6293 16581 -6283
rect 16529 -6327 16538 -6293
rect 16538 -6327 16572 -6293
rect 16572 -6327 16581 -6293
rect 16529 -6335 16581 -6327
rect 16721 -6293 16773 -6283
rect 16721 -6327 16730 -6293
rect 16730 -6327 16764 -6293
rect 16764 -6327 16773 -6293
rect 16721 -6335 16773 -6327
rect 16912 -6293 16964 -6283
rect 16912 -6327 16922 -6293
rect 16922 -6327 16956 -6293
rect 16956 -6327 16964 -6293
rect 16912 -6335 16964 -6327
rect 17105 -6293 17157 -6283
rect 17105 -6327 17114 -6293
rect 17114 -6327 17148 -6293
rect 17148 -6327 17157 -6293
rect 17105 -6335 17157 -6327
rect 7145 -7101 7197 -7091
rect 7145 -7135 7154 -7101
rect 7154 -7135 7188 -7101
rect 7188 -7135 7197 -7101
rect 7145 -7143 7197 -7135
rect 7337 -7101 7389 -7091
rect 7337 -7135 7346 -7101
rect 7346 -7135 7380 -7101
rect 7380 -7135 7389 -7101
rect 7337 -7143 7389 -7135
rect 7530 -7101 7582 -7090
rect 7530 -7135 7538 -7101
rect 7538 -7135 7572 -7101
rect 7572 -7135 7582 -7101
rect 7530 -7142 7582 -7135
rect 7722 -7101 7774 -7090
rect 7722 -7135 7730 -7101
rect 7730 -7135 7764 -7101
rect 7764 -7135 7774 -7101
rect 7722 -7142 7774 -7135
rect 7914 -7101 7966 -7090
rect 7914 -7135 7922 -7101
rect 7922 -7135 7956 -7101
rect 7956 -7135 7966 -7101
rect 7914 -7142 7966 -7135
rect 8105 -7101 8157 -7090
rect 8105 -7135 8114 -7101
rect 8114 -7135 8148 -7101
rect 8148 -7135 8157 -7101
rect 8105 -7142 8157 -7135
rect 8600 -6834 8664 -6770
rect 15820 -6832 15884 -6768
rect 8382 -7142 8434 -7090
rect 17382 -6335 17434 -6283
rect 17831 -6585 17895 -6521
rect 16145 -7101 16197 -7091
rect 16145 -7135 16154 -7101
rect 16154 -7135 16188 -7101
rect 16188 -7135 16197 -7101
rect 16145 -7143 16197 -7135
rect 16337 -7101 16389 -7091
rect 16337 -7135 16346 -7101
rect 16346 -7135 16380 -7101
rect 16380 -7135 16389 -7101
rect 16337 -7143 16389 -7135
rect 16530 -7101 16582 -7090
rect 16530 -7135 16538 -7101
rect 16538 -7135 16572 -7101
rect 16572 -7135 16582 -7101
rect 16530 -7142 16582 -7135
rect 16722 -7101 16774 -7090
rect 16722 -7135 16730 -7101
rect 16730 -7135 16764 -7101
rect 16764 -7135 16774 -7101
rect 16722 -7142 16774 -7135
rect 16914 -7101 16966 -7090
rect 16914 -7135 16922 -7101
rect 16922 -7135 16956 -7101
rect 16956 -7135 16966 -7101
rect 16914 -7142 16966 -7135
rect 17105 -7101 17157 -7090
rect 17105 -7135 17114 -7101
rect 17114 -7135 17148 -7101
rect 17148 -7135 17157 -7101
rect 17105 -7142 17157 -7135
rect 17382 -7142 17434 -7090
rect -3873 -7743 -3821 -7691
rect -3731 -7837 -3679 -7785
rect -3541 -7840 -3489 -7788
rect -5502 -12324 -5449 -12271
rect -6077 -12565 -6024 -12512
rect -5626 -12565 -5573 -12512
rect -6223 -13115 -6170 -13062
rect -6426 -13905 -6373 -13852
rect -5000 -12325 -4947 -12272
rect -4502 -12324 -4449 -12271
rect -5376 -12441 -5323 -12388
rect -5127 -12441 -5074 -12388
rect -4877 -12565 -4824 -12512
rect -4627 -12565 -4574 -12512
rect -4377 -12441 -4324 -12388
rect -3928 -12442 -3875 -12389
rect -5751 -13115 -5698 -13062
rect -5251 -13242 -5198 -13189
rect -4752 -13115 -4699 -13062
rect -4251 -13242 -4198 -13189
rect -6077 -13798 -6024 -13745
rect -5376 -13798 -5323 -13745
rect -5626 -13905 -5573 -13852
rect -5730 -14010 -5677 -13957
rect -5126 -13798 -5073 -13745
rect -4877 -13905 -4824 -13852
rect -4376 -13798 -4323 -13745
rect -4627 -13905 -4574 -13852
rect -4752 -14010 -4699 -13957
rect -3788 -13242 -3735 -13189
rect -3928 -13905 -3875 -13852
rect -3788 -14010 -3735 -13957
rect -6223 -14108 -6170 -14055
rect -5250 -14108 -5197 -14055
rect -4250 -14108 -4197 -14055
rect -6159 -14848 -6106 -14795
rect -5860 -14848 -5807 -14795
rect -5504 -14954 -5451 -14901
rect -5147 -14848 -5094 -14795
rect -4791 -14954 -4738 -14901
rect -4436 -14848 -4383 -14795
rect 4771 -7907 4824 -7854
rect 4906 -7905 4959 -7852
rect 5037 -7903 5090 -7850
rect -3382 -7986 -3329 -7933
rect -1382 -7975 -1329 -7922
rect -3542 -13242 -3489 -13189
rect -1203 -7976 -1150 -7923
rect -1025 -7975 -972 -7922
rect -848 -7975 -795 -7922
rect -670 -7975 -617 -7922
rect -490 -7975 -437 -7922
rect 755 -7975 808 -7922
rect 932 -7975 985 -7922
rect 1112 -7975 1165 -7922
rect 1289 -7976 1342 -7923
rect 1467 -7975 1520 -7922
rect 1644 -7975 1697 -7922
rect 2890 -7975 2943 -7922
rect 3069 -7975 3122 -7922
rect 3247 -7975 3300 -7922
rect 3424 -7975 3477 -7922
rect 3603 -7976 3656 -7923
rect 3778 -7975 3831 -7922
rect 4208 -7976 4261 -7923
rect -1916 -8587 -1863 -8534
rect -1739 -8587 -1686 -8534
rect -1826 -8706 -1773 -8653
rect -2447 -8820 -2394 -8767
rect -2005 -8820 -1952 -8767
rect -1558 -8587 -1505 -8534
rect -1382 -8587 -1329 -8534
rect -1470 -8706 -1417 -8653
rect -1648 -8820 -1595 -8767
rect -1203 -8587 -1150 -8534
rect -1293 -8820 -1240 -8767
rect -1026 -8587 -973 -8534
rect -1115 -8706 -1062 -8653
rect -848 -8587 -795 -8534
rect -936 -8820 -883 -8767
rect -670 -8587 -617 -8534
rect -758 -8706 -705 -8653
rect -491 -8587 -438 -8534
rect -580 -8819 -527 -8766
rect -314 -8587 -261 -8534
rect -402 -8706 -349 -8653
rect -136 -8587 -83 -8534
rect 42 -8587 95 -8534
rect -47 -8706 6 -8653
rect -225 -8820 -172 -8767
rect 221 -8587 274 -8534
rect 398 -8587 451 -8534
rect 310 -8706 363 -8653
rect 132 -8821 185 -8768
rect 577 -8587 630 -8534
rect 754 -8587 807 -8534
rect 666 -8706 719 -8653
rect 489 -8819 542 -8766
rect 932 -8587 985 -8534
rect 843 -8819 896 -8766
rect 1111 -8587 1164 -8534
rect 1022 -8706 1075 -8653
rect 1289 -8587 1342 -8534
rect 1201 -8820 1254 -8767
rect 1466 -8587 1519 -8534
rect 1377 -8706 1430 -8653
rect 1644 -8587 1697 -8534
rect 1556 -8820 1609 -8767
rect 1822 -8587 1875 -8534
rect 1733 -8706 1786 -8653
rect 2000 -8587 2053 -8534
rect 2178 -8587 2231 -8534
rect 2090 -8706 2143 -8653
rect 1911 -8820 1964 -8767
rect 2357 -8587 2410 -8534
rect 2534 -8587 2587 -8534
rect 2446 -8706 2499 -8653
rect 2267 -8820 2320 -8767
rect 2712 -8587 2765 -8534
rect 2890 -8587 2943 -8534
rect 2802 -8706 2855 -8653
rect 2624 -8820 2677 -8767
rect 3068 -8587 3121 -8534
rect 2980 -8820 3033 -8767
rect 3246 -8587 3299 -8534
rect 3158 -8706 3211 -8653
rect 3424 -8587 3477 -8534
rect 3336 -8820 3389 -8767
rect 3602 -8587 3655 -8534
rect 3513 -8706 3566 -8653
rect 3781 -8587 3834 -8534
rect 3692 -8820 3745 -8767
rect 3869 -8706 3922 -8653
rect -2315 -9978 -2262 -9925
rect -2447 -12325 -2394 -12272
rect -3382 -14108 -3329 -14055
rect -3936 -14954 -3883 -14901
rect -6159 -15535 -6106 -15482
rect -5860 -15641 -5807 -15588
rect -5504 -15534 -5451 -15481
rect -5148 -15642 -5095 -15589
rect -4792 -15534 -4739 -15481
rect -4435 -15641 -4383 -15589
rect -3935 -15641 -3883 -15589
rect -6159 -16246 -6106 -16193
rect -5860 -16347 -5807 -16294
rect -5504 -16246 -5451 -16193
rect -5148 -16347 -5095 -16294
rect -4792 -16246 -4739 -16193
rect -4436 -16347 -4383 -16294
rect -1916 -9599 -1863 -9546
rect -1916 -9978 -1863 -9925
rect -1738 -9599 -1685 -9546
rect -1738 -9979 -1685 -9926
rect -1558 -9599 -1505 -9546
rect -1560 -9978 -1507 -9925
rect -1382 -9977 -1329 -9924
rect -312 -9599 -259 -9546
rect -314 -9978 -261 -9925
rect -136 -9598 -83 -9545
rect -136 -9979 -83 -9926
rect 42 -9599 95 -9546
rect 43 -9978 96 -9925
rect 222 -9598 275 -9545
rect 220 -9978 273 -9925
rect 399 -9599 452 -9546
rect 398 -9978 451 -9925
rect 577 -9599 630 -9546
rect 576 -9978 629 -9925
rect 2178 -9600 2231 -9547
rect 2357 -9599 2410 -9546
rect 2356 -9978 2409 -9925
rect 2534 -9599 2587 -9546
rect 2534 -9978 2587 -9925
rect 2713 -9599 2766 -9546
rect 2712 -9979 2765 -9926
rect 2891 -9978 2944 -9925
rect 3069 -9978 3122 -9925
rect 3246 -9978 3299 -9925
rect 4771 -9367 4824 -9314
rect 4208 -9599 4261 -9546
rect -1827 -10961 -1774 -10908
rect -1470 -10961 -1417 -10908
rect -1114 -10961 -1061 -10908
rect -758 -10961 -705 -10908
rect -402 -10961 -349 -10908
rect -46 -10961 7 -10908
rect 309 -10961 362 -10908
rect 665 -10961 718 -10908
rect 931 -10961 984 -10908
rect 1199 -10961 1252 -10908
rect 1556 -10961 1609 -10908
rect 1913 -10961 1966 -10908
rect 2268 -10961 2321 -10908
rect 2623 -10961 2676 -10908
rect 2980 -10961 3033 -10908
rect 3335 -10961 3388 -10908
rect 3692 -10961 3745 -10908
rect -2004 -11690 -1951 -11637
rect -1915 -11972 -1862 -11919
rect -1649 -11581 -1596 -11528
rect -1738 -11972 -1685 -11919
rect -1559 -11972 -1506 -11919
rect -1293 -11581 -1240 -11528
rect -1381 -11972 -1328 -11919
rect -1203 -11972 -1150 -11919
rect -937 -11581 -884 -11528
rect -1025 -11972 -972 -11919
rect -848 -11972 -795 -11919
rect -580 -11690 -527 -11637
rect -670 -11972 -617 -11919
rect -492 -11972 -439 -11919
rect -224 -11810 -171 -11757
rect -314 -11972 -261 -11919
rect -136 -11972 -83 -11919
rect 131 -11810 184 -11757
rect 42 -11972 95 -11919
rect 220 -11972 273 -11919
rect 487 -11810 540 -11757
rect 399 -11972 452 -11919
rect 577 -11972 630 -11919
rect 1377 -11581 1430 -11528
rect 1288 -11972 1341 -11919
rect 1468 -11972 1521 -11919
rect 1733 -11581 1786 -11528
rect 1644 -11973 1697 -11920
rect 1823 -11972 1876 -11919
rect 2089 -11581 2142 -11528
rect 2000 -11972 2053 -11919
rect 2178 -11972 2231 -11919
rect 2446 -11690 2499 -11637
rect 2357 -11972 2410 -11919
rect 2534 -11972 2587 -11919
rect 2800 -11810 2853 -11757
rect 2713 -11972 2766 -11919
rect 2890 -11972 2943 -11919
rect 3157 -11810 3210 -11757
rect 3068 -11972 3121 -11919
rect 3247 -11972 3300 -11919
rect 3513 -11810 3566 -11757
rect 3425 -11972 3478 -11919
rect 3603 -11972 3656 -11919
rect 3871 -11691 3924 -11638
rect 3781 -11972 3834 -11919
rect -2005 -12595 -1952 -12542
rect -1649 -12595 -1596 -12542
rect -1294 -12707 -1241 -12654
rect -937 -12836 -884 -12783
rect -582 -12706 -529 -12653
rect -224 -12836 -171 -12783
rect 130 -12706 183 -12653
rect 486 -12837 539 -12784
rect 1378 -12836 1431 -12783
rect 1735 -12707 1788 -12654
rect 2088 -12835 2141 -12782
rect 2445 -12706 2498 -12653
rect 2801 -12835 2854 -12782
rect 3158 -12705 3211 -12652
rect 3514 -12595 3567 -12542
rect 3871 -12595 3924 -12542
rect -2004 -13598 -1951 -13545
rect -1648 -13725 -1595 -13672
rect -581 -13598 -528 -13545
rect -1291 -13725 -1238 -13672
rect -937 -13725 -884 -13672
rect -225 -13847 -172 -13794
rect 133 -13847 186 -13794
rect 487 -13848 540 -13795
rect 1379 -13725 1432 -13672
rect 1732 -13725 1785 -13672
rect 2091 -13725 2144 -13672
rect 2446 -13598 2499 -13545
rect 2802 -13847 2855 -13794
rect 3157 -13848 3210 -13795
rect 3870 -13598 3923 -13545
rect 3512 -13847 3565 -13794
rect -2315 -14596 -2262 -14543
rect -1381 -14596 -1328 -14543
rect -1204 -14596 -1151 -14543
rect -1026 -14596 -973 -14543
rect -848 -14596 -795 -14543
rect -847 -14979 -794 -14926
rect -669 -14596 -616 -14543
rect -669 -14979 -616 -14926
rect -491 -14596 -438 -14543
rect -491 -14979 -438 -14926
rect -314 -14980 -261 -14927
rect -137 -14979 -84 -14926
rect 43 -14979 96 -14926
rect 1288 -14596 1341 -14543
rect 1289 -14980 1342 -14927
rect 1466 -14596 1519 -14543
rect 1467 -14979 1520 -14926
rect 1644 -14596 1697 -14543
rect 1644 -14979 1697 -14926
rect 1823 -14595 1876 -14542
rect 1822 -14979 1875 -14926
rect 2000 -14596 2053 -14543
rect 1999 -14979 2052 -14926
rect 2178 -14596 2231 -14543
rect 2180 -14979 2233 -14926
rect 3246 -14597 3299 -14544
rect 3424 -14596 3477 -14543
rect 3425 -14979 3478 -14926
rect 3602 -14596 3655 -14543
rect 3603 -14979 3656 -14926
rect 3781 -14596 3834 -14543
rect 3780 -14979 3833 -14926
rect 5184 -7908 5237 -7855
rect 5337 -7903 5390 -7850
rect 5185 -8687 5237 -8635
rect 11054 -8769 11107 -8716
rect 11345 -8769 11398 -8716
rect 11638 -8769 11691 -8716
rect 11932 -8769 11985 -8716
rect 12222 -8769 12275 -8716
rect 6769 -9367 6822 -9314
rect 6679 -9598 6732 -9545
rect 6947 -9368 7000 -9315
rect 7126 -9368 7179 -9315
rect 7303 -9366 7356 -9313
rect 7482 -9366 7535 -9313
rect 7659 -9368 7712 -9315
rect 7837 -9367 7890 -9314
rect 8015 -9368 8068 -9315
rect 8194 -9367 8247 -9314
rect 8371 -9367 8424 -9314
rect 8549 -9367 8602 -9314
rect 8727 -9368 8780 -9315
rect 8906 -9367 8959 -9314
rect 11144 -9427 11197 -9374
rect 11436 -9428 11489 -9375
rect 11728 -9428 11781 -9375
rect 12020 -9429 12073 -9376
rect 12312 -9428 12365 -9375
rect 5337 -9978 5390 -9925
rect 6680 -10366 6733 -10313
rect 6858 -10520 6911 -10467
rect 7214 -10519 7267 -10466
rect 7571 -10519 7624 -10466
rect 7927 -10519 7980 -10466
rect 8283 -10520 8336 -10467
rect 8638 -10519 8691 -10466
rect 9171 -10367 9224 -10314
rect 8995 -10520 9048 -10467
rect 7037 -11419 7090 -11366
rect 7393 -11419 7446 -11366
rect 7748 -11420 7801 -11367
rect 8103 -11419 8156 -11366
rect 8461 -11419 8514 -11366
rect 8817 -11419 8870 -11366
rect 11053 -11727 11106 -11674
rect 11347 -11728 11400 -11675
rect 11638 -11727 11691 -11674
rect 11931 -11727 11984 -11674
rect 12223 -11727 12276 -11674
rect 13022 -11726 13075 -11673
rect 5037 -13349 5090 -13296
rect 5534 -13349 5587 -13296
rect 5031 -13486 5084 -13433
rect 4905 -14598 4958 -14545
rect 4239 -14979 4292 -14926
rect -2447 -15874 -2394 -15821
rect -2005 -15875 -1952 -15822
rect -1915 -15986 -1862 -15933
rect -1649 -15875 -1596 -15822
rect -1738 -15986 -1685 -15933
rect -1560 -15986 -1507 -15933
rect -1293 -15875 -1240 -15822
rect -1382 -15986 -1329 -15933
rect -1204 -15986 -1151 -15933
rect -937 -15875 -884 -15822
rect -1025 -15986 -972 -15933
rect -847 -15986 -794 -15933
rect -581 -15875 -528 -15822
rect -670 -15986 -617 -15933
rect -491 -15986 -438 -15933
rect -225 -15875 -172 -15822
rect -313 -15986 -260 -15933
rect -136 -15986 -83 -15933
rect 132 -15874 185 -15821
rect 43 -15986 96 -15933
rect 221 -15986 274 -15933
rect 487 -15875 540 -15822
rect 398 -15986 451 -15933
rect 575 -15986 628 -15933
rect 843 -15875 896 -15822
rect 755 -15986 808 -15933
rect 931 -15986 984 -15933
rect 1201 -15875 1254 -15822
rect 1110 -15986 1163 -15933
rect 1289 -15986 1342 -15933
rect 1555 -15875 1608 -15822
rect 1466 -15986 1519 -15933
rect 1643 -15986 1696 -15933
rect 1910 -15875 1963 -15822
rect 1822 -15986 1875 -15933
rect 2000 -15986 2053 -15933
rect 2267 -15875 2320 -15822
rect 2179 -15986 2232 -15933
rect 2356 -15986 2409 -15933
rect 2624 -15875 2677 -15822
rect 2534 -15986 2587 -15933
rect 2712 -15986 2765 -15933
rect 2979 -15875 3032 -15822
rect 2891 -15986 2944 -15933
rect 3068 -15986 3121 -15933
rect 3335 -15875 3388 -15822
rect 3247 -15986 3300 -15933
rect 3424 -15986 3477 -15933
rect 3692 -15875 3745 -15822
rect 3603 -15986 3656 -15933
rect 3780 -15986 3833 -15933
rect 4238 -15592 4291 -15539
rect 5400 -13598 5453 -13545
rect 5142 -13847 5195 -13794
rect 5143 -14711 5196 -14658
rect -3935 -16347 -3883 -16295
rect -5682 -16939 -5629 -16886
rect -6159 -17060 -6106 -17007
rect -5859 -17060 -5806 -17007
rect -5326 -16939 -5273 -16886
rect -4970 -16939 -4917 -16886
rect -5148 -17060 -5095 -17007
rect -5504 -17171 -5451 -17118
rect -4614 -16939 -4561 -16886
rect -4258 -16939 -4205 -16886
rect -4437 -17060 -4384 -17007
rect -1917 -16595 -1864 -16542
rect -1738 -16595 -1685 -16542
rect -1561 -16594 -1508 -16541
rect -1827 -16718 -1774 -16665
rect -1381 -16596 -1328 -16543
rect -1204 -16595 -1151 -16542
rect -1026 -16595 -973 -16542
rect -1471 -16719 -1418 -16666
rect -1114 -16718 -1061 -16665
rect -759 -16717 -706 -16664
rect 220 -16595 273 -16542
rect -403 -16718 -350 -16665
rect -47 -16718 6 -16665
rect 397 -16595 450 -16542
rect 576 -16595 629 -16542
rect 755 -16595 808 -16542
rect 933 -16595 986 -16542
rect 1111 -16595 1164 -16542
rect 2356 -16595 2409 -16542
rect 309 -16719 362 -16666
rect 665 -16718 718 -16665
rect 845 -16718 898 -16665
rect 1021 -16718 1074 -16665
rect 1377 -16718 1430 -16665
rect 1735 -16718 1788 -16665
rect 2090 -16717 2143 -16664
rect 2534 -16595 2587 -16542
rect 2713 -16594 2766 -16541
rect 2891 -16595 2944 -16542
rect 3070 -16595 3123 -16542
rect 3249 -16595 3302 -16542
rect 2445 -16718 2498 -16665
rect 2801 -16718 2854 -16665
rect 3157 -16717 3210 -16664
rect 5031 -15593 5084 -15540
rect 4238 -16595 4291 -16542
rect -4792 -17171 -4739 -17118
rect -3935 -17170 -3883 -17118
rect 3514 -16719 3567 -16666
rect 3868 -16718 3921 -16665
rect 5534 -13725 5587 -13672
rect 8950 -13486 9003 -13433
rect 9305 -13486 9358 -13433
rect 8772 -13609 8825 -13556
rect 7526 -13725 7579 -13672
rect 7348 -13849 7401 -13796
rect 5833 -13975 5886 -13922
rect 6013 -13975 6066 -13922
rect 6190 -13976 6243 -13923
rect 6369 -13975 6422 -13922
rect 6547 -13976 6600 -13923
rect 6725 -13975 6778 -13922
rect 6902 -13975 6955 -13922
rect 7437 -13975 7490 -13922
rect 7882 -13726 7935 -13673
rect 8238 -13724 8291 -13671
rect 7704 -13848 7757 -13795
rect 7615 -13975 7668 -13922
rect 7793 -13976 7846 -13923
rect 8061 -13849 8114 -13796
rect 7970 -13975 8023 -13922
rect 8148 -13975 8201 -13922
rect 8415 -13849 8468 -13796
rect 8326 -13975 8379 -13922
rect 8861 -13975 8914 -13922
rect 9127 -13609 9180 -13556
rect 9038 -13975 9091 -13922
rect 9217 -13975 9270 -13922
rect 9483 -13609 9536 -13556
rect 9394 -13975 9447 -13922
rect 11442 -13725 11495 -13672
rect 11798 -13725 11851 -13672
rect 11264 -13849 11317 -13796
rect 9929 -13976 9982 -13923
rect 10108 -13975 10161 -13922
rect 10284 -13976 10337 -13923
rect 10462 -13976 10515 -13923
rect 10640 -13975 10693 -13922
rect 10819 -13976 10872 -13923
rect 11353 -13975 11406 -13922
rect 11620 -13850 11673 -13797
rect 11530 -13975 11583 -13922
rect 11709 -13975 11762 -13922
rect 12152 -13726 12205 -13673
rect 12509 -13725 12562 -13672
rect 11977 -13849 12030 -13796
rect 11886 -13976 11939 -13923
rect 12064 -13975 12117 -13922
rect 12334 -13849 12387 -13796
rect 12242 -13976 12295 -13923
rect 12420 -13975 12473 -13922
rect 5746 -14598 5799 -14545
rect 5924 -14711 5977 -14658
rect 6101 -14598 6154 -14545
rect 6279 -14711 6332 -14658
rect 6459 -14598 6512 -14545
rect 6813 -14598 6866 -14545
rect 6636 -14711 6689 -14658
rect 6991 -14711 7044 -14658
rect 6993 -14877 7046 -14824
rect 7347 -14877 7400 -14824
rect 7080 -14976 7133 -14923
rect 7260 -14977 7313 -14924
rect 7439 -14976 7492 -14923
rect 7704 -14878 7757 -14825
rect 8236 -14598 8289 -14545
rect 8060 -14874 8113 -14821
rect 8417 -14710 8470 -14657
rect 8327 -14976 8380 -14923
rect 8595 -14598 8648 -14545
rect 8504 -14859 8557 -14806
rect 8505 -14977 8558 -14924
rect 8772 -14711 8825 -14658
rect 8683 -14977 8736 -14924
rect 8950 -14599 9003 -14546
rect 9127 -14712 9180 -14659
rect 9304 -14598 9357 -14545
rect 9661 -14598 9714 -14545
rect 9483 -14711 9536 -14658
rect 9572 -14976 9625 -14923
rect 9837 -14712 9890 -14659
rect 9753 -14859 9806 -14806
rect 9750 -14976 9803 -14923
rect 10016 -14598 10069 -14545
rect 9929 -14976 9982 -14923
rect 10373 -14599 10426 -14546
rect 10196 -14711 10249 -14658
rect 10195 -14875 10248 -14822
rect 10550 -14711 10603 -14658
rect 10552 -14868 10605 -14815
rect 10729 -14598 10782 -14545
rect 10908 -14711 10961 -14658
rect 11087 -14711 11140 -14658
rect 10908 -14866 10961 -14813
rect 11440 -14709 11493 -14656
rect 10819 -14976 10872 -14923
rect 11264 -14868 11317 -14815
rect 10996 -14976 11049 -14923
rect 11175 -14976 11228 -14923
rect 5745 -15592 5798 -15539
rect 5400 -15706 5453 -15653
rect 5747 -15803 5800 -15750
rect 5923 -15705 5976 -15652
rect 5921 -16001 5974 -15948
rect 6101 -15592 6154 -15539
rect 6101 -15802 6154 -15749
rect 6279 -15705 6332 -15652
rect 6279 -16001 6332 -15948
rect 6458 -15592 6511 -15539
rect 6456 -15803 6509 -15750
rect 6635 -15705 6688 -15652
rect 6713 -15804 6766 -15751
rect 6634 -16001 6687 -15948
rect 6813 -15904 6866 -15851
rect 7169 -15803 7222 -15750
rect 7169 -15905 7222 -15852
rect 6994 -16004 7047 -15951
rect 7526 -15802 7579 -15749
rect 7526 -16006 7579 -15953
rect 7882 -15802 7935 -15749
rect 8060 -15904 8113 -15851
rect 7881 -16005 7934 -15952
rect 8237 -16005 8290 -15952
rect 8593 -15905 8646 -15852
rect 9663 -15905 9716 -15852
rect 10373 -15804 10426 -15751
rect 10194 -15905 10247 -15852
rect 10730 -15803 10783 -15750
rect 11086 -15803 11139 -15750
rect 11619 -15705 11672 -15652
rect 11084 -15905 11137 -15852
rect 11440 -15894 11493 -15841
rect 11441 -16005 11494 -15952
rect 11798 -15593 11851 -15540
rect 11797 -16005 11850 -15952
rect 11975 -15705 12028 -15652
rect 12155 -15592 12208 -15539
rect 12154 -16005 12207 -15952
rect 12332 -15705 12385 -15652
rect 12511 -15592 12564 -15539
rect 12511 -16005 12564 -15952
rect 6548 -16597 6601 -16544
rect 6726 -16597 6779 -16544
rect 6903 -16598 6956 -16545
rect 5399 -16720 5452 -16667
rect 5031 -16835 5084 -16782
rect 7970 -16598 8023 -16545
rect 8149 -16597 8202 -16544
rect 8771 -16719 8824 -16666
rect 9128 -16719 9181 -16666
rect 9484 -16719 9537 -16666
rect 8950 -16835 9003 -16782
rect 9305 -16835 9358 -16782
rect 7347 -16943 7400 -16890
rect 7704 -16943 7757 -16890
rect 8060 -16943 8113 -16890
rect 8416 -16943 8469 -16890
rect 9929 -16597 9982 -16544
rect 9838 -16719 9891 -16666
rect 10107 -16598 10160 -16545
rect 10287 -16598 10340 -16545
rect 10195 -16718 10248 -16665
rect 10550 -16718 10603 -16665
rect 10907 -16718 10960 -16665
rect 10017 -16834 10070 -16781
rect 10374 -16834 10427 -16781
rect 10731 -16832 10784 -16779
rect 11352 -16598 11405 -16545
rect 11530 -16599 11583 -16546
rect 11709 -16598 11762 -16545
rect 11263 -16943 11316 -16890
rect 11620 -16943 11673 -16890
rect 11975 -16942 12028 -16889
rect 12331 -16942 12384 -16889
rect 18337 -13496 18412 -13421
<< metal2 >>
rect 6451 2729 6515 2739
rect 17950 2729 18014 2739
rect 7145 2717 7197 2727
rect 7337 2717 7389 2727
rect 7529 2717 7581 2727
rect 7721 2717 7773 2727
rect 7912 2717 7964 2727
rect 8105 2717 8157 2727
rect 8382 2717 8434 2727
rect 16145 2717 16197 2727
rect 16337 2717 16389 2727
rect 16529 2717 16581 2727
rect 16721 2717 16773 2727
rect 16912 2717 16964 2727
rect 17105 2717 17157 2727
rect 17382 2717 17434 2727
rect 6515 2665 7145 2717
rect 7197 2665 7337 2717
rect 7389 2665 7529 2717
rect 7581 2665 7721 2717
rect 7773 2665 7912 2717
rect 7964 2665 8105 2717
rect 8157 2665 8382 2717
rect 16138 2665 16145 2717
rect 16197 2665 16337 2717
rect 16389 2665 16529 2717
rect 16581 2665 16721 2717
rect 16773 2665 16912 2717
rect 16964 2665 17105 2717
rect 17157 2665 17382 2717
rect 17434 2665 17950 2717
rect 6451 2655 6515 2665
rect 7145 2655 7197 2665
rect 7337 2655 7389 2665
rect 7529 2655 7581 2665
rect 7721 2655 7773 2665
rect 7912 2655 7964 2665
rect 8105 2655 8157 2665
rect 8382 2655 8434 2665
rect 16145 2655 16197 2665
rect 16337 2655 16389 2665
rect 16529 2655 16581 2665
rect 16721 2655 16773 2665
rect 16912 2655 16964 2665
rect 17105 2655 17157 2665
rect 17382 2655 17434 2665
rect 17950 2655 18014 2665
rect 8080 2386 11162 2450
rect 8080 2226 8144 2386
rect 8080 2152 8144 2162
rect 6704 1921 6768 1931
rect 7145 1910 7197 1919
rect 7337 1910 7389 1919
rect 7530 1910 7582 1920
rect 7722 1910 7774 1920
rect 7914 1910 7966 1920
rect 8105 1910 8157 1920
rect 8382 1910 8434 1920
rect 7138 1909 7530 1910
rect 6768 1857 7145 1909
rect 7197 1858 7337 1909
rect 6704 1847 6768 1857
rect 7145 1847 7197 1857
rect 7389 1858 7530 1909
rect 7582 1858 7722 1910
rect 7774 1858 7914 1910
rect 7966 1858 8105 1910
rect 8157 1858 8382 1910
rect 7337 1847 7389 1857
rect 7530 1848 7582 1858
rect 7722 1848 7774 1858
rect 7914 1848 7966 1858
rect 8105 1848 8157 1858
rect 8382 1848 8434 1858
rect 11098 1287 11162 2386
rect 15793 2228 15857 2238
rect 15793 2154 15857 2164
rect 17697 1922 17761 1932
rect 16145 1910 16197 1919
rect 16337 1910 16389 1919
rect 16530 1910 16582 1920
rect 16722 1910 16774 1920
rect 16914 1910 16966 1920
rect 17105 1910 17157 1920
rect 17382 1910 17434 1920
rect 16138 1909 16530 1910
rect 16138 1858 16145 1909
rect 16197 1858 16337 1909
rect 16145 1847 16197 1857
rect 16389 1858 16530 1909
rect 16582 1858 16722 1910
rect 16774 1858 16914 1910
rect 16966 1858 17105 1910
rect 17157 1858 17382 1910
rect 17434 1858 17697 1910
rect 16337 1847 16389 1857
rect 16530 1848 16582 1858
rect 16722 1848 16774 1858
rect 16914 1848 16966 1858
rect 17105 1848 17157 1858
rect 17382 1848 17434 1858
rect 17697 1848 17761 1858
rect 11098 1213 11162 1223
rect 10730 1007 10794 1017
rect 6451 929 6515 939
rect 10730 933 10794 943
rect 17950 929 18014 939
rect 7145 917 7197 927
rect 7337 917 7389 927
rect 7529 917 7581 927
rect 7721 917 7773 927
rect 7912 917 7964 927
rect 8105 917 8157 927
rect 8382 917 8434 927
rect 16145 917 16197 927
rect 16337 917 16389 927
rect 16529 917 16581 927
rect 16721 917 16773 927
rect 16912 917 16964 927
rect 17105 917 17157 927
rect 17382 917 17434 927
rect 6515 865 7145 917
rect 7197 865 7337 917
rect 7389 865 7529 917
rect 7581 865 7721 917
rect 7773 865 7912 917
rect 7964 865 8105 917
rect 8157 865 8382 917
rect 16138 865 16145 917
rect 16197 865 16337 917
rect 16389 865 16529 917
rect 16581 865 16721 917
rect 16773 865 16912 917
rect 16964 865 17105 917
rect 17157 865 17382 917
rect 17434 865 17950 917
rect 6451 855 6515 865
rect 7145 855 7197 865
rect 7337 855 7389 865
rect 7529 855 7581 865
rect 7721 855 7773 865
rect 7912 855 7964 865
rect 8105 855 8157 865
rect 8382 855 8434 865
rect 16145 855 16197 865
rect 16337 855 16389 865
rect 16529 855 16581 865
rect 16721 855 16773 865
rect 16912 855 16964 865
rect 17105 855 17157 865
rect 17382 855 17434 865
rect 17950 855 18014 865
rect 8074 426 8138 436
rect 8074 257 8138 362
rect 8625 424 8689 434
rect 8625 350 8689 360
rect 15806 426 15870 436
rect 15806 352 15870 362
rect 12512 312 12576 322
rect 8074 193 8969 257
rect 6704 121 6768 131
rect 7145 110 7197 119
rect 7337 110 7389 119
rect 7530 110 7582 120
rect 7722 110 7774 120
rect 7914 110 7966 120
rect 8105 110 8157 120
rect 8382 110 8434 120
rect 7138 109 7530 110
rect 6768 57 7145 109
rect 7197 58 7337 109
rect 6704 47 6768 57
rect 7145 47 7197 57
rect 7389 58 7530 109
rect 7582 58 7722 110
rect 7774 58 7914 110
rect 7966 58 8105 110
rect 8157 58 8382 110
rect 7337 47 7389 57
rect 7530 48 7582 58
rect 7722 48 7774 58
rect 7914 48 7966 58
rect 8105 48 8157 58
rect 8382 48 8434 58
rect 8905 -299 8969 193
rect 8905 -373 8969 -363
rect 10384 143 10448 153
rect 6451 -871 6515 -861
rect 7145 -883 7197 -873
rect 7337 -883 7389 -873
rect 7529 -883 7581 -873
rect 7721 -883 7773 -873
rect 7912 -883 7964 -873
rect 8105 -883 8157 -873
rect 8382 -883 8434 -873
rect 6515 -935 7145 -883
rect 7197 -935 7337 -883
rect 7389 -935 7529 -883
rect 7581 -935 7721 -883
rect 7773 -935 7912 -883
rect 7964 -935 8105 -883
rect 8157 -935 8382 -883
rect 6451 -945 6515 -935
rect 7145 -945 7197 -935
rect 7337 -945 7389 -935
rect 7529 -945 7581 -935
rect 7721 -945 7773 -935
rect 7912 -945 7964 -935
rect 8105 -945 8157 -935
rect 8382 -945 8434 -935
rect 10384 -1250 10448 79
rect 10732 144 10796 154
rect 10530 -1250 10594 -1240
rect 8668 -1314 10530 -1250
rect 8078 -1374 8142 -1364
rect 8078 -1546 8142 -1438
rect 8668 -1375 8732 -1314
rect 10530 -1324 10594 -1314
rect 8668 -1449 8732 -1439
rect 8078 -1610 8733 -1546
rect 6704 -1679 6768 -1669
rect 7145 -1690 7197 -1681
rect 7337 -1690 7389 -1681
rect 7530 -1690 7582 -1680
rect 7722 -1690 7774 -1680
rect 7914 -1690 7966 -1680
rect 8105 -1690 8157 -1680
rect 8382 -1690 8434 -1680
rect 7138 -1691 7530 -1690
rect 6768 -1743 7145 -1691
rect 7197 -1742 7337 -1691
rect 6704 -1753 6768 -1743
rect 7145 -1753 7197 -1743
rect 7389 -1742 7530 -1691
rect 7582 -1742 7722 -1690
rect 7774 -1742 7914 -1690
rect 7966 -1742 8105 -1690
rect 8157 -1742 8382 -1690
rect 7337 -1753 7389 -1743
rect 7530 -1752 7582 -1742
rect 7722 -1752 7774 -1742
rect 7914 -1752 7966 -1742
rect 8105 -1752 8157 -1742
rect 8382 -1752 8434 -1742
rect -5867 -1910 -5814 -1900
rect -5689 -1910 -5636 -1900
rect -5510 -1910 -5457 -1900
rect -5333 -1910 -5280 -1900
rect -5155 -1910 -5102 -1900
rect -4976 -1910 -4923 -1900
rect -4799 -1910 -4746 -1900
rect -4621 -1910 -4568 -1900
rect -4443 -1910 -4390 -1900
rect -4265 -1910 -4212 -1900
rect -4086 -1910 -4033 -1900
rect -3909 -1910 -3856 -1900
rect -1109 -1910 -1056 -1900
rect -5814 -1963 -5689 -1910
rect -5636 -1963 -5510 -1910
rect -5457 -1963 -5333 -1910
rect -5280 -1963 -5155 -1910
rect -5102 -1963 -4976 -1910
rect -4923 -1963 -4799 -1910
rect -4746 -1963 -4621 -1910
rect -4568 -1963 -4443 -1910
rect -4390 -1963 -4265 -1910
rect -4212 -1963 -4086 -1910
rect -4033 -1963 -3909 -1910
rect -3856 -1963 -1109 -1910
rect -5867 -1973 -5814 -1963
rect -5689 -1973 -5636 -1963
rect -5510 -1973 -5457 -1963
rect -5333 -1973 -5280 -1963
rect -5155 -1973 -5102 -1963
rect -4976 -1973 -4923 -1963
rect -4799 -1973 -4746 -1963
rect -4621 -1973 -4568 -1963
rect -4443 -1973 -4390 -1963
rect -4265 -1973 -4212 -1963
rect -4086 -1973 -4033 -1963
rect -3909 -1973 -3856 -1963
rect -1109 -1973 -1056 -1963
rect 8669 -2142 8733 -1610
rect 10732 -1626 10796 80
rect 12259 89 12323 99
rect 12259 15 12323 25
rect 12512 -300 12576 248
rect 17697 122 17761 132
rect 16145 110 16197 119
rect 16337 110 16389 119
rect 16530 110 16582 120
rect 16722 110 16774 120
rect 16914 110 16966 120
rect 17105 110 17157 120
rect 17382 110 17434 120
rect 16138 109 16530 110
rect 16138 58 16145 109
rect 16197 58 16337 109
rect 16145 47 16197 57
rect 16389 58 16530 109
rect 16582 58 16722 110
rect 16774 58 16914 110
rect 16966 58 17105 110
rect 17157 58 17382 110
rect 17434 58 17697 110
rect 16337 47 16389 57
rect 16530 48 16582 58
rect 16722 48 16774 58
rect 16914 48 16966 58
rect 17105 48 17157 58
rect 17382 48 17434 58
rect 17697 48 17761 58
rect 12512 -374 12576 -364
rect 13760 -363 13824 -353
rect 14520 -363 14584 -353
rect 12259 -385 12323 -375
rect 13824 -427 14520 -363
rect 13760 -437 13824 -427
rect 14520 -437 14584 -427
rect 12259 -459 12323 -449
rect 12870 -541 12934 -531
rect 12870 -615 12934 -605
rect 13186 -541 13250 -531
rect 14808 -541 14872 -531
rect 13250 -605 14808 -541
rect 13186 -615 13250 -605
rect 14808 -615 14872 -605
rect 15268 -537 15332 -527
rect 15268 -611 15332 -601
rect 17950 -871 18014 -861
rect 16145 -883 16197 -873
rect 16337 -883 16389 -873
rect 16529 -883 16581 -873
rect 16721 -883 16773 -873
rect 16912 -883 16964 -873
rect 17105 -883 17157 -873
rect 17382 -883 17434 -873
rect 12208 -906 12272 -896
rect 16138 -935 16145 -883
rect 16197 -935 16337 -883
rect 16389 -935 16529 -883
rect 16581 -935 16721 -883
rect 16773 -935 16912 -883
rect 16964 -935 17105 -883
rect 17157 -935 17382 -883
rect 17434 -935 17950 -883
rect 16145 -945 16197 -935
rect 16337 -945 16389 -935
rect 16529 -945 16581 -935
rect 16721 -945 16773 -935
rect 16912 -945 16964 -935
rect 17105 -945 17157 -935
rect 17382 -945 17434 -935
rect 17950 -945 18014 -935
rect 12208 -980 12272 -970
rect 14309 -1079 14373 -1069
rect 14309 -1153 14373 -1143
rect 12410 -1257 12474 -1247
rect 12410 -1331 12474 -1321
rect 15861 -1374 15925 -1364
rect 15054 -1438 15861 -1374
rect 13978 -1489 14042 -1479
rect 14308 -1489 14372 -1479
rect 14042 -1553 14308 -1489
rect 13978 -1563 14042 -1553
rect 14308 -1563 14372 -1553
rect 12408 -1607 12472 -1597
rect 10732 -1690 10968 -1626
rect 9435 -1986 9499 -1976
rect 9435 -2060 9499 -2050
rect 9867 -1986 9931 -1976
rect 10510 -1986 10574 -1976
rect 9931 -2050 10510 -1986
rect 9867 -2060 9931 -2050
rect 10510 -2060 10574 -2050
rect 10733 -1986 10797 -1976
rect 10733 -2060 10797 -2050
rect 9435 -2142 9499 -2132
rect 8669 -2162 9435 -2142
rect 5337 -2205 5390 -2195
rect 6680 -2199 6744 -2189
rect 5390 -2258 6680 -2205
rect 5337 -2268 5390 -2258
rect 6744 -2258 6748 -2205
rect 8668 -2206 9435 -2162
rect 9499 -2206 9504 -2142
rect 6680 -2273 6744 -2263
rect -1109 -2425 -1056 -2415
rect -752 -2425 -699 -2415
rect -1056 -2478 -752 -2425
rect -1109 -2488 -1056 -2478
rect -752 -2488 -699 -2478
rect 1919 -2426 1972 -2416
rect 2275 -2426 2328 -2416
rect 3193 -2426 3246 -2417
rect 1972 -2479 2275 -2426
rect 2328 -2427 3246 -2426
rect 2328 -2479 3193 -2427
rect 1919 -2489 1972 -2479
rect 2275 -2489 2328 -2479
rect 3193 -2490 3246 -2480
rect -6498 -2529 -6445 -2519
rect -5777 -2529 -5724 -2520
rect -6445 -2530 -5724 -2529
rect -5066 -2530 -5013 -2520
rect -4354 -2530 -4301 -2520
rect -6445 -2582 -5777 -2530
rect -6498 -2592 -6445 -2582
rect -5724 -2583 -5066 -2530
rect -5013 -2583 -4354 -2530
rect -5777 -2593 -5724 -2583
rect -5066 -2593 -5013 -2583
rect -4354 -2593 -4301 -2583
rect -2624 -2558 -2571 -2548
rect -1285 -2558 -1232 -2548
rect -930 -2558 -877 -2548
rect -2571 -2611 -1285 -2558
rect -1232 -2611 -930 -2558
rect -2624 -2621 -2571 -2611
rect -1285 -2621 -1232 -2611
rect -930 -2621 -877 -2611
rect 2097 -2554 2150 -2544
rect 2453 -2554 2506 -2544
rect 2150 -2607 2453 -2554
rect 2097 -2617 2150 -2607
rect 2453 -2617 2506 -2607
rect -5421 -2668 -5368 -2658
rect -4710 -2668 -4657 -2658
rect -3998 -2668 -3945 -2658
rect -3298 -2668 -3245 -2658
rect -5368 -2721 -4710 -2668
rect -4657 -2721 -3998 -2668
rect -3945 -2721 -3298 -2668
rect -5421 -2731 -5368 -2721
rect -4710 -2731 -4657 -2721
rect -3998 -2731 -3945 -2721
rect -3298 -2731 -3245 -2721
rect -1197 -2665 -1144 -2655
rect -1019 -2665 -966 -2655
rect -841 -2665 -788 -2655
rect -129 -2665 -76 -2655
rect 50 -2665 103 -2655
rect 227 -2665 280 -2655
rect 940 -2665 993 -2655
rect 1117 -2665 1170 -2655
rect 1295 -2665 1348 -2655
rect 2007 -2665 2060 -2655
rect 2186 -2665 2239 -2655
rect 2363 -2665 2416 -2655
rect -1144 -2718 -1019 -2665
rect -966 -2718 -841 -2665
rect -788 -2718 -129 -2665
rect -76 -2718 50 -2665
rect 103 -2718 227 -2665
rect 280 -2718 940 -2665
rect 993 -2718 1117 -2665
rect 1170 -2718 1295 -2665
rect 1348 -2718 2007 -2665
rect 2060 -2718 2186 -2665
rect 2239 -2718 2363 -2665
rect -1197 -2728 -1144 -2718
rect -1019 -2728 -966 -2718
rect -841 -2728 -788 -2718
rect -129 -2728 -76 -2718
rect 50 -2728 103 -2718
rect 227 -2728 280 -2718
rect 940 -2728 993 -2718
rect 1117 -2728 1170 -2718
rect 1295 -2728 1348 -2718
rect 2007 -2728 2060 -2718
rect 2186 -2728 2239 -2718
rect 2363 -2728 2416 -2718
rect 6451 -2671 6515 -2661
rect 7145 -2683 7197 -2673
rect 7337 -2683 7389 -2673
rect 7529 -2683 7581 -2673
rect 7721 -2683 7773 -2673
rect 7912 -2683 7964 -2673
rect 8105 -2683 8157 -2673
rect 8382 -2683 8434 -2673
rect 6515 -2735 7145 -2683
rect 7197 -2735 7337 -2683
rect 7389 -2735 7529 -2683
rect 7581 -2735 7721 -2683
rect 7773 -2735 7912 -2683
rect 7964 -2735 8105 -2683
rect 8157 -2735 8382 -2683
rect 6451 -2745 6515 -2735
rect 7145 -2745 7197 -2735
rect 7337 -2745 7389 -2735
rect 7529 -2745 7581 -2735
rect 7721 -2745 7773 -2735
rect 7912 -2745 7964 -2735
rect 8105 -2745 8157 -2735
rect 8382 -2745 8434 -2735
rect -6044 -2780 -5991 -2770
rect -5866 -2780 -5813 -2770
rect -5991 -2833 -5866 -2780
rect -6044 -2843 -5991 -2833
rect -5866 -2843 -5813 -2833
rect -3908 -2780 -3855 -2770
rect -3731 -2780 -3678 -2770
rect -3855 -2833 -3731 -2780
rect -3908 -2843 -3855 -2833
rect -3731 -2843 -3678 -2833
rect 8668 -2933 8732 -2206
rect 9435 -2216 9499 -2206
rect 9435 -2315 9499 -2305
rect 9435 -2389 9499 -2379
rect 9866 -2316 9930 -2306
rect 10904 -2316 10968 -1690
rect 9930 -2380 10968 -2316
rect 9866 -2390 9930 -2380
rect 12408 -2846 12472 -1671
rect 13976 -1827 14040 -1817
rect 13976 -1901 14040 -1891
rect 13612 -2007 13676 -1997
rect 15054 -2007 15118 -1438
rect 15861 -1448 15925 -1438
rect 17697 -1678 17761 -1668
rect 16145 -1690 16197 -1681
rect 16337 -1690 16389 -1681
rect 16530 -1690 16582 -1680
rect 16722 -1690 16774 -1680
rect 16914 -1690 16966 -1680
rect 17105 -1690 17157 -1680
rect 17382 -1690 17434 -1680
rect 16138 -1691 16530 -1690
rect 16138 -1742 16145 -1691
rect 16197 -1742 16337 -1691
rect 16145 -1753 16197 -1743
rect 16389 -1742 16530 -1691
rect 16582 -1742 16722 -1690
rect 16774 -1742 16914 -1690
rect 16966 -1742 17105 -1690
rect 17157 -1742 17382 -1690
rect 17434 -1742 17697 -1690
rect 16337 -1753 16389 -1743
rect 16530 -1752 16582 -1742
rect 16722 -1752 16774 -1742
rect 16914 -1752 16966 -1742
rect 17105 -1752 17157 -1742
rect 17382 -1752 17434 -1742
rect 17697 -1752 17761 -1742
rect 13676 -2071 15118 -2007
rect 13612 -2081 13676 -2071
rect 13610 -2318 13674 -2308
rect 13674 -2382 15113 -2318
rect 13610 -2392 13674 -2382
rect 12408 -2920 12472 -2910
rect 8075 -2997 8732 -2933
rect 8075 -3174 8139 -2997
rect 8075 -3248 8139 -3238
rect 8668 -3178 8732 -3168
rect 15049 -3172 15113 -2382
rect 17950 -2671 18014 -2661
rect 16145 -2683 16197 -2673
rect 16337 -2683 16389 -2673
rect 16529 -2683 16581 -2673
rect 16721 -2683 16773 -2673
rect 16912 -2683 16964 -2673
rect 17105 -2683 17157 -2673
rect 17382 -2683 17434 -2673
rect 16138 -2735 16145 -2683
rect 16197 -2735 16337 -2683
rect 16389 -2735 16529 -2683
rect 16581 -2735 16721 -2683
rect 16773 -2735 16912 -2683
rect 16964 -2735 17105 -2683
rect 17157 -2735 17382 -2683
rect 17434 -2735 17950 -2683
rect 16145 -2745 16197 -2735
rect 16337 -2745 16389 -2735
rect 16529 -2745 16581 -2735
rect 16721 -2745 16773 -2735
rect 16912 -2745 16964 -2735
rect 17105 -2745 17157 -2735
rect 17382 -2745 17434 -2735
rect 17950 -2745 18014 -2735
rect 15866 -3172 15930 -3162
rect 15049 -3236 15866 -3172
rect -484 -3301 -431 -3291
rect 583 -3301 636 -3291
rect 1654 -3301 1707 -3291
rect -431 -3354 583 -3301
rect 636 -3354 1654 -3301
rect -484 -3364 -431 -3354
rect 583 -3364 636 -3354
rect 1654 -3364 1707 -3354
rect -6625 -3401 -6572 -3391
rect -6134 -3401 -6081 -3391
rect -5066 -3401 -5013 -3391
rect -6572 -3454 -6134 -3401
rect -6081 -3454 -5066 -3401
rect -6625 -3464 -6572 -3454
rect -6134 -3464 -6081 -3454
rect -5066 -3464 -5013 -3454
rect -4710 -3401 -4657 -3391
rect -3642 -3401 -3589 -3391
rect -3131 -3401 -3078 -3391
rect -4657 -3454 -3642 -3401
rect -3589 -3454 -3131 -3401
rect -4710 -3464 -4657 -3454
rect -3642 -3464 -3589 -3454
rect -3131 -3464 -3078 -3454
rect -1645 -3449 -1584 -3439
rect -5777 -3516 -5724 -3506
rect -3998 -3516 -3945 -3506
rect -3298 -3516 -3245 -3506
rect -5724 -3569 -3998 -3516
rect -3945 -3569 -3298 -3516
rect -1108 -3456 -1055 -3446
rect -750 -3456 -697 -3446
rect -396 -3456 -343 -3446
rect -39 -3456 14 -3446
rect 317 -3456 370 -3446
rect -1584 -3509 -1108 -3456
rect -1055 -3509 -750 -3456
rect -697 -3509 -396 -3456
rect -343 -3509 -39 -3456
rect 14 -3509 317 -3456
rect -1645 -3520 -1584 -3510
rect -1108 -3519 -1055 -3509
rect -750 -3519 -697 -3509
rect -396 -3519 -343 -3509
rect -39 -3519 14 -3509
rect 317 -3519 370 -3509
rect 850 -3456 903 -3446
rect 1206 -3456 1259 -3446
rect 1562 -3456 1615 -3446
rect 1919 -3456 1972 -3446
rect 2275 -3456 2328 -3446
rect 3019 -3452 3080 -3442
rect 903 -3509 1206 -3456
rect 1259 -3509 1562 -3456
rect 1615 -3509 1919 -3456
rect 1972 -3509 2275 -3456
rect 2328 -3509 3019 -3456
rect 850 -3519 903 -3509
rect 1206 -3519 1259 -3509
rect 1562 -3519 1615 -3509
rect 1919 -3519 1972 -3509
rect 2275 -3519 2328 -3509
rect 6222 -3451 6286 -3441
rect 3080 -3509 6222 -3456
rect 3019 -3523 3080 -3513
rect 6286 -3509 6297 -3456
rect 6704 -3479 6768 -3469
rect 6222 -3525 6286 -3515
rect 7145 -3490 7197 -3481
rect 7337 -3490 7389 -3481
rect 7530 -3490 7582 -3480
rect 7722 -3490 7774 -3480
rect 7914 -3490 7966 -3480
rect 8105 -3490 8157 -3480
rect 8382 -3490 8434 -3480
rect 7138 -3491 7530 -3490
rect 6768 -3543 7145 -3491
rect 7197 -3542 7337 -3491
rect 6704 -3553 6768 -3543
rect 7145 -3553 7197 -3543
rect 7389 -3542 7530 -3491
rect 7582 -3542 7722 -3490
rect 7774 -3542 7914 -3490
rect 7966 -3542 8105 -3490
rect 8157 -3542 8382 -3490
rect 7337 -3553 7389 -3543
rect 7530 -3552 7582 -3542
rect 7722 -3552 7774 -3542
rect 7914 -3552 7966 -3542
rect 8105 -3552 8157 -3542
rect 8382 -3552 8434 -3542
rect -5777 -3579 -5724 -3569
rect -3998 -3579 -3945 -3569
rect -3298 -3579 -3245 -3569
rect -1286 -3571 -1233 -3561
rect -929 -3571 -876 -3561
rect -573 -3571 -520 -3561
rect -217 -3571 -164 -3561
rect -1702 -3624 -1286 -3571
rect -1233 -3624 -929 -3571
rect -876 -3624 -573 -3571
rect -520 -3624 -217 -3571
rect -6498 -3640 -6445 -3630
rect -5422 -3640 -5369 -3630
rect -4353 -3640 -4300 -3630
rect -1702 -3640 -1649 -3624
rect -1286 -3634 -1233 -3624
rect -929 -3634 -876 -3624
rect -573 -3634 -520 -3624
rect -217 -3634 -164 -3624
rect 1384 -3564 1437 -3554
rect 1741 -3564 1794 -3554
rect 2097 -3564 2150 -3554
rect 2451 -3564 2504 -3554
rect 1437 -3617 1741 -3564
rect 1794 -3617 2097 -3564
rect 2150 -3617 2451 -3564
rect 1384 -3627 1437 -3617
rect 1741 -3627 1794 -3617
rect 2097 -3627 2150 -3617
rect 2451 -3627 2504 -3617
rect -6445 -3693 -5422 -3640
rect -5369 -3693 -4353 -3640
rect -4300 -3693 -1649 -3640
rect -6498 -3703 -6445 -3693
rect -5422 -3703 -5369 -3693
rect -4353 -3703 -4300 -3693
rect -2546 -3928 -2485 -3693
rect 8668 -3795 8732 -3242
rect 12410 -3246 12474 -3236
rect 15866 -3246 15930 -3236
rect 12410 -3320 12474 -3310
rect 17697 -3478 17761 -3468
rect 16145 -3490 16197 -3481
rect 16337 -3490 16389 -3481
rect 16530 -3490 16582 -3480
rect 16722 -3490 16774 -3480
rect 16914 -3490 16966 -3480
rect 17105 -3490 17157 -3480
rect 17382 -3490 17434 -3480
rect 16138 -3491 16530 -3490
rect 16138 -3542 16145 -3491
rect 16197 -3542 16337 -3491
rect 16145 -3553 16197 -3543
rect 16389 -3542 16530 -3491
rect 16582 -3542 16722 -3490
rect 16774 -3542 16914 -3490
rect 16966 -3542 17105 -3490
rect 17157 -3542 17382 -3490
rect 17434 -3542 17697 -3490
rect 16337 -3553 16389 -3543
rect 16530 -3552 16582 -3542
rect 16722 -3552 16774 -3542
rect 16914 -3552 16966 -3542
rect 17105 -3552 17157 -3542
rect 17382 -3552 17434 -3542
rect 17697 -3552 17761 -3542
rect 13539 -3765 13603 -3755
rect 14528 -3765 14592 -3755
rect 9642 -3795 9706 -3785
rect 10932 -3795 10996 -3785
rect 8668 -3859 9642 -3795
rect 9706 -3859 10932 -3795
rect 9642 -3869 9706 -3859
rect 10932 -3869 10996 -3859
rect 11432 -3829 11496 -3819
rect 13603 -3829 14528 -3765
rect 13539 -3839 13603 -3829
rect 14528 -3839 14592 -3829
rect 11432 -3903 11496 -3893
rect -2546 -3999 -2485 -3989
rect 12704 -3943 12768 -3933
rect 12704 -4017 12768 -4007
rect 12996 -3947 13060 -3937
rect 14838 -3947 14902 -3937
rect 13060 -4011 14838 -3947
rect 12996 -4021 13060 -4011
rect 14838 -4021 14902 -4011
rect 15254 -3943 15318 -3933
rect 15254 -4017 15318 -4007
rect 9272 -4128 9336 -4118
rect -841 -4192 -788 -4182
rect -662 -4192 -609 -4182
rect -483 -4192 -430 -4182
rect -306 -4192 -253 -4182
rect 407 -4192 460 -4182
rect 583 -4192 636 -4182
rect 761 -4192 814 -4182
rect 1474 -4192 1527 -4182
rect 1652 -4192 1705 -4182
rect 1830 -4192 1883 -4182
rect 2008 -4192 2061 -4182
rect -788 -4245 -662 -4192
rect -609 -4245 -483 -4192
rect -430 -4245 -306 -4192
rect -253 -4245 407 -4192
rect 460 -4245 583 -4192
rect 636 -4245 761 -4192
rect 814 -4245 1474 -4192
rect 1527 -4245 1652 -4192
rect 1705 -4245 1830 -4192
rect 1883 -4245 2008 -4192
rect 9272 -4202 9336 -4192
rect 10032 -4128 10096 -4118
rect 13045 -4128 13109 -4118
rect 10096 -4192 13045 -4128
rect 10032 -4202 10096 -4192
rect 13045 -4202 13109 -4192
rect 13428 -4128 13492 -4118
rect 13428 -4202 13492 -4192
rect -841 -4255 -788 -4245
rect -662 -4255 -609 -4245
rect -483 -4255 -430 -4245
rect -306 -4255 -253 -4245
rect 407 -4255 460 -4245
rect 583 -4255 636 -4245
rect 761 -4255 814 -4245
rect 1474 -4255 1527 -4245
rect 1652 -4255 1705 -4245
rect 1830 -4255 1883 -4245
rect 2008 -4255 2061 -4245
rect -6498 -4271 -6445 -4261
rect -5778 -4271 -5725 -4261
rect -3998 -4271 -3945 -4261
rect -6445 -4324 -5778 -4271
rect -5725 -4324 -3998 -4271
rect 2538 -4266 2599 -4256
rect 317 -4304 370 -4294
rect 673 -4304 726 -4294
rect -6498 -4334 -6445 -4324
rect -5778 -4334 -5725 -4324
rect -3998 -4334 -3945 -4324
rect -2357 -4357 317 -4304
rect 370 -4357 673 -4304
rect 2538 -4337 2599 -4327
rect -6134 -4390 -6081 -4380
rect -5066 -4390 -5013 -4380
rect -4709 -4390 -4656 -4380
rect -3642 -4390 -3589 -4380
rect -2357 -4390 -2304 -4357
rect 317 -4367 370 -4357
rect 673 -4367 726 -4357
rect -6081 -4443 -5066 -4390
rect -5013 -4443 -4709 -4390
rect -4656 -4443 -3642 -4390
rect -3589 -4443 -2304 -4390
rect -2004 -4412 -1951 -4402
rect 495 -4412 548 -4402
rect 850 -4412 903 -4402
rect -6134 -4453 -6081 -4443
rect -5066 -4453 -5013 -4443
rect -4709 -4453 -4656 -4443
rect -3642 -4453 -3589 -4443
rect -1951 -4465 495 -4412
rect 548 -4465 850 -4412
rect -2004 -4475 -1951 -4465
rect 495 -4475 548 -4465
rect 850 -4475 903 -4465
rect 2746 -4446 2807 -4436
rect -5422 -4506 -5369 -4496
rect -4353 -4506 -4300 -4496
rect -3298 -4506 -3245 -4496
rect -2385 -4505 -2324 -4495
rect -5369 -4559 -4353 -4506
rect -4300 -4559 -3298 -4506
rect -3245 -4559 -2385 -4506
rect -5422 -4569 -5369 -4559
rect -4353 -4569 -4300 -4559
rect -3298 -4569 -3245 -4559
rect 2746 -4517 2807 -4507
rect 6451 -4471 6515 -4461
rect 17950 -4471 18014 -4461
rect 7145 -4483 7197 -4473
rect 7337 -4483 7389 -4473
rect 7529 -4483 7581 -4473
rect 7721 -4483 7773 -4473
rect 7912 -4483 7964 -4473
rect 8105 -4483 8157 -4473
rect 8382 -4483 8434 -4473
rect 16145 -4483 16197 -4473
rect 16337 -4483 16389 -4473
rect 16529 -4483 16581 -4473
rect 16721 -4483 16773 -4473
rect 16912 -4483 16964 -4473
rect 17105 -4483 17157 -4473
rect 17382 -4483 17434 -4473
rect 6515 -4535 7145 -4483
rect 7197 -4535 7337 -4483
rect 7389 -4535 7529 -4483
rect 7581 -4535 7721 -4483
rect 7773 -4535 7912 -4483
rect 7964 -4535 8105 -4483
rect 8157 -4535 8382 -4483
rect 16138 -4535 16145 -4483
rect 16197 -4535 16337 -4483
rect 16389 -4535 16529 -4483
rect 16581 -4535 16721 -4483
rect 16773 -4535 16912 -4483
rect 16964 -4535 17105 -4483
rect 17157 -4535 17382 -4483
rect 17434 -4535 17950 -4483
rect 6451 -4545 6515 -4535
rect 7145 -4545 7197 -4535
rect 7337 -4545 7389 -4535
rect 7529 -4545 7581 -4535
rect 7721 -4545 7773 -4535
rect 7912 -4545 7964 -4535
rect 8105 -4545 8157 -4535
rect 8382 -4545 8434 -4535
rect 16145 -4545 16197 -4535
rect 16337 -4545 16389 -4535
rect 16529 -4545 16581 -4535
rect 16721 -4545 16773 -4535
rect 16912 -4545 16964 -4535
rect 17105 -4545 17157 -4535
rect 17382 -4545 17434 -4535
rect 17950 -4545 18014 -4535
rect -2385 -4576 -2324 -4566
rect 3194 -4805 3246 -4795
rect 4771 -4805 4823 -4795
rect 3246 -4857 4771 -4805
rect 3194 -4867 3246 -4857
rect 4771 -4867 4823 -4857
rect 8082 -4972 8146 -4962
rect 3021 -5002 3082 -4992
rect 5037 -5006 5090 -4996
rect 4985 -5007 5037 -5006
rect 3082 -5059 5037 -5007
rect 3021 -5073 3082 -5063
rect 5037 -5069 5090 -5059
rect -2385 -5093 -2324 -5083
rect -6498 -5141 -6445 -5131
rect -5422 -5141 -5369 -5131
rect -6445 -5187 -5422 -5147
rect -6498 -5204 -6445 -5194
rect -4353 -5141 -4300 -5131
rect -5369 -5188 -4353 -5148
rect -5422 -5204 -5369 -5194
rect -1287 -5097 -1234 -5087
rect -929 -5097 -876 -5087
rect -572 -5097 -519 -5087
rect -218 -5097 -165 -5087
rect -2324 -5150 -1287 -5097
rect -1234 -5150 -929 -5097
rect -876 -5150 -572 -5097
rect -519 -5150 -218 -5097
rect 1385 -5093 1438 -5083
rect 1740 -5093 1793 -5083
rect 2096 -5093 2149 -5083
rect 2453 -5093 2506 -5083
rect -2385 -5164 -2324 -5154
rect -1287 -5160 -1234 -5150
rect -929 -5160 -876 -5150
rect -572 -5160 -519 -5150
rect -218 -5160 -165 -5150
rect 311 -5148 372 -5138
rect -4353 -5204 -4300 -5194
rect -1105 -5213 -1052 -5203
rect -751 -5213 -698 -5203
rect -396 -5213 -343 -5203
rect -41 -5213 12 -5203
rect 1438 -5146 1740 -5093
rect 1793 -5146 2096 -5093
rect 2149 -5146 2453 -5093
rect 1385 -5156 1438 -5146
rect 1740 -5156 1793 -5146
rect 2096 -5156 2149 -5146
rect 2453 -5156 2506 -5146
rect 8082 -5121 8146 -5036
rect 15802 -4976 15866 -4966
rect 15802 -5050 15866 -5040
rect 10525 -5120 10589 -5110
rect 8082 -5184 10525 -5121
rect 8082 -5185 10589 -5184
rect 10525 -5194 10589 -5185
rect 311 -5213 372 -5209
rect -6134 -5232 -6081 -5222
rect -5066 -5233 -5013 -5223
rect -6081 -5279 -5066 -5239
rect -6134 -5295 -6081 -5285
rect -3130 -5233 -3077 -5223
rect -5013 -5279 -3130 -5239
rect -5066 -5296 -5013 -5286
rect -1876 -5232 -1823 -5222
rect -3077 -5279 -1876 -5239
rect -3130 -5296 -3077 -5286
rect -1052 -5266 -751 -5213
rect -698 -5266 -396 -5213
rect -343 -5266 -41 -5213
rect 12 -5266 316 -5213
rect 369 -5219 372 -5213
rect 846 -5213 903 -5203
rect 1207 -5213 1260 -5203
rect 1563 -5213 1616 -5203
rect 1917 -5213 1970 -5203
rect 2274 -5213 2327 -5203
rect 4905 -5212 4958 -5202
rect -1876 -5295 -1823 -5285
rect -1646 -5278 -1585 -5268
rect -1105 -5276 -1052 -5266
rect -751 -5276 -698 -5266
rect -396 -5276 -343 -5266
rect -41 -5276 12 -5266
rect 316 -5276 369 -5266
rect 846 -5266 850 -5213
rect 903 -5266 1207 -5213
rect 1260 -5266 1563 -5213
rect 1616 -5266 1917 -5213
rect 1970 -5266 2274 -5213
rect 2327 -5265 4905 -5213
rect 5614 -5207 5678 -5197
rect 4958 -5265 5614 -5213
rect 2327 -5266 5614 -5265
rect -6625 -5322 -6572 -5312
rect -4710 -5322 -4657 -5312
rect -6572 -5369 -4710 -5329
rect -6625 -5385 -6572 -5375
rect -3642 -5319 -3589 -5309
rect -4657 -5369 -3642 -5329
rect -4710 -5385 -4657 -5375
rect -2624 -5324 -2571 -5314
rect -3589 -5369 -2624 -5329
rect -3642 -5382 -3589 -5372
rect -1646 -5349 -1585 -5339
rect 846 -5278 907 -5266
rect 1207 -5276 1260 -5266
rect 1563 -5276 1616 -5266
rect 1917 -5276 1970 -5266
rect 2274 -5276 2327 -5266
rect 4905 -5275 4958 -5266
rect 5678 -5266 5685 -5213
rect 5614 -5281 5678 -5271
rect 6704 -5279 6768 -5269
rect 846 -5349 907 -5339
rect 17697 -5278 17761 -5268
rect 7145 -5290 7197 -5281
rect 7337 -5290 7389 -5281
rect 7530 -5290 7582 -5280
rect 7722 -5290 7774 -5280
rect 7914 -5290 7966 -5280
rect 8105 -5290 8157 -5280
rect 8382 -5290 8434 -5280
rect 16145 -5290 16197 -5281
rect 16337 -5290 16389 -5281
rect 16530 -5290 16582 -5280
rect 16722 -5290 16774 -5280
rect 16914 -5290 16966 -5280
rect 17105 -5290 17157 -5280
rect 17382 -5290 17434 -5280
rect 7138 -5291 7530 -5290
rect 6768 -5343 7145 -5291
rect 7197 -5342 7337 -5291
rect 6704 -5353 6768 -5343
rect 7145 -5353 7197 -5343
rect 7389 -5342 7530 -5291
rect 7582 -5342 7722 -5290
rect 7774 -5342 7914 -5290
rect 7966 -5342 8105 -5290
rect 8157 -5342 8382 -5290
rect 16138 -5291 16530 -5290
rect 16138 -5342 16145 -5291
rect 7337 -5353 7389 -5343
rect 7530 -5352 7582 -5342
rect 7722 -5352 7774 -5342
rect 7914 -5352 7966 -5342
rect 8105 -5352 8157 -5342
rect 8382 -5352 8434 -5342
rect 16197 -5342 16337 -5291
rect 16145 -5353 16197 -5343
rect 16389 -5342 16530 -5291
rect 16582 -5342 16722 -5290
rect 16774 -5342 16914 -5290
rect 16966 -5342 17105 -5290
rect 17157 -5342 17382 -5290
rect 17434 -5342 17697 -5290
rect 16337 -5353 16389 -5343
rect 16530 -5352 16582 -5342
rect 16722 -5352 16774 -5342
rect 16914 -5352 16966 -5342
rect 17105 -5352 17157 -5342
rect 17382 -5352 17434 -5342
rect 17697 -5352 17761 -5342
rect -2624 -5387 -2571 -5377
rect -128 -5380 -75 -5370
rect 50 -5380 103 -5370
rect 228 -5380 281 -5370
rect 940 -5380 993 -5371
rect 1119 -5380 1172 -5370
rect 1296 -5380 1349 -5370
rect -5777 -5415 -5724 -5405
rect -3997 -5415 -3944 -5405
rect -5724 -5462 -3997 -5422
rect -5777 -5478 -5724 -5468
rect -3298 -5416 -3245 -5406
rect -3944 -5462 -3298 -5422
rect -3997 -5478 -3944 -5468
rect -75 -5433 50 -5380
rect 103 -5433 228 -5380
rect 281 -5381 1119 -5380
rect 281 -5433 940 -5381
rect -128 -5443 -75 -5433
rect 50 -5443 103 -5433
rect 228 -5443 281 -5433
rect 993 -5433 1119 -5381
rect 1172 -5433 1296 -5380
rect 940 -5444 993 -5434
rect 1119 -5443 1172 -5433
rect 1296 -5443 1349 -5433
rect -3298 -5479 -3245 -5469
rect 5337 -5527 5390 -5517
rect -5956 -6016 -5903 -6006
rect -5601 -6016 -5548 -6006
rect -5244 -6016 -5191 -6006
rect -4888 -6016 -4835 -6006
rect -4532 -6016 -4479 -6006
rect -4175 -6016 -4122 -6006
rect -3820 -6016 -3767 -6006
rect -5903 -6069 -5601 -6016
rect -5548 -6069 -5244 -6016
rect -5191 -6069 -4888 -6016
rect -4835 -6069 -4532 -6016
rect -4479 -6069 -4175 -6016
rect -4122 -6069 -3820 -6016
rect -5956 -6079 -5903 -6069
rect -5601 -6079 -5548 -6069
rect -5244 -6079 -5191 -6069
rect -4888 -6079 -4835 -6069
rect -4532 -6079 -4479 -6069
rect -4175 -6079 -4122 -6069
rect -3820 -6079 -3767 -6069
rect -2624 -6007 -2571 -5997
rect 2096 -6007 2149 -5997
rect 2452 -6007 2505 -5997
rect -2571 -6060 2096 -6007
rect 2149 -6060 2452 -6007
rect -2624 -6070 -2571 -6060
rect 2096 -6070 2149 -6060
rect 2452 -6070 2505 -6060
rect -5778 -6131 -5725 -6121
rect -5065 -6131 -5012 -6121
rect -4354 -6131 -4301 -6121
rect -3298 -6131 -3245 -6121
rect 1918 -6124 1971 -6114
rect 2275 -6124 2328 -6114
rect -2821 -6125 1918 -6124
rect -5725 -6184 -5065 -6131
rect -5012 -6184 -4354 -6131
rect -4301 -6184 -3298 -6131
rect -5778 -6194 -5725 -6184
rect -5065 -6194 -5012 -6184
rect -4354 -6194 -4301 -6184
rect -3298 -6194 -3245 -6184
rect -2856 -6177 1918 -6125
rect 1971 -6177 2275 -6124
rect -6498 -6248 -6445 -6238
rect -5421 -6248 -5368 -6238
rect -4710 -6248 -4657 -6238
rect -3998 -6247 -3945 -6237
rect -6445 -6301 -5421 -6248
rect -5368 -6301 -4710 -6248
rect -4657 -6300 -3998 -6248
rect -4657 -6301 -3945 -6300
rect -6498 -6311 -6445 -6301
rect -5421 -6311 -5368 -6301
rect -4710 -6311 -4657 -6301
rect -3998 -6310 -3945 -6301
rect -4786 -6378 -4733 -6368
rect -2856 -6401 -2803 -6177
rect 1918 -6187 1971 -6177
rect 2275 -6187 2328 -6177
rect -3874 -6408 -2803 -6401
rect -4733 -6431 -2803 -6408
rect -4786 -6454 -2803 -6431
rect -2702 -6250 -2649 -6249
rect 227 -6250 280 -6240
rect 942 -6250 995 -6240
rect -2702 -6303 227 -6250
rect 280 -6303 942 -6250
rect -4786 -6461 -3820 -6454
rect -3874 -7691 -3821 -6461
rect -2702 -6542 -2649 -6303
rect 227 -6313 280 -6303
rect 942 -6313 995 -6303
rect -1876 -6364 -1823 -6354
rect -1282 -6364 -1229 -6354
rect -1823 -6417 -1282 -6364
rect -1229 -6365 -1177 -6364
rect -928 -6365 -876 -6355
rect 2879 -6365 2931 -6355
rect -1229 -6417 -928 -6365
rect -876 -6417 2879 -6365
rect -1876 -6427 -1823 -6417
rect -1282 -6427 -1229 -6417
rect -928 -6427 -876 -6417
rect 2879 -6427 2931 -6417
rect -1110 -6479 -1057 -6469
rect -752 -6479 -699 -6469
rect -1057 -6532 -752 -6479
rect -1110 -6542 -1057 -6532
rect -752 -6542 -699 -6532
rect -3874 -7743 -3873 -7691
rect -3873 -7753 -3821 -7743
rect -3731 -6595 -2649 -6542
rect -3731 -7785 -3678 -6595
rect -753 -6598 -700 -6588
rect 4772 -6597 4825 -6587
rect -700 -6650 4772 -6598
rect -700 -6651 4825 -6650
rect -753 -6661 -700 -6651
rect 4772 -6660 4825 -6651
rect -2003 -6714 -1950 -6704
rect -1950 -6767 5237 -6714
rect -2003 -6777 -1950 -6767
rect -3545 -6806 -3484 -6796
rect -3545 -6877 -3484 -6867
rect -3679 -7837 -3678 -7785
rect -3541 -7788 -3489 -6877
rect 4770 -6891 4823 -6881
rect -3386 -6979 -3325 -6969
rect 4770 -6996 4823 -6944
rect 4906 -6889 4959 -6879
rect 4906 -6994 4959 -6942
rect -3386 -7050 -3325 -7040
rect -3731 -7847 -3679 -7837
rect -3541 -7850 -3489 -7840
rect -3382 -7933 -3329 -7050
rect 4771 -7844 4823 -6996
rect 4907 -7842 4959 -6994
rect 5038 -6887 5091 -6877
rect 5038 -7840 5091 -6940
rect 4771 -7854 4824 -7844
rect -1382 -7922 -1329 -7912
rect -1203 -7922 -1150 -7913
rect -1025 -7922 -972 -7912
rect -848 -7922 -795 -7912
rect -670 -7922 -617 -7912
rect -490 -7922 -437 -7912
rect 755 -7922 808 -7912
rect 932 -7922 985 -7912
rect 1112 -7922 1165 -7912
rect 1289 -7922 1342 -7913
rect 1467 -7922 1520 -7912
rect 1644 -7922 1697 -7912
rect 2890 -7922 2943 -7912
rect 3069 -7922 3122 -7912
rect 3247 -7922 3300 -7912
rect 3424 -7922 3477 -7912
rect 3603 -7922 3656 -7913
rect 3778 -7922 3831 -7912
rect -1329 -7923 -1025 -7922
rect -1329 -7975 -1203 -7923
rect -1382 -7985 -1329 -7975
rect -1150 -7975 -1025 -7923
rect -972 -7975 -848 -7922
rect -795 -7975 -670 -7922
rect -617 -7975 -490 -7922
rect -437 -7975 755 -7922
rect 808 -7975 932 -7922
rect 985 -7975 1112 -7922
rect 1165 -7923 1467 -7922
rect 1165 -7975 1289 -7923
rect -1203 -7986 -1150 -7976
rect -1025 -7985 -972 -7975
rect -848 -7985 -795 -7975
rect -670 -7985 -617 -7975
rect -490 -7985 -437 -7975
rect 755 -7985 808 -7975
rect 932 -7985 985 -7975
rect 1112 -7985 1165 -7975
rect 1342 -7975 1467 -7923
rect 1520 -7975 1644 -7922
rect 1697 -7975 2890 -7922
rect 2943 -7975 3069 -7922
rect 3122 -7975 3247 -7922
rect 3300 -7975 3424 -7922
rect 3477 -7923 3778 -7922
rect 3477 -7975 3603 -7923
rect 1289 -7986 1342 -7976
rect 1467 -7985 1520 -7975
rect 1644 -7985 1697 -7975
rect 2890 -7985 2943 -7975
rect 3069 -7985 3122 -7975
rect 3247 -7985 3300 -7975
rect 3424 -7985 3477 -7975
rect 3656 -7975 3778 -7923
rect 4208 -7923 4261 -7913
rect 4771 -7917 4824 -7907
rect 4906 -7852 4959 -7842
rect 4906 -7915 4959 -7905
rect 5037 -7850 5091 -7840
rect 5090 -7898 5091 -7850
rect 5184 -7855 5237 -6767
rect 5037 -7913 5090 -7903
rect 5184 -7918 5237 -7908
rect 5337 -7850 5390 -5580
rect 9262 -5687 9326 -5677
rect 6451 -6271 6515 -6261
rect 7145 -6283 7197 -6273
rect 7337 -6283 7389 -6273
rect 7529 -6283 7581 -6273
rect 7721 -6283 7773 -6273
rect 7912 -6283 7964 -6273
rect 8105 -6283 8157 -6273
rect 8382 -6283 8434 -6273
rect 6515 -6335 7145 -6283
rect 7197 -6335 7337 -6283
rect 7389 -6335 7529 -6283
rect 7581 -6335 7721 -6283
rect 7773 -6335 7912 -6283
rect 7964 -6335 8105 -6283
rect 8157 -6335 8382 -6283
rect 6451 -6345 6515 -6335
rect 7145 -6345 7197 -6335
rect 7337 -6345 7389 -6335
rect 7529 -6345 7581 -6335
rect 7721 -6345 7773 -6335
rect 7912 -6345 7964 -6335
rect 8105 -6345 8157 -6335
rect 8382 -6345 8434 -6335
rect 8738 -6543 8802 -6533
rect 8083 -6607 8738 -6543
rect 8083 -6773 8147 -6607
rect 8738 -6617 8802 -6607
rect 8083 -6847 8147 -6837
rect 8600 -6770 8664 -6760
rect 9262 -6770 9326 -5751
rect 17950 -6271 18014 -6261
rect 16145 -6283 16197 -6273
rect 16337 -6283 16389 -6273
rect 16529 -6283 16581 -6273
rect 16721 -6283 16773 -6273
rect 16912 -6283 16964 -6273
rect 17105 -6283 17157 -6273
rect 17382 -6283 17434 -6273
rect 16138 -6335 16145 -6283
rect 16197 -6335 16337 -6283
rect 16389 -6335 16529 -6283
rect 16581 -6335 16721 -6283
rect 16773 -6335 16912 -6283
rect 16964 -6335 17105 -6283
rect 17157 -6335 17382 -6283
rect 17434 -6335 17950 -6283
rect 16145 -6345 16197 -6335
rect 16337 -6345 16389 -6335
rect 16529 -6345 16581 -6335
rect 16721 -6345 16773 -6335
rect 16912 -6345 16964 -6335
rect 17105 -6345 17157 -6335
rect 17382 -6345 17434 -6335
rect 17950 -6345 18014 -6335
rect 17831 -6521 17895 -6511
rect 8664 -6834 9326 -6770
rect 15820 -6768 15884 -6758
rect 8600 -6844 8664 -6834
rect 15820 -6842 15884 -6832
rect 6704 -7079 6768 -7069
rect 17697 -7078 17761 -7068
rect 7145 -7090 7197 -7081
rect 7337 -7090 7389 -7081
rect 7530 -7090 7582 -7080
rect 7722 -7090 7774 -7080
rect 7914 -7090 7966 -7080
rect 8105 -7090 8157 -7080
rect 8382 -7090 8434 -7080
rect 16145 -7090 16197 -7081
rect 16337 -7090 16389 -7081
rect 16530 -7090 16582 -7080
rect 16722 -7090 16774 -7080
rect 16914 -7090 16966 -7080
rect 17105 -7090 17157 -7080
rect 17382 -7090 17434 -7080
rect 7138 -7091 7530 -7090
rect 6768 -7143 7145 -7091
rect 7197 -7142 7337 -7091
rect 6704 -7153 6768 -7143
rect 7145 -7153 7197 -7143
rect 7389 -7142 7530 -7091
rect 7582 -7142 7722 -7090
rect 7774 -7142 7914 -7090
rect 7966 -7142 8105 -7090
rect 8157 -7142 8382 -7090
rect 16138 -7091 16530 -7090
rect 16138 -7142 16145 -7091
rect 7337 -7153 7389 -7143
rect 7530 -7152 7582 -7142
rect 7722 -7152 7774 -7142
rect 7914 -7152 7966 -7142
rect 8105 -7152 8157 -7142
rect 8382 -7152 8434 -7142
rect 16197 -7142 16337 -7091
rect 16145 -7153 16197 -7143
rect 16389 -7142 16530 -7091
rect 16582 -7142 16722 -7090
rect 16774 -7142 16914 -7090
rect 16966 -7142 17105 -7090
rect 17157 -7142 17382 -7090
rect 17434 -7142 17697 -7090
rect 16337 -7153 16389 -7143
rect 16530 -7152 16582 -7142
rect 16722 -7152 16774 -7142
rect 16914 -7152 16966 -7142
rect 17105 -7152 17157 -7142
rect 17382 -7152 17434 -7142
rect 17697 -7152 17761 -7142
rect 5337 -7913 5390 -7903
rect 3831 -7975 4208 -7923
rect 3603 -7986 3656 -7976
rect 3778 -7976 4208 -7975
rect 3778 -7985 3831 -7976
rect 4208 -7986 4261 -7976
rect -3382 -7996 -3329 -7986
rect -1916 -8534 -1863 -8524
rect -1739 -8534 -1686 -8524
rect -1558 -8534 -1505 -8524
rect -1382 -8534 -1329 -8524
rect -1203 -8534 -1150 -8524
rect -1026 -8534 -973 -8524
rect -848 -8534 -795 -8524
rect -670 -8534 -617 -8524
rect -491 -8534 -438 -8524
rect -314 -8534 -261 -8524
rect -136 -8534 -83 -8524
rect 42 -8534 95 -8524
rect 221 -8534 274 -8524
rect 398 -8534 451 -8524
rect 577 -8534 630 -8524
rect 754 -8534 807 -8524
rect 932 -8534 985 -8524
rect 1111 -8534 1164 -8524
rect 1289 -8534 1342 -8524
rect 1466 -8534 1519 -8524
rect 1644 -8534 1697 -8524
rect 1822 -8534 1875 -8524
rect 2000 -8534 2053 -8524
rect 2178 -8534 2231 -8524
rect 2357 -8534 2410 -8524
rect 2534 -8534 2587 -8524
rect 2712 -8534 2765 -8524
rect 2890 -8534 2943 -8524
rect 3068 -8534 3121 -8524
rect 3246 -8534 3299 -8524
rect 3424 -8534 3477 -8524
rect 3602 -8534 3655 -8524
rect 3781 -8534 3834 -8524
rect -1863 -8587 -1739 -8534
rect -1686 -8587 -1558 -8534
rect -1505 -8587 -1382 -8534
rect -1329 -8587 -1203 -8534
rect -1150 -8587 -1026 -8534
rect -973 -8587 -848 -8534
rect -795 -8587 -670 -8534
rect -617 -8587 -491 -8534
rect -438 -8587 -314 -8534
rect -261 -8587 -136 -8534
rect -83 -8587 42 -8534
rect 95 -8587 221 -8534
rect 274 -8587 398 -8534
rect 451 -8587 577 -8534
rect 630 -8587 754 -8534
rect 807 -8587 932 -8534
rect 985 -8587 1111 -8534
rect 1164 -8587 1289 -8534
rect 1342 -8587 1466 -8534
rect 1519 -8587 1644 -8534
rect 1697 -8587 1822 -8534
rect 1875 -8587 2000 -8534
rect 2053 -8587 2178 -8534
rect 2231 -8587 2357 -8534
rect 2410 -8587 2534 -8534
rect 2587 -8587 2712 -8534
rect 2765 -8587 2890 -8534
rect 2943 -8587 3068 -8534
rect 3121 -8587 3246 -8534
rect 3299 -8587 3424 -8534
rect 3477 -8587 3602 -8534
rect 3655 -8587 3781 -8534
rect -1916 -8597 -1863 -8587
rect -1739 -8597 -1686 -8587
rect -1558 -8597 -1505 -8587
rect -1382 -8597 -1329 -8587
rect -1203 -8597 -1150 -8587
rect -1026 -8597 -973 -8587
rect -848 -8597 -795 -8587
rect -670 -8597 -617 -8587
rect -491 -8597 -438 -8587
rect -314 -8597 -261 -8587
rect -136 -8597 -83 -8587
rect 42 -8597 95 -8587
rect 221 -8597 274 -8587
rect 398 -8597 451 -8587
rect 577 -8597 630 -8587
rect 754 -8597 807 -8587
rect 932 -8597 985 -8587
rect 1111 -8597 1164 -8587
rect 1289 -8597 1342 -8587
rect 1466 -8597 1519 -8587
rect 1644 -8597 1697 -8587
rect 1822 -8597 1875 -8587
rect 2000 -8597 2053 -8587
rect 2178 -8597 2231 -8587
rect 2357 -8597 2410 -8587
rect 2534 -8597 2587 -8587
rect 2712 -8597 2765 -8587
rect 2890 -8597 2943 -8587
rect 3068 -8597 3121 -8587
rect 3246 -8597 3299 -8587
rect 3424 -8597 3477 -8587
rect 3602 -8597 3655 -8587
rect 3781 -8597 3834 -8587
rect 5185 -8633 5237 -8625
rect 5185 -8635 10564 -8633
rect -1826 -8653 -1773 -8643
rect -1470 -8653 -1417 -8643
rect -1115 -8653 -1062 -8643
rect -758 -8653 -705 -8643
rect -402 -8653 -349 -8643
rect -47 -8653 6 -8643
rect 310 -8653 363 -8643
rect 666 -8653 719 -8643
rect 1022 -8653 1075 -8643
rect 1377 -8653 1430 -8643
rect 1733 -8653 1786 -8643
rect 2090 -8653 2143 -8643
rect 2446 -8653 2499 -8643
rect 2802 -8653 2855 -8643
rect 3158 -8653 3211 -8643
rect 3513 -8653 3566 -8643
rect 3869 -8653 3922 -8643
rect -1773 -8706 -1470 -8653
rect -1417 -8706 -1115 -8653
rect -1062 -8706 -758 -8653
rect -705 -8706 -402 -8653
rect -349 -8706 -47 -8653
rect 6 -8706 310 -8653
rect 363 -8706 666 -8653
rect 719 -8706 1022 -8653
rect 1075 -8706 1377 -8653
rect 1430 -8706 1733 -8653
rect 1786 -8706 2090 -8653
rect 2143 -8706 2446 -8653
rect 2499 -8706 2802 -8653
rect 2855 -8706 3158 -8653
rect 3211 -8706 3513 -8653
rect 3566 -8706 3869 -8653
rect 5237 -8685 10564 -8635
rect 5185 -8697 5237 -8687
rect -1826 -8716 -1773 -8706
rect -1470 -8716 -1417 -8706
rect -1115 -8716 -1062 -8706
rect -758 -8716 -705 -8706
rect -402 -8716 -349 -8706
rect -47 -8716 6 -8706
rect 310 -8716 363 -8706
rect 666 -8716 719 -8706
rect 1022 -8716 1075 -8706
rect 1377 -8716 1430 -8706
rect 1733 -8716 1786 -8706
rect 2090 -8716 2143 -8706
rect 2446 -8716 2499 -8706
rect 2802 -8716 2855 -8706
rect 3158 -8716 3211 -8706
rect 3513 -8716 3566 -8706
rect 3869 -8716 3922 -8706
rect 10512 -8716 10564 -8685
rect 11054 -8716 11107 -8706
rect 11345 -8716 11398 -8706
rect 11638 -8716 11691 -8706
rect 11932 -8716 11985 -8706
rect 12222 -8716 12275 -8706
rect 17831 -8716 17895 -6585
rect -2447 -8767 -2394 -8757
rect -2005 -8767 -1952 -8757
rect -1648 -8767 -1595 -8757
rect -1293 -8767 -1240 -8757
rect -936 -8767 -883 -8757
rect -580 -8766 -527 -8756
rect -2394 -8820 -2005 -8767
rect -1952 -8820 -1648 -8767
rect -1595 -8820 -1293 -8767
rect -1240 -8820 -936 -8767
rect -883 -8819 -580 -8767
rect -225 -8767 -172 -8757
rect 132 -8767 185 -8758
rect 489 -8766 542 -8756
rect -527 -8819 -225 -8767
rect -883 -8820 -225 -8819
rect -172 -8768 489 -8767
rect -172 -8820 132 -8768
rect -2447 -8830 -2394 -8820
rect -2005 -8830 -1952 -8820
rect -1648 -8830 -1595 -8820
rect -1293 -8830 -1240 -8820
rect -936 -8830 -883 -8820
rect -580 -8829 -527 -8820
rect -225 -8830 -172 -8820
rect 185 -8819 489 -8768
rect 843 -8766 896 -8756
rect 542 -8819 843 -8767
rect 1201 -8767 1254 -8757
rect 1556 -8767 1609 -8757
rect 1911 -8767 1964 -8757
rect 2267 -8767 2320 -8757
rect 2624 -8767 2677 -8757
rect 2980 -8767 3033 -8757
rect 3336 -8767 3389 -8757
rect 3692 -8767 3745 -8757
rect 896 -8819 1201 -8767
rect 185 -8820 1201 -8819
rect 1254 -8820 1556 -8767
rect 1609 -8820 1911 -8767
rect 1964 -8820 2267 -8767
rect 2320 -8820 2624 -8767
rect 2677 -8820 2980 -8767
rect 3033 -8820 3336 -8767
rect 3389 -8820 3692 -8767
rect 10512 -8768 11054 -8716
rect 10584 -8769 11054 -8768
rect 11107 -8769 11345 -8716
rect 11398 -8769 11638 -8716
rect 11691 -8769 11932 -8716
rect 11985 -8769 12222 -8716
rect 12275 -8769 17895 -8716
rect 11054 -8779 11107 -8769
rect 11345 -8779 11398 -8769
rect 11638 -8779 11691 -8769
rect 11932 -8779 11985 -8769
rect 12222 -8779 12275 -8769
rect 132 -8831 185 -8821
rect 489 -8829 542 -8820
rect 843 -8829 896 -8820
rect 1201 -8830 1254 -8820
rect 1556 -8830 1609 -8820
rect 1911 -8830 1964 -8820
rect 2267 -8830 2320 -8820
rect 2624 -8830 2677 -8820
rect 2980 -8830 3033 -8820
rect 3336 -8830 3389 -8820
rect 3692 -8830 3745 -8820
rect 4771 -9314 4824 -9304
rect 6769 -9314 6822 -9304
rect 6947 -9314 7000 -9305
rect 7126 -9314 7179 -9305
rect 7303 -9313 7356 -9303
rect 4824 -9367 6769 -9314
rect 6822 -9315 7303 -9314
rect 6822 -9367 6947 -9315
rect 4771 -9377 4824 -9367
rect 6769 -9377 6822 -9367
rect 7000 -9367 7126 -9315
rect 6947 -9378 7000 -9368
rect 7179 -9366 7303 -9315
rect 7482 -9313 7535 -9303
rect 7356 -9366 7482 -9314
rect 7659 -9314 7712 -9305
rect 7837 -9314 7890 -9304
rect 8015 -9314 8068 -9305
rect 8194 -9314 8247 -9304
rect 8371 -9314 8424 -9304
rect 8549 -9314 8602 -9304
rect 8727 -9314 8780 -9305
rect 8906 -9314 8959 -9304
rect 7535 -9315 7837 -9314
rect 7535 -9366 7659 -9315
rect 7179 -9367 7659 -9366
rect 7126 -9378 7179 -9368
rect 7303 -9376 7356 -9367
rect 7482 -9376 7535 -9367
rect 7712 -9367 7837 -9315
rect 7890 -9315 8194 -9314
rect 7890 -9367 8015 -9315
rect 7659 -9378 7712 -9368
rect 7837 -9377 7890 -9367
rect 8068 -9367 8194 -9315
rect 8247 -9367 8371 -9314
rect 8424 -9367 8549 -9314
rect 8602 -9315 8906 -9314
rect 8602 -9367 8727 -9315
rect 8015 -9378 8068 -9368
rect 8194 -9377 8247 -9367
rect 8371 -9377 8424 -9367
rect 8549 -9377 8602 -9367
rect 8780 -9367 8906 -9315
rect 8727 -9378 8780 -9368
rect 8906 -9377 8959 -9367
rect 11144 -9374 11197 -9364
rect 11436 -9375 11489 -9365
rect 11728 -9375 11781 -9365
rect 12020 -9375 12073 -9366
rect 12312 -9375 12365 -9365
rect 11197 -9427 11436 -9375
rect 11144 -9428 11436 -9427
rect 11489 -9428 11728 -9375
rect 11781 -9376 12312 -9375
rect 11781 -9428 12020 -9376
rect 11144 -9437 11197 -9428
rect 11436 -9438 11489 -9428
rect 11728 -9438 11781 -9428
rect 12073 -9428 12312 -9376
rect 12020 -9439 12073 -9429
rect 12312 -9438 12365 -9428
rect -1916 -9546 -1863 -9536
rect -1738 -9546 -1685 -9536
rect -1558 -9546 -1505 -9536
rect -312 -9546 -259 -9536
rect -136 -9545 -83 -9535
rect -1863 -9599 -1738 -9546
rect -1685 -9599 -1558 -9546
rect -1505 -9599 -312 -9546
rect -259 -9598 -136 -9546
rect 42 -9546 95 -9536
rect 222 -9545 275 -9535
rect -83 -9598 42 -9546
rect -259 -9599 42 -9598
rect 95 -9598 222 -9546
rect 399 -9546 452 -9536
rect 577 -9546 630 -9536
rect 2178 -9546 2231 -9537
rect 2357 -9546 2410 -9536
rect 2534 -9546 2587 -9536
rect 2713 -9546 2766 -9536
rect 4208 -9546 4261 -9536
rect 6679 -9545 6732 -9535
rect 275 -9598 399 -9546
rect 95 -9599 399 -9598
rect 452 -9599 577 -9546
rect 630 -9547 2357 -9546
rect 630 -9599 2178 -9547
rect -1916 -9609 -1863 -9599
rect -1738 -9609 -1685 -9599
rect -1558 -9609 -1505 -9599
rect -312 -9609 -259 -9599
rect -136 -9608 -83 -9599
rect 42 -9609 95 -9599
rect 222 -9608 275 -9599
rect 399 -9609 452 -9599
rect 577 -9609 630 -9599
rect 2231 -9599 2357 -9547
rect 2410 -9599 2534 -9546
rect 2587 -9599 2713 -9546
rect 2766 -9599 4208 -9546
rect 4261 -9598 6679 -9546
rect 4261 -9599 6732 -9598
rect 2178 -9610 2231 -9600
rect 2357 -9609 2410 -9599
rect 2534 -9609 2587 -9599
rect 2713 -9609 2766 -9599
rect 4208 -9609 4261 -9599
rect 6679 -9608 6732 -9599
rect -2315 -9925 -2262 -9915
rect -1916 -9925 -1863 -9915
rect -1738 -9925 -1685 -9916
rect -1560 -9925 -1507 -9915
rect -1382 -9924 -1329 -9914
rect -2262 -9978 -1916 -9925
rect -1863 -9926 -1560 -9925
rect -1863 -9978 -1738 -9926
rect -2315 -9988 -2262 -9978
rect -1916 -9988 -1863 -9978
rect -1685 -9978 -1560 -9926
rect -1507 -9977 -1382 -9925
rect -314 -9925 -261 -9915
rect -136 -9925 -83 -9916
rect 43 -9925 96 -9915
rect 220 -9925 273 -9915
rect 398 -9925 451 -9915
rect 576 -9925 629 -9915
rect 2356 -9925 2409 -9915
rect 2534 -9925 2587 -9915
rect 2712 -9925 2765 -9916
rect 2891 -9925 2944 -9915
rect 3069 -9925 3122 -9915
rect 3246 -9925 3299 -9915
rect 5337 -9925 5390 -9915
rect -1329 -9977 -314 -9925
rect -1507 -9978 -314 -9977
rect -261 -9926 43 -9925
rect -261 -9978 -136 -9926
rect -1738 -9989 -1685 -9979
rect -1560 -9988 -1507 -9978
rect -1382 -9987 -1329 -9978
rect -314 -9988 -261 -9978
rect -83 -9978 43 -9926
rect 96 -9978 220 -9925
rect 273 -9978 398 -9925
rect 451 -9978 576 -9925
rect 629 -9978 2356 -9925
rect 2409 -9978 2534 -9925
rect 2587 -9926 2891 -9925
rect 2587 -9978 2712 -9926
rect -136 -9989 -83 -9979
rect 43 -9988 96 -9978
rect 220 -9988 273 -9978
rect 398 -9988 451 -9978
rect 576 -9988 629 -9978
rect 2356 -9988 2409 -9978
rect 2534 -9988 2587 -9978
rect 2765 -9978 2891 -9926
rect 2944 -9978 3069 -9925
rect 3122 -9978 3246 -9925
rect 3299 -9978 5337 -9925
rect 2712 -9989 2765 -9979
rect 2891 -9988 2944 -9978
rect 3069 -9988 3122 -9978
rect 3246 -9988 3299 -9978
rect 5337 -9988 5390 -9978
rect 6680 -10313 6733 -10303
rect 9171 -10313 9224 -10304
rect 6733 -10314 9224 -10313
rect 6733 -10366 9171 -10314
rect 6680 -10376 6733 -10366
rect 9171 -10377 9224 -10367
rect 6858 -10466 6911 -10457
rect 7214 -10466 7267 -10456
rect 7571 -10466 7624 -10456
rect 7927 -10466 7980 -10456
rect 8283 -10466 8336 -10457
rect 8638 -10466 8691 -10456
rect 8995 -10466 9048 -10457
rect 6858 -10467 7214 -10466
rect 6911 -10519 7214 -10467
rect 7267 -10519 7571 -10466
rect 7624 -10519 7927 -10466
rect 7980 -10467 8638 -10466
rect 7980 -10519 8283 -10467
rect 6858 -10530 6911 -10520
rect 7214 -10529 7267 -10519
rect 7571 -10529 7624 -10519
rect 7927 -10529 7980 -10519
rect 8336 -10519 8638 -10467
rect 8691 -10467 9048 -10466
rect 8691 -10519 8995 -10467
rect 8283 -10530 8336 -10520
rect 8638 -10529 8691 -10519
rect 8995 -10530 9048 -10520
rect -1827 -10908 -1774 -10898
rect -1470 -10908 -1417 -10898
rect -1114 -10908 -1061 -10898
rect -758 -10908 -705 -10898
rect -402 -10908 -349 -10898
rect -46 -10908 7 -10898
rect 309 -10908 362 -10898
rect 665 -10908 718 -10898
rect 931 -10908 984 -10898
rect 1199 -10908 1252 -10898
rect 1556 -10908 1609 -10898
rect 1913 -10908 1966 -10898
rect 2268 -10908 2321 -10898
rect 2623 -10908 2676 -10898
rect 2980 -10908 3033 -10898
rect 3335 -10908 3388 -10898
rect 3692 -10908 3745 -10898
rect -1774 -10961 -1470 -10908
rect -1417 -10961 -1114 -10908
rect -1061 -10961 -758 -10908
rect -705 -10961 -402 -10908
rect -349 -10961 -46 -10908
rect 7 -10961 309 -10908
rect 362 -10961 665 -10908
rect 718 -10961 931 -10908
rect 984 -10961 1199 -10908
rect 1252 -10961 1556 -10908
rect 1609 -10961 1913 -10908
rect 1966 -10961 2268 -10908
rect 2321 -10961 2623 -10908
rect 2676 -10961 2980 -10908
rect 3033 -10961 3335 -10908
rect 3388 -10961 3692 -10908
rect -1827 -10971 -1774 -10961
rect -1470 -10971 -1417 -10961
rect -1114 -10971 -1061 -10961
rect -758 -10971 -705 -10961
rect -402 -10971 -349 -10961
rect -46 -10971 7 -10961
rect 309 -10971 362 -10961
rect 665 -10971 718 -10961
rect 931 -10971 984 -10961
rect 1199 -10971 1252 -10961
rect 1556 -10971 1609 -10961
rect 1913 -10971 1966 -10961
rect 2268 -10971 2321 -10961
rect 2623 -10971 2676 -10961
rect 2980 -10971 3033 -10961
rect 3335 -10971 3388 -10961
rect 3692 -10971 3745 -10961
rect 7037 -11366 7090 -11356
rect 7393 -11366 7446 -11356
rect 7748 -11366 7801 -11357
rect 8103 -11366 8156 -11356
rect 8461 -11366 8514 -11356
rect 8817 -11366 8870 -11356
rect 7090 -11419 7393 -11366
rect 7446 -11367 8103 -11366
rect 7446 -11419 7748 -11367
rect 7037 -11429 7090 -11419
rect 7393 -11429 7446 -11419
rect 7801 -11419 8103 -11367
rect 8156 -11419 8461 -11366
rect 8514 -11419 8817 -11366
rect 7748 -11430 7801 -11420
rect 8103 -11429 8156 -11419
rect 8461 -11429 8514 -11419
rect 8817 -11429 8870 -11419
rect -1649 -11528 -1596 -11518
rect -1293 -11528 -1240 -11518
rect -937 -11528 -884 -11518
rect 1377 -11528 1430 -11518
rect 1733 -11528 1786 -11518
rect 2089 -11528 2142 -11518
rect -1596 -11581 -1293 -11528
rect -1240 -11581 -937 -11528
rect -884 -11581 1377 -11528
rect 1430 -11581 1733 -11528
rect 1786 -11581 2089 -11528
rect -1649 -11591 -1596 -11581
rect -1293 -11591 -1240 -11581
rect -937 -11591 -884 -11581
rect 1377 -11591 1430 -11581
rect 1733 -11591 1786 -11581
rect 2089 -11591 2142 -11581
rect -2004 -11637 -1951 -11627
rect -580 -11637 -527 -11627
rect 2446 -11637 2499 -11627
rect 3871 -11637 3924 -11628
rect -1951 -11690 -580 -11637
rect -527 -11690 2446 -11637
rect 2499 -11638 3924 -11637
rect 2499 -11690 3871 -11638
rect -2004 -11700 -1951 -11690
rect -580 -11700 -527 -11690
rect 2446 -11700 2499 -11690
rect 3871 -11701 3924 -11691
rect 11053 -11674 11106 -11664
rect 11347 -11674 11400 -11665
rect 11638 -11674 11691 -11664
rect 11931 -11674 11984 -11664
rect 12223 -11674 12276 -11664
rect 13022 -11673 13075 -11663
rect 11106 -11675 11638 -11674
rect 11106 -11727 11347 -11675
rect 11053 -11737 11106 -11727
rect 11400 -11727 11638 -11675
rect 11691 -11727 11931 -11674
rect 11984 -11727 12223 -11674
rect 12276 -11726 13022 -11674
rect 12276 -11727 13075 -11726
rect 11347 -11738 11400 -11728
rect 11638 -11737 11691 -11727
rect 11931 -11737 11984 -11727
rect 12223 -11737 12276 -11727
rect 13022 -11736 13075 -11727
rect -224 -11757 -171 -11747
rect 131 -11757 184 -11747
rect 487 -11757 540 -11747
rect 2800 -11757 2853 -11747
rect 3157 -11757 3210 -11747
rect 3513 -11757 3566 -11747
rect -171 -11810 131 -11757
rect 184 -11810 487 -11757
rect 540 -11810 2800 -11757
rect 2853 -11810 3157 -11757
rect 3210 -11810 3513 -11757
rect -224 -11820 -171 -11810
rect 131 -11820 184 -11810
rect 487 -11820 540 -11810
rect 2800 -11820 2853 -11810
rect 3157 -11820 3210 -11810
rect 3513 -11820 3566 -11810
rect -1915 -11919 -1862 -11909
rect -1738 -11919 -1685 -11909
rect -1559 -11919 -1506 -11909
rect -1381 -11919 -1328 -11909
rect -1203 -11919 -1150 -11909
rect -1025 -11919 -972 -11909
rect -848 -11919 -795 -11909
rect -670 -11919 -617 -11909
rect -492 -11919 -439 -11909
rect -314 -11919 -261 -11909
rect -136 -11919 -83 -11909
rect 42 -11919 95 -11909
rect 220 -11919 273 -11909
rect 399 -11919 452 -11909
rect 577 -11919 630 -11909
rect 1288 -11919 1341 -11909
rect 1468 -11919 1521 -11909
rect 1644 -11919 1697 -11910
rect 1823 -11919 1876 -11909
rect 2000 -11919 2053 -11909
rect 2178 -11919 2231 -11909
rect 2357 -11919 2410 -11909
rect 2534 -11919 2587 -11909
rect 2713 -11919 2766 -11909
rect 2890 -11919 2943 -11909
rect 3068 -11919 3121 -11909
rect 3247 -11919 3300 -11909
rect 3425 -11919 3478 -11909
rect 3603 -11919 3656 -11909
rect 3781 -11919 3834 -11909
rect -1862 -11972 -1738 -11919
rect -1685 -11972 -1559 -11919
rect -1506 -11972 -1381 -11919
rect -1328 -11972 -1203 -11919
rect -1150 -11972 -1025 -11919
rect -972 -11972 -848 -11919
rect -795 -11972 -670 -11919
rect -617 -11972 -492 -11919
rect -439 -11972 -314 -11919
rect -261 -11972 -136 -11919
rect -83 -11972 42 -11919
rect 95 -11972 220 -11919
rect 273 -11972 399 -11919
rect 452 -11972 577 -11919
rect 630 -11972 1288 -11919
rect 1341 -11972 1468 -11919
rect 1521 -11920 1823 -11919
rect 1521 -11972 1644 -11920
rect -1915 -11982 -1862 -11972
rect -1738 -11982 -1685 -11972
rect -1559 -11982 -1506 -11972
rect -1381 -11982 -1328 -11972
rect -1203 -11982 -1150 -11972
rect -1025 -11982 -972 -11972
rect -848 -11982 -795 -11972
rect -670 -11982 -617 -11972
rect -492 -11982 -439 -11972
rect -314 -11982 -261 -11972
rect -136 -11982 -83 -11972
rect 42 -11982 95 -11972
rect 220 -11982 273 -11972
rect 399 -11982 452 -11972
rect 577 -11982 630 -11972
rect 1288 -11982 1341 -11972
rect 1468 -11982 1521 -11972
rect 1697 -11972 1823 -11920
rect 1876 -11972 2000 -11919
rect 2053 -11972 2178 -11919
rect 2231 -11972 2357 -11919
rect 2410 -11972 2534 -11919
rect 2587 -11972 2713 -11919
rect 2766 -11972 2890 -11919
rect 2943 -11972 3068 -11919
rect 3121 -11972 3247 -11919
rect 3300 -11972 3425 -11919
rect 3478 -11972 3603 -11919
rect 3656 -11972 3781 -11919
rect 1644 -11983 1697 -11973
rect 1823 -11982 1876 -11972
rect 2000 -11982 2053 -11972
rect 2178 -11982 2231 -11972
rect 2357 -11982 2410 -11972
rect 2534 -11982 2587 -11972
rect 2713 -11982 2766 -11972
rect 2890 -11982 2943 -11972
rect 3068 -11982 3121 -11972
rect 3247 -11982 3300 -11972
rect 3425 -11982 3478 -11972
rect 3603 -11982 3656 -11972
rect 3781 -11982 3834 -11972
rect -5502 -12271 -5449 -12261
rect -5000 -12271 -4947 -12262
rect -4502 -12271 -4449 -12261
rect -5449 -12272 -4502 -12271
rect -5449 -12324 -5000 -12272
rect -5502 -12334 -5449 -12324
rect -4947 -12324 -4502 -12272
rect -2447 -12272 -2394 -12262
rect -4449 -12324 -2447 -12272
rect -5000 -12335 -4947 -12325
rect -4502 -12325 -2447 -12324
rect -4502 -12334 -4449 -12325
rect -2447 -12335 -2394 -12325
rect -5376 -12388 -5323 -12378
rect -5127 -12388 -5074 -12378
rect -4377 -12388 -4324 -12378
rect -3928 -12388 -3875 -12379
rect -5323 -12441 -5127 -12388
rect -5074 -12441 -4377 -12388
rect -4324 -12389 -3875 -12388
rect -4324 -12441 -3928 -12389
rect -5376 -12451 -5323 -12441
rect -5127 -12451 -5074 -12441
rect -4377 -12451 -4324 -12441
rect -3928 -12452 -3875 -12442
rect -6077 -12512 -6024 -12502
rect -5626 -12512 -5573 -12502
rect -4877 -12512 -4824 -12502
rect -4627 -12512 -4574 -12502
rect -6024 -12565 -5626 -12512
rect -5573 -12565 -4877 -12512
rect -4824 -12565 -4627 -12512
rect -6077 -12575 -6024 -12565
rect -5626 -12575 -5573 -12565
rect -4877 -12575 -4824 -12565
rect -4627 -12575 -4574 -12565
rect -2005 -12542 -1952 -12532
rect -1649 -12542 -1596 -12532
rect 3514 -12542 3567 -12532
rect 3871 -12542 3924 -12532
rect -1952 -12595 -1649 -12542
rect -1596 -12544 -1284 -12542
rect -1250 -12544 3514 -12542
rect -1596 -12595 3514 -12544
rect 3567 -12595 3871 -12542
rect -2005 -12605 -1952 -12595
rect -1649 -12605 -1596 -12595
rect 3514 -12605 3567 -12595
rect 3871 -12605 3924 -12595
rect -1294 -12653 -1241 -12644
rect -582 -12653 -529 -12643
rect 130 -12653 183 -12643
rect 1735 -12653 1788 -12644
rect 2445 -12653 2498 -12643
rect 3158 -12652 3211 -12642
rect -1294 -12654 -582 -12653
rect -1241 -12706 -582 -12654
rect -529 -12706 130 -12653
rect 183 -12654 2445 -12653
rect 183 -12706 1735 -12654
rect -1294 -12717 -1241 -12707
rect -582 -12716 -529 -12706
rect 130 -12716 183 -12706
rect 1788 -12706 2445 -12654
rect 2498 -12705 3158 -12653
rect 2498 -12706 3211 -12705
rect 1735 -12717 1788 -12707
rect 2445 -12716 2498 -12706
rect 3158 -12715 3211 -12706
rect -937 -12783 -884 -12773
rect -224 -12783 -171 -12773
rect 486 -12783 539 -12774
rect 1378 -12783 1431 -12773
rect 2088 -12782 2141 -12772
rect -884 -12836 -224 -12783
rect -171 -12784 1378 -12783
rect -171 -12836 486 -12784
rect -937 -12846 -884 -12836
rect -224 -12846 -171 -12836
rect 539 -12836 1378 -12784
rect 1431 -12835 2088 -12783
rect 2801 -12782 2854 -12772
rect 2141 -12835 2801 -12783
rect 1431 -12836 2854 -12835
rect 486 -12847 539 -12837
rect 1378 -12846 1431 -12836
rect 2088 -12845 2141 -12836
rect 2801 -12845 2854 -12836
rect -6223 -13062 -6170 -13052
rect -5751 -13062 -5698 -13052
rect -4752 -13062 -4699 -13052
rect -6170 -13115 -5751 -13062
rect -5698 -13115 -4752 -13062
rect -6223 -13125 -6170 -13115
rect -5751 -13125 -5698 -13115
rect -4752 -13125 -4699 -13115
rect -5251 -13189 -5198 -13179
rect -4251 -13189 -4198 -13179
rect -3788 -13189 -3735 -13179
rect -3542 -13189 -3489 -13179
rect -5198 -13242 -4251 -13189
rect -4198 -13242 -3788 -13189
rect -3735 -13242 -3542 -13189
rect -5251 -13252 -5198 -13242
rect -4251 -13252 -4198 -13242
rect -3788 -13252 -3735 -13242
rect -3542 -13252 -3489 -13242
rect 5037 -13296 5090 -13286
rect 5534 -13296 5587 -13286
rect 5090 -13349 5534 -13296
rect 5037 -13359 5090 -13349
rect 5534 -13359 5587 -13349
rect 18337 -13421 18412 -13411
rect 5031 -13433 5084 -13423
rect 8950 -13433 9003 -13423
rect 9305 -13433 9358 -13423
rect 5084 -13486 8950 -13433
rect 9003 -13486 9305 -13433
rect 9358 -13486 18337 -13433
rect 5031 -13496 5084 -13486
rect 8950 -13496 9003 -13486
rect 9305 -13496 9358 -13486
rect 18412 -13486 18422 -13433
rect 18337 -13506 18412 -13496
rect -2004 -13545 -1951 -13535
rect -581 -13545 -528 -13535
rect 2446 -13545 2499 -13535
rect 3870 -13545 3923 -13535
rect 5400 -13545 5453 -13535
rect -1951 -13598 -581 -13545
rect -528 -13598 2446 -13545
rect 2499 -13598 3870 -13545
rect 3923 -13598 5400 -13545
rect 5453 -13556 8828 -13545
rect 9127 -13556 9180 -13546
rect 9483 -13556 9536 -13546
rect 5453 -13598 8772 -13556
rect -2004 -13608 -1951 -13598
rect -581 -13608 -528 -13598
rect 2446 -13608 2499 -13598
rect 3870 -13608 3923 -13598
rect 5400 -13608 5453 -13598
rect 8825 -13609 9127 -13556
rect 9180 -13609 9483 -13556
rect 8772 -13619 8825 -13609
rect 9127 -13619 9180 -13609
rect 9483 -13619 9536 -13609
rect -1648 -13672 -1595 -13662
rect -1291 -13672 -1238 -13662
rect -937 -13672 -884 -13662
rect 1379 -13672 1432 -13662
rect 1732 -13672 1785 -13662
rect 2091 -13672 2144 -13662
rect 5534 -13672 5587 -13662
rect 7526 -13672 7579 -13662
rect 7882 -13672 7935 -13663
rect 8238 -13671 8291 -13661
rect -1595 -13725 -1291 -13672
rect -1238 -13725 -937 -13672
rect -884 -13725 1379 -13672
rect 1432 -13725 1732 -13672
rect 1785 -13725 2091 -13672
rect 2144 -13725 5323 -13672
rect -1648 -13735 -1595 -13725
rect -1291 -13735 -1238 -13725
rect -937 -13735 -884 -13725
rect 1379 -13735 1432 -13725
rect 1732 -13735 1785 -13725
rect 2091 -13735 2144 -13725
rect -6077 -13745 -6024 -13735
rect -5376 -13745 -5323 -13735
rect -5126 -13745 -5073 -13735
rect -4376 -13745 -4323 -13735
rect -6024 -13798 -5376 -13745
rect -5323 -13798 -5126 -13745
rect -5073 -13798 -4376 -13745
rect -6077 -13808 -6024 -13798
rect -5376 -13808 -5323 -13798
rect -5126 -13808 -5073 -13798
rect -4376 -13808 -4323 -13798
rect -225 -13794 -172 -13784
rect 133 -13794 186 -13784
rect 487 -13794 540 -13785
rect 2802 -13794 2855 -13784
rect 3157 -13794 3210 -13785
rect 3512 -13794 3565 -13784
rect 5142 -13794 5195 -13784
rect -6426 -13852 -6373 -13842
rect -5626 -13852 -5573 -13842
rect -4877 -13852 -4824 -13842
rect -4627 -13852 -4574 -13842
rect -3928 -13852 -3875 -13842
rect -6373 -13905 -5626 -13852
rect -5573 -13905 -4877 -13852
rect -4824 -13905 -4627 -13852
rect -4574 -13905 -3928 -13852
rect -172 -13847 133 -13794
rect 186 -13795 2802 -13794
rect 186 -13847 487 -13795
rect -225 -13857 -172 -13847
rect 133 -13857 186 -13847
rect 540 -13847 2802 -13795
rect 2855 -13795 3512 -13794
rect 2855 -13847 3157 -13795
rect 487 -13858 540 -13848
rect 2802 -13857 2855 -13847
rect 3210 -13847 3512 -13795
rect 3565 -13847 5142 -13794
rect 3157 -13858 3210 -13848
rect 3512 -13857 3565 -13847
rect 5142 -13857 5195 -13847
rect 5270 -13796 5323 -13725
rect 5587 -13725 7526 -13672
rect 7579 -13673 8238 -13672
rect 7579 -13725 7882 -13673
rect 5534 -13735 5587 -13725
rect 7526 -13735 7579 -13725
rect 7935 -13724 8238 -13673
rect 11442 -13672 11495 -13662
rect 11798 -13672 11851 -13662
rect 12152 -13672 12205 -13663
rect 12509 -13672 12562 -13662
rect 8291 -13724 11442 -13672
rect 7935 -13725 11442 -13724
rect 11495 -13725 11798 -13672
rect 11851 -13673 12509 -13672
rect 11851 -13725 12152 -13673
rect 7882 -13736 7935 -13726
rect 8238 -13734 8291 -13725
rect 11442 -13735 11495 -13725
rect 11798 -13735 11851 -13725
rect 12205 -13725 12509 -13673
rect 12152 -13736 12205 -13726
rect 12509 -13735 12562 -13725
rect 7348 -13796 7401 -13786
rect 7704 -13795 7757 -13785
rect 5270 -13849 7348 -13796
rect 7401 -13848 7704 -13796
rect 8061 -13796 8114 -13786
rect 8415 -13796 8468 -13786
rect 11264 -13796 11317 -13786
rect 11620 -13796 11673 -13787
rect 11977 -13796 12030 -13786
rect 12334 -13796 12387 -13786
rect 7757 -13848 8061 -13796
rect 7401 -13849 8061 -13848
rect 8114 -13849 8415 -13796
rect 8468 -13849 11264 -13796
rect 11317 -13797 11977 -13796
rect 11317 -13849 11620 -13797
rect 7348 -13859 7401 -13849
rect 7704 -13858 7757 -13849
rect 8061 -13859 8114 -13849
rect 8415 -13859 8468 -13849
rect 11264 -13859 11317 -13849
rect 11673 -13849 11977 -13797
rect 12030 -13849 12334 -13796
rect 11620 -13860 11673 -13850
rect 11977 -13859 12030 -13849
rect 12334 -13859 12387 -13849
rect -6426 -13915 -6373 -13905
rect -5626 -13915 -5573 -13905
rect -4877 -13915 -4824 -13905
rect -4627 -13915 -4574 -13905
rect -3928 -13915 -3875 -13905
rect 5833 -13922 5886 -13912
rect 6013 -13922 6066 -13912
rect 6190 -13922 6243 -13913
rect 6369 -13922 6422 -13912
rect 6547 -13922 6600 -13913
rect 6725 -13922 6778 -13912
rect 6902 -13922 6955 -13912
rect 7437 -13922 7490 -13912
rect 7615 -13922 7668 -13912
rect 7793 -13922 7846 -13913
rect 7970 -13922 8023 -13912
rect 8148 -13922 8201 -13912
rect 8326 -13922 8379 -13912
rect 8861 -13922 8914 -13912
rect 9038 -13922 9091 -13912
rect 9217 -13922 9270 -13912
rect 9394 -13922 9447 -13912
rect 9929 -13922 9982 -13913
rect 10108 -13922 10161 -13912
rect 10284 -13922 10337 -13913
rect 10462 -13922 10515 -13913
rect 10640 -13922 10693 -13912
rect 10819 -13922 10872 -13913
rect 11353 -13922 11406 -13912
rect 11530 -13922 11583 -13912
rect 11709 -13922 11762 -13912
rect 11886 -13922 11939 -13913
rect 12064 -13922 12117 -13912
rect 12242 -13922 12295 -13913
rect 12420 -13922 12473 -13912
rect -5730 -13957 -5677 -13947
rect -4752 -13957 -4699 -13947
rect -3788 -13957 -3735 -13947
rect -5677 -14010 -4752 -13957
rect -4699 -14010 -3788 -13957
rect 5886 -13975 6013 -13922
rect 6066 -13923 6369 -13922
rect 6066 -13975 6190 -13923
rect 5833 -13985 5886 -13975
rect 6013 -13985 6066 -13975
rect 6243 -13975 6369 -13923
rect 6422 -13923 6725 -13922
rect 6422 -13975 6547 -13923
rect 6190 -13986 6243 -13976
rect 6369 -13985 6422 -13975
rect 6600 -13975 6725 -13923
rect 6778 -13975 6902 -13922
rect 6955 -13975 7437 -13922
rect 7490 -13975 7615 -13922
rect 7668 -13923 7970 -13922
rect 7668 -13975 7793 -13923
rect 6547 -13986 6600 -13976
rect 6725 -13985 6778 -13975
rect 6902 -13985 6955 -13975
rect 7437 -13985 7490 -13975
rect 7615 -13985 7668 -13975
rect 7846 -13975 7970 -13923
rect 8023 -13975 8148 -13922
rect 8201 -13975 8326 -13922
rect 8379 -13975 8861 -13922
rect 8914 -13975 9038 -13922
rect 9091 -13975 9217 -13922
rect 9270 -13975 9394 -13922
rect 9447 -13923 10108 -13922
rect 9447 -13975 9929 -13923
rect 7793 -13986 7846 -13976
rect 7970 -13985 8023 -13975
rect 8148 -13985 8201 -13975
rect 8326 -13985 8379 -13975
rect 8861 -13985 8914 -13975
rect 9038 -13985 9091 -13975
rect 9217 -13985 9270 -13975
rect 9394 -13985 9447 -13975
rect 9982 -13975 10108 -13923
rect 10161 -13923 10640 -13922
rect 10161 -13975 10284 -13923
rect 9929 -13986 9982 -13976
rect 10108 -13985 10161 -13975
rect 10337 -13975 10462 -13923
rect 10284 -13986 10337 -13976
rect 10515 -13975 10640 -13923
rect 10693 -13923 11353 -13922
rect 10693 -13975 10819 -13923
rect 10462 -13986 10515 -13976
rect 10640 -13985 10693 -13975
rect 10872 -13975 11353 -13923
rect 11406 -13975 11530 -13922
rect 11583 -13975 11709 -13922
rect 11762 -13923 12064 -13922
rect 11762 -13975 11886 -13923
rect 10819 -13986 10872 -13976
rect 11353 -13985 11406 -13975
rect 11530 -13985 11583 -13975
rect 11709 -13985 11762 -13975
rect 11939 -13975 12064 -13923
rect 12117 -13923 12420 -13922
rect 12117 -13975 12242 -13923
rect 11886 -13986 11939 -13976
rect 12064 -13985 12117 -13975
rect 12295 -13975 12420 -13923
rect 12242 -13986 12295 -13976
rect 12420 -13985 12473 -13975
rect -5730 -14020 -5677 -14010
rect -4752 -14020 -4699 -14010
rect -3788 -14020 -3735 -14010
rect -6223 -14055 -6170 -14045
rect -5250 -14055 -5197 -14045
rect -4250 -14055 -4197 -14045
rect -3382 -14055 -3329 -14045
rect -6170 -14108 -5250 -14055
rect -5197 -14108 -4250 -14055
rect -4197 -14108 -3382 -14055
rect -6223 -14118 -6170 -14108
rect -5250 -14118 -5197 -14108
rect -4250 -14118 -4197 -14108
rect -3382 -14118 -3329 -14108
rect -2315 -14543 -2262 -14533
rect -1381 -14543 -1328 -14533
rect -1204 -14543 -1151 -14533
rect -1026 -14543 -973 -14533
rect -848 -14543 -795 -14533
rect -669 -14543 -616 -14533
rect -491 -14543 -438 -14533
rect 1288 -14543 1341 -14533
rect 1466 -14543 1519 -14533
rect 1644 -14543 1697 -14533
rect 1823 -14542 1876 -14532
rect -2262 -14596 -1381 -14543
rect -1328 -14596 -1204 -14543
rect -1151 -14596 -1026 -14543
rect -973 -14596 -848 -14543
rect -795 -14596 -669 -14543
rect -616 -14596 -491 -14543
rect -438 -14596 1288 -14543
rect 1341 -14596 1466 -14543
rect 1519 -14596 1644 -14543
rect 1697 -14595 1823 -14543
rect 2000 -14543 2053 -14533
rect 2178 -14543 2231 -14533
rect 3246 -14543 3299 -14534
rect 3424 -14543 3477 -14533
rect 3602 -14543 3655 -14533
rect 3781 -14543 3834 -14533
rect 1876 -14595 2000 -14543
rect 1697 -14596 2000 -14595
rect 2053 -14596 2178 -14543
rect 2231 -14544 3424 -14543
rect 2231 -14596 3246 -14544
rect -2315 -14606 -2262 -14596
rect -1381 -14606 -1328 -14596
rect -1204 -14606 -1151 -14596
rect -1026 -14606 -973 -14596
rect -848 -14606 -795 -14596
rect -669 -14606 -616 -14596
rect -491 -14606 -438 -14596
rect 1288 -14606 1341 -14596
rect 1466 -14606 1519 -14596
rect 1644 -14606 1697 -14596
rect 1823 -14605 1876 -14596
rect 2000 -14606 2053 -14596
rect 2178 -14606 2231 -14596
rect 3299 -14596 3424 -14544
rect 3477 -14596 3602 -14543
rect 3655 -14596 3781 -14543
rect 3246 -14607 3299 -14597
rect 3424 -14606 3477 -14596
rect 3602 -14606 3655 -14596
rect 3781 -14606 3834 -14596
rect 4905 -14545 4958 -14535
rect 5746 -14545 5799 -14535
rect 6101 -14545 6154 -14535
rect 6459 -14545 6512 -14535
rect 6813 -14545 6866 -14535
rect 8236 -14545 8289 -14535
rect 8595 -14545 8648 -14535
rect 8950 -14545 9003 -14536
rect 9304 -14545 9357 -14535
rect 9661 -14545 9714 -14535
rect 10016 -14545 10069 -14535
rect 10373 -14545 10426 -14536
rect 10729 -14545 10782 -14535
rect 4958 -14598 5746 -14545
rect 5799 -14598 6101 -14545
rect 6154 -14598 6459 -14545
rect 6512 -14598 6813 -14545
rect 6866 -14598 8236 -14545
rect 8289 -14598 8595 -14545
rect 8648 -14546 9304 -14545
rect 8648 -14598 8950 -14546
rect 4905 -14608 4958 -14598
rect 5746 -14608 5799 -14598
rect 6101 -14608 6154 -14598
rect 6459 -14608 6512 -14598
rect 6813 -14608 6866 -14598
rect 8236 -14608 8289 -14598
rect 8595 -14608 8648 -14598
rect 9003 -14598 9304 -14546
rect 9357 -14598 9661 -14545
rect 9714 -14598 10016 -14545
rect 10069 -14546 10729 -14545
rect 10069 -14598 10373 -14546
rect 8950 -14609 9003 -14599
rect 9304 -14608 9357 -14598
rect 9661 -14608 9714 -14598
rect 10016 -14608 10069 -14598
rect 10426 -14598 10729 -14546
rect 10373 -14609 10426 -14599
rect 10729 -14608 10782 -14598
rect 5143 -14658 5196 -14648
rect 5924 -14658 5977 -14648
rect 6279 -14658 6332 -14648
rect 6636 -14658 6689 -14648
rect 6991 -14658 7044 -14648
rect 8417 -14657 8470 -14647
rect 5196 -14711 5924 -14658
rect 5977 -14711 6279 -14658
rect 6332 -14711 6636 -14658
rect 6689 -14711 6991 -14658
rect 7044 -14710 8417 -14658
rect 8772 -14658 8825 -14648
rect 9127 -14658 9180 -14649
rect 9483 -14658 9536 -14648
rect 9837 -14658 9890 -14649
rect 10196 -14658 10249 -14648
rect 10550 -14658 10603 -14648
rect 10908 -14658 10961 -14648
rect 8470 -14710 8772 -14658
rect 7044 -14711 8772 -14710
rect 8825 -14659 9483 -14658
rect 8825 -14711 9127 -14659
rect 5143 -14721 5196 -14711
rect 5924 -14721 5977 -14711
rect 6279 -14721 6332 -14711
rect 6636 -14721 6689 -14711
rect 6991 -14721 7044 -14711
rect 8417 -14720 8470 -14711
rect 8772 -14721 8825 -14711
rect 9180 -14711 9483 -14659
rect 9536 -14659 10196 -14658
rect 9536 -14711 9837 -14659
rect 9127 -14722 9180 -14712
rect 9483 -14721 9536 -14711
rect 9890 -14711 10196 -14659
rect 10249 -14711 10550 -14658
rect 10603 -14711 10908 -14658
rect 9837 -14722 9890 -14712
rect 10196 -14721 10249 -14711
rect 10550 -14721 10603 -14711
rect 10908 -14721 10961 -14711
rect 11087 -14656 11140 -14648
rect 11440 -14656 11493 -14646
rect 11087 -14658 11440 -14656
rect 11140 -14708 11440 -14658
rect 11140 -14709 11192 -14708
rect 11087 -14721 11140 -14711
rect 11440 -14719 11493 -14709
rect -6159 -14795 -6106 -14785
rect -5860 -14795 -5807 -14785
rect -5147 -14795 -5094 -14785
rect -4436 -14795 -4383 -14785
rect -6106 -14848 -5860 -14795
rect -5807 -14848 -5147 -14795
rect -5094 -14848 -4436 -14795
rect 8504 -14806 8557 -14796
rect -6159 -14858 -6106 -14848
rect -5860 -14858 -5807 -14848
rect -5147 -14858 -5094 -14848
rect -4436 -14858 -4383 -14848
rect 6993 -14824 7046 -14814
rect 7347 -14824 7400 -14814
rect 7704 -14824 7757 -14815
rect 7046 -14877 7347 -14824
rect 7400 -14825 7757 -14824
rect 7400 -14877 7704 -14825
rect 6993 -14887 7046 -14877
rect 7347 -14887 7400 -14877
rect 7704 -14888 7757 -14878
rect 8060 -14821 8113 -14811
rect 8113 -14859 8504 -14821
rect 9753 -14806 9806 -14796
rect 8557 -14859 9753 -14821
rect 10195 -14821 10248 -14812
rect 9806 -14822 10248 -14821
rect 9806 -14859 10195 -14822
rect 8113 -14874 10195 -14859
rect 8060 -14884 8113 -14874
rect 10195 -14885 10248 -14875
rect 10552 -14814 10605 -14805
rect 10908 -14813 10961 -14803
rect 10552 -14815 10908 -14814
rect 10605 -14866 10908 -14815
rect 10961 -14814 11013 -14813
rect 11264 -14814 11317 -14805
rect 10961 -14815 11317 -14814
rect 10961 -14866 11264 -14815
rect 10552 -14878 10605 -14868
rect 10908 -14876 10961 -14866
rect 11264 -14878 11317 -14868
rect -5504 -14901 -5451 -14891
rect -4791 -14901 -4738 -14891
rect -3936 -14901 -3883 -14891
rect -5451 -14954 -4791 -14901
rect -4738 -14954 -3936 -14901
rect -5504 -14964 -5451 -14954
rect -4791 -14964 -4738 -14954
rect -3936 -14964 -3883 -14954
rect -847 -14926 -794 -14916
rect -669 -14926 -616 -14916
rect -491 -14926 -438 -14916
rect -314 -14926 -261 -14917
rect -137 -14926 -84 -14916
rect 43 -14926 96 -14916
rect 1289 -14926 1342 -14917
rect 1467 -14926 1520 -14916
rect 1644 -14926 1697 -14916
rect 1822 -14926 1875 -14916
rect 1999 -14926 2052 -14916
rect 2180 -14926 2233 -14916
rect 3425 -14926 3478 -14916
rect 3603 -14926 3656 -14916
rect 3780 -14926 3833 -14916
rect 4239 -14926 4292 -14916
rect -794 -14979 -669 -14926
rect -616 -14979 -491 -14926
rect -438 -14927 -137 -14926
rect -438 -14979 -314 -14927
rect -847 -14989 -794 -14979
rect -669 -14989 -616 -14979
rect -491 -14989 -438 -14979
rect -261 -14979 -137 -14927
rect -84 -14979 43 -14926
rect 96 -14927 1467 -14926
rect 96 -14979 1289 -14927
rect -314 -14990 -261 -14980
rect -137 -14989 -84 -14979
rect 43 -14989 96 -14979
rect 1342 -14979 1467 -14927
rect 1520 -14979 1644 -14926
rect 1697 -14979 1822 -14926
rect 1875 -14979 1999 -14926
rect 2052 -14979 2180 -14926
rect 2233 -14979 3425 -14926
rect 3478 -14979 3603 -14926
rect 3656 -14979 3780 -14926
rect 3833 -14979 4239 -14926
rect 1289 -14990 1342 -14980
rect 1467 -14989 1520 -14979
rect 1644 -14989 1697 -14979
rect 1822 -14989 1875 -14979
rect 1999 -14989 2052 -14979
rect 2180 -14989 2233 -14979
rect 3425 -14989 3478 -14979
rect 3603 -14989 3656 -14979
rect 3780 -14989 3833 -14979
rect 4239 -14989 4292 -14979
rect 7080 -14923 7133 -14913
rect 7260 -14923 7313 -14914
rect 7439 -14923 7492 -14913
rect 8327 -14923 8380 -14913
rect 8505 -14923 8558 -14914
rect 8683 -14923 8736 -14914
rect 9572 -14923 9625 -14913
rect 9750 -14923 9803 -14913
rect 9929 -14923 9982 -14913
rect 10819 -14923 10872 -14913
rect 10996 -14923 11049 -14913
rect 11175 -14923 11228 -14913
rect 7133 -14924 7439 -14923
rect 7133 -14976 7260 -14924
rect 7080 -14986 7133 -14976
rect 7313 -14976 7439 -14924
rect 7492 -14976 8327 -14923
rect 8380 -14924 9572 -14923
rect 8380 -14976 8505 -14924
rect 7260 -14987 7313 -14977
rect 7439 -14986 7492 -14976
rect 8327 -14986 8380 -14976
rect 8558 -14976 8683 -14924
rect 8505 -14987 8558 -14977
rect 8736 -14976 9572 -14924
rect 9625 -14976 9750 -14923
rect 9803 -14976 9929 -14923
rect 9982 -14976 10819 -14923
rect 10872 -14976 10996 -14923
rect 11049 -14976 11175 -14923
rect 8683 -14987 8736 -14977
rect 9572 -14986 9625 -14976
rect 9750 -14986 9803 -14976
rect 9929 -14986 9982 -14976
rect 10819 -14986 10872 -14976
rect 10996 -14986 11049 -14976
rect 11175 -14986 11228 -14976
rect -6159 -15481 -6106 -15472
rect -5504 -15481 -5451 -15471
rect -4792 -15481 -4739 -15471
rect -6159 -15482 -5504 -15481
rect -6106 -15534 -5504 -15482
rect -5451 -15534 -4792 -15481
rect -6159 -15545 -6106 -15535
rect -5504 -15544 -5451 -15534
rect -4792 -15544 -4739 -15534
rect 4238 -15539 4291 -15529
rect 5031 -15539 5084 -15530
rect 5745 -15539 5798 -15529
rect 6101 -15539 6154 -15529
rect 6458 -15539 6511 -15529
rect 11798 -15539 11851 -15530
rect 12155 -15539 12208 -15529
rect 12511 -15539 12564 -15529
rect -5860 -15588 -5807 -15578
rect -5148 -15589 -5095 -15579
rect -4435 -15589 -4383 -15579
rect -3935 -15589 -3883 -15579
rect -5807 -15641 -5148 -15589
rect -5860 -15651 -5807 -15641
rect -5095 -15641 -4435 -15589
rect -4383 -15641 -3935 -15589
rect 4291 -15540 5745 -15539
rect 4291 -15592 5031 -15540
rect 4238 -15602 4291 -15592
rect 5084 -15592 5745 -15540
rect 5798 -15592 6101 -15539
rect 6154 -15592 6458 -15539
rect 6511 -15540 12155 -15539
rect 6511 -15592 11798 -15540
rect 5031 -15603 5084 -15593
rect 5745 -15602 5798 -15592
rect 6101 -15602 6154 -15592
rect 6458 -15602 6511 -15592
rect 11851 -15592 12155 -15540
rect 12208 -15592 12511 -15539
rect 11798 -15603 11851 -15593
rect 12155 -15602 12208 -15592
rect 12511 -15602 12564 -15592
rect -5148 -15652 -5095 -15642
rect -4435 -15651 -4383 -15641
rect -3935 -15651 -3883 -15641
rect 5400 -15652 5453 -15643
rect 5923 -15652 5976 -15642
rect 6279 -15652 6332 -15642
rect 6635 -15652 6688 -15642
rect 11619 -15652 11672 -15642
rect 11975 -15652 12028 -15642
rect 12332 -15652 12385 -15642
rect 5400 -15653 5923 -15652
rect 5453 -15705 5923 -15653
rect 5976 -15705 6279 -15652
rect 6332 -15705 6635 -15652
rect 6688 -15705 11619 -15652
rect 11672 -15705 11975 -15652
rect 12028 -15705 12332 -15652
rect 5400 -15716 5453 -15706
rect 5923 -15715 5976 -15705
rect 6279 -15715 6332 -15705
rect 6635 -15715 6688 -15705
rect 11619 -15715 11672 -15705
rect 11975 -15715 12028 -15705
rect 12332 -15715 12385 -15705
rect 5747 -15750 5800 -15740
rect 6101 -15749 6154 -15739
rect 5800 -15802 6101 -15750
rect 6456 -15750 6509 -15740
rect 6713 -15750 6766 -15741
rect 7169 -15750 7222 -15740
rect 7526 -15749 7579 -15739
rect 6154 -15802 6456 -15750
rect 5800 -15803 6456 -15802
rect 6509 -15751 7169 -15750
rect 6509 -15803 6713 -15751
rect -2447 -15821 -2394 -15811
rect -2005 -15821 -1952 -15812
rect -2394 -15822 -1952 -15821
rect -1649 -15822 -1596 -15812
rect -1293 -15822 -1240 -15812
rect -937 -15822 -884 -15812
rect -581 -15822 -528 -15812
rect -225 -15822 -172 -15812
rect 132 -15821 185 -15811
rect -2394 -15874 -2005 -15822
rect -2447 -15884 -2394 -15874
rect -1952 -15875 -1649 -15822
rect -1596 -15875 -1293 -15822
rect -1240 -15875 -937 -15822
rect -884 -15875 -581 -15822
rect -528 -15875 -225 -15822
rect -172 -15874 132 -15822
rect 487 -15822 540 -15812
rect 843 -15822 896 -15812
rect 1201 -15822 1254 -15812
rect 1555 -15822 1608 -15812
rect 1910 -15822 1963 -15812
rect 2267 -15822 2320 -15812
rect 2624 -15822 2677 -15812
rect 2979 -15822 3032 -15812
rect 3335 -15822 3388 -15812
rect 3692 -15822 3745 -15812
rect 5747 -15813 5800 -15803
rect 6101 -15812 6154 -15803
rect 6456 -15813 6509 -15803
rect 6766 -15803 7169 -15751
rect 7222 -15802 7526 -15750
rect 7882 -15749 7935 -15739
rect 7579 -15802 7882 -15750
rect 10373 -15750 10426 -15741
rect 10730 -15750 10783 -15740
rect 11086 -15750 11139 -15740
rect 7935 -15751 10730 -15750
rect 7935 -15802 10373 -15751
rect 7222 -15803 10373 -15802
rect 6713 -15814 6766 -15804
rect 7169 -15813 7222 -15803
rect 7526 -15812 7579 -15803
rect 7882 -15812 7935 -15803
rect 10426 -15803 10730 -15751
rect 10783 -15803 11086 -15750
rect 10373 -15814 10426 -15804
rect 10730 -15813 10783 -15803
rect 11086 -15813 11139 -15803
rect 185 -15874 487 -15822
rect -172 -15875 487 -15874
rect 540 -15875 843 -15822
rect 896 -15875 1201 -15822
rect 1254 -15875 1555 -15822
rect 1608 -15875 1910 -15822
rect 1963 -15875 2267 -15822
rect 2320 -15875 2624 -15822
rect 2677 -15875 2979 -15822
rect 3032 -15875 3335 -15822
rect 3388 -15875 3692 -15822
rect 11440 -15841 11493 -15831
rect -2005 -15885 -1952 -15875
rect -1649 -15885 -1596 -15875
rect -1293 -15885 -1240 -15875
rect -937 -15885 -884 -15875
rect -581 -15885 -528 -15875
rect -225 -15885 -172 -15875
rect 132 -15884 185 -15875
rect 487 -15885 540 -15875
rect 843 -15885 896 -15875
rect 1201 -15885 1254 -15875
rect 1555 -15885 1608 -15875
rect 1910 -15885 1963 -15875
rect 2267 -15885 2320 -15875
rect 2624 -15885 2677 -15875
rect 2979 -15885 3032 -15875
rect 3335 -15885 3388 -15875
rect 3692 -15885 3745 -15875
rect 6813 -15851 6866 -15841
rect 7169 -15851 7222 -15842
rect 8060 -15851 8113 -15841
rect 8593 -15851 8646 -15842
rect 9663 -15851 9716 -15842
rect 10194 -15851 10247 -15842
rect 11084 -15851 11137 -15842
rect 6866 -15852 8060 -15851
rect 6866 -15904 7169 -15852
rect 6813 -15914 6866 -15904
rect 7222 -15904 8060 -15852
rect 8113 -15852 11440 -15851
rect 8113 -15904 8593 -15852
rect 7169 -15915 7222 -15905
rect 8060 -15914 8113 -15904
rect 8646 -15904 9663 -15852
rect 8593 -15915 8646 -15905
rect 9716 -15904 10194 -15852
rect 9663 -15915 9716 -15905
rect 10247 -15904 11084 -15852
rect 10194 -15915 10247 -15905
rect 11137 -15894 11440 -15852
rect 11137 -15904 11493 -15894
rect 11084 -15915 11137 -15905
rect -1915 -15933 -1862 -15923
rect -1738 -15933 -1685 -15923
rect -1560 -15933 -1507 -15923
rect -1382 -15933 -1329 -15923
rect -1204 -15933 -1151 -15923
rect -1025 -15933 -972 -15923
rect -847 -15933 -794 -15923
rect -670 -15933 -617 -15923
rect -491 -15933 -438 -15923
rect -313 -15933 -260 -15923
rect -136 -15933 -83 -15923
rect 43 -15933 96 -15923
rect 221 -15933 274 -15923
rect 398 -15933 451 -15923
rect 575 -15933 628 -15923
rect 755 -15933 808 -15923
rect 931 -15933 984 -15923
rect 1110 -15933 1163 -15923
rect 1289 -15933 1342 -15923
rect 1466 -15933 1519 -15923
rect 1643 -15933 1696 -15923
rect 1822 -15933 1875 -15923
rect 2000 -15933 2053 -15923
rect 2179 -15933 2232 -15923
rect 2356 -15933 2409 -15923
rect 2534 -15933 2587 -15923
rect 2712 -15933 2765 -15923
rect 2891 -15933 2944 -15923
rect 3068 -15933 3121 -15923
rect 3247 -15933 3300 -15923
rect 3424 -15933 3477 -15923
rect 3603 -15933 3656 -15923
rect 3780 -15933 3833 -15923
rect -1862 -15986 -1738 -15933
rect -1685 -15986 -1560 -15933
rect -1507 -15986 -1382 -15933
rect -1329 -15986 -1204 -15933
rect -1151 -15986 -1025 -15933
rect -972 -15986 -847 -15933
rect -794 -15986 -670 -15933
rect -617 -15986 -491 -15933
rect -438 -15986 -313 -15933
rect -260 -15986 -136 -15933
rect -83 -15986 43 -15933
rect 96 -15986 221 -15933
rect 274 -15986 398 -15933
rect 451 -15986 575 -15933
rect 628 -15986 755 -15933
rect 808 -15986 931 -15933
rect 984 -15986 1110 -15933
rect 1163 -15986 1289 -15933
rect 1342 -15986 1466 -15933
rect 1519 -15986 1643 -15933
rect 1696 -15986 1822 -15933
rect 1875 -15986 2000 -15933
rect 2053 -15986 2179 -15933
rect 2232 -15986 2356 -15933
rect 2409 -15986 2534 -15933
rect 2587 -15986 2712 -15933
rect 2765 -15986 2891 -15933
rect 2944 -15986 3068 -15933
rect 3121 -15986 3247 -15933
rect 3300 -15986 3424 -15933
rect 3477 -15986 3603 -15933
rect 3656 -15986 3780 -15933
rect -1915 -15996 -1862 -15986
rect -1738 -15996 -1685 -15986
rect -1560 -15996 -1507 -15986
rect -1382 -15996 -1329 -15986
rect -1204 -15996 -1151 -15986
rect -1025 -15996 -972 -15986
rect -847 -15996 -794 -15986
rect -670 -15996 -617 -15986
rect -491 -15996 -438 -15986
rect -313 -15996 -260 -15986
rect -136 -15996 -83 -15986
rect 43 -15996 96 -15986
rect 221 -15996 274 -15986
rect 398 -15996 451 -15986
rect 575 -15996 628 -15986
rect 755 -15996 808 -15986
rect 931 -15996 984 -15986
rect 1110 -15996 1163 -15986
rect 1289 -15996 1342 -15986
rect 1466 -15996 1519 -15986
rect 1643 -15996 1696 -15986
rect 1822 -15996 1875 -15986
rect 2000 -15996 2053 -15986
rect 2179 -15996 2232 -15986
rect 2356 -15996 2409 -15986
rect 2534 -15996 2587 -15986
rect 2712 -15996 2765 -15986
rect 2891 -15996 2944 -15986
rect 3068 -15996 3121 -15986
rect 3247 -15996 3300 -15986
rect 3424 -15996 3477 -15986
rect 3603 -15996 3656 -15986
rect 3780 -15996 3833 -15986
rect 5921 -15947 5974 -15938
rect 6279 -15947 6332 -15938
rect 6634 -15947 6687 -15938
rect 6994 -15947 7047 -15941
rect 5921 -15948 7047 -15947
rect 5974 -16000 6279 -15948
rect 5921 -16011 5974 -16001
rect 6332 -16000 6634 -15948
rect 6279 -16011 6332 -16001
rect 6687 -15951 7047 -15948
rect 6687 -16000 6994 -15951
rect 6634 -16011 6687 -16001
rect 6994 -16014 7047 -16004
rect 7526 -15952 7579 -15943
rect 7881 -15952 7934 -15942
rect 8237 -15952 8290 -15942
rect 11441 -15952 11494 -15942
rect 11797 -15952 11850 -15942
rect 12154 -15952 12207 -15942
rect 12511 -15952 12564 -15942
rect 7526 -15953 7881 -15952
rect 7579 -16005 7881 -15953
rect 7934 -16005 8237 -15952
rect 8290 -16005 11441 -15952
rect 11494 -16005 11797 -15952
rect 11850 -16005 12154 -15952
rect 12207 -16005 12511 -15952
rect 7526 -16016 7579 -16006
rect 7881 -16015 7934 -16005
rect 8237 -16015 8290 -16005
rect 11441 -16015 11494 -16005
rect 11797 -16015 11850 -16005
rect 12154 -16015 12207 -16005
rect 12511 -16015 12564 -16005
rect -6159 -16193 -6106 -16183
rect -5504 -16193 -5451 -16183
rect -4792 -16193 -4739 -16183
rect -6106 -16246 -5504 -16193
rect -5451 -16246 -4792 -16193
rect -6159 -16256 -6106 -16246
rect -5504 -16256 -5451 -16246
rect -4792 -16256 -4739 -16246
rect -5860 -16294 -5807 -16284
rect -5148 -16294 -5095 -16284
rect -4436 -16294 -4383 -16284
rect -3935 -16294 -3883 -16285
rect -5807 -16347 -5148 -16294
rect -5095 -16346 -4436 -16294
rect -5860 -16357 -5807 -16347
rect -5148 -16357 -5095 -16347
rect -4383 -16295 -3883 -16294
rect -4383 -16346 -3935 -16295
rect -4436 -16357 -4383 -16347
rect -3935 -16357 -3883 -16347
rect -1917 -16542 -1864 -16532
rect -1738 -16542 -1685 -16532
rect -1561 -16541 -1508 -16531
rect -1864 -16595 -1738 -16542
rect -1685 -16594 -1561 -16542
rect -1381 -16542 -1328 -16533
rect -1204 -16542 -1151 -16532
rect -1026 -16542 -973 -16532
rect 220 -16542 273 -16532
rect 397 -16542 450 -16532
rect 576 -16542 629 -16532
rect 755 -16542 808 -16532
rect 933 -16542 986 -16532
rect 1111 -16542 1164 -16532
rect 2356 -16542 2409 -16532
rect 2534 -16542 2587 -16532
rect 2713 -16541 2766 -16531
rect -1508 -16543 -1204 -16542
rect -1508 -16594 -1381 -16543
rect -1685 -16595 -1381 -16594
rect -1917 -16605 -1864 -16595
rect -1738 -16605 -1685 -16595
rect -1561 -16604 -1508 -16595
rect -1328 -16595 -1204 -16543
rect -1151 -16595 -1026 -16542
rect -973 -16595 220 -16542
rect 273 -16595 397 -16542
rect 450 -16595 576 -16542
rect 629 -16595 755 -16542
rect 808 -16595 933 -16542
rect 986 -16595 1111 -16542
rect 1164 -16595 2356 -16542
rect 2409 -16595 2534 -16542
rect 2587 -16594 2713 -16542
rect 2891 -16542 2944 -16532
rect 3070 -16542 3123 -16532
rect 3249 -16542 3302 -16532
rect 4238 -16542 4291 -16532
rect 2766 -16594 2891 -16542
rect 2587 -16595 2891 -16594
rect 2944 -16595 3070 -16542
rect 3123 -16595 3249 -16542
rect 3302 -16595 4238 -16542
rect -1381 -16606 -1328 -16596
rect -1204 -16605 -1151 -16595
rect -1026 -16605 -973 -16595
rect 220 -16605 273 -16595
rect 397 -16605 450 -16595
rect 576 -16605 629 -16595
rect 755 -16605 808 -16595
rect 933 -16605 986 -16595
rect 1111 -16605 1164 -16595
rect 2356 -16605 2409 -16595
rect 2534 -16605 2587 -16595
rect 2713 -16604 2766 -16595
rect 2891 -16605 2944 -16595
rect 3070 -16605 3123 -16595
rect 3249 -16605 3302 -16595
rect 4238 -16605 4291 -16595
rect 6548 -16544 6601 -16534
rect 6726 -16544 6779 -16534
rect 6601 -16597 6726 -16545
rect 6903 -16545 6956 -16535
rect 7970 -16545 8023 -16535
rect 8149 -16544 8202 -16534
rect 6779 -16597 6903 -16545
rect 6548 -16598 6903 -16597
rect 6956 -16598 7970 -16545
rect 8023 -16597 8149 -16545
rect 9929 -16544 9982 -16534
rect 8202 -16597 9929 -16545
rect 10107 -16545 10160 -16535
rect 10287 -16545 10340 -16535
rect 11352 -16545 11405 -16535
rect 11530 -16545 11583 -16536
rect 11709 -16545 11762 -16535
rect 9982 -16597 10107 -16545
rect 8023 -16598 10107 -16597
rect 10160 -16598 10287 -16545
rect 10340 -16598 11352 -16545
rect 11405 -16546 11709 -16545
rect 11405 -16598 11530 -16546
rect 6548 -16607 6601 -16598
rect 6726 -16607 6779 -16598
rect 6903 -16608 6956 -16598
rect 7970 -16608 8023 -16598
rect 8149 -16607 8202 -16598
rect 9929 -16607 9982 -16598
rect 10107 -16608 10160 -16598
rect 10287 -16608 10340 -16598
rect 11352 -16608 11405 -16598
rect 11583 -16598 11709 -16546
rect 11530 -16609 11583 -16599
rect 11709 -16608 11762 -16598
rect -1827 -16665 -1774 -16655
rect -1471 -16665 -1418 -16656
rect -1114 -16665 -1061 -16655
rect -759 -16664 -706 -16654
rect -1774 -16666 -1114 -16665
rect -1774 -16718 -1471 -16666
rect -1827 -16728 -1774 -16718
rect -1418 -16718 -1114 -16666
rect -1061 -16717 -759 -16665
rect -403 -16665 -350 -16655
rect -47 -16665 6 -16655
rect 309 -16665 362 -16656
rect 665 -16665 718 -16655
rect 845 -16665 898 -16655
rect 1021 -16665 1074 -16655
rect 1377 -16665 1430 -16655
rect 1735 -16665 1788 -16655
rect 2090 -16664 2143 -16654
rect -706 -16717 -403 -16665
rect -1061 -16718 -403 -16717
rect -350 -16718 -47 -16665
rect 6 -16666 665 -16665
rect 6 -16718 309 -16666
rect -1471 -16729 -1418 -16719
rect -1114 -16728 -1061 -16718
rect -759 -16727 -706 -16718
rect -403 -16728 -350 -16718
rect -47 -16728 6 -16718
rect 362 -16718 665 -16666
rect 718 -16718 845 -16665
rect 898 -16718 1021 -16665
rect 1074 -16718 1377 -16665
rect 1430 -16718 1735 -16665
rect 1788 -16717 2090 -16665
rect 2445 -16665 2498 -16655
rect 2801 -16665 2854 -16655
rect 3157 -16664 3210 -16654
rect 2143 -16717 2445 -16665
rect 1788 -16718 2445 -16717
rect 2498 -16718 2801 -16665
rect 2854 -16717 3157 -16665
rect 3514 -16665 3567 -16656
rect 3868 -16665 3921 -16655
rect 3210 -16666 3868 -16665
rect 3210 -16717 3514 -16666
rect 2854 -16718 3514 -16717
rect 309 -16729 362 -16719
rect 665 -16728 718 -16718
rect 845 -16728 898 -16718
rect 1021 -16728 1074 -16718
rect 1377 -16728 1430 -16718
rect 1735 -16728 1788 -16718
rect 2090 -16727 2143 -16718
rect 2445 -16728 2498 -16718
rect 2801 -16728 2854 -16718
rect 3157 -16727 3210 -16718
rect 3567 -16718 3868 -16666
rect 3514 -16729 3567 -16719
rect 3868 -16728 3921 -16718
rect 5399 -16666 5452 -16657
rect 8771 -16666 8824 -16656
rect 9128 -16666 9181 -16656
rect 9484 -16666 9537 -16656
rect 5399 -16667 8771 -16666
rect 5452 -16719 8771 -16667
rect 8824 -16719 9128 -16666
rect 9181 -16719 9484 -16666
rect 5399 -16730 5452 -16720
rect 8771 -16729 8824 -16719
rect 9128 -16729 9181 -16719
rect 9484 -16729 9537 -16719
rect 9838 -16665 9891 -16656
rect 10195 -16665 10248 -16655
rect 10550 -16665 10603 -16655
rect 10907 -16665 10960 -16655
rect 9838 -16666 10195 -16665
rect 9891 -16718 10195 -16666
rect 10248 -16718 10550 -16665
rect 10603 -16718 10907 -16665
rect 9838 -16729 9891 -16719
rect 10195 -16728 10248 -16718
rect 10550 -16728 10603 -16718
rect 10907 -16728 10960 -16718
rect 5031 -16782 5084 -16772
rect 8950 -16782 9003 -16772
rect 9305 -16782 9358 -16772
rect 5084 -16835 8950 -16782
rect 9003 -16835 9305 -16782
rect 5031 -16845 5084 -16835
rect 8950 -16845 9003 -16835
rect 9305 -16845 9358 -16835
rect 10017 -16780 10070 -16771
rect 10374 -16780 10427 -16771
rect 10731 -16779 10784 -16769
rect 10017 -16781 10731 -16780
rect 10070 -16833 10374 -16781
rect 10017 -16844 10070 -16834
rect 10427 -16832 10731 -16781
rect 10427 -16833 10784 -16832
rect 10374 -16844 10427 -16834
rect 10731 -16842 10784 -16833
rect -5682 -16886 -5629 -16876
rect -5326 -16886 -5273 -16876
rect -4970 -16886 -4917 -16876
rect -4614 -16886 -4561 -16876
rect -4258 -16886 -4205 -16876
rect -5629 -16939 -5326 -16886
rect -5273 -16939 -4970 -16886
rect -4917 -16939 -4614 -16886
rect -4561 -16939 -4258 -16886
rect -5682 -16949 -5629 -16939
rect -5326 -16949 -5273 -16939
rect -4970 -16949 -4917 -16939
rect -4614 -16949 -4561 -16939
rect -4258 -16949 -4205 -16939
rect 7347 -16890 7400 -16880
rect 7704 -16890 7757 -16880
rect 8060 -16890 8113 -16880
rect 8416 -16890 8469 -16880
rect 11263 -16890 11316 -16880
rect 11620 -16890 11673 -16880
rect 11975 -16889 12028 -16879
rect 7400 -16943 7704 -16890
rect 7757 -16943 8060 -16890
rect 8113 -16943 8416 -16890
rect 8469 -16943 11263 -16890
rect 11316 -16943 11620 -16890
rect 11673 -16942 11975 -16890
rect 12331 -16889 12384 -16879
rect 12028 -16942 12331 -16890
rect 11673 -16943 12384 -16942
rect 7347 -16953 7400 -16943
rect 7704 -16953 7757 -16943
rect 8060 -16953 8113 -16943
rect 8416 -16953 8469 -16943
rect 11263 -16953 11316 -16943
rect 11620 -16953 11673 -16943
rect 11975 -16952 12028 -16943
rect 12331 -16952 12384 -16943
rect -6159 -17007 -6106 -16997
rect -5859 -17007 -5806 -16997
rect -5148 -17007 -5095 -16997
rect -4437 -17007 -4384 -16997
rect -6106 -17060 -5859 -17007
rect -5806 -17060 -5148 -17007
rect -5095 -17060 -4437 -17007
rect -6159 -17070 -6106 -17060
rect -5859 -17070 -5806 -17060
rect -5148 -17070 -5095 -17060
rect -4437 -17070 -4384 -17060
rect -5504 -17118 -5451 -17108
rect -4792 -17118 -4739 -17108
rect -3935 -17118 -3883 -17108
rect -5451 -17170 -4792 -17118
rect -5504 -17181 -5451 -17171
rect -4739 -17170 -3935 -17118
rect -4792 -17181 -4739 -17171
rect -3935 -17180 -3883 -17170
<< via2 >>
rect 6451 2665 6515 2729
rect 17950 2665 18014 2729
rect 6704 1857 6768 1921
rect 15793 2164 15857 2228
rect 17697 1858 17761 1922
rect 11098 1223 11162 1287
rect 10730 943 10794 1007
rect 6451 865 6515 929
rect 17950 865 18014 929
rect 8625 360 8689 424
rect 15806 362 15870 426
rect 6704 57 6768 121
rect 12512 248 12576 312
rect 8905 -363 8969 -299
rect 10384 79 10448 143
rect 6451 -935 6515 -871
rect 10732 80 10796 144
rect 10530 -1314 10594 -1250
rect 6704 -1743 6768 -1679
rect 12259 25 12323 89
rect 17697 58 17761 122
rect 12512 -364 12576 -300
rect 12259 -449 12323 -385
rect 13760 -427 13824 -363
rect 14520 -427 14584 -363
rect 12870 -605 12934 -541
rect 13186 -605 13250 -541
rect 14808 -605 14872 -541
rect 15268 -601 15332 -537
rect 12208 -970 12272 -906
rect 17950 -935 18014 -871
rect 14309 -1143 14373 -1079
rect 12410 -1321 12474 -1257
rect 13978 -1553 14042 -1489
rect 14308 -1553 14372 -1489
rect 9435 -2050 9499 -1986
rect 9867 -2050 9931 -1986
rect 10510 -2050 10574 -1986
rect 10733 -2050 10797 -1986
rect 9435 -2206 9499 -2142
rect 6451 -2735 6515 -2671
rect 9435 -2379 9499 -2315
rect 9866 -2380 9930 -2316
rect 12408 -1671 12472 -1607
rect 13976 -1891 14040 -1827
rect 17697 -1742 17761 -1678
rect 13612 -2071 13676 -2007
rect 13610 -2382 13674 -2318
rect 12408 -2910 12472 -2846
rect 17950 -2735 18014 -2671
rect 3019 -3513 3080 -3452
rect 6704 -3543 6768 -3479
rect 12410 -3310 12474 -3246
rect 17697 -3542 17761 -3478
rect 9642 -3859 9706 -3795
rect 10932 -3859 10996 -3795
rect 11432 -3893 11496 -3829
rect 13539 -3829 13603 -3765
rect 14528 -3829 14592 -3765
rect -2546 -3989 -2485 -3928
rect 12704 -4007 12768 -3943
rect 12996 -4011 13060 -3947
rect 14838 -4011 14902 -3947
rect 15254 -4007 15318 -3943
rect 9272 -4192 9336 -4128
rect 10032 -4192 10096 -4128
rect 13045 -4192 13109 -4128
rect 13428 -4192 13492 -4128
rect 2538 -4327 2599 -4266
rect -2385 -4566 -2324 -4505
rect 2746 -4507 2807 -4446
rect 6451 -4535 6515 -4471
rect 17950 -4535 18014 -4471
rect 3021 -5063 3082 -5002
rect -2385 -5154 -2324 -5093
rect 311 -5209 372 -5148
rect 15802 -5040 15866 -4976
rect 10525 -5184 10589 -5120
rect -1646 -5339 -1585 -5278
rect 846 -5339 907 -5278
rect 6704 -5343 6768 -5279
rect 17697 -5342 17761 -5278
rect -3545 -6867 -3484 -6806
rect -3386 -7040 -3325 -6979
rect 9262 -5751 9326 -5687
rect 6451 -6335 6515 -6271
rect 8738 -6607 8802 -6543
rect 17950 -6335 18014 -6271
rect 15820 -6832 15884 -6768
rect 6704 -7143 6768 -7079
rect 17697 -7142 17761 -7078
<< metal3 >>
rect 6451 2734 6515 2739
rect 6441 2729 6525 2734
rect 6441 2665 6451 2729
rect 6515 2665 6525 2729
rect 6441 2660 6525 2665
rect 6451 934 6515 2660
rect 6704 1926 6768 1931
rect 6694 1921 6778 1926
rect 6694 1857 6704 1921
rect 6768 1857 6778 1921
rect 6694 1852 6778 1857
rect 6441 929 6525 934
rect 6441 865 6451 929
rect 6515 865 6525 929
rect 6441 860 6525 865
rect 6451 -866 6515 860
rect 6704 126 6768 1852
rect 7302 1731 8460 2891
rect 9102 1731 10260 2891
rect 10902 1731 12060 2891
rect 12702 1731 13860 2891
rect 14502 1731 15660 2891
rect 15783 2228 15867 2233
rect 15783 2164 15793 2228
rect 15857 2164 15867 2228
rect 15783 2159 15867 2164
rect 11077 1287 11182 1311
rect 15793 1310 15857 2159
rect 16302 1731 17460 2891
rect 17950 2734 18014 2739
rect 17940 2729 18024 2734
rect 17940 2665 17950 2729
rect 18014 2665 18024 2729
rect 17940 2660 18024 2665
rect 17697 1927 17761 1932
rect 17687 1922 17771 1927
rect 17687 1858 17697 1922
rect 17761 1858 17771 1922
rect 17687 1853 17771 1858
rect 11077 1223 11098 1287
rect 11162 1223 11182 1287
rect 11077 1200 11182 1223
rect 15293 1246 15857 1310
rect 15293 1091 15357 1246
rect 6694 121 6778 126
rect 6694 57 6704 121
rect 6768 57 6778 121
rect 6694 52 6778 57
rect 6441 -871 6525 -866
rect 6441 -935 6451 -871
rect 6515 -935 6525 -871
rect 6441 -940 6525 -935
rect 6451 -945 6515 -940
rect 6704 -1674 6768 52
rect 7302 -69 8460 1091
rect 8605 424 8711 446
rect 8605 360 8625 424
rect 8689 360 8711 424
rect 8605 339 8711 360
rect 9102 143 10260 1091
rect 10720 1007 10804 1012
rect 10902 1007 12060 1091
rect 10720 943 10730 1007
rect 10794 943 12060 1007
rect 10720 938 10804 943
rect 10374 143 10458 148
rect 9102 79 10384 143
rect 10448 79 10458 143
rect 9102 -69 10260 79
rect 10374 74 10458 79
rect 10718 144 10810 177
rect 10718 80 10732 144
rect 10796 80 10810 144
rect 10718 55 10810 80
rect 10902 -69 12060 943
rect 12702 728 13860 1091
rect 12259 664 13860 728
rect 12259 94 12323 664
rect 12502 312 12586 341
rect 12502 248 12512 312
rect 12576 248 12586 312
rect 12502 224 12586 248
rect 12249 89 12333 94
rect 12249 25 12259 89
rect 12323 25 12333 89
rect 12249 20 12333 25
rect 12702 -69 13860 664
rect 14502 -69 15660 1091
rect 15788 426 15886 445
rect 15788 362 15806 426
rect 15870 362 15886 426
rect 15788 345 15886 362
rect 16302 -69 17460 1091
rect 17697 127 17761 1853
rect 17950 934 18014 2660
rect 17940 929 18024 934
rect 17940 865 17950 929
rect 18014 865 18024 929
rect 17940 860 18024 865
rect 17687 122 17771 127
rect 17687 58 17697 122
rect 17761 58 17771 122
rect 17687 53 17771 58
rect 9646 -158 9710 -69
rect 9646 -222 14207 -158
rect 8864 -299 9004 -268
rect 8864 -363 8905 -299
rect 8969 -363 9004 -299
rect 8864 -397 9004 -363
rect 12481 -300 12610 -292
rect 12481 -364 12512 -300
rect 12576 -364 12610 -300
rect 12481 -372 12610 -364
rect 13750 -363 13834 -358
rect 12249 -385 12333 -380
rect 9856 -449 12259 -385
rect 12323 -449 12333 -385
rect 13750 -427 13760 -363
rect 13824 -427 13834 -363
rect 13750 -432 13834 -427
rect 9856 -709 9920 -449
rect 12249 -454 12333 -449
rect 12860 -541 12944 -536
rect 10343 -605 12870 -541
rect 12934 -605 12944 -541
rect 6694 -1679 6778 -1674
rect 6694 -1743 6704 -1679
rect 6768 -1743 6778 -1679
rect 6694 -1748 6778 -1743
rect 7302 -1869 8460 -709
rect 9102 -1869 10260 -709
rect 9435 -1981 9499 -1869
rect 9425 -1986 9509 -1981
rect 9425 -2050 9435 -1986
rect 9499 -2050 9509 -1986
rect 9425 -2055 9509 -2050
rect 9845 -1986 9951 -1968
rect 9845 -2050 9867 -1986
rect 9931 -2050 9951 -1986
rect 9435 -2137 9499 -2055
rect 9845 -2065 9951 -2050
rect 9425 -2142 9509 -2137
rect 9425 -2206 9435 -2142
rect 9499 -2206 9509 -2142
rect 9425 -2211 9509 -2206
rect 9435 -2310 9499 -2211
rect 9425 -2315 9509 -2310
rect 9425 -2379 9435 -2315
rect 9499 -2379 9509 -2315
rect 9425 -2384 9509 -2379
rect 9847 -2311 9939 -2286
rect 9847 -2316 9940 -2311
rect 9847 -2380 9866 -2316
rect 9930 -2380 9940 -2316
rect 9435 -2509 9499 -2384
rect 9847 -2385 9940 -2380
rect 9847 -2408 9939 -2385
rect 6451 -2666 6515 -2661
rect 6441 -2671 6525 -2666
rect 6441 -2735 6451 -2671
rect 6515 -2735 6525 -2671
rect 6441 -2740 6525 -2735
rect 3009 -3452 3090 -3447
rect 3009 -3513 3019 -3452
rect 3080 -3513 3090 -3452
rect 3009 -3518 3090 -3513
rect -2556 -3928 -2475 -3923
rect -2556 -3989 -2546 -3928
rect -2485 -3989 -2475 -3928
rect -2556 -3994 -2475 -3989
rect -2546 -4266 -2485 -3994
rect 2528 -4266 2609 -4261
rect -2546 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect -2546 -6637 -2485 -4327
rect 2528 -4332 2609 -4327
rect 2736 -4446 2817 -4441
rect -2385 -4500 2746 -4446
rect -2395 -4505 2746 -4500
rect -2395 -4566 -2385 -4505
rect -2324 -4507 2746 -4505
rect 2807 -4507 2817 -4446
rect -2324 -4566 -2314 -4507
rect 2736 -4512 2817 -4507
rect -2395 -4571 -2314 -4566
rect -2385 -5088 -2324 -4571
rect 3021 -4997 3082 -3518
rect 6451 -4466 6515 -2740
rect 6704 -3474 6768 -3469
rect 6694 -3479 6778 -3474
rect 6694 -3543 6704 -3479
rect 6768 -3543 6778 -3479
rect 6694 -3548 6778 -3543
rect 6441 -4471 6525 -4466
rect 6441 -4535 6451 -4471
rect 6515 -4535 6525 -4471
rect 6441 -4540 6525 -4535
rect 3011 -5002 3092 -4997
rect 3011 -5063 3021 -5002
rect 3082 -5063 3092 -5002
rect 3011 -5068 3092 -5063
rect -2395 -5093 -2314 -5088
rect -2395 -5154 -2385 -5093
rect -2324 -5154 -2314 -5093
rect -2395 -5159 -2314 -5154
rect 301 -5147 382 -5143
rect 3021 -5147 3082 -5068
rect 301 -5148 3082 -5147
rect -3545 -6698 -2485 -6637
rect -3545 -6801 -3484 -6698
rect -2385 -6786 -2324 -5159
rect 301 -5209 311 -5148
rect 372 -5208 3082 -5148
rect 372 -5209 382 -5208
rect 301 -5214 382 -5209
rect -1656 -5278 -1575 -5273
rect 836 -5278 917 -5273
rect -1656 -5339 -1646 -5278
rect -1585 -5339 846 -5278
rect 907 -5339 917 -5278
rect -1656 -5344 -1575 -5339
rect 836 -5344 917 -5339
rect 6451 -6266 6515 -4540
rect 6704 -5274 6768 -3548
rect 7302 -3669 8460 -2509
rect 9102 -3669 10260 -2509
rect 9272 -4123 9336 -3669
rect 9632 -3795 9716 -3790
rect 9632 -3859 9642 -3795
rect 9706 -3859 9716 -3795
rect 9632 -3864 9716 -3859
rect 9262 -4128 9346 -4123
rect 9262 -4192 9272 -4128
rect 9336 -4192 9346 -4128
rect 9262 -4197 9346 -4192
rect 9642 -4309 9706 -3864
rect 10012 -4128 10113 -4112
rect 10012 -4192 10032 -4128
rect 10096 -4192 10113 -4128
rect 10012 -4210 10113 -4192
rect 6694 -5279 6778 -5274
rect 6694 -5343 6704 -5279
rect 6768 -5343 6778 -5279
rect 6694 -5348 6778 -5343
rect 6441 -6271 6525 -6266
rect 6441 -6335 6451 -6271
rect 6515 -6335 6525 -6271
rect 6441 -6340 6525 -6335
rect 6451 -6345 6515 -6340
rect -3555 -6806 -3474 -6801
rect -3555 -6867 -3545 -6806
rect -3484 -6867 -3474 -6806
rect -3555 -6872 -3474 -6867
rect -3386 -6847 -2324 -6786
rect -3386 -6974 -3325 -6847
rect -3396 -6979 -3315 -6974
rect -3396 -7040 -3386 -6979
rect -3325 -7040 -3315 -6979
rect -3396 -7045 -3315 -7040
rect 6704 -7074 6768 -5348
rect 7302 -5469 8460 -4309
rect 9102 -5115 10260 -4309
rect 10343 -5115 10407 -605
rect 12860 -610 12944 -605
rect 13163 -541 13273 -525
rect 13163 -605 13186 -541
rect 13250 -605 13273 -541
rect 13163 -619 13273 -605
rect 13760 -709 13824 -432
rect 10520 -1250 10604 -1245
rect 10902 -1250 12060 -709
rect 12183 -906 12292 -883
rect 12183 -970 12208 -906
rect 12272 -970 12292 -906
rect 12183 -990 12292 -970
rect 10520 -1314 10530 -1250
rect 10594 -1314 12060 -1250
rect 10520 -1319 10604 -1314
rect 10902 -1869 12060 -1314
rect 12400 -1257 12484 -1252
rect 12702 -1257 13860 -709
rect 12400 -1321 12410 -1257
rect 12474 -1321 13860 -1257
rect 12400 -1326 12484 -1321
rect 12385 -1607 12491 -1584
rect 12385 -1671 12408 -1607
rect 12472 -1671 12491 -1607
rect 12385 -1691 12491 -1671
rect 12702 -1869 13860 -1321
rect 13964 -1489 14055 -1450
rect 13964 -1553 13978 -1489
rect 14042 -1553 14055 -1489
rect 13964 -1590 14055 -1553
rect 13966 -1827 14050 -1822
rect 10499 -1986 10586 -1952
rect 10499 -2050 10510 -1986
rect 10574 -2050 10586 -1986
rect 10499 -2081 10586 -2050
rect 10723 -1986 10807 -1981
rect 10723 -2050 10733 -1986
rect 10797 -2050 10807 -1986
rect 10723 -2055 10807 -2050
rect 11450 -2037 11514 -1869
rect 13966 -1891 13976 -1827
rect 14040 -1891 14050 -1827
rect 13966 -1896 14050 -1891
rect 13581 -2007 13706 -1977
rect 9102 -5179 10407 -5115
rect 10507 -5120 10605 -5089
rect 9102 -5469 10260 -5179
rect 10507 -5184 10525 -5120
rect 10589 -5184 10605 -5120
rect 10733 -5104 10797 -2055
rect 11450 -2101 13014 -2037
rect 13581 -2071 13612 -2007
rect 13676 -2071 13706 -2007
rect 13581 -2098 13706 -2071
rect 12950 -2509 13014 -2101
rect 13588 -2318 13692 -2298
rect 13588 -2382 13610 -2318
rect 13674 -2382 13692 -2318
rect 13588 -2398 13692 -2382
rect 10902 -3246 12060 -2509
rect 12386 -2846 12492 -2824
rect 12386 -2910 12408 -2846
rect 12472 -2910 12492 -2846
rect 12386 -2931 12492 -2910
rect 12400 -3246 12484 -3241
rect 10902 -3310 12410 -3246
rect 12474 -3310 12484 -3246
rect 10902 -3669 12060 -3310
rect 12400 -3315 12484 -3310
rect 12702 -3669 13860 -2509
rect 10932 -3790 10996 -3669
rect 13539 -3760 13603 -3669
rect 13529 -3765 13613 -3760
rect 10922 -3795 11006 -3790
rect 10922 -3859 10932 -3795
rect 10996 -3859 11006 -3795
rect 10922 -3864 11006 -3859
rect 11409 -3829 11517 -3803
rect 11409 -3893 11432 -3829
rect 11496 -3893 11517 -3829
rect 13529 -3829 13539 -3765
rect 13603 -3829 13613 -3765
rect 13529 -3834 13613 -3829
rect 11409 -3916 11517 -3893
rect 12694 -3943 12778 -3938
rect 12185 -4007 12704 -3943
rect 12768 -4007 12778 -3943
rect 10902 -5104 12060 -4309
rect 10733 -5106 12060 -5104
rect 12185 -5106 12249 -4007
rect 12694 -4012 12778 -4007
rect 12975 -3947 13080 -3923
rect 12975 -4011 12996 -3947
rect 13060 -4011 13080 -3947
rect 12975 -4032 13080 -4011
rect 13025 -4128 13126 -4109
rect 13025 -4192 13045 -4128
rect 13109 -4192 13126 -4128
rect 13025 -4207 13126 -4192
rect 13418 -4128 13502 -4123
rect 13418 -4192 13428 -4128
rect 13492 -4192 13502 -4128
rect 13418 -4197 13502 -4192
rect 13428 -4309 13492 -4197
rect 10733 -5168 12249 -5106
rect 10507 -5209 10605 -5184
rect 10902 -5170 12249 -5168
rect 12702 -5021 13860 -4309
rect 13976 -5021 14040 -1896
rect 14143 -4853 14207 -222
rect 14520 -358 14584 -69
rect 14510 -363 14594 -358
rect 14510 -427 14520 -363
rect 14584 -427 14594 -363
rect 14510 -432 14594 -427
rect 14785 -541 14895 -526
rect 15268 -532 15332 -69
rect 14785 -605 14808 -541
rect 14872 -605 14895 -541
rect 14785 -620 14895 -605
rect 15258 -537 15342 -532
rect 15258 -601 15268 -537
rect 15332 -601 15342 -537
rect 15258 -606 15342 -601
rect 14299 -1079 14383 -1074
rect 14502 -1079 15660 -709
rect 14299 -1143 14309 -1079
rect 14373 -1143 15660 -1079
rect 14299 -1148 14383 -1143
rect 14295 -1489 14386 -1451
rect 14295 -1553 14308 -1489
rect 14372 -1553 14386 -1489
rect 14295 -1591 14386 -1553
rect 14502 -1869 15660 -1143
rect 16302 -1869 17460 -709
rect 17697 -1673 17761 53
rect 17950 -866 18014 860
rect 17940 -871 18024 -866
rect 17940 -935 17950 -871
rect 18014 -935 18024 -871
rect 17940 -940 18024 -935
rect 17687 -1678 17771 -1673
rect 17687 -1742 17697 -1678
rect 17761 -1742 17771 -1678
rect 17687 -1747 17771 -1742
rect 17697 -1752 17761 -1747
rect 14502 -3669 15660 -2509
rect 16302 -3669 17460 -2509
rect 17950 -2666 18014 -2661
rect 17940 -2671 18024 -2666
rect 17940 -2735 17950 -2671
rect 18014 -2735 18024 -2671
rect 17940 -2740 18024 -2735
rect 17697 -3473 17761 -3468
rect 17687 -3478 17771 -3473
rect 17687 -3542 17697 -3478
rect 17761 -3542 17771 -3478
rect 17687 -3547 17771 -3542
rect 14518 -3765 14602 -3760
rect 14518 -3829 14528 -3765
rect 14592 -3829 14602 -3765
rect 14518 -3834 14602 -3829
rect 14528 -4309 14592 -3834
rect 14817 -3947 14922 -3925
rect 15254 -3938 15318 -3669
rect 14817 -4011 14838 -3947
rect 14902 -4011 14922 -3947
rect 14817 -4034 14922 -4011
rect 15244 -3943 15328 -3938
rect 15244 -4007 15254 -3943
rect 15318 -4007 15328 -3943
rect 15244 -4012 15328 -4007
rect 14502 -4853 15660 -4309
rect 14143 -4917 15660 -4853
rect 12702 -5085 14043 -5021
rect 10902 -5469 12060 -5170
rect 12702 -5469 13860 -5085
rect 14502 -5469 15660 -4917
rect 15785 -4976 15887 -4955
rect 15785 -5040 15802 -4976
rect 15866 -5040 15887 -4976
rect 15785 -5058 15887 -5040
rect 16302 -5469 17460 -4309
rect 17697 -5273 17761 -3547
rect 17950 -4466 18014 -2740
rect 17940 -4471 18024 -4466
rect 17940 -4535 17950 -4471
rect 18014 -4535 18024 -4471
rect 17940 -4540 18024 -4535
rect 17687 -5278 17771 -5273
rect 17687 -5342 17697 -5278
rect 17761 -5342 17771 -5278
rect 17687 -5347 17771 -5342
rect 9241 -5687 9347 -5664
rect 9241 -5751 9262 -5687
rect 9326 -5751 9347 -5687
rect 9241 -5768 9347 -5751
rect 15281 -5911 15345 -5469
rect 15281 -5975 15884 -5911
rect 6694 -7079 6778 -7074
rect 6694 -7143 6704 -7079
rect 6768 -7143 6778 -7079
rect 6694 -7148 6778 -7143
rect 6704 -7153 6768 -7148
rect 7302 -7269 8460 -6109
rect 8724 -6543 8822 -6525
rect 8724 -6607 8738 -6543
rect 8802 -6607 8822 -6543
rect 8724 -6628 8822 -6607
rect 9102 -7269 10260 -6109
rect 10902 -7269 12060 -6109
rect 12702 -7269 13860 -6109
rect 14502 -7269 15660 -6109
rect 15820 -6763 15884 -5975
rect 15810 -6768 15894 -6763
rect 15810 -6832 15820 -6768
rect 15884 -6832 15894 -6768
rect 15810 -6837 15894 -6832
rect 15820 -6841 15884 -6837
rect 16302 -7269 17460 -6109
rect 17697 -7073 17761 -5347
rect 17950 -6266 18014 -4540
rect 17940 -6271 18024 -6266
rect 17940 -6335 17950 -6271
rect 18014 -6335 18024 -6271
rect 17940 -6340 18024 -6335
rect 17687 -7078 17771 -7073
rect 17687 -7142 17697 -7078
rect 17761 -7142 17771 -7078
rect 17687 -7147 17771 -7142
rect 17697 -7152 17761 -7147
<< via3 >>
rect 11098 1223 11162 1287
rect 8625 360 8689 424
rect 10732 80 10796 144
rect 12512 248 12576 312
rect 15806 362 15870 426
rect 8905 -363 8969 -299
rect 12512 -364 12576 -300
rect 9867 -2050 9931 -1986
rect 9866 -2380 9930 -2316
rect 10032 -4192 10096 -4128
rect 13186 -605 13250 -541
rect 12208 -970 12272 -906
rect 12408 -1671 12472 -1607
rect 13978 -1553 14042 -1489
rect 10510 -2050 10574 -1986
rect 10525 -5184 10589 -5120
rect 13612 -2071 13676 -2007
rect 13610 -2382 13674 -2318
rect 12408 -2910 12472 -2846
rect 11432 -3893 11496 -3829
rect 12996 -4011 13060 -3947
rect 13045 -4192 13109 -4128
rect 14808 -605 14872 -541
rect 14308 -1553 14372 -1489
rect 14838 -4011 14902 -3947
rect 15802 -5040 15866 -4976
rect 9262 -5751 9326 -5687
rect 8738 -6607 8802 -6543
<< mimcap >>
rect 7402 2751 8362 2791
rect 7402 1871 7442 2751
rect 8322 1871 8362 2751
rect 7402 1831 8362 1871
rect 9202 2751 10162 2791
rect 9202 1871 9242 2751
rect 10122 1871 10162 2751
rect 9202 1831 10162 1871
rect 11002 2751 11962 2791
rect 11002 1871 11042 2751
rect 11922 1871 11962 2751
rect 11002 1831 11962 1871
rect 12802 2751 13762 2791
rect 12802 1871 12842 2751
rect 13722 1871 13762 2751
rect 12802 1831 13762 1871
rect 14602 2751 15562 2791
rect 14602 1871 14642 2751
rect 15522 1871 15562 2751
rect 14602 1831 15562 1871
rect 16402 2751 17362 2791
rect 16402 1871 16442 2751
rect 17322 1871 17362 2751
rect 16402 1831 17362 1871
rect 7402 951 8362 991
rect 7402 71 7442 951
rect 8322 71 8362 951
rect 7402 31 8362 71
rect 9202 951 10162 991
rect 9202 71 9242 951
rect 10122 71 10162 951
rect 9202 31 10162 71
rect 11002 951 11962 991
rect 11002 71 11042 951
rect 11922 71 11962 951
rect 11002 31 11962 71
rect 12802 951 13762 991
rect 12802 71 12842 951
rect 13722 71 13762 951
rect 12802 31 13762 71
rect 14602 951 15562 991
rect 14602 71 14642 951
rect 15522 71 15562 951
rect 14602 31 15562 71
rect 16402 951 17362 991
rect 16402 71 16442 951
rect 17322 71 17362 951
rect 16402 31 17362 71
rect 7402 -849 8362 -809
rect 7402 -1729 7442 -849
rect 8322 -1729 8362 -849
rect 7402 -1769 8362 -1729
rect 9202 -849 10162 -809
rect 9202 -1729 9242 -849
rect 10122 -1729 10162 -849
rect 9202 -1769 10162 -1729
rect 11002 -849 11962 -809
rect 11002 -1729 11042 -849
rect 11922 -1729 11962 -849
rect 11002 -1769 11962 -1729
rect 12802 -849 13762 -809
rect 12802 -1729 12842 -849
rect 13722 -1729 13762 -849
rect 12802 -1769 13762 -1729
rect 14602 -849 15562 -809
rect 14602 -1729 14642 -849
rect 15522 -1729 15562 -849
rect 14602 -1769 15562 -1729
rect 16402 -849 17362 -809
rect 16402 -1729 16442 -849
rect 17322 -1729 17362 -849
rect 16402 -1769 17362 -1729
rect 7402 -2649 8362 -2609
rect 7402 -3529 7442 -2649
rect 8322 -3529 8362 -2649
rect 7402 -3569 8362 -3529
rect 9202 -2649 10162 -2609
rect 9202 -3529 9242 -2649
rect 10122 -3529 10162 -2649
rect 9202 -3569 10162 -3529
rect 11002 -2649 11962 -2609
rect 11002 -3529 11042 -2649
rect 11922 -3529 11962 -2649
rect 11002 -3569 11962 -3529
rect 12802 -2649 13762 -2609
rect 12802 -3529 12842 -2649
rect 13722 -3529 13762 -2649
rect 12802 -3569 13762 -3529
rect 14602 -2649 15562 -2609
rect 14602 -3529 14642 -2649
rect 15522 -3529 15562 -2649
rect 14602 -3569 15562 -3529
rect 16402 -2649 17362 -2609
rect 16402 -3529 16442 -2649
rect 17322 -3529 17362 -2649
rect 16402 -3569 17362 -3529
rect 7402 -4449 8362 -4409
rect 7402 -5329 7442 -4449
rect 8322 -5329 8362 -4449
rect 7402 -5369 8362 -5329
rect 9202 -4449 10162 -4409
rect 9202 -5329 9242 -4449
rect 10122 -5329 10162 -4449
rect 9202 -5369 10162 -5329
rect 11002 -4449 11962 -4409
rect 11002 -5329 11042 -4449
rect 11922 -5329 11962 -4449
rect 11002 -5369 11962 -5329
rect 12802 -4449 13762 -4409
rect 12802 -5329 12842 -4449
rect 13722 -5329 13762 -4449
rect 12802 -5369 13762 -5329
rect 14602 -4449 15562 -4409
rect 14602 -5329 14642 -4449
rect 15522 -5329 15562 -4449
rect 14602 -5369 15562 -5329
rect 16402 -4449 17362 -4409
rect 16402 -5329 16442 -4449
rect 17322 -5329 17362 -4449
rect 16402 -5369 17362 -5329
rect 7402 -6249 8362 -6209
rect 7402 -7129 7442 -6249
rect 8322 -7129 8362 -6249
rect 7402 -7169 8362 -7129
rect 9202 -6249 10162 -6209
rect 9202 -7129 9242 -6249
rect 10122 -7129 10162 -6249
rect 9202 -7169 10162 -7129
rect 11002 -6249 11962 -6209
rect 11002 -7129 11042 -6249
rect 11922 -7129 11962 -6249
rect 11002 -7169 11962 -7129
rect 12802 -6249 13762 -6209
rect 12802 -7129 12842 -6249
rect 13722 -7129 13762 -6249
rect 12802 -7169 13762 -7129
rect 14602 -6249 15562 -6209
rect 14602 -7129 14642 -6249
rect 15522 -7129 15562 -6249
rect 14602 -7169 15562 -7129
rect 16402 -6249 17362 -6209
rect 16402 -7129 16442 -6249
rect 17322 -7129 17362 -6249
rect 16402 -7169 17362 -7129
<< mimcapcontact >>
rect 7442 1871 8322 2751
rect 9242 1871 10122 2751
rect 11042 1871 11922 2751
rect 12842 1871 13722 2751
rect 14642 1871 15522 2751
rect 16442 1871 17322 2751
rect 7442 71 8322 951
rect 9242 71 10122 951
rect 11042 71 11922 951
rect 12842 71 13722 951
rect 14642 71 15522 951
rect 16442 71 17322 951
rect 7442 -1729 8322 -849
rect 9242 -1729 10122 -849
rect 11042 -1729 11922 -849
rect 12842 -1729 13722 -849
rect 14642 -1729 15522 -849
rect 16442 -1729 17322 -849
rect 7442 -3529 8322 -2649
rect 9242 -3529 10122 -2649
rect 11042 -3529 11922 -2649
rect 12842 -3529 13722 -2649
rect 14642 -3529 15522 -2649
rect 16442 -3529 17322 -2649
rect 7442 -5329 8322 -4449
rect 9242 -5329 10122 -4449
rect 11042 -5329 11922 -4449
rect 12842 -5329 13722 -4449
rect 14642 -5329 15522 -4449
rect 16442 -5329 17322 -4449
rect 7442 -7129 8322 -6249
rect 9242 -7129 10122 -6249
rect 11042 -7129 11922 -6249
rect 12842 -7129 13722 -6249
rect 14642 -7129 15522 -6249
rect 16442 -7129 17322 -6249
<< metal4 >>
rect 7441 2751 8323 2752
rect 7441 1871 7442 2751
rect 8322 1871 8323 2751
rect 7441 1870 8323 1871
rect 9241 2751 10123 2752
rect 9241 1871 9242 2751
rect 10122 1871 10123 2751
rect 9241 1870 10123 1871
rect 11041 2751 11923 2752
rect 11041 1871 11042 2751
rect 11922 1871 11923 2751
rect 11041 1870 11923 1871
rect 12841 2751 13723 2752
rect 12841 1871 12842 2751
rect 13722 1871 13723 2751
rect 12841 1870 13723 1871
rect 14641 2751 15523 2752
rect 14641 1871 14642 2751
rect 15522 1871 15523 2751
rect 14641 1870 15523 1871
rect 16441 2751 17323 2752
rect 16441 1871 16442 2751
rect 17322 1871 17323 2751
rect 16441 1870 17323 1871
rect 11097 1287 11163 1288
rect 11097 1223 11098 1287
rect 11162 1223 11163 1287
rect 11097 1222 11163 1223
rect 11098 952 11162 1222
rect 7441 951 8323 952
rect 7441 71 7442 951
rect 8322 71 8323 951
rect 9241 951 10123 952
rect 8624 424 8690 425
rect 9241 424 9242 951
rect 8624 360 8625 424
rect 8689 360 9242 424
rect 8624 359 8690 360
rect 7441 70 8323 71
rect 9241 71 9242 360
rect 10122 71 10123 951
rect 11041 951 11923 952
rect 10731 144 10797 145
rect 11041 144 11042 951
rect 10731 80 10732 144
rect 10796 80 11042 144
rect 10731 79 10797 80
rect 9241 70 10123 71
rect 11041 71 11042 80
rect 11922 71 11923 951
rect 12841 951 13723 952
rect 12511 312 12577 313
rect 12841 312 12842 951
rect 12511 248 12512 312
rect 12576 248 12842 312
rect 12511 247 12577 248
rect 11041 70 11923 71
rect 12841 71 12842 248
rect 13722 71 13723 951
rect 12841 70 13723 71
rect 14641 951 15523 952
rect 14641 71 14642 951
rect 15522 426 15523 951
rect 16441 951 17323 952
rect 15805 426 15871 427
rect 15522 362 15806 426
rect 15870 362 15871 426
rect 15522 71 15523 362
rect 15805 361 15871 362
rect 14641 70 15523 71
rect 16441 71 16442 951
rect 17322 71 17323 951
rect 16441 70 17323 71
rect 9646 -158 9710 70
rect 9646 -222 14207 -158
rect 8904 -299 8970 -298
rect 8904 -363 8905 -299
rect 8969 -300 8970 -299
rect 12511 -300 12577 -299
rect 8969 -363 12512 -300
rect 8904 -364 12512 -363
rect 12576 -364 12577 -300
rect 9422 -848 9486 -364
rect 12511 -365 12577 -364
rect 13185 -541 13251 -540
rect 10344 -605 13186 -541
rect 13250 -605 13252 -541
rect 7441 -849 8323 -848
rect 7441 -1729 7442 -849
rect 8322 -1729 8323 -849
rect 7441 -1730 8323 -1729
rect 9241 -849 10123 -848
rect 9241 -1729 9242 -849
rect 10122 -1729 10123 -849
rect 9241 -1730 10123 -1729
rect 9867 -1985 9931 -1730
rect 9866 -1986 9932 -1985
rect 9866 -2050 9867 -1986
rect 9931 -2050 9932 -1986
rect 9866 -2051 9932 -2050
rect 9865 -2316 9931 -2315
rect 9865 -2380 9866 -2316
rect 9930 -2380 9931 -2316
rect 9865 -2381 9931 -2380
rect 9866 -2648 9930 -2381
rect 7441 -2649 8323 -2648
rect 7441 -3529 7442 -2649
rect 8322 -3529 8323 -2649
rect 9241 -2649 10123 -2648
rect 9241 -3420 9242 -2649
rect 7441 -3530 8323 -3529
rect 8738 -3484 9242 -3420
rect 7441 -4449 8323 -4448
rect 7441 -5329 7442 -4449
rect 8322 -5329 8323 -4449
rect 7441 -5330 8323 -5329
rect 7441 -6249 8323 -6248
rect 7441 -7129 7442 -6249
rect 8322 -7129 8323 -6249
rect 8738 -6542 8802 -3484
rect 9241 -3529 9242 -3484
rect 10122 -3529 10123 -2649
rect 9241 -3530 10123 -3529
rect 10032 -4127 10096 -3530
rect 10031 -4128 10097 -4127
rect 10031 -4192 10032 -4128
rect 10096 -4192 10097 -4128
rect 10031 -4193 10097 -4192
rect 9241 -4449 10123 -4448
rect 9241 -5329 9242 -4449
rect 10122 -4610 10123 -4449
rect 10344 -4610 10408 -605
rect 13185 -606 13251 -605
rect 11041 -849 11923 -848
rect 11041 -1729 11042 -849
rect 11922 -906 11923 -849
rect 12841 -849 13723 -848
rect 12207 -906 12273 -905
rect 11922 -970 12208 -906
rect 12272 -970 12273 -906
rect 11922 -1729 11923 -970
rect 12207 -971 12273 -970
rect 12407 -1607 12473 -1606
rect 12841 -1607 12842 -849
rect 12407 -1671 12408 -1607
rect 12472 -1671 12842 -1607
rect 12407 -1672 12473 -1671
rect 11041 -1730 11923 -1729
rect 12841 -1729 12842 -1671
rect 13722 -1729 13723 -849
rect 13977 -1489 14043 -1488
rect 13977 -1553 13978 -1489
rect 14042 -1553 14043 -1489
rect 13977 -1554 14043 -1553
rect 12841 -1730 13723 -1729
rect 10509 -1986 10575 -1985
rect 10509 -2050 10510 -1986
rect 10574 -2050 10575 -1986
rect 10509 -2051 10575 -2050
rect 11450 -2037 11514 -1730
rect 13612 -2006 13676 -1730
rect 13611 -2007 13677 -2006
rect 10122 -4674 10408 -4610
rect 10510 -4656 10574 -2051
rect 11450 -2101 13014 -2037
rect 13611 -2071 13612 -2007
rect 13676 -2071 13677 -2007
rect 13611 -2072 13677 -2071
rect 12950 -2648 13014 -2101
rect 13609 -2318 13675 -2317
rect 13609 -2382 13610 -2318
rect 13674 -2382 13675 -2318
rect 13609 -2383 13675 -2382
rect 13610 -2648 13674 -2383
rect 11041 -2649 11923 -2648
rect 11041 -3529 11042 -2649
rect 11922 -2846 11923 -2649
rect 12841 -2649 13723 -2648
rect 12407 -2846 12473 -2845
rect 11922 -2910 12408 -2846
rect 12472 -2910 12473 -2846
rect 11922 -3529 11923 -2910
rect 12407 -2911 12473 -2910
rect 11041 -3530 11923 -3529
rect 12841 -3529 12842 -2649
rect 13722 -3529 13723 -2649
rect 12841 -3530 13723 -3529
rect 11432 -3828 11496 -3530
rect 11431 -3829 11497 -3828
rect 11431 -3893 11432 -3829
rect 11496 -3893 11497 -3829
rect 11431 -3894 11497 -3893
rect 12995 -3947 13061 -3946
rect 12185 -4011 12996 -3947
rect 13060 -4011 13061 -3947
rect 11041 -4449 11923 -4448
rect 11041 -4656 11042 -4449
rect 10122 -5329 10123 -4674
rect 10510 -4720 11042 -4656
rect 10524 -5120 10590 -5119
rect 11041 -5120 11042 -4720
rect 10522 -5184 10525 -5120
rect 10589 -5184 11042 -5120
rect 10524 -5185 10590 -5184
rect 9241 -5330 10123 -5329
rect 11041 -5329 11042 -5184
rect 11922 -4657 11923 -4449
rect 12185 -4657 12249 -4011
rect 12995 -4012 13061 -4011
rect 13045 -4127 13109 -4124
rect 13044 -4128 13110 -4127
rect 13044 -4192 13045 -4128
rect 13109 -4192 13110 -4128
rect 13044 -4193 13110 -4192
rect 13045 -4448 13109 -4193
rect 11922 -4721 12249 -4657
rect 12841 -4449 13723 -4448
rect 11922 -5329 11923 -4721
rect 11041 -5330 11923 -5329
rect 12841 -5329 12842 -4449
rect 13722 -4625 13723 -4449
rect 13978 -4625 14042 -1554
rect 13722 -4689 14042 -4625
rect 13722 -5329 13723 -4689
rect 14143 -4853 14207 -222
rect 14808 -540 14872 70
rect 14807 -541 14873 -540
rect 14807 -605 14808 -541
rect 14872 -605 14873 -541
rect 14807 -606 14873 -605
rect 14641 -849 15523 -848
rect 14307 -1489 14373 -1488
rect 14641 -1489 14642 -849
rect 14307 -1553 14308 -1489
rect 14372 -1553 14642 -1489
rect 14307 -1554 14373 -1553
rect 14641 -1729 14642 -1553
rect 15522 -1729 15523 -849
rect 14641 -1730 15523 -1729
rect 16441 -849 17323 -848
rect 16441 -1729 16442 -849
rect 17322 -1729 17323 -849
rect 16441 -1730 17323 -1729
rect 14641 -2649 15523 -2648
rect 14641 -3529 14642 -2649
rect 15522 -3529 15523 -2649
rect 14641 -3530 15523 -3529
rect 16441 -2649 17323 -2648
rect 16441 -3529 16442 -2649
rect 17322 -3529 17323 -2649
rect 16441 -3530 17323 -3529
rect 14838 -3946 14902 -3530
rect 14837 -3947 14903 -3946
rect 14837 -4011 14838 -3947
rect 14902 -4011 14903 -3947
rect 14837 -4012 14903 -4011
rect 14641 -4449 15523 -4448
rect 14641 -4853 14642 -4449
rect 14143 -4917 14642 -4853
rect 12841 -5330 13723 -5329
rect 14641 -5329 14642 -4917
rect 15522 -4976 15523 -4449
rect 16441 -4449 17323 -4448
rect 15801 -4976 15867 -4975
rect 15522 -5040 15802 -4976
rect 15866 -5040 15868 -4976
rect 15522 -5329 15523 -5040
rect 15801 -5041 15867 -5040
rect 14641 -5330 15523 -5329
rect 16441 -5329 16442 -4449
rect 17322 -5329 17323 -4449
rect 16441 -5330 17323 -5329
rect 9262 -5686 9326 -5330
rect 9261 -5687 9327 -5686
rect 9261 -5751 9262 -5687
rect 9326 -5751 9327 -5687
rect 9261 -5752 9327 -5751
rect 9241 -6249 10123 -6248
rect 8737 -6543 8803 -6542
rect 8737 -6607 8738 -6543
rect 8802 -6607 8803 -6543
rect 8737 -6608 8803 -6607
rect 7441 -7130 8323 -7129
rect 9241 -7129 9242 -6249
rect 10122 -7129 10123 -6249
rect 9241 -7130 10123 -7129
rect 11041 -6249 11923 -6248
rect 11041 -7129 11042 -6249
rect 11922 -7129 11923 -6249
rect 11041 -7130 11923 -7129
rect 12841 -6249 13723 -6248
rect 12841 -7129 12842 -6249
rect 13722 -7129 13723 -6249
rect 12841 -7130 13723 -7129
rect 14641 -6249 15523 -6248
rect 14641 -7129 14642 -6249
rect 15522 -7129 15523 -6249
rect 14641 -7130 15523 -7129
rect 16441 -6249 17323 -6248
rect 16441 -7129 16442 -6249
rect 17322 -7129 17323 -6249
rect 16441 -7130 17323 -7129
<< labels >>
flabel metal2 3147 -3484 3147 -3484 1 FreeSans 1200 0 0 0 on
port 8 n
flabel metal2 3431 -5243 3431 -5243 1 FreeSans 1200 0 0 0 op
port 7 n
flabel metal2 5049 -9956 5049 -9956 1 FreeSans 1200 0 0 0 cmc
flabel metal1 4262 -15741 4262 -15741 1 FreeSans 1200 0 0 0 bias_a
flabel metal1 6929 -13167 6929 -13167 1 FreeSans 1200 0 0 0 bias_d
flabel metal1 -7420 -1403 -7420 -1403 1 FreeSans 1200 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 -7407 -17402 -7407 -17402 1 FreeSans 1200 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 -6957 -14245 -6957 -14245 1 FreeSans 1200 0 0 0 i_bias
port 9 n
flabel metal1 -3636 -12323 -3636 -12323 1 FreeSans 1200 0 0 0 bias_c
flabel metal1 -6950 -12541 -6950 -12541 1 FreeSans 1200 0 0 0 ip
port 1 n
flabel metal1 -6952 -13880 -6952 -13880 1 FreeSans 1200 0 0 0 in
port 2 n
flabel metal1 -4277 -7715 -4277 -7715 1 FreeSans 1200 0 0 0 bias_b
flabel viali 10071 -9280 10071 -9280 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali 10071 -11280 10071 -11280 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali 11526 -12643 11526 -12643 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali 8526 -12643 8526 -12643 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali 5775 -11240 5775 -11240 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali -2896 -9365 -2896 -9365 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali -2896 -11365 -2896 -11365 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali -2896 -13365 -2896 -13365 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali -2896 -15365 -2896 -15365 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali 4632 -14958 4632 -14958 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel viali -2097 -3132 -2097 -3132 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel viali -2945 -5751 -2945 -5751 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 7057 2874 7057 2874 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 7057 1707 7057 1707 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 7058 -83 7058 -83 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 7058 -739 7058 -739 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 7058 -1885 7058 -1885 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 7058 -2537 7058 -2537 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 7051 -4329 7051 -4329 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 7054 -5489 7054 -5489 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 7054 -7288 7054 -7288 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16056 -7290 16056 -7290 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16057 -6136 16057 -6136 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 16055 -5482 16055 -5482 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16057 -2529 16057 -2529 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 16055 -1886 16055 -1886 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16057 -86 16057 -86 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16057 1070 16057 1070 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 16057 1716 16057 1716 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16057 2870 16057 2870 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal3 6479 2585 6479 2585 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal3 6738 1807 6738 1807 1 FreeSans 400 0 0 0 p2
port 5 n
flabel metal3 6486 -6211 6486 -6211 1 FreeSans 400 0 0 0 p1_b
port 4 n
flabel metal3 6735 -5207 6735 -5207 1 FreeSans 400 0 0 0 p1
port 3 n
flabel metal3 17730 1821 17730 1821 1 FreeSans 400 0 0 0 p2
port 5 n
flabel metal3 17980 2631 17980 2631 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal3 17727 -7023 17727 -7023 1 FreeSans 400 0 0 0 p1
port 3 n
flabel metal3 17984 -6236 17984 -6236 1 FreeSans 400 0 0 0 p1_b
port 4 n
flabel metal2 17862 -8732 17862 -8732 1 FreeSans 800 0 0 0 cm
port 10 n
flabel metal1 7058 1058 7058 1058 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 7058 -3672 7058 -3672 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 7058 -6144 7058 -6144 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 16056 -4338 16056 -4338 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal1 16056 -3678 16056 -3678 1 FreeSans 400 0 0 0 VSS
port 12 n power bidirectional
flabel metal1 16056 -738 16056 -738 1 FreeSans 400 0 0 0 VDD
port 11 n power bidirectional
flabel metal3 6460 2550 6460 2550 1 FreeSans 400 0 0 0 sc_cmfb_0/p2_b
flabel metal3 6713 1767 6713 1767 1 FreeSans 400 0 0 0 sc_cmfb_0/p2
flabel metal3 6463 -2843 6463 -2843 1 FreeSans 400 0 0 0 sc_cmfb_0/p1_b
flabel metal3 6713 -3629 6713 -3629 1 FreeSans 400 0 0 0 sc_cmfb_0/p1
flabel metal3 17747 -7006 17747 -7006 1 FreeSans 400 0 0 0 sc_cmfb_0/p1
flabel metal3 18000 -6139 18000 -6139 1 FreeSans 400 0 0 0 sc_cmfb_0/p1_b
flabel metal3 17750 1777 17750 1777 1 FreeSans 400 0 0 0 sc_cmfb_0/p2
flabel metal3 18006 2547 18006 2547 1 FreeSans 400 0 0 0 sc_cmfb_0/p2_b
flabel metal1 5618 -2100 5618 -2100 1 FreeSans 400 0 0 0 sc_cmfb_0/op
flabel metal1 6230 -2101 6230 -2101 1 FreeSans 400 0 0 0 sc_cmfb_0/on
flabel metal1 6690 -2098 6690 -2098 1 FreeSans 400 0 0 0 sc_cmfb_0/cmc
flabel metal1 17892 -2174 17892 -2174 1 FreeSans 400 0 0 0 sc_cmfb_0/cm
flabel metal1 18394 -2171 18394 -2171 1 FreeSans 400 0 0 0 sc_cmfb_0/bias_a
flabel metal1 7056 2881 7056 2881 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 7057 1709 7057 1709 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 7059 1074 7059 1074 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 7057 -99 7057 -99 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 7059 -726 7059 -726 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 7055 -1895 7055 -1895 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 7055 -2527 7055 -2527 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 7057 -3693 7057 -3693 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 7059 -4323 7059 -4323 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 7055 -5496 7055 -5496 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 7057 -6128 7057 -6128 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 7057 -7291 7057 -7291 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16059 -7291 16059 -7291 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16056 -6128 16056 -6128 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 16059 -5495 16059 -5495 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16054 -4328 16054 -4328 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 16054 -3693 16054 -3693 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16056 -2525 16056 -2525 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 16056 -1890 16056 -1890 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16059 -729 16059 -729 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 16056 -94 16056 -94 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16054 1078 16054 1078 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 16056 1711 16056 1711 1 FreeSans 400 0 0 0 sc_cmfb_0/VSS
flabel metal1 16056 2876 16056 2876 1 FreeSans 400 0 0 0 sc_cmfb_0/VDD
flabel metal1 8456 -6309 8456 -6309 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/en_b
flabel metal1 8457 -6805 8457 -6805 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/in
flabel metal1 8457 -7116 8457 -7116 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/en
flabel metal1 6966 -6806 6966 -6806 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/out
flabel metal1 7057 -6160 7057 -6160 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/VDD
flabel metal1 7057 -7266 7057 -7266 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_11/VSS
flabel metal1 17456 -6309 17456 -6309 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/en_b
flabel metal1 17457 -6805 17457 -6805 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/in
flabel metal1 17457 -7116 17457 -7116 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/en
flabel metal1 15966 -6806 15966 -6806 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/out
flabel metal1 16057 -6160 16057 -6160 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/VDD
flabel metal1 16057 -7266 16057 -7266 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_2/VSS
flabel metal1 8456 -4509 8456 -4509 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/en_b
flabel metal1 8457 -5005 8457 -5005 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/in
flabel metal1 8457 -5316 8457 -5316 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/en
flabel metal1 6966 -5006 6966 -5006 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/out
flabel metal1 7057 -4360 7057 -4360 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/VDD
flabel metal1 7057 -5466 7057 -5466 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_10/VSS
flabel metal1 17456 -4509 17456 -4509 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/en_b
flabel metal1 17457 -5005 17457 -5005 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/in
flabel metal1 17457 -5316 17457 -5316 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/en
flabel metal1 15966 -5006 15966 -5006 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/out
flabel metal1 16057 -4360 16057 -4360 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/VDD
flabel metal1 16057 -5466 16057 -5466 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_0/VSS
flabel metal1 8456 -2709 8456 -2709 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/en_b
flabel metal1 8457 -3205 8457 -3205 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/in
flabel metal1 8457 -3516 8457 -3516 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/en
flabel metal1 6966 -3206 6966 -3206 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/out
flabel metal1 7057 -2560 7057 -2560 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/VDD
flabel metal1 7057 -3666 7057 -3666 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_9/VSS
flabel metal1 17456 -2709 17456 -2709 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/en_b
flabel metal1 17457 -3205 17457 -3205 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/in
flabel metal1 17457 -3516 17457 -3516 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/en
flabel metal1 15966 -3206 15966 -3206 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/out
flabel metal1 16057 -2560 16057 -2560 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/VDD
flabel metal1 16057 -3666 16057 -3666 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_1/VSS
flabel metal1 8456 -909 8456 -909 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/en_b
flabel metal1 8457 -1405 8457 -1405 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/in
flabel metal1 8457 -1716 8457 -1716 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/en
flabel metal1 6966 -1406 6966 -1406 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/out
flabel metal1 7057 -760 7057 -760 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/VDD
flabel metal1 7057 -1866 7057 -1866 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_8/VSS
flabel metal1 17456 -909 17456 -909 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/en_b
flabel metal1 17457 -1405 17457 -1405 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/in
flabel metal1 17457 -1716 17457 -1716 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/en
flabel metal1 15966 -1406 15966 -1406 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/out
flabel metal1 16057 -760 16057 -760 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/VDD
flabel metal1 16057 -1866 16057 -1866 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_3/VSS
flabel metal1 8456 891 8456 891 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/en_b
flabel metal1 8457 395 8457 395 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/in
flabel metal1 8457 84 8457 84 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/en
flabel metal1 6966 394 6966 394 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/out
flabel metal1 7057 1040 7057 1040 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/VDD
flabel metal1 7057 -66 7057 -66 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_7/VSS
flabel metal1 17456 891 17456 891 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/en_b
flabel metal1 17457 395 17457 395 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/in
flabel metal1 17457 84 17457 84 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/en
flabel metal1 15966 394 15966 394 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/out
flabel metal1 16057 1040 16057 1040 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/VDD
flabel metal1 16057 -66 16057 -66 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_4/VSS
flabel metal1 8456 2691 8456 2691 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/en_b
flabel metal1 8457 2195 8457 2195 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/in
flabel metal1 8457 1884 8457 1884 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/en
flabel metal1 6966 2194 6966 2194 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/out
flabel metal1 7057 2840 7057 2840 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/VDD
flabel metal1 7057 1734 7057 1734 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_6/VSS
flabel metal1 17456 2691 17456 2691 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/en_b
flabel metal1 17457 2195 17457 2195 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/in
flabel metal1 17457 1884 17457 1884 7 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/en
flabel metal1 15966 2194 15966 2194 3 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/out
flabel metal1 16057 2840 16057 2840 5 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/VDD
flabel metal1 16057 1734 16057 1734 1 FreeSans 400 0 0 0 sc_cmfb_0/transmission_gate_5/VSS
<< end >>
