magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< error_p >>
rect -749 181 -691 187
rect -557 181 -499 187
rect -365 181 -307 187
rect -173 181 -115 187
rect 19 181 77 187
rect 211 181 269 187
rect 403 181 461 187
rect 595 181 653 187
rect -749 147 -737 181
rect -557 147 -545 181
rect -365 147 -353 181
rect -173 147 -161 181
rect 19 147 31 181
rect 211 147 223 181
rect 403 147 415 181
rect 595 147 607 181
rect -749 141 -691 147
rect -557 141 -499 147
rect -365 141 -307 147
rect -173 141 -115 147
rect 19 141 77 147
rect 211 141 269 147
rect 403 141 461 147
rect 595 141 653 147
rect -653 -147 -595 -141
rect -461 -147 -403 -141
rect -269 -147 -211 -141
rect -77 -147 -19 -141
rect 115 -147 173 -141
rect 307 -147 365 -141
rect 499 -147 557 -141
rect 691 -147 749 -141
rect -653 -181 -641 -147
rect -461 -181 -449 -147
rect -269 -181 -257 -147
rect -77 -181 -65 -147
rect 115 -181 127 -147
rect 307 -181 319 -147
rect 499 -181 511 -147
rect 691 -181 703 -147
rect -653 -187 -595 -181
rect -461 -187 -403 -181
rect -269 -187 -211 -181
rect -77 -187 -19 -181
rect 115 -187 173 -181
rect 307 -187 365 -181
rect 499 -187 557 -181
rect 691 -187 749 -181
<< nwell >>
rect -1031 -319 1031 319
<< pmos >>
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
<< pdiff >>
rect -893 85 -831 100
rect -893 51 -881 85
rect -847 51 -831 85
rect -893 17 -831 51
rect -893 -17 -881 17
rect -847 -17 -831 17
rect -893 -51 -831 -17
rect -893 -85 -881 -51
rect -847 -85 -831 -51
rect -893 -100 -831 -85
rect -801 85 -735 100
rect -801 51 -785 85
rect -751 51 -735 85
rect -801 17 -735 51
rect -801 -17 -785 17
rect -751 -17 -735 17
rect -801 -51 -735 -17
rect -801 -85 -785 -51
rect -751 -85 -735 -51
rect -801 -100 -735 -85
rect -705 85 -639 100
rect -705 51 -689 85
rect -655 51 -639 85
rect -705 17 -639 51
rect -705 -17 -689 17
rect -655 -17 -639 17
rect -705 -51 -639 -17
rect -705 -85 -689 -51
rect -655 -85 -639 -51
rect -705 -100 -639 -85
rect -609 85 -543 100
rect -609 51 -593 85
rect -559 51 -543 85
rect -609 17 -543 51
rect -609 -17 -593 17
rect -559 -17 -543 17
rect -609 -51 -543 -17
rect -609 -85 -593 -51
rect -559 -85 -543 -51
rect -609 -100 -543 -85
rect -513 85 -447 100
rect -513 51 -497 85
rect -463 51 -447 85
rect -513 17 -447 51
rect -513 -17 -497 17
rect -463 -17 -447 17
rect -513 -51 -447 -17
rect -513 -85 -497 -51
rect -463 -85 -447 -51
rect -513 -100 -447 -85
rect -417 85 -351 100
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -100 -351 -85
rect -321 85 -255 100
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -100 -255 -85
rect -225 85 -159 100
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 225 100
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -100 225 -85
rect 255 85 321 100
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -100 321 -85
rect 351 85 417 100
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -100 417 -85
rect 447 85 513 100
rect 447 51 463 85
rect 497 51 513 85
rect 447 17 513 51
rect 447 -17 463 17
rect 497 -17 513 17
rect 447 -51 513 -17
rect 447 -85 463 -51
rect 497 -85 513 -51
rect 447 -100 513 -85
rect 543 85 609 100
rect 543 51 559 85
rect 593 51 609 85
rect 543 17 609 51
rect 543 -17 559 17
rect 593 -17 609 17
rect 543 -51 609 -17
rect 543 -85 559 -51
rect 593 -85 609 -51
rect 543 -100 609 -85
rect 639 85 705 100
rect 639 51 655 85
rect 689 51 705 85
rect 639 17 705 51
rect 639 -17 655 17
rect 689 -17 705 17
rect 639 -51 705 -17
rect 639 -85 655 -51
rect 689 -85 705 -51
rect 639 -100 705 -85
rect 735 85 801 100
rect 735 51 751 85
rect 785 51 801 85
rect 735 17 801 51
rect 735 -17 751 17
rect 785 -17 801 17
rect 735 -51 801 -17
rect 735 -85 751 -51
rect 785 -85 801 -51
rect 735 -100 801 -85
rect 831 85 893 100
rect 831 51 847 85
rect 881 51 893 85
rect 831 17 893 51
rect 831 -17 847 17
rect 881 -17 893 17
rect 831 -51 893 -17
rect 831 -85 847 -51
rect 881 -85 893 -51
rect 831 -100 893 -85
<< pdiffc >>
rect -881 51 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -51
rect -785 51 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -51
rect -689 51 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -51
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
rect 655 51 689 85
rect 655 -17 689 17
rect 655 -85 689 -51
rect 751 51 785 85
rect 751 -17 785 17
rect 751 -85 785 -51
rect 847 51 881 85
rect 847 -17 881 17
rect 847 -85 881 -51
<< nsubdiff >>
rect -995 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 995 283
rect -995 187 -961 249
rect -995 119 -961 153
rect 961 187 995 249
rect 961 119 995 153
rect -995 51 -961 85
rect -995 -17 -961 17
rect -995 -85 -961 -51
rect 961 51 995 85
rect 961 -17 995 17
rect 961 -85 995 -51
rect -995 -153 -961 -119
rect -995 -249 -961 -187
rect 961 -153 995 -119
rect 961 -249 995 -187
rect -995 -283 -867 -249
rect -833 -283 -799 -249
rect -765 -283 -731 -249
rect -697 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 697 -249
rect 731 -283 765 -249
rect 799 -283 833 -249
rect 867 -283 995 -249
<< nsubdiffcont >>
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect -995 153 -961 187
rect 961 153 995 187
rect -995 85 -961 119
rect -995 17 -961 51
rect -995 -51 -961 -17
rect -995 -119 -961 -85
rect 961 85 995 119
rect 961 17 995 51
rect 961 -51 995 -17
rect 961 -119 995 -85
rect -995 -187 -961 -153
rect 961 -187 995 -153
rect -867 -283 -833 -249
rect -799 -283 -765 -249
rect -731 -283 -697 -249
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
rect 697 -283 731 -249
rect 765 -283 799 -249
rect 833 -283 867 -249
<< poly >>
rect -753 181 -687 197
rect -753 147 -737 181
rect -703 147 -687 181
rect -753 131 -687 147
rect -561 181 -495 197
rect -561 147 -545 181
rect -511 147 -495 181
rect -561 131 -495 147
rect -369 181 -303 197
rect -369 147 -353 181
rect -319 147 -303 181
rect -369 131 -303 147
rect -177 181 -111 197
rect -177 147 -161 181
rect -127 147 -111 181
rect -177 131 -111 147
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect 207 181 273 197
rect 207 147 223 181
rect 257 147 273 181
rect 207 131 273 147
rect 399 181 465 197
rect 399 147 415 181
rect 449 147 465 181
rect 399 131 465 147
rect 591 181 657 197
rect 591 147 607 181
rect 641 147 657 181
rect 591 131 657 147
rect 783 181 849 197
rect 783 147 799 181
rect 833 147 849 181
rect 783 131 849 147
rect -831 100 -801 127
rect -735 100 -705 131
rect -639 100 -609 127
rect -543 100 -513 131
rect -447 100 -417 127
rect -351 100 -321 131
rect -255 100 -225 127
rect -159 100 -129 131
rect -63 100 -33 127
rect 33 100 63 131
rect 129 100 159 127
rect 225 100 255 131
rect 321 100 351 127
rect 417 100 447 131
rect 513 100 543 127
rect 609 100 639 131
rect 705 100 735 127
rect 801 100 831 131
rect -831 -131 -801 -100
rect -735 -127 -705 -100
rect -639 -131 -609 -100
rect -543 -127 -513 -100
rect -447 -131 -417 -100
rect -351 -127 -321 -100
rect -255 -131 -225 -100
rect -159 -127 -129 -100
rect -63 -131 -33 -100
rect 33 -127 63 -100
rect 129 -131 159 -100
rect 225 -127 255 -100
rect 321 -131 351 -100
rect 417 -127 447 -100
rect 513 -131 543 -100
rect 609 -127 639 -100
rect 705 -131 735 -100
rect 801 -127 831 -100
rect -849 -147 -783 -131
rect -849 -181 -833 -147
rect -799 -181 -783 -147
rect -849 -197 -783 -181
rect -657 -147 -591 -131
rect -657 -181 -641 -147
rect -607 -181 -591 -147
rect -657 -197 -591 -181
rect -465 -147 -399 -131
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -465 -197 -399 -181
rect -273 -147 -207 -131
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -273 -197 -207 -181
rect -81 -147 -15 -131
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect -81 -197 -15 -181
rect 111 -147 177 -131
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 111 -197 177 -181
rect 303 -147 369 -131
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 303 -197 369 -181
rect 495 -147 561 -131
rect 495 -181 511 -147
rect 545 -181 561 -147
rect 495 -197 561 -181
rect 687 -147 753 -131
rect 687 -181 703 -147
rect 737 -181 753 -147
rect 687 -197 753 -181
<< polycont >>
rect -737 147 -703 181
rect -545 147 -511 181
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect 607 147 641 181
rect 799 147 833 181
rect -833 -181 -799 -147
rect -641 -181 -607 -147
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
rect 511 -181 545 -147
rect 703 -181 737 -147
<< locali >>
rect -995 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 995 283
rect -995 187 -961 249
rect 847 181 881 249
rect -995 119 -961 153
rect -753 147 -737 181
rect -703 147 -687 181
rect -561 147 -545 181
rect -511 147 -495 181
rect -369 147 -353 181
rect -319 147 -303 181
rect -177 147 -161 181
rect -127 147 -111 181
rect 15 147 31 181
rect 65 147 81 181
rect 207 147 223 181
rect 257 147 273 181
rect 399 147 415 181
rect 449 147 465 181
rect 591 147 607 181
rect 641 147 657 181
rect 783 147 799 181
rect 833 147 881 181
rect -995 51 -961 85
rect -995 -17 -961 17
rect -995 -85 -961 -51
rect -995 -153 -961 -119
rect -995 -249 -961 -187
rect -881 85 -847 104
rect -881 17 -847 51
rect -881 -51 -847 -17
rect -881 -147 -847 -85
rect -785 85 -751 104
rect -785 17 -751 51
rect -785 -51 -751 -17
rect -785 -104 -751 -85
rect -689 85 -655 104
rect -689 17 -655 51
rect -689 -51 -655 -17
rect -689 -104 -655 -85
rect -593 85 -559 104
rect -593 17 -559 51
rect -593 -51 -559 -17
rect -593 -104 -559 -85
rect -497 85 -463 104
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -104 -463 -85
rect -401 85 -367 104
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -104 -367 -85
rect -305 85 -271 104
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -104 -271 -85
rect -209 85 -175 104
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -104 209 -85
rect 271 85 305 104
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -104 305 -85
rect 367 85 401 104
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -104 401 -85
rect 463 85 497 104
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -104 497 -85
rect 559 85 593 104
rect 559 17 593 51
rect 559 -51 593 -17
rect 559 -104 593 -85
rect 655 85 689 104
rect 655 17 689 51
rect 655 -51 689 -17
rect 655 -104 689 -85
rect 751 85 785 104
rect 751 17 785 51
rect 751 -51 785 -17
rect 751 -104 785 -85
rect 847 85 881 147
rect 847 17 881 51
rect 847 -51 881 -17
rect 847 -104 881 -85
rect 961 187 995 249
rect 961 119 995 153
rect 961 51 995 85
rect 961 -17 995 17
rect 961 -85 995 -51
rect -881 -181 -833 -147
rect -799 -181 -783 -147
rect -657 -181 -641 -147
rect -607 -181 -591 -147
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 495 -181 511 -147
rect 545 -181 561 -147
rect 687 -181 703 -147
rect 737 -181 753 -147
rect 961 -153 995 -119
rect -881 -249 -847 -181
rect 961 -249 995 -187
rect -995 -283 -867 -249
rect -833 -283 -799 -249
rect -765 -283 -731 -249
rect -697 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 697 -249
rect 731 -283 765 -249
rect 799 -283 833 -249
rect 867 -283 995 -249
<< viali >>
rect -737 147 -703 181
rect -545 147 -511 181
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect 607 147 641 181
rect -641 -181 -607 -147
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
rect 511 -181 545 -147
rect 703 -181 737 -147
<< metal1 >>
rect -749 181 -691 187
rect -749 147 -737 181
rect -703 147 -691 181
rect -749 141 -691 147
rect -557 181 -499 187
rect -557 147 -545 181
rect -511 147 -499 181
rect -557 141 -499 147
rect -365 181 -307 187
rect -365 147 -353 181
rect -319 147 -307 181
rect -365 141 -307 147
rect -173 181 -115 187
rect -173 147 -161 181
rect -127 147 -115 181
rect -173 141 -115 147
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect 211 181 269 187
rect 211 147 223 181
rect 257 147 269 181
rect 211 141 269 147
rect 403 181 461 187
rect 403 147 415 181
rect 449 147 461 181
rect 403 141 461 147
rect 595 181 653 187
rect 595 147 607 181
rect 641 147 653 181
rect 595 141 653 147
rect -653 -147 -595 -141
rect -653 -181 -641 -147
rect -607 -181 -595 -147
rect -653 -187 -595 -181
rect -461 -147 -403 -141
rect -461 -181 -449 -147
rect -415 -181 -403 -147
rect -461 -187 -403 -181
rect -269 -147 -211 -141
rect -269 -181 -257 -147
rect -223 -181 -211 -147
rect -269 -187 -211 -181
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
rect 115 -147 173 -141
rect 115 -181 127 -147
rect 161 -181 173 -147
rect 115 -187 173 -181
rect 307 -147 365 -141
rect 307 -181 319 -147
rect 353 -181 365 -147
rect 307 -187 365 -181
rect 499 -147 557 -141
rect 499 -181 511 -147
rect 545 -181 557 -147
rect 499 -187 557 -181
rect 691 -147 749 -141
rect 691 -181 703 -147
rect 737 -181 749 -147
rect 691 -187 749 -181
<< properties >>
string FIXED_BBOX -978 -266 978 266
<< end >>
