magic
tech sky130A
magscale 1 2
timestamp 1654720150
<< nmos >>
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
<< ndiff >>
rect -1008 128 -950 140
rect -1008 -128 -996 128
rect -962 -128 -950 128
rect -1008 -140 -950 -128
rect -830 128 -772 140
rect -830 -128 -818 128
rect -784 -128 -772 128
rect -830 -140 -772 -128
rect -652 128 -594 140
rect -652 -128 -640 128
rect -606 -128 -594 128
rect -652 -140 -594 -128
rect -474 128 -416 140
rect -474 -128 -462 128
rect -428 -128 -416 128
rect -474 -140 -416 -128
rect -296 128 -238 140
rect -296 -128 -284 128
rect -250 -128 -238 128
rect -296 -140 -238 -128
rect -118 128 -60 140
rect -118 -128 -106 128
rect -72 -128 -60 128
rect -118 -140 -60 -128
rect 60 128 118 140
rect 60 -128 72 128
rect 106 -128 118 128
rect 60 -140 118 -128
rect 238 128 296 140
rect 238 -128 250 128
rect 284 -128 296 128
rect 238 -140 296 -128
rect 416 128 474 140
rect 416 -128 428 128
rect 462 -128 474 128
rect 416 -140 474 -128
rect 594 128 652 140
rect 594 -128 606 128
rect 640 -128 652 128
rect 594 -140 652 -128
rect 772 128 830 140
rect 772 -128 784 128
rect 818 -128 830 128
rect 772 -140 830 -128
rect 950 128 1008 140
rect 950 -128 962 128
rect 996 -128 1008 128
rect 950 -140 1008 -128
<< ndiffc >>
rect -996 -128 -962 128
rect -818 -128 -784 128
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect 784 -128 818 128
rect 962 -128 996 128
<< poly >>
rect -932 212 -848 228
rect -932 195 -916 212
rect -950 178 -916 195
rect -864 195 -848 212
rect -754 212 -670 228
rect -754 195 -738 212
rect -864 178 -830 195
rect -950 140 -830 178
rect -772 178 -738 195
rect -686 195 -670 212
rect -576 212 -492 228
rect -576 195 -560 212
rect -686 178 -652 195
rect -772 140 -652 178
rect -594 178 -560 195
rect -508 195 -492 212
rect -398 212 -314 228
rect -398 195 -382 212
rect -508 178 -474 195
rect -594 140 -474 178
rect -416 178 -382 195
rect -330 195 -314 212
rect -220 212 -136 228
rect -220 195 -204 212
rect -330 178 -296 195
rect -416 140 -296 178
rect -238 178 -204 195
rect -152 195 -136 212
rect -42 212 42 228
rect -42 195 -26 212
rect -152 178 -118 195
rect -238 140 -118 178
rect -60 178 -26 195
rect 26 195 42 212
rect 136 212 220 228
rect 136 195 152 212
rect 26 178 60 195
rect -60 140 60 178
rect 118 178 152 195
rect 204 195 220 212
rect 314 212 398 228
rect 314 195 330 212
rect 204 178 238 195
rect 118 140 238 178
rect 296 178 330 195
rect 382 195 398 212
rect 492 212 576 228
rect 492 195 508 212
rect 382 178 416 195
rect 296 140 416 178
rect 474 178 508 195
rect 560 195 576 212
rect 670 212 754 228
rect 670 195 686 212
rect 560 178 594 195
rect 474 140 594 178
rect 652 178 686 195
rect 738 195 754 212
rect 848 212 932 228
rect 848 195 864 212
rect 738 178 772 195
rect 652 140 772 178
rect 830 178 864 195
rect 916 195 932 212
rect 916 178 950 195
rect 830 140 950 178
rect -950 -178 -830 -140
rect -950 -195 -916 -178
rect -932 -212 -916 -195
rect -864 -195 -830 -178
rect -772 -178 -652 -140
rect -772 -195 -738 -178
rect -864 -212 -848 -195
rect -932 -228 -848 -212
rect -754 -212 -738 -195
rect -686 -195 -652 -178
rect -594 -178 -474 -140
rect -594 -195 -560 -178
rect -686 -212 -670 -195
rect -754 -228 -670 -212
rect -576 -212 -560 -195
rect -508 -195 -474 -178
rect -416 -178 -296 -140
rect -416 -195 -382 -178
rect -508 -212 -492 -195
rect -576 -228 -492 -212
rect -398 -212 -382 -195
rect -330 -195 -296 -178
rect -238 -178 -118 -140
rect -238 -195 -204 -178
rect -330 -212 -314 -195
rect -398 -228 -314 -212
rect -220 -212 -204 -195
rect -152 -195 -118 -178
rect -60 -178 60 -140
rect -60 -195 -26 -178
rect -152 -212 -136 -195
rect -220 -228 -136 -212
rect -42 -212 -26 -195
rect 26 -195 60 -178
rect 118 -178 238 -140
rect 118 -195 152 -178
rect 26 -212 42 -195
rect -42 -228 42 -212
rect 136 -212 152 -195
rect 204 -195 238 -178
rect 296 -178 416 -140
rect 296 -195 330 -178
rect 204 -212 220 -195
rect 136 -228 220 -212
rect 314 -212 330 -195
rect 382 -195 416 -178
rect 474 -178 594 -140
rect 474 -195 508 -178
rect 382 -212 398 -195
rect 314 -228 398 -212
rect 492 -212 508 -195
rect 560 -195 594 -178
rect 652 -178 772 -140
rect 652 -195 686 -178
rect 560 -212 576 -195
rect 492 -228 576 -212
rect 670 -212 686 -195
rect 738 -195 772 -178
rect 830 -178 950 -140
rect 830 -195 864 -178
rect 738 -212 754 -195
rect 670 -228 754 -212
rect 848 -212 864 -195
rect 916 -195 950 -178
rect 916 -212 932 -195
rect 848 -228 932 -212
<< polycont >>
rect -916 178 -864 212
rect -738 178 -686 212
rect -560 178 -508 212
rect -382 178 -330 212
rect -204 178 -152 212
rect -26 178 26 212
rect 152 178 204 212
rect 330 178 382 212
rect 508 178 560 212
rect 686 178 738 212
rect 864 178 916 212
rect -916 -212 -864 -178
rect -738 -212 -686 -178
rect -560 -212 -508 -178
rect -382 -212 -330 -178
rect -204 -212 -152 -178
rect -26 -212 26 -178
rect 152 -212 204 -178
rect 330 -212 382 -178
rect 508 -212 560 -178
rect 686 -212 738 -178
rect 864 -212 916 -178
<< locali >>
rect -996 178 -916 212
rect -864 178 -848 212
rect -754 178 -738 212
rect -686 178 -670 212
rect -576 178 -560 212
rect -508 178 -492 212
rect -398 178 -382 212
rect -330 178 -314 212
rect -220 178 -204 212
rect -152 178 -136 212
rect -42 178 -26 212
rect 26 178 42 212
rect 136 178 152 212
rect 204 178 220 212
rect 314 178 330 212
rect 382 178 398 212
rect 492 178 508 212
rect 560 178 576 212
rect 670 178 686 212
rect 738 178 754 212
rect 848 178 864 212
rect 916 178 996 212
rect -996 128 -962 178
rect -996 -178 -962 -128
rect -818 128 -784 144
rect -818 -144 -784 -128
rect -640 128 -606 144
rect -640 -144 -606 -128
rect -462 128 -428 144
rect -462 -144 -428 -128
rect -284 128 -250 144
rect -284 -144 -250 -128
rect -106 128 -72 144
rect -106 -144 -72 -128
rect 72 128 106 144
rect 72 -144 106 -128
rect 250 128 284 144
rect 250 -144 284 -128
rect 428 128 462 144
rect 428 -144 462 -128
rect 606 128 640 144
rect 606 -144 640 -128
rect 784 128 818 144
rect 784 -144 818 -128
rect 962 128 996 178
rect 962 -178 996 -128
rect -996 -212 -916 -178
rect -864 -212 -848 -178
rect -754 -212 -738 -178
rect -686 -212 -670 -178
rect -576 -212 -560 -178
rect -508 -212 -492 -178
rect -398 -212 -382 -178
rect -330 -212 -314 -178
rect -220 -212 -204 -178
rect -152 -212 -136 -178
rect -42 -212 -26 -178
rect 26 -212 42 -178
rect 136 -212 152 -178
rect 204 -212 220 -178
rect 314 -212 330 -178
rect 382 -212 398 -178
rect 492 -212 508 -178
rect 560 -212 576 -178
rect 670 -212 686 -178
rect 738 -212 754 -178
rect 848 -212 864 -178
rect 916 -212 996 -178
<< viali >>
rect -738 178 -686 212
rect -560 178 -508 212
rect -382 178 -330 212
rect -204 178 -152 212
rect -26 178 26 212
rect 152 178 204 212
rect 330 178 382 212
rect 508 178 560 212
rect 686 178 738 212
rect -738 -212 -686 -178
rect -560 -212 -508 -178
rect -382 -212 -330 -178
rect -204 -212 -152 -178
rect -26 -212 26 -178
rect 152 -212 204 -178
rect 330 -212 382 -178
rect 508 -212 560 -178
rect 686 -212 738 -178
<< metal1 >>
rect -750 212 -674 218
rect -750 178 -738 212
rect -686 178 -674 212
rect -750 172 -674 178
rect -572 212 -496 218
rect -572 178 -560 212
rect -508 178 -496 212
rect -572 172 -496 178
rect -394 212 -318 218
rect -394 178 -382 212
rect -330 178 -318 212
rect -394 172 -318 178
rect -216 212 -140 218
rect -216 178 -204 212
rect -152 178 -140 212
rect -216 172 -140 178
rect -38 212 38 218
rect -38 178 -26 212
rect 26 178 38 212
rect -38 172 38 178
rect 140 212 216 218
rect 140 178 152 212
rect 204 178 216 212
rect 140 172 216 178
rect 318 212 394 218
rect 318 178 330 212
rect 382 178 394 212
rect 318 172 394 178
rect 496 212 572 218
rect 496 178 508 212
rect 560 178 572 212
rect 496 172 572 178
rect 674 212 750 218
rect 674 178 686 212
rect 738 178 750 212
rect 674 172 750 178
rect -750 -178 -674 -172
rect -750 -212 -738 -178
rect -686 -212 -674 -178
rect -750 -218 -674 -212
rect -572 -178 -496 -172
rect -572 -212 -560 -178
rect -508 -212 -496 -178
rect -572 -218 -496 -212
rect -394 -178 -318 -172
rect -394 -212 -382 -178
rect -330 -212 -318 -178
rect -394 -218 -318 -212
rect -216 -178 -140 -172
rect -216 -212 -204 -178
rect -152 -212 -140 -178
rect -216 -218 -140 -212
rect -38 -178 38 -172
rect -38 -212 -26 -178
rect 26 -212 38 -178
rect -38 -218 38 -212
rect 140 -178 216 -172
rect 140 -212 152 -178
rect 204 -212 216 -178
rect 140 -218 216 -212
rect 318 -178 394 -172
rect 318 -212 330 -178
rect 382 -212 394 -178
rect 318 -218 394 -212
rect 496 -178 572 -172
rect 496 -212 508 -178
rect 560 -212 572 -178
rect 496 -218 572 -212
rect 674 -178 750 -172
rect 674 -212 686 -178
rect 738 -212 750 -178
rect 674 -218 750 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 11 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
