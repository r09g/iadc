magic
tech sky130A
magscale 1 2
timestamp 1652838679
<< nwell >>
rect 163 464 1457 1114
rect 157 -688 1451 -38
<< pwell >>
rect 163 0 1457 464
rect 157 -1152 1451 -688
<< nmos >>
rect 363 210 393 316
rect 459 210 489 316
rect 555 210 585 316
rect 651 210 681 316
rect 747 210 777 316
rect 843 210 873 316
rect 939 210 969 316
rect 1035 210 1065 316
rect 1131 210 1161 316
rect 1227 210 1257 316
rect 357 -942 387 -836
rect 453 -942 483 -836
rect 549 -942 579 -836
rect 645 -942 675 -836
rect 741 -942 771 -836
rect 837 -942 867 -836
rect 933 -942 963 -836
rect 1029 -942 1059 -836
rect 1125 -942 1155 -836
rect 1221 -942 1251 -836
<< pmos >>
rect 363 621 393 895
rect 459 621 489 895
rect 555 621 585 895
rect 651 621 681 895
rect 747 621 777 895
rect 843 621 873 895
rect 939 621 969 895
rect 1035 621 1065 895
rect 1131 621 1161 895
rect 1227 621 1257 895
rect 357 -531 387 -257
rect 453 -531 483 -257
rect 549 -531 579 -257
rect 645 -531 675 -257
rect 741 -531 771 -257
rect 837 -531 867 -257
rect 933 -531 963 -257
rect 1029 -531 1059 -257
rect 1125 -531 1155 -257
rect 1221 -531 1251 -257
<< ndiff >>
rect 301 304 363 316
rect 301 222 313 304
rect 347 222 363 304
rect 301 210 363 222
rect 393 304 459 316
rect 393 222 409 304
rect 443 222 459 304
rect 393 210 459 222
rect 489 304 555 316
rect 489 222 505 304
rect 539 222 555 304
rect 489 210 555 222
rect 585 304 651 316
rect 585 222 601 304
rect 635 222 651 304
rect 585 210 651 222
rect 681 304 747 316
rect 681 222 697 304
rect 731 222 747 304
rect 681 210 747 222
rect 777 304 843 316
rect 777 222 793 304
rect 827 222 843 304
rect 777 210 843 222
rect 873 304 939 316
rect 873 222 889 304
rect 923 222 939 304
rect 873 210 939 222
rect 969 304 1035 316
rect 969 222 985 304
rect 1019 222 1035 304
rect 969 210 1035 222
rect 1065 304 1131 316
rect 1065 222 1081 304
rect 1115 222 1131 304
rect 1065 210 1131 222
rect 1161 304 1227 316
rect 1161 222 1177 304
rect 1211 222 1227 304
rect 1161 210 1227 222
rect 1257 304 1319 316
rect 1257 222 1273 304
rect 1307 222 1319 304
rect 1257 210 1319 222
rect 295 -848 357 -836
rect 295 -930 307 -848
rect 341 -930 357 -848
rect 295 -942 357 -930
rect 387 -848 453 -836
rect 387 -930 403 -848
rect 437 -930 453 -848
rect 387 -942 453 -930
rect 483 -848 549 -836
rect 483 -930 499 -848
rect 533 -930 549 -848
rect 483 -942 549 -930
rect 579 -848 645 -836
rect 579 -930 595 -848
rect 629 -930 645 -848
rect 579 -942 645 -930
rect 675 -848 741 -836
rect 675 -930 691 -848
rect 725 -930 741 -848
rect 675 -942 741 -930
rect 771 -848 837 -836
rect 771 -930 787 -848
rect 821 -930 837 -848
rect 771 -942 837 -930
rect 867 -848 933 -836
rect 867 -930 883 -848
rect 917 -930 933 -848
rect 867 -942 933 -930
rect 963 -848 1029 -836
rect 963 -930 979 -848
rect 1013 -930 1029 -848
rect 963 -942 1029 -930
rect 1059 -848 1125 -836
rect 1059 -930 1075 -848
rect 1109 -930 1125 -848
rect 1059 -942 1125 -930
rect 1155 -848 1221 -836
rect 1155 -930 1171 -848
rect 1205 -930 1221 -848
rect 1155 -942 1221 -930
rect 1251 -848 1313 -836
rect 1251 -930 1267 -848
rect 1301 -930 1313 -848
rect 1251 -942 1313 -930
<< pdiff >>
rect 301 883 363 895
rect 301 633 313 883
rect 347 633 363 883
rect 301 621 363 633
rect 393 883 459 895
rect 393 633 409 883
rect 443 633 459 883
rect 393 621 459 633
rect 489 883 555 895
rect 489 633 505 883
rect 539 633 555 883
rect 489 621 555 633
rect 585 883 651 895
rect 585 633 601 883
rect 635 633 651 883
rect 585 621 651 633
rect 681 883 747 895
rect 681 633 697 883
rect 731 633 747 883
rect 681 621 747 633
rect 777 883 843 895
rect 777 633 793 883
rect 827 633 843 883
rect 777 621 843 633
rect 873 883 939 895
rect 873 633 889 883
rect 923 633 939 883
rect 873 621 939 633
rect 969 883 1035 895
rect 969 633 985 883
rect 1019 633 1035 883
rect 969 621 1035 633
rect 1065 883 1131 895
rect 1065 633 1081 883
rect 1115 633 1131 883
rect 1065 621 1131 633
rect 1161 883 1227 895
rect 1161 633 1177 883
rect 1211 633 1227 883
rect 1161 621 1227 633
rect 1257 883 1319 895
rect 1257 633 1273 883
rect 1307 633 1319 883
rect 1257 621 1319 633
rect 295 -269 357 -257
rect 295 -519 307 -269
rect 341 -519 357 -269
rect 295 -531 357 -519
rect 387 -269 453 -257
rect 387 -519 403 -269
rect 437 -519 453 -269
rect 387 -531 453 -519
rect 483 -269 549 -257
rect 483 -519 499 -269
rect 533 -519 549 -269
rect 483 -531 549 -519
rect 579 -269 645 -257
rect 579 -519 595 -269
rect 629 -519 645 -269
rect 579 -531 645 -519
rect 675 -269 741 -257
rect 675 -519 691 -269
rect 725 -519 741 -269
rect 675 -531 741 -519
rect 771 -269 837 -257
rect 771 -519 787 -269
rect 821 -519 837 -269
rect 771 -531 837 -519
rect 867 -269 933 -257
rect 867 -519 883 -269
rect 917 -519 933 -269
rect 867 -531 933 -519
rect 963 -269 1029 -257
rect 963 -519 979 -269
rect 1013 -519 1029 -269
rect 963 -531 1029 -519
rect 1059 -269 1125 -257
rect 1059 -519 1075 -269
rect 1109 -519 1125 -269
rect 1059 -531 1125 -519
rect 1155 -269 1221 -257
rect 1155 -519 1171 -269
rect 1205 -519 1221 -269
rect 1155 -531 1221 -519
rect 1251 -269 1313 -257
rect 1251 -519 1267 -269
rect 1301 -519 1313 -269
rect 1251 -531 1313 -519
<< ndiffc >>
rect 313 222 347 304
rect 409 222 443 304
rect 505 222 539 304
rect 601 222 635 304
rect 697 222 731 304
rect 793 222 827 304
rect 889 222 923 304
rect 985 222 1019 304
rect 1081 222 1115 304
rect 1177 222 1211 304
rect 1273 222 1307 304
rect 307 -930 341 -848
rect 403 -930 437 -848
rect 499 -930 533 -848
rect 595 -930 629 -848
rect 691 -930 725 -848
rect 787 -930 821 -848
rect 883 -930 917 -848
rect 979 -930 1013 -848
rect 1075 -930 1109 -848
rect 1171 -930 1205 -848
rect 1267 -930 1301 -848
<< pdiffc >>
rect 313 633 347 883
rect 409 633 443 883
rect 505 633 539 883
rect 601 633 635 883
rect 697 633 731 883
rect 793 633 827 883
rect 889 633 923 883
rect 985 633 1019 883
rect 1081 633 1115 883
rect 1177 633 1211 883
rect 1273 633 1307 883
rect 307 -519 341 -269
rect 403 -519 437 -269
rect 499 -519 533 -269
rect 595 -519 629 -269
rect 691 -519 725 -269
rect 787 -519 821 -269
rect 883 -519 917 -269
rect 979 -519 1013 -269
rect 1075 -519 1109 -269
rect 1171 -519 1205 -269
rect 1267 -519 1301 -269
<< psubdiff >>
rect 199 394 295 428
rect 1325 394 1421 428
rect 199 332 233 394
rect 1387 332 1421 394
rect 199 70 233 132
rect 1387 70 1421 132
rect 199 36 295 70
rect 1325 36 1421 70
rect 193 -758 289 -724
rect 1319 -758 1415 -724
rect 193 -820 227 -758
rect 1381 -820 1415 -758
rect 193 -1082 227 -1020
rect 1381 -1082 1415 -1020
rect 193 -1116 289 -1082
rect 1319 -1116 1415 -1082
<< nsubdiff >>
rect 199 1044 295 1078
rect 1325 1044 1421 1078
rect 199 982 233 1044
rect 1387 982 1421 1044
rect 199 534 233 596
rect 1387 534 1421 596
rect 199 500 295 534
rect 1325 500 1421 534
rect 193 -108 289 -74
rect 1319 -108 1415 -74
rect 193 -170 227 -108
rect 1381 -170 1415 -108
rect 193 -618 227 -556
rect 1381 -618 1415 -556
rect 193 -652 289 -618
rect 1319 -652 1415 -618
<< psubdiffcont >>
rect 295 394 1325 428
rect 199 132 233 332
rect 1387 132 1421 332
rect 295 36 1325 70
rect 289 -758 1319 -724
rect 193 -1020 227 -820
rect 1381 -1020 1415 -820
rect 289 -1116 1319 -1082
<< nsubdiffcont >>
rect 295 1044 1325 1078
rect 199 596 233 982
rect 1387 596 1421 982
rect 295 500 1325 534
rect 289 -108 1319 -74
rect 193 -556 227 -170
rect 1381 -556 1415 -170
rect 289 -652 1319 -618
<< poly >>
rect 297 976 1323 992
rect 297 942 313 976
rect 347 942 505 976
rect 539 942 697 976
rect 731 942 889 976
rect 923 942 1081 976
rect 1115 942 1273 976
rect 1307 942 1323 976
rect 297 926 1323 942
rect 363 895 393 926
rect 459 895 489 926
rect 555 895 585 926
rect 651 895 681 926
rect 747 895 777 926
rect 843 895 873 926
rect 939 895 969 926
rect 1035 895 1065 926
rect 1131 895 1161 926
rect 1227 895 1257 926
rect 363 595 393 621
rect 459 595 489 621
rect 555 595 585 621
rect 651 595 681 621
rect 747 595 777 621
rect 843 595 873 621
rect 939 595 969 621
rect 1035 595 1065 621
rect 1131 595 1161 621
rect 1227 595 1257 621
rect 363 316 393 342
rect 459 316 489 342
rect 555 316 585 342
rect 651 316 681 342
rect 747 316 777 342
rect 843 316 873 342
rect 939 316 969 342
rect 1035 316 1065 342
rect 1131 316 1161 342
rect 1227 316 1257 342
rect 363 188 393 210
rect 459 188 489 210
rect 555 188 585 210
rect 651 188 681 210
rect 747 188 777 210
rect 843 188 873 210
rect 939 188 969 210
rect 1035 188 1065 210
rect 1131 188 1161 210
rect 1227 188 1257 210
rect 297 169 1323 188
rect 297 135 313 169
rect 347 135 505 169
rect 539 135 697 169
rect 731 135 889 169
rect 923 135 1081 169
rect 1115 135 1273 169
rect 1307 135 1323 169
rect 297 122 1323 135
rect 291 -176 1317 -160
rect 291 -210 307 -176
rect 341 -210 499 -176
rect 533 -210 691 -176
rect 725 -210 883 -176
rect 917 -210 1075 -176
rect 1109 -210 1267 -176
rect 1301 -210 1317 -176
rect 291 -226 1317 -210
rect 357 -257 387 -226
rect 453 -257 483 -226
rect 549 -257 579 -226
rect 645 -257 675 -226
rect 741 -257 771 -226
rect 837 -257 867 -226
rect 933 -257 963 -226
rect 1029 -257 1059 -226
rect 1125 -257 1155 -226
rect 1221 -257 1251 -226
rect 357 -557 387 -531
rect 453 -557 483 -531
rect 549 -557 579 -531
rect 645 -557 675 -531
rect 741 -557 771 -531
rect 837 -557 867 -531
rect 933 -557 963 -531
rect 1029 -557 1059 -531
rect 1125 -557 1155 -531
rect 1221 -557 1251 -531
rect 357 -836 387 -810
rect 453 -836 483 -810
rect 549 -836 579 -810
rect 645 -836 675 -810
rect 741 -836 771 -810
rect 837 -836 867 -810
rect 933 -836 963 -810
rect 1029 -836 1059 -810
rect 1125 -836 1155 -810
rect 1221 -836 1251 -810
rect 357 -964 387 -942
rect 453 -964 483 -942
rect 549 -964 579 -942
rect 645 -964 675 -942
rect 741 -964 771 -942
rect 837 -964 867 -942
rect 933 -964 963 -942
rect 1029 -964 1059 -942
rect 1125 -964 1155 -942
rect 1221 -964 1251 -942
rect 291 -983 1317 -964
rect 291 -1017 307 -983
rect 341 -1017 499 -983
rect 533 -1017 691 -983
rect 725 -1017 883 -983
rect 917 -1017 1075 -983
rect 1109 -1017 1267 -983
rect 1301 -1017 1317 -983
rect 291 -1030 1317 -1017
<< polycont >>
rect 313 942 347 976
rect 505 942 539 976
rect 697 942 731 976
rect 889 942 923 976
rect 1081 942 1115 976
rect 1273 942 1307 976
rect 313 135 347 169
rect 505 135 539 169
rect 697 135 731 169
rect 889 135 923 169
rect 1081 135 1115 169
rect 1273 135 1307 169
rect 307 -210 341 -176
rect 499 -210 533 -176
rect 691 -210 725 -176
rect 883 -210 917 -176
rect 1075 -210 1109 -176
rect 1267 -210 1301 -176
rect 307 -1017 341 -983
rect 499 -1017 533 -983
rect 691 -1017 725 -983
rect 883 -1017 917 -983
rect 1075 -1017 1109 -983
rect 1267 -1017 1301 -983
<< locali >>
rect 199 1044 295 1078
rect 1325 1044 1421 1078
rect 199 982 233 1044
rect 1387 982 1421 1044
rect 297 942 313 976
rect 347 942 363 976
rect 489 942 505 976
rect 539 942 555 976
rect 681 942 697 976
rect 731 942 747 976
rect 873 942 889 976
rect 923 942 939 976
rect 1065 942 1081 976
rect 1115 942 1131 976
rect 1257 942 1273 976
rect 1307 942 1323 976
rect 313 883 347 899
rect 313 617 347 633
rect 409 883 443 899
rect 409 617 443 633
rect 505 883 539 899
rect 505 617 539 633
rect 601 883 635 899
rect 601 617 635 633
rect 697 883 731 899
rect 697 617 731 633
rect 793 883 827 899
rect 793 617 827 633
rect 889 883 923 899
rect 889 617 923 633
rect 985 883 1019 899
rect 985 617 1019 633
rect 1081 883 1115 899
rect 1081 617 1115 633
rect 1177 883 1211 899
rect 1177 617 1211 633
rect 1273 883 1307 899
rect 1273 617 1307 633
rect 199 534 233 596
rect 1387 534 1421 596
rect 199 500 295 534
rect 1325 500 1421 534
rect 199 394 295 428
rect 1325 394 1421 428
rect 199 332 233 394
rect 1387 332 1421 394
rect 313 304 347 320
rect 313 206 347 222
rect 409 304 443 320
rect 409 206 443 222
rect 505 304 539 320
rect 505 206 539 222
rect 601 304 635 320
rect 601 206 635 222
rect 697 304 731 320
rect 697 206 731 222
rect 793 304 827 320
rect 793 206 827 222
rect 889 304 923 320
rect 889 206 923 222
rect 985 304 1019 320
rect 985 206 1019 222
rect 1081 304 1115 320
rect 1081 206 1115 222
rect 1177 304 1211 320
rect 1177 206 1211 222
rect 1273 304 1307 320
rect 1273 206 1307 222
rect 297 135 313 169
rect 347 135 363 169
rect 489 135 505 169
rect 539 135 555 169
rect 681 135 697 169
rect 731 135 747 169
rect 873 135 889 169
rect 923 135 939 169
rect 1065 135 1081 169
rect 1115 135 1131 169
rect 1257 135 1273 169
rect 1307 135 1323 169
rect 199 70 233 132
rect 1387 70 1421 132
rect 199 36 295 70
rect 1325 36 1421 70
rect 193 -108 289 -74
rect 1319 -108 1415 -74
rect 193 -170 227 -108
rect 1381 -170 1415 -108
rect 291 -210 307 -176
rect 341 -210 357 -176
rect 483 -210 499 -176
rect 533 -210 549 -176
rect 675 -210 691 -176
rect 725 -210 741 -176
rect 867 -210 883 -176
rect 917 -210 933 -176
rect 1059 -210 1075 -176
rect 1109 -210 1125 -176
rect 1251 -210 1267 -176
rect 1301 -210 1317 -176
rect 307 -269 341 -253
rect 307 -535 341 -519
rect 403 -269 437 -253
rect 403 -535 437 -519
rect 499 -269 533 -253
rect 499 -535 533 -519
rect 595 -269 629 -253
rect 595 -535 629 -519
rect 691 -269 725 -253
rect 691 -535 725 -519
rect 787 -269 821 -253
rect 787 -535 821 -519
rect 883 -269 917 -253
rect 883 -535 917 -519
rect 979 -269 1013 -253
rect 979 -535 1013 -519
rect 1075 -269 1109 -253
rect 1075 -535 1109 -519
rect 1171 -269 1205 -253
rect 1171 -535 1205 -519
rect 1267 -269 1301 -253
rect 1267 -535 1301 -519
rect 193 -618 227 -556
rect 1381 -618 1415 -556
rect 193 -652 289 -618
rect 1319 -652 1415 -618
rect 193 -758 289 -724
rect 1319 -758 1415 -724
rect 193 -820 227 -758
rect 1381 -820 1415 -758
rect 307 -848 341 -832
rect 307 -946 341 -930
rect 403 -848 437 -832
rect 403 -946 437 -930
rect 499 -848 533 -832
rect 499 -946 533 -930
rect 595 -848 629 -832
rect 595 -946 629 -930
rect 691 -848 725 -832
rect 691 -946 725 -930
rect 787 -848 821 -832
rect 787 -946 821 -930
rect 883 -848 917 -832
rect 883 -946 917 -930
rect 979 -848 1013 -832
rect 979 -946 1013 -930
rect 1075 -848 1109 -832
rect 1075 -946 1109 -930
rect 1171 -848 1205 -832
rect 1171 -946 1205 -930
rect 1267 -848 1301 -832
rect 1267 -946 1301 -930
rect 291 -1017 307 -983
rect 341 -1017 357 -983
rect 483 -1017 499 -983
rect 533 -1017 549 -983
rect 675 -1017 691 -983
rect 725 -1017 741 -983
rect 867 -1017 883 -983
rect 917 -1017 933 -983
rect 1059 -1017 1075 -983
rect 1109 -1017 1125 -983
rect 1251 -1017 1267 -983
rect 1301 -1017 1317 -983
rect 193 -1082 227 -1020
rect 1381 -1082 1415 -1020
rect 193 -1116 289 -1082
rect 1319 -1116 1415 -1082
<< viali >>
rect 313 942 347 976
rect 505 942 539 976
rect 697 942 731 976
rect 889 942 923 976
rect 1081 942 1115 976
rect 1273 942 1307 976
rect 313 633 347 883
rect 409 633 443 883
rect 505 633 539 883
rect 601 633 635 883
rect 697 633 731 883
rect 793 633 827 883
rect 889 633 923 883
rect 985 633 1019 883
rect 1081 633 1115 883
rect 1177 633 1211 883
rect 1273 633 1307 883
rect 1387 596 1421 982
rect 313 222 347 304
rect 409 222 443 304
rect 505 222 539 304
rect 601 222 635 304
rect 697 222 731 304
rect 793 222 827 304
rect 889 222 923 304
rect 985 222 1019 304
rect 1081 222 1115 304
rect 1177 222 1211 304
rect 1273 222 1307 304
rect 313 135 347 169
rect 505 135 539 169
rect 697 135 731 169
rect 889 135 923 169
rect 1081 135 1115 169
rect 1273 135 1307 169
rect 1387 132 1421 332
rect 307 -210 341 -176
rect 499 -210 533 -176
rect 691 -210 725 -176
rect 883 -210 917 -176
rect 1075 -210 1109 -176
rect 1267 -210 1301 -176
rect 307 -519 341 -269
rect 403 -519 437 -269
rect 499 -519 533 -269
rect 595 -519 629 -269
rect 691 -519 725 -269
rect 787 -519 821 -269
rect 883 -519 917 -269
rect 979 -519 1013 -269
rect 1075 -519 1109 -269
rect 1171 -519 1205 -269
rect 1267 -519 1301 -269
rect 1381 -556 1415 -170
rect 307 -930 341 -848
rect 403 -930 437 -848
rect 499 -930 533 -848
rect 595 -930 629 -848
rect 691 -930 725 -848
rect 787 -930 821 -848
rect 883 -930 917 -848
rect 979 -930 1013 -848
rect 1075 -930 1109 -848
rect 1171 -930 1205 -848
rect 1267 -930 1301 -848
rect 307 -1017 341 -983
rect 499 -1017 533 -983
rect 691 -1017 725 -983
rect 883 -1017 917 -983
rect 1075 -1017 1109 -983
rect 1267 -1017 1301 -983
rect 1381 -1020 1415 -820
<< metal1 >>
rect 129 1044 1211 1078
rect -133 934 27 986
rect 79 934 89 986
rect -300 438 -238 490
rect -186 438 -176 490
rect -298 -38 -236 14
rect -184 -38 -174 14
rect -133 -326 -81 934
rect -10 438 0 490
rect 52 481 62 490
rect 129 481 163 1044
rect 294 934 304 986
rect 356 934 366 986
rect 409 895 443 1044
rect 487 934 497 986
rect 549 934 559 986
rect 601 895 635 1044
rect 678 934 688 986
rect 740 934 750 986
rect 793 895 827 1044
rect 870 934 880 986
rect 932 934 942 986
rect 985 895 1019 1044
rect 1062 934 1072 986
rect 1124 934 1134 986
rect 1177 895 1211 1044
rect 1381 1062 1892 1114
rect 1254 934 1264 986
rect 1316 934 1326 986
rect 1381 982 1427 1062
rect 307 883 353 895
rect 307 633 313 883
rect 347 633 353 883
rect 307 621 353 633
rect 403 883 449 895
rect 403 633 409 883
rect 443 633 449 883
rect 403 621 449 633
rect 499 883 545 895
rect 499 633 505 883
rect 539 633 545 883
rect 499 621 545 633
rect 595 883 641 895
rect 595 633 601 883
rect 635 633 641 883
rect 595 621 641 633
rect 691 883 737 895
rect 691 633 697 883
rect 731 633 737 883
rect 691 621 737 633
rect 787 883 833 895
rect 787 633 793 883
rect 827 633 833 883
rect 787 621 833 633
rect 883 883 929 895
rect 883 633 889 883
rect 923 633 929 883
rect 883 621 929 633
rect 979 883 1025 895
rect 979 633 985 883
rect 1019 633 1025 883
rect 979 621 1025 633
rect 1075 883 1121 895
rect 1075 633 1081 883
rect 1115 633 1121 883
rect 1075 621 1121 633
rect 1171 883 1217 895
rect 1171 633 1177 883
rect 1211 633 1217 883
rect 1171 621 1217 633
rect 1267 883 1313 895
rect 1267 633 1273 883
rect 1307 633 1313 883
rect 1267 621 1313 633
rect 52 447 163 481
rect 52 438 62 447
rect -31 127 27 179
rect 79 127 89 179
rect -31 14 21 127
rect 129 70 163 447
rect 313 481 347 621
rect 505 481 539 621
rect 697 481 731 621
rect 889 481 923 621
rect 1081 481 1115 621
rect 1273 481 1307 621
rect 1381 596 1387 982
rect 1421 630 1427 982
rect 1421 596 1727 630
rect 1381 584 1427 596
rect 313 447 1530 481
rect 313 316 347 447
rect 505 316 539 447
rect 697 316 731 447
rect 889 316 923 447
rect 1081 316 1115 447
rect 1273 316 1307 447
rect 1381 333 1427 344
rect 307 304 353 316
rect 307 222 313 304
rect 347 222 353 304
rect 307 210 353 222
rect 403 304 449 316
rect 403 222 409 304
rect 443 222 449 304
rect 403 210 449 222
rect 499 304 545 316
rect 499 222 505 304
rect 539 222 545 304
rect 499 210 545 222
rect 595 304 641 316
rect 595 222 601 304
rect 635 222 641 304
rect 595 210 641 222
rect 691 304 737 316
rect 691 222 697 304
rect 731 222 737 304
rect 691 210 737 222
rect 787 304 833 316
rect 787 222 793 304
rect 827 222 833 304
rect 787 210 833 222
rect 883 304 929 316
rect 883 222 889 304
rect 923 222 929 304
rect 883 210 929 222
rect 979 304 1025 316
rect 979 222 985 304
rect 1019 222 1025 304
rect 979 210 1025 222
rect 1075 304 1121 316
rect 1075 222 1081 304
rect 1115 222 1121 304
rect 1075 210 1121 222
rect 1171 304 1217 316
rect 1171 222 1177 304
rect 1211 222 1217 304
rect 1171 210 1217 222
rect 1267 304 1313 316
rect 1267 222 1273 304
rect 1307 222 1313 304
rect 1368 281 1378 333
rect 1430 281 1440 333
rect 1267 210 1313 222
rect 297 179 363 182
rect 294 127 304 179
rect 356 127 366 179
rect 297 122 363 127
rect 409 70 443 210
rect 489 179 555 182
rect 485 127 495 179
rect 547 127 557 179
rect 489 122 555 127
rect 601 70 635 210
rect 681 179 747 182
rect 677 127 687 179
rect 739 127 749 179
rect 681 122 747 127
rect 793 70 827 210
rect 873 179 939 182
rect 869 127 879 179
rect 931 127 941 179
rect 873 122 939 127
rect 985 70 1019 210
rect 1065 178 1131 182
rect 1062 126 1072 178
rect 1124 126 1134 178
rect 1065 122 1131 126
rect 1177 70 1211 210
rect 1257 178 1323 182
rect 1254 126 1264 178
rect 1316 126 1326 178
rect 1381 132 1387 281
rect 1421 132 1427 281
rect 1257 122 1323 126
rect 129 36 1211 70
rect -41 -38 -31 14
rect 21 -38 31 14
rect 1381 0 1427 132
rect 1496 5 1530 447
rect 1571 281 1581 333
rect 1633 281 1643 333
rect -31 -218 21 -38
rect 123 -108 1205 -74
rect 73 -218 83 -166
rect -313 -378 -81 -326
rect -300 -715 -238 -663
rect -186 -715 -176 -663
rect -133 -973 -81 -378
rect -17 -715 -7 -663
rect 45 -671 55 -663
rect 123 -671 157 -108
rect 288 -218 298 -166
rect 350 -218 360 -166
rect 403 -257 437 -108
rect 481 -218 491 -166
rect 543 -218 553 -166
rect 595 -257 629 -108
rect 672 -218 682 -166
rect 734 -218 744 -166
rect 787 -257 821 -108
rect 864 -218 874 -166
rect 926 -218 936 -166
rect 979 -257 1013 -108
rect 1056 -218 1066 -166
rect 1118 -218 1128 -166
rect 1171 -257 1205 -108
rect 1248 -218 1258 -166
rect 1310 -218 1320 -166
rect 1375 -170 1421 -38
rect 1477 -47 1487 5
rect 1539 -47 1549 5
rect 301 -269 347 -257
rect 301 -519 307 -269
rect 341 -519 347 -269
rect 301 -531 347 -519
rect 397 -269 443 -257
rect 397 -519 403 -269
rect 437 -519 443 -269
rect 397 -531 443 -519
rect 493 -269 539 -257
rect 493 -519 499 -269
rect 533 -519 539 -269
rect 493 -531 539 -519
rect 589 -269 635 -257
rect 589 -519 595 -269
rect 629 -519 635 -269
rect 589 -531 635 -519
rect 685 -269 731 -257
rect 685 -519 691 -269
rect 725 -519 731 -269
rect 685 -531 731 -519
rect 781 -269 827 -257
rect 781 -519 787 -269
rect 821 -519 827 -269
rect 781 -531 827 -519
rect 877 -269 923 -257
rect 877 -519 883 -269
rect 917 -519 923 -269
rect 877 -531 923 -519
rect 973 -269 1019 -257
rect 973 -519 979 -269
rect 1013 -519 1019 -269
rect 973 -531 1019 -519
rect 1069 -269 1115 -257
rect 1069 -519 1075 -269
rect 1109 -519 1115 -269
rect 1069 -531 1115 -519
rect 1165 -269 1211 -257
rect 1165 -519 1171 -269
rect 1205 -519 1211 -269
rect 1165 -531 1211 -519
rect 1261 -269 1307 -257
rect 1261 -519 1267 -269
rect 1301 -519 1307 -269
rect 1375 -505 1381 -170
rect 1415 -505 1421 -170
rect 1261 -531 1307 -519
rect 45 -705 157 -671
rect 45 -715 55 -705
rect -133 -1025 21 -973
rect 73 -1025 83 -973
rect 123 -1082 157 -705
rect 307 -671 341 -531
rect 499 -671 533 -531
rect 691 -671 725 -531
rect 883 -671 917 -531
rect 1075 -671 1109 -531
rect 1267 -671 1301 -531
rect 1362 -557 1372 -505
rect 1424 -557 1434 -505
rect 1375 -568 1421 -557
rect 1496 -671 1530 -47
rect 307 -705 1530 -671
rect 307 -836 341 -705
rect 499 -836 533 -705
rect 691 -836 725 -705
rect 883 -836 917 -705
rect 1075 -836 1109 -705
rect 1267 -836 1301 -705
rect 1375 -820 1421 -808
rect 1590 -820 1624 281
rect 1693 -505 1727 596
rect 1782 -47 1792 5
rect 1844 -47 1895 5
rect 1674 -557 1684 -505
rect 1736 -557 1746 -505
rect 301 -848 347 -836
rect 301 -930 307 -848
rect 341 -930 347 -848
rect 301 -942 347 -930
rect 397 -848 443 -836
rect 397 -930 403 -848
rect 437 -930 443 -848
rect 397 -942 443 -930
rect 493 -848 539 -836
rect 493 -930 499 -848
rect 533 -930 539 -848
rect 493 -942 539 -930
rect 589 -848 635 -836
rect 589 -930 595 -848
rect 629 -930 635 -848
rect 589 -942 635 -930
rect 685 -848 731 -836
rect 685 -930 691 -848
rect 725 -930 731 -848
rect 685 -942 731 -930
rect 781 -848 827 -836
rect 781 -930 787 -848
rect 821 -930 827 -848
rect 781 -942 827 -930
rect 877 -848 923 -836
rect 877 -930 883 -848
rect 917 -930 923 -848
rect 877 -942 923 -930
rect 973 -848 1019 -836
rect 973 -930 979 -848
rect 1013 -930 1019 -848
rect 973 -942 1019 -930
rect 1069 -848 1115 -836
rect 1069 -930 1075 -848
rect 1109 -930 1115 -848
rect 1069 -942 1115 -930
rect 1165 -848 1211 -836
rect 1165 -930 1171 -848
rect 1205 -930 1211 -848
rect 1165 -942 1211 -930
rect 1261 -848 1307 -836
rect 1261 -930 1267 -848
rect 1301 -930 1307 -848
rect 1261 -942 1307 -930
rect 291 -973 357 -970
rect 288 -1025 298 -973
rect 350 -1025 360 -973
rect 291 -1030 357 -1025
rect 403 -1082 437 -942
rect 483 -973 549 -970
rect 479 -1025 489 -973
rect 541 -1025 551 -973
rect 483 -1030 549 -1025
rect 595 -1082 629 -942
rect 675 -973 741 -970
rect 671 -1025 681 -973
rect 733 -1025 743 -973
rect 675 -1030 741 -1025
rect 787 -1082 821 -942
rect 867 -973 933 -970
rect 863 -1025 873 -973
rect 925 -1025 935 -973
rect 867 -1030 933 -1025
rect 979 -1082 1013 -942
rect 1059 -974 1125 -970
rect 1056 -1026 1066 -974
rect 1118 -1026 1128 -974
rect 1059 -1030 1125 -1026
rect 1171 -1082 1205 -942
rect 1251 -974 1317 -970
rect 1248 -1026 1258 -974
rect 1310 -1026 1320 -974
rect 1375 -1020 1381 -820
rect 1415 -854 1624 -820
rect 1415 -1020 1421 -854
rect 1251 -1030 1317 -1026
rect 123 -1116 1205 -1082
rect 1375 -1102 1421 -1020
rect 1374 -1154 1885 -1102
<< via1 >>
rect 27 934 79 986
rect -238 438 -186 490
rect -236 -38 -184 14
rect 0 438 52 490
rect 304 976 356 986
rect 304 942 313 976
rect 313 942 347 976
rect 347 942 356 976
rect 304 934 356 942
rect 497 976 549 986
rect 497 942 505 976
rect 505 942 539 976
rect 539 942 549 976
rect 497 934 549 942
rect 688 976 740 986
rect 688 942 697 976
rect 697 942 731 976
rect 731 942 740 976
rect 688 934 740 942
rect 880 976 932 986
rect 880 942 889 976
rect 889 942 923 976
rect 923 942 932 976
rect 880 934 932 942
rect 1072 976 1124 986
rect 1072 942 1081 976
rect 1081 942 1115 976
rect 1115 942 1124 976
rect 1072 934 1124 942
rect 1264 976 1316 986
rect 1264 942 1273 976
rect 1273 942 1307 976
rect 1307 942 1316 976
rect 1264 934 1316 942
rect 27 127 79 179
rect 1378 332 1430 333
rect 1378 281 1387 332
rect 1387 281 1421 332
rect 1421 281 1430 332
rect 304 169 356 179
rect 304 135 313 169
rect 313 135 347 169
rect 347 135 356 169
rect 304 127 356 135
rect 495 169 547 179
rect 495 135 505 169
rect 505 135 539 169
rect 539 135 547 169
rect 495 127 547 135
rect 687 169 739 179
rect 687 135 697 169
rect 697 135 731 169
rect 731 135 739 169
rect 687 127 739 135
rect 879 169 931 179
rect 879 135 889 169
rect 889 135 923 169
rect 923 135 931 169
rect 879 127 931 135
rect 1072 169 1124 178
rect 1072 135 1081 169
rect 1081 135 1115 169
rect 1115 135 1124 169
rect 1072 126 1124 135
rect 1264 169 1316 178
rect 1264 135 1273 169
rect 1273 135 1307 169
rect 1307 135 1316 169
rect 1264 126 1316 135
rect -31 -38 21 14
rect 1581 281 1633 333
rect 21 -218 73 -166
rect -238 -715 -186 -663
rect -7 -715 45 -663
rect 298 -176 350 -166
rect 298 -210 307 -176
rect 307 -210 341 -176
rect 341 -210 350 -176
rect 298 -218 350 -210
rect 491 -176 543 -166
rect 491 -210 499 -176
rect 499 -210 533 -176
rect 533 -210 543 -176
rect 491 -218 543 -210
rect 682 -176 734 -166
rect 682 -210 691 -176
rect 691 -210 725 -176
rect 725 -210 734 -176
rect 682 -218 734 -210
rect 874 -176 926 -166
rect 874 -210 883 -176
rect 883 -210 917 -176
rect 917 -210 926 -176
rect 874 -218 926 -210
rect 1066 -176 1118 -166
rect 1066 -210 1075 -176
rect 1075 -210 1109 -176
rect 1109 -210 1118 -176
rect 1066 -218 1118 -210
rect 1258 -176 1310 -166
rect 1258 -210 1267 -176
rect 1267 -210 1301 -176
rect 1301 -210 1310 -176
rect 1258 -218 1310 -210
rect 1487 -47 1539 5
rect 21 -1025 73 -973
rect 1372 -556 1381 -505
rect 1381 -556 1415 -505
rect 1415 -556 1424 -505
rect 1372 -557 1424 -556
rect 1792 -47 1844 5
rect 1684 -557 1736 -505
rect 298 -983 350 -973
rect 298 -1017 307 -983
rect 307 -1017 341 -983
rect 341 -1017 350 -983
rect 298 -1025 350 -1017
rect 489 -983 541 -973
rect 489 -1017 499 -983
rect 499 -1017 533 -983
rect 533 -1017 541 -983
rect 489 -1025 541 -1017
rect 681 -983 733 -973
rect 681 -1017 691 -983
rect 691 -1017 725 -983
rect 725 -1017 733 -983
rect 681 -1025 733 -1017
rect 873 -983 925 -973
rect 873 -1017 883 -983
rect 883 -1017 917 -983
rect 917 -1017 925 -983
rect 873 -1025 925 -1017
rect 1066 -983 1118 -974
rect 1066 -1017 1075 -983
rect 1075 -1017 1109 -983
rect 1109 -1017 1118 -983
rect 1066 -1026 1118 -1017
rect 1258 -983 1310 -974
rect 1258 -1017 1267 -983
rect 1267 -1017 1301 -983
rect 1301 -1017 1310 -983
rect 1258 -1026 1310 -1017
<< metal2 >>
rect 27 986 79 996
rect 304 986 356 996
rect 497 986 549 996
rect 688 986 740 996
rect 880 986 932 996
rect 1072 986 1124 996
rect 1264 986 1316 996
rect 79 934 304 986
rect 356 934 497 986
rect 549 934 688 986
rect 740 934 880 986
rect 932 934 1072 986
rect 1124 934 1264 986
rect 1316 934 1323 986
rect 27 924 79 934
rect 304 924 356 934
rect 497 924 549 934
rect 688 924 740 934
rect 880 924 932 934
rect 1072 924 1124 934
rect 1264 924 1316 934
rect -238 490 -186 500
rect 0 490 52 500
rect -186 438 0 490
rect -238 428 -186 438
rect 0 428 52 438
rect 1378 333 1430 343
rect 1581 333 1633 343
rect 1430 281 1581 333
rect 1378 271 1430 281
rect 1581 271 1633 281
rect 27 179 79 189
rect 304 179 356 189
rect 495 179 547 189
rect 687 179 739 189
rect 879 179 931 189
rect 1072 179 1124 188
rect 1264 179 1316 188
rect 79 127 304 179
rect 356 127 495 179
rect 547 127 687 179
rect 739 127 879 179
rect 931 178 1323 179
rect 931 127 1072 178
rect 27 117 79 127
rect 304 117 356 127
rect 495 117 547 127
rect 687 117 739 127
rect 879 117 931 127
rect 1124 127 1264 178
rect 1072 116 1124 126
rect 1316 127 1323 178
rect 1264 116 1316 126
rect -236 14 -184 24
rect -31 14 21 24
rect -184 -38 -31 14
rect -236 -48 -184 -38
rect -31 -48 21 -38
rect 1487 5 1539 15
rect 1792 5 1844 15
rect 1539 -47 1792 5
rect 1487 -57 1539 -47
rect 1792 -57 1844 -47
rect 21 -166 73 -156
rect 298 -166 350 -156
rect 491 -166 543 -156
rect 682 -166 734 -156
rect 874 -166 926 -156
rect 1066 -166 1118 -156
rect 1258 -166 1310 -156
rect 73 -218 298 -166
rect 350 -218 491 -166
rect 543 -218 682 -166
rect 734 -218 874 -166
rect 926 -218 1066 -166
rect 1118 -218 1258 -166
rect 1310 -218 1317 -166
rect 21 -228 73 -218
rect 298 -228 350 -218
rect 491 -228 543 -218
rect 682 -228 734 -218
rect 874 -228 926 -218
rect 1066 -228 1118 -218
rect 1258 -228 1310 -218
rect 1372 -505 1424 -495
rect 1684 -505 1736 -495
rect 1424 -557 1684 -505
rect 1372 -567 1424 -557
rect 1684 -567 1736 -557
rect -238 -663 -186 -653
rect -7 -663 45 -653
rect -186 -715 -7 -663
rect -238 -725 -186 -715
rect -7 -725 45 -715
rect 21 -973 73 -963
rect 298 -973 350 -963
rect 489 -973 541 -963
rect 681 -973 733 -963
rect 873 -973 925 -963
rect 1066 -973 1118 -964
rect 1258 -973 1310 -964
rect 73 -1025 298 -973
rect 350 -1025 489 -973
rect 541 -1025 681 -973
rect 733 -1025 873 -973
rect 925 -974 1317 -973
rect 925 -1025 1066 -974
rect 21 -1035 73 -1025
rect 298 -1035 350 -1025
rect 489 -1035 541 -1025
rect 681 -1035 733 -1025
rect 873 -1035 925 -1025
rect 1118 -1025 1258 -974
rect 1066 -1036 1118 -1026
rect 1310 -1025 1317 -974
rect 1258 -1036 1310 -1026
<< labels >>
flabel metal1 -285 464 -285 464 1 FreeSans 400 0 0 0 v_hi
port 1 n
flabel metal1 -280 -690 -280 -690 1 FreeSans 400 0 0 0 v_lo
port 2 n
flabel metal1 -275 -14 -275 -14 1 FreeSans 400 0 0 0 v
port 3 n
flabel metal1 -286 -352 -286 -352 1 FreeSans 400 0 0 0 v_b
port 4 n
flabel metal1 1879 -24 1879 -24 1 FreeSans 400 0 0 0 out
port 5 n
flabel metal1 1868 1086 1868 1086 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 1867 -1131 1867 -1131 1 FreeSans 400 0 0 0 VSS
port 7 n ground bidirectional
flabel metal1 1398 -1149 1398 -1149 1 FreeSans 400 0 0 0 transmission_gate_1/VSS
flabel metal1 1398 -43 1398 -43 5 FreeSans 400 0 0 0 transmission_gate_1/VDD
flabel metal1 -1 -192 -1 -192 3 FreeSans 400 0 0 0 transmission_gate_1/en_b
flabel metal1 -2 -688 -2 -688 3 FreeSans 400 0 0 0 transmission_gate_1/in
flabel metal1 -2 -999 -2 -999 3 FreeSans 400 0 0 0 transmission_gate_1/en
flabel metal1 1489 -689 1489 -689 7 FreeSans 400 0 0 0 transmission_gate_1/out
flabel metal1 1404 3 1404 3 1 FreeSans 400 0 0 0 transmission_gate_0/VSS
flabel metal1 1404 1109 1404 1109 5 FreeSans 400 0 0 0 transmission_gate_0/VDD
flabel metal1 5 960 5 960 3 FreeSans 400 0 0 0 transmission_gate_0/en_b
flabel metal1 4 464 4 464 3 FreeSans 400 0 0 0 transmission_gate_0/in
flabel metal1 4 153 4 153 3 FreeSans 400 0 0 0 transmission_gate_0/en
flabel metal1 1495 463 1495 463 7 FreeSans 400 0 0 0 transmission_gate_0/out
<< end >>
