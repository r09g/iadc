magic
tech sky130A
magscale 1 2
timestamp 1654894986
<< error_p >>
rect -6387 18944 -6327 25142
rect -6307 18944 -6247 25142
rect -70 18944 -10 25142
rect 10 18944 70 25142
rect 6247 18944 6307 25142
rect 6327 18944 6387 25142
rect -6387 12646 -6327 18844
rect -6307 12646 -6247 18844
rect -70 12646 -10 18844
rect 10 12646 70 18844
rect 6247 12646 6307 18844
rect 6327 12646 6387 18844
rect -6387 6348 -6327 12546
rect -6307 6348 -6247 12546
rect -70 6348 -10 12546
rect 10 6348 70 12546
rect 6247 6348 6307 12546
rect 6327 6348 6387 12546
rect -6387 50 -6327 6248
rect -6307 50 -6247 6248
rect -70 50 -10 6248
rect 10 50 70 6248
rect 6247 50 6307 6248
rect 6327 50 6387 6248
rect -6387 -6248 -6327 -50
rect -6307 -6248 -6247 -50
rect -70 -6248 -10 -50
rect 10 -6248 70 -50
rect 6247 -6248 6307 -50
rect 6327 -6248 6387 -50
rect -6387 -12546 -6327 -6348
rect -6307 -12546 -6247 -6348
rect -70 -12546 -10 -6348
rect 10 -12546 70 -6348
rect 6247 -12546 6307 -6348
rect 6327 -12546 6387 -6348
rect -6387 -18844 -6327 -12646
rect -6307 -18844 -6247 -12646
rect -70 -18844 -10 -12646
rect 10 -18844 70 -12646
rect 6247 -18844 6307 -12646
rect 6327 -18844 6387 -12646
rect -6387 -25142 -6327 -18944
rect -6307 -25142 -6247 -18944
rect -70 -25142 -10 -18944
rect 10 -25142 70 -18944
rect 6247 -25142 6307 -18944
rect 6327 -25142 6387 -18944
<< metal3 >>
rect -12624 25114 -6327 25142
rect -12624 18972 -6411 25114
rect -6347 18972 -6327 25114
rect -12624 18944 -6327 18972
rect -6307 25114 -10 25142
rect -6307 18972 -94 25114
rect -30 18972 -10 25114
rect -6307 18944 -10 18972
rect 10 25114 6307 25142
rect 10 18972 6223 25114
rect 6287 18972 6307 25114
rect 10 18944 6307 18972
rect 6327 25114 12624 25142
rect 6327 18972 12540 25114
rect 12604 18972 12624 25114
rect 6327 18944 12624 18972
rect -12624 18816 -6327 18844
rect -12624 12674 -6411 18816
rect -6347 12674 -6327 18816
rect -12624 12646 -6327 12674
rect -6307 18816 -10 18844
rect -6307 12674 -94 18816
rect -30 12674 -10 18816
rect -6307 12646 -10 12674
rect 10 18816 6307 18844
rect 10 12674 6223 18816
rect 6287 12674 6307 18816
rect 10 12646 6307 12674
rect 6327 18816 12624 18844
rect 6327 12674 12540 18816
rect 12604 12674 12624 18816
rect 6327 12646 12624 12674
rect -12624 12518 -6327 12546
rect -12624 6376 -6411 12518
rect -6347 6376 -6327 12518
rect -12624 6348 -6327 6376
rect -6307 12518 -10 12546
rect -6307 6376 -94 12518
rect -30 6376 -10 12518
rect -6307 6348 -10 6376
rect 10 12518 6307 12546
rect 10 6376 6223 12518
rect 6287 6376 6307 12518
rect 10 6348 6307 6376
rect 6327 12518 12624 12546
rect 6327 6376 12540 12518
rect 12604 6376 12624 12518
rect 6327 6348 12624 6376
rect -12624 6220 -6327 6248
rect -12624 78 -6411 6220
rect -6347 78 -6327 6220
rect -12624 50 -6327 78
rect -6307 6220 -10 6248
rect -6307 78 -94 6220
rect -30 78 -10 6220
rect -6307 50 -10 78
rect 10 6220 6307 6248
rect 10 78 6223 6220
rect 6287 78 6307 6220
rect 10 50 6307 78
rect 6327 6220 12624 6248
rect 6327 78 12540 6220
rect 12604 78 12624 6220
rect 6327 50 12624 78
rect -12624 -78 -6327 -50
rect -12624 -6220 -6411 -78
rect -6347 -6220 -6327 -78
rect -12624 -6248 -6327 -6220
rect -6307 -78 -10 -50
rect -6307 -6220 -94 -78
rect -30 -6220 -10 -78
rect -6307 -6248 -10 -6220
rect 10 -78 6307 -50
rect 10 -6220 6223 -78
rect 6287 -6220 6307 -78
rect 10 -6248 6307 -6220
rect 6327 -78 12624 -50
rect 6327 -6220 12540 -78
rect 12604 -6220 12624 -78
rect 6327 -6248 12624 -6220
rect -12624 -6376 -6327 -6348
rect -12624 -12518 -6411 -6376
rect -6347 -12518 -6327 -6376
rect -12624 -12546 -6327 -12518
rect -6307 -6376 -10 -6348
rect -6307 -12518 -94 -6376
rect -30 -12518 -10 -6376
rect -6307 -12546 -10 -12518
rect 10 -6376 6307 -6348
rect 10 -12518 6223 -6376
rect 6287 -12518 6307 -6376
rect 10 -12546 6307 -12518
rect 6327 -6376 12624 -6348
rect 6327 -12518 12540 -6376
rect 12604 -12518 12624 -6376
rect 6327 -12546 12624 -12518
rect -12624 -12674 -6327 -12646
rect -12624 -18816 -6411 -12674
rect -6347 -18816 -6327 -12674
rect -12624 -18844 -6327 -18816
rect -6307 -12674 -10 -12646
rect -6307 -18816 -94 -12674
rect -30 -18816 -10 -12674
rect -6307 -18844 -10 -18816
rect 10 -12674 6307 -12646
rect 10 -18816 6223 -12674
rect 6287 -18816 6307 -12674
rect 10 -18844 6307 -18816
rect 6327 -12674 12624 -12646
rect 6327 -18816 12540 -12674
rect 12604 -18816 12624 -12674
rect 6327 -18844 12624 -18816
rect -12624 -18972 -6327 -18944
rect -12624 -25114 -6411 -18972
rect -6347 -25114 -6327 -18972
rect -12624 -25142 -6327 -25114
rect -6307 -18972 -10 -18944
rect -6307 -25114 -94 -18972
rect -30 -25114 -10 -18972
rect -6307 -25142 -10 -25114
rect 10 -18972 6307 -18944
rect 10 -25114 6223 -18972
rect 6287 -25114 6307 -18972
rect 10 -25142 6307 -25114
rect 6327 -18972 12624 -18944
rect 6327 -25114 12540 -18972
rect 12604 -25114 12624 -18972
rect 6327 -25142 12624 -25114
<< via3 >>
rect -6411 18972 -6347 25114
rect -94 18972 -30 25114
rect 6223 18972 6287 25114
rect 12540 18972 12604 25114
rect -6411 12674 -6347 18816
rect -94 12674 -30 18816
rect 6223 12674 6287 18816
rect 12540 12674 12604 18816
rect -6411 6376 -6347 12518
rect -94 6376 -30 12518
rect 6223 6376 6287 12518
rect 12540 6376 12604 12518
rect -6411 78 -6347 6220
rect -94 78 -30 6220
rect 6223 78 6287 6220
rect 12540 78 12604 6220
rect -6411 -6220 -6347 -78
rect -94 -6220 -30 -78
rect 6223 -6220 6287 -78
rect 12540 -6220 12604 -78
rect -6411 -12518 -6347 -6376
rect -94 -12518 -30 -6376
rect 6223 -12518 6287 -6376
rect 12540 -12518 12604 -6376
rect -6411 -18816 -6347 -12674
rect -94 -18816 -30 -12674
rect 6223 -18816 6287 -12674
rect 12540 -18816 12604 -12674
rect -6411 -25114 -6347 -18972
rect -94 -25114 -30 -18972
rect 6223 -25114 6287 -18972
rect 12540 -25114 12604 -18972
<< mimcap >>
rect -12524 25002 -6526 25042
rect -12524 19084 -12484 25002
rect -6566 19084 -6526 25002
rect -12524 19044 -6526 19084
rect -6207 25002 -209 25042
rect -6207 19084 -6167 25002
rect -249 19084 -209 25002
rect -6207 19044 -209 19084
rect 110 25002 6108 25042
rect 110 19084 150 25002
rect 6068 19084 6108 25002
rect 110 19044 6108 19084
rect 6427 25002 12425 25042
rect 6427 19084 6467 25002
rect 12385 19084 12425 25002
rect 6427 19044 12425 19084
rect -12524 18704 -6526 18744
rect -12524 12786 -12484 18704
rect -6566 12786 -6526 18704
rect -12524 12746 -6526 12786
rect -6207 18704 -209 18744
rect -6207 12786 -6167 18704
rect -249 12786 -209 18704
rect -6207 12746 -209 12786
rect 110 18704 6108 18744
rect 110 12786 150 18704
rect 6068 12786 6108 18704
rect 110 12746 6108 12786
rect 6427 18704 12425 18744
rect 6427 12786 6467 18704
rect 12385 12786 12425 18704
rect 6427 12746 12425 12786
rect -12524 12406 -6526 12446
rect -12524 6488 -12484 12406
rect -6566 6488 -6526 12406
rect -12524 6448 -6526 6488
rect -6207 12406 -209 12446
rect -6207 6488 -6167 12406
rect -249 6488 -209 12406
rect -6207 6448 -209 6488
rect 110 12406 6108 12446
rect 110 6488 150 12406
rect 6068 6488 6108 12406
rect 110 6448 6108 6488
rect 6427 12406 12425 12446
rect 6427 6488 6467 12406
rect 12385 6488 12425 12406
rect 6427 6448 12425 6488
rect -12524 6108 -6526 6148
rect -12524 190 -12484 6108
rect -6566 190 -6526 6108
rect -12524 150 -6526 190
rect -6207 6108 -209 6148
rect -6207 190 -6167 6108
rect -249 190 -209 6108
rect -6207 150 -209 190
rect 110 6108 6108 6148
rect 110 190 150 6108
rect 6068 190 6108 6108
rect 110 150 6108 190
rect 6427 6108 12425 6148
rect 6427 190 6467 6108
rect 12385 190 12425 6108
rect 6427 150 12425 190
rect -12524 -190 -6526 -150
rect -12524 -6108 -12484 -190
rect -6566 -6108 -6526 -190
rect -12524 -6148 -6526 -6108
rect -6207 -190 -209 -150
rect -6207 -6108 -6167 -190
rect -249 -6108 -209 -190
rect -6207 -6148 -209 -6108
rect 110 -190 6108 -150
rect 110 -6108 150 -190
rect 6068 -6108 6108 -190
rect 110 -6148 6108 -6108
rect 6427 -190 12425 -150
rect 6427 -6108 6467 -190
rect 12385 -6108 12425 -190
rect 6427 -6148 12425 -6108
rect -12524 -6488 -6526 -6448
rect -12524 -12406 -12484 -6488
rect -6566 -12406 -6526 -6488
rect -12524 -12446 -6526 -12406
rect -6207 -6488 -209 -6448
rect -6207 -12406 -6167 -6488
rect -249 -12406 -209 -6488
rect -6207 -12446 -209 -12406
rect 110 -6488 6108 -6448
rect 110 -12406 150 -6488
rect 6068 -12406 6108 -6488
rect 110 -12446 6108 -12406
rect 6427 -6488 12425 -6448
rect 6427 -12406 6467 -6488
rect 12385 -12406 12425 -6488
rect 6427 -12446 12425 -12406
rect -12524 -12786 -6526 -12746
rect -12524 -18704 -12484 -12786
rect -6566 -18704 -6526 -12786
rect -12524 -18744 -6526 -18704
rect -6207 -12786 -209 -12746
rect -6207 -18704 -6167 -12786
rect -249 -18704 -209 -12786
rect -6207 -18744 -209 -18704
rect 110 -12786 6108 -12746
rect 110 -18704 150 -12786
rect 6068 -18704 6108 -12786
rect 110 -18744 6108 -18704
rect 6427 -12786 12425 -12746
rect 6427 -18704 6467 -12786
rect 12385 -18704 12425 -12786
rect 6427 -18744 12425 -18704
rect -12524 -19084 -6526 -19044
rect -12524 -25002 -12484 -19084
rect -6566 -25002 -6526 -19084
rect -12524 -25042 -6526 -25002
rect -6207 -19084 -209 -19044
rect -6207 -25002 -6167 -19084
rect -249 -25002 -209 -19084
rect -6207 -25042 -209 -25002
rect 110 -19084 6108 -19044
rect 110 -25002 150 -19084
rect 6068 -25002 6108 -19084
rect 110 -25042 6108 -25002
rect 6427 -19084 12425 -19044
rect 6427 -25002 6467 -19084
rect 12385 -25002 12425 -19084
rect 6427 -25042 12425 -25002
<< mimcapcontact >>
rect -12484 19084 -6566 25002
rect -6167 19084 -249 25002
rect 150 19084 6068 25002
rect 6467 19084 12385 25002
rect -12484 12786 -6566 18704
rect -6167 12786 -249 18704
rect 150 12786 6068 18704
rect 6467 12786 12385 18704
rect -12484 6488 -6566 12406
rect -6167 6488 -249 12406
rect 150 6488 6068 12406
rect 6467 6488 12385 12406
rect -12484 190 -6566 6108
rect -6167 190 -249 6108
rect 150 190 6068 6108
rect 6467 190 12385 6108
rect -12484 -6108 -6566 -190
rect -6167 -6108 -249 -190
rect 150 -6108 6068 -190
rect 6467 -6108 12385 -190
rect -12484 -12406 -6566 -6488
rect -6167 -12406 -249 -6488
rect 150 -12406 6068 -6488
rect 6467 -12406 12385 -6488
rect -12484 -18704 -6566 -12786
rect -6167 -18704 -249 -12786
rect 150 -18704 6068 -12786
rect 6467 -18704 12385 -12786
rect -12484 -25002 -6566 -19084
rect -6167 -25002 -249 -19084
rect 150 -25002 6068 -19084
rect 6467 -25002 12385 -19084
<< metal4 >>
rect -9577 25003 -9473 25192
rect -6458 25130 -6354 25192
rect -6458 25114 -6331 25130
rect -12485 25002 -6565 25003
rect -12485 19084 -12484 25002
rect -6566 19084 -6565 25002
rect -12485 19083 -6565 19084
rect -9577 18705 -9473 19083
rect -6458 18972 -6411 25114
rect -6347 18972 -6331 25114
rect -3260 25003 -3156 25192
rect -141 25130 -37 25192
rect -141 25114 -14 25130
rect -6168 25002 -248 25003
rect -6168 19084 -6167 25002
rect -249 19084 -248 25002
rect -6168 19083 -248 19084
rect -6458 18956 -6331 18972
rect -6458 18832 -6354 18956
rect -6458 18816 -6331 18832
rect -12485 18704 -6565 18705
rect -12485 12786 -12484 18704
rect -6566 12786 -6565 18704
rect -12485 12785 -6565 12786
rect -9577 12407 -9473 12785
rect -6458 12674 -6411 18816
rect -6347 12674 -6331 18816
rect -3260 18705 -3156 19083
rect -141 18972 -94 25114
rect -30 18972 -14 25114
rect 3057 25003 3161 25192
rect 6176 25130 6280 25192
rect 6176 25114 6303 25130
rect 149 25002 6069 25003
rect 149 19084 150 25002
rect 6068 19084 6069 25002
rect 149 19083 6069 19084
rect -141 18956 -14 18972
rect -141 18832 -37 18956
rect -141 18816 -14 18832
rect -6168 18704 -248 18705
rect -6168 12786 -6167 18704
rect -249 12786 -248 18704
rect -6168 12785 -248 12786
rect -6458 12658 -6331 12674
rect -6458 12534 -6354 12658
rect -6458 12518 -6331 12534
rect -12485 12406 -6565 12407
rect -12485 6488 -12484 12406
rect -6566 6488 -6565 12406
rect -12485 6487 -6565 6488
rect -9577 6109 -9473 6487
rect -6458 6376 -6411 12518
rect -6347 6376 -6331 12518
rect -3260 12407 -3156 12785
rect -141 12674 -94 18816
rect -30 12674 -14 18816
rect 3057 18705 3161 19083
rect 6176 18972 6223 25114
rect 6287 18972 6303 25114
rect 9374 25003 9478 25192
rect 12493 25130 12597 25192
rect 12493 25114 12620 25130
rect 6466 25002 12386 25003
rect 6466 19084 6467 25002
rect 12385 19084 12386 25002
rect 6466 19083 12386 19084
rect 6176 18956 6303 18972
rect 6176 18832 6280 18956
rect 6176 18816 6303 18832
rect 149 18704 6069 18705
rect 149 12786 150 18704
rect 6068 12786 6069 18704
rect 149 12785 6069 12786
rect -141 12658 -14 12674
rect -141 12534 -37 12658
rect -141 12518 -14 12534
rect -6168 12406 -248 12407
rect -6168 6488 -6167 12406
rect -249 6488 -248 12406
rect -6168 6487 -248 6488
rect -6458 6360 -6331 6376
rect -6458 6236 -6354 6360
rect -6458 6220 -6331 6236
rect -12485 6108 -6565 6109
rect -12485 190 -12484 6108
rect -6566 190 -6565 6108
rect -12485 189 -6565 190
rect -9577 -189 -9473 189
rect -6458 78 -6411 6220
rect -6347 78 -6331 6220
rect -3260 6109 -3156 6487
rect -141 6376 -94 12518
rect -30 6376 -14 12518
rect 3057 12407 3161 12785
rect 6176 12674 6223 18816
rect 6287 12674 6303 18816
rect 9374 18705 9478 19083
rect 12493 18972 12540 25114
rect 12604 18972 12620 25114
rect 12493 18956 12620 18972
rect 12493 18832 12597 18956
rect 12493 18816 12620 18832
rect 6466 18704 12386 18705
rect 6466 12786 6467 18704
rect 12385 12786 12386 18704
rect 6466 12785 12386 12786
rect 6176 12658 6303 12674
rect 6176 12534 6280 12658
rect 6176 12518 6303 12534
rect 149 12406 6069 12407
rect 149 6488 150 12406
rect 6068 6488 6069 12406
rect 149 6487 6069 6488
rect -141 6360 -14 6376
rect -141 6236 -37 6360
rect -141 6220 -14 6236
rect -6168 6108 -248 6109
rect -6168 190 -6167 6108
rect -249 190 -248 6108
rect -6168 189 -248 190
rect -6458 62 -6331 78
rect -6458 -62 -6354 62
rect -6458 -78 -6331 -62
rect -12485 -190 -6565 -189
rect -12485 -6108 -12484 -190
rect -6566 -6108 -6565 -190
rect -12485 -6109 -6565 -6108
rect -9577 -6487 -9473 -6109
rect -6458 -6220 -6411 -78
rect -6347 -6220 -6331 -78
rect -3260 -189 -3156 189
rect -141 78 -94 6220
rect -30 78 -14 6220
rect 3057 6109 3161 6487
rect 6176 6376 6223 12518
rect 6287 6376 6303 12518
rect 9374 12407 9478 12785
rect 12493 12674 12540 18816
rect 12604 12674 12620 18816
rect 12493 12658 12620 12674
rect 12493 12534 12597 12658
rect 12493 12518 12620 12534
rect 6466 12406 12386 12407
rect 6466 6488 6467 12406
rect 12385 6488 12386 12406
rect 6466 6487 12386 6488
rect 6176 6360 6303 6376
rect 6176 6236 6280 6360
rect 6176 6220 6303 6236
rect 149 6108 6069 6109
rect 149 190 150 6108
rect 6068 190 6069 6108
rect 149 189 6069 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -6168 -190 -248 -189
rect -6168 -6108 -6167 -190
rect -249 -6108 -248 -190
rect -6168 -6109 -248 -6108
rect -6458 -6236 -6331 -6220
rect -6458 -6360 -6354 -6236
rect -6458 -6376 -6331 -6360
rect -12485 -6488 -6565 -6487
rect -12485 -12406 -12484 -6488
rect -6566 -12406 -6565 -6488
rect -12485 -12407 -6565 -12406
rect -9577 -12785 -9473 -12407
rect -6458 -12518 -6411 -6376
rect -6347 -12518 -6331 -6376
rect -3260 -6487 -3156 -6109
rect -141 -6220 -94 -78
rect -30 -6220 -14 -78
rect 3057 -189 3161 189
rect 6176 78 6223 6220
rect 6287 78 6303 6220
rect 9374 6109 9478 6487
rect 12493 6376 12540 12518
rect 12604 6376 12620 12518
rect 12493 6360 12620 6376
rect 12493 6236 12597 6360
rect 12493 6220 12620 6236
rect 6466 6108 12386 6109
rect 6466 190 6467 6108
rect 12385 190 12386 6108
rect 6466 189 12386 190
rect 6176 62 6303 78
rect 6176 -62 6280 62
rect 6176 -78 6303 -62
rect 149 -190 6069 -189
rect 149 -6108 150 -190
rect 6068 -6108 6069 -190
rect 149 -6109 6069 -6108
rect -141 -6236 -14 -6220
rect -141 -6360 -37 -6236
rect -141 -6376 -14 -6360
rect -6168 -6488 -248 -6487
rect -6168 -12406 -6167 -6488
rect -249 -12406 -248 -6488
rect -6168 -12407 -248 -12406
rect -6458 -12534 -6331 -12518
rect -6458 -12658 -6354 -12534
rect -6458 -12674 -6331 -12658
rect -12485 -12786 -6565 -12785
rect -12485 -18704 -12484 -12786
rect -6566 -18704 -6565 -12786
rect -12485 -18705 -6565 -18704
rect -9577 -19083 -9473 -18705
rect -6458 -18816 -6411 -12674
rect -6347 -18816 -6331 -12674
rect -3260 -12785 -3156 -12407
rect -141 -12518 -94 -6376
rect -30 -12518 -14 -6376
rect 3057 -6487 3161 -6109
rect 6176 -6220 6223 -78
rect 6287 -6220 6303 -78
rect 9374 -189 9478 189
rect 12493 78 12540 6220
rect 12604 78 12620 6220
rect 12493 62 12620 78
rect 12493 -62 12597 62
rect 12493 -78 12620 -62
rect 6466 -190 12386 -189
rect 6466 -6108 6467 -190
rect 12385 -6108 12386 -190
rect 6466 -6109 12386 -6108
rect 6176 -6236 6303 -6220
rect 6176 -6360 6280 -6236
rect 6176 -6376 6303 -6360
rect 149 -6488 6069 -6487
rect 149 -12406 150 -6488
rect 6068 -12406 6069 -6488
rect 149 -12407 6069 -12406
rect -141 -12534 -14 -12518
rect -141 -12658 -37 -12534
rect -141 -12674 -14 -12658
rect -6168 -12786 -248 -12785
rect -6168 -18704 -6167 -12786
rect -249 -18704 -248 -12786
rect -6168 -18705 -248 -18704
rect -6458 -18832 -6331 -18816
rect -6458 -18956 -6354 -18832
rect -6458 -18972 -6331 -18956
rect -12485 -19084 -6565 -19083
rect -12485 -25002 -12484 -19084
rect -6566 -25002 -6565 -19084
rect -12485 -25003 -6565 -25002
rect -9577 -25192 -9473 -25003
rect -6458 -25114 -6411 -18972
rect -6347 -25114 -6331 -18972
rect -3260 -19083 -3156 -18705
rect -141 -18816 -94 -12674
rect -30 -18816 -14 -12674
rect 3057 -12785 3161 -12407
rect 6176 -12518 6223 -6376
rect 6287 -12518 6303 -6376
rect 9374 -6487 9478 -6109
rect 12493 -6220 12540 -78
rect 12604 -6220 12620 -78
rect 12493 -6236 12620 -6220
rect 12493 -6360 12597 -6236
rect 12493 -6376 12620 -6360
rect 6466 -6488 12386 -6487
rect 6466 -12406 6467 -6488
rect 12385 -12406 12386 -6488
rect 6466 -12407 12386 -12406
rect 6176 -12534 6303 -12518
rect 6176 -12658 6280 -12534
rect 6176 -12674 6303 -12658
rect 149 -12786 6069 -12785
rect 149 -18704 150 -12786
rect 6068 -18704 6069 -12786
rect 149 -18705 6069 -18704
rect -141 -18832 -14 -18816
rect -141 -18956 -37 -18832
rect -141 -18972 -14 -18956
rect -6168 -19084 -248 -19083
rect -6168 -25002 -6167 -19084
rect -249 -25002 -248 -19084
rect -6168 -25003 -248 -25002
rect -6458 -25130 -6331 -25114
rect -6458 -25192 -6354 -25130
rect -3260 -25192 -3156 -25003
rect -141 -25114 -94 -18972
rect -30 -25114 -14 -18972
rect 3057 -19083 3161 -18705
rect 6176 -18816 6223 -12674
rect 6287 -18816 6303 -12674
rect 9374 -12785 9478 -12407
rect 12493 -12518 12540 -6376
rect 12604 -12518 12620 -6376
rect 12493 -12534 12620 -12518
rect 12493 -12658 12597 -12534
rect 12493 -12674 12620 -12658
rect 6466 -12786 12386 -12785
rect 6466 -18704 6467 -12786
rect 12385 -18704 12386 -12786
rect 6466 -18705 12386 -18704
rect 6176 -18832 6303 -18816
rect 6176 -18956 6280 -18832
rect 6176 -18972 6303 -18956
rect 149 -19084 6069 -19083
rect 149 -25002 150 -19084
rect 6068 -25002 6069 -19084
rect 149 -25003 6069 -25002
rect -141 -25130 -14 -25114
rect -141 -25192 -37 -25130
rect 3057 -25192 3161 -25003
rect 6176 -25114 6223 -18972
rect 6287 -25114 6303 -18972
rect 9374 -19083 9478 -18705
rect 12493 -18816 12540 -12674
rect 12604 -18816 12620 -12674
rect 12493 -18832 12620 -18816
rect 12493 -18956 12597 -18832
rect 12493 -18972 12620 -18956
rect 6466 -19084 12386 -19083
rect 6466 -25002 6467 -19084
rect 12385 -25002 12386 -19084
rect 6466 -25003 12386 -25002
rect 6176 -25130 6303 -25114
rect 6176 -25192 6280 -25130
rect 9374 -25192 9478 -25003
rect 12493 -25114 12540 -18972
rect 12604 -25114 12620 -18972
rect 12493 -25130 12620 -25114
rect 12493 -25192 12597 -25130
<< properties >>
string FIXED_BBOX 6327 18944 12525 25142
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 29.993 l 29.993 val 1.821k carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
