* NGSPICE file created from esd_cell.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_BRTJC6 a_n345_n500# a_1135_n588# a_n603_n588#
+ a_n1393_n588# a_n1609_n500# a_661_n588# a_n1135_n500# a_n977_n500# a_1293_n588#
+ a_n761_n588# a_n503_n500# a_n1551_n588# a_129_n500# a_n1293_n500# a_287_n500# a_n661_n500#
+ a_1451_n588# a_n1451_n500# a_919_n500# a_445_n500# a_1077_n500# a_29_n588# a_n129_n588#
+ a_603_n500# a_187_n588# a_1235_n500# a_n287_n588# a_761_n500# a_819_n588# a_345_n588#
+ a_n1077_n588# a_n29_n500# a_1393_n500# a_n919_n588# a_n1743_n722# a_n187_n500# a_977_n588#
+ a_n445_n588# a_503_n588# a_n1235_n588# a_1551_n500# a_n819_n500#
X0 a_n819_n500# a_n919_n588# a_n977_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n588# a_n819_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n588# a_761_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n588# a_n345_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n588# a_603_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n588# a_129_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n588# a_n1451_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n588# a_1235_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n588# a_n503_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n588# a_n29_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n588# a_287_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n588# a_n1609_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n588# a_1393_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n588# a_n1135_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_n503_n500# a_n603_n588# a_n661_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_1077_n500# a_977_n588# a_919_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n588# a_n187_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n588# a_445_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n588# a_n1293_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n588# a_1077_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_1551_n500# a_1393_n500# 0.56fF
C1 a_1551_n500# a_1235_n500# 0.24fF
C2 a_1235_n500# a_1393_n500# 0.56fF
C3 a_1551_n500# a_1077_n500# 0.15fF
C4 a_1077_n500# a_1393_n500# 0.24fF
C5 a_1551_n500# a_919_n500# 0.11fF
C6 a_1393_n500# a_919_n500# 0.15fF
C7 a_1235_n500# a_1077_n500# 0.56fF
C8 a_1235_n500# a_919_n500# 0.24fF
C9 a_603_n500# a_1551_n500# 0.07fF
C10 a_761_n500# a_1551_n500# 0.09fF
C11 a_1077_n500# a_919_n500# 0.56fF
C12 a_603_n500# a_1393_n500# 0.09fF
C13 a_761_n500# a_1393_n500# 0.11fF
C14 a_445_n500# a_1551_n500# 0.06fF
C15 a_445_n500# a_1393_n500# 0.07fF
C16 a_603_n500# a_1235_n500# 0.11fF
C17 a_761_n500# a_1235_n500# 0.15fF
C18 a_445_n500# a_1235_n500# 0.09fF
C19 a_1551_n500# a_287_n500# 0.05fF
C20 a_287_n500# a_1393_n500# 0.06fF
C21 a_603_n500# a_1077_n500# 0.15fF
C22 a_761_n500# a_1077_n500# 0.24fF
C23 a_1551_n500# a_n29_n500# 0.04fF
C24 a_445_n500# a_1077_n500# 0.11fF
C25 a_n29_n500# a_1393_n500# 0.05fF
C26 a_603_n500# a_919_n500# 0.24fF
C27 a_129_n500# a_1551_n500# 0.05fF
C28 a_761_n500# a_919_n500# 0.56fF
C29 a_129_n500# a_1393_n500# 0.05fF
C30 a_1235_n500# a_287_n500# 0.07fF
C31 a_445_n500# a_919_n500# 0.15fF
C32 a_n187_n500# a_1393_n500# 0.04fF
C33 a_n29_n500# a_1235_n500# 0.05fF
C34 a_287_n500# a_1077_n500# 0.09fF
C35 a_129_n500# a_1235_n500# 0.06fF
C36 a_287_n500# a_919_n500# 0.11fF
C37 a_n187_n500# a_1235_n500# 0.05fF
C38 a_n29_n500# a_1077_n500# 0.06fF
C39 a_n345_n500# a_1235_n500# 0.04fF
C40 a_761_n500# a_603_n500# 0.56fF
C41 a_129_n500# a_1077_n500# 0.07fF
C42 a_n29_n500# a_919_n500# 0.07fF
C43 a_445_n500# a_603_n500# 0.56fF
C44 a_761_n500# a_445_n500# 0.24fF
C45 a_n187_n500# a_1077_n500# 0.05fF
C46 a_129_n500# a_919_n500# 0.09fF
C47 a_n345_n500# a_1077_n500# 0.05fF
C48 a_n503_n500# a_1077_n500# 0.04fF
C49 a_n187_n500# a_919_n500# 0.06fF
C50 a_n345_n500# a_919_n500# 0.05fF
C51 a_n503_n500# a_919_n500# 0.05fF
C52 a_603_n500# a_287_n500# 0.24fF
C53 a_761_n500# a_287_n500# 0.15fF
C54 a_445_n500# a_287_n500# 0.56fF
C55 a_603_n500# a_n29_n500# 0.11fF
C56 a_761_n500# a_n29_n500# 0.09fF
C57 a_603_n500# a_129_n500# 0.15fF
C58 a_445_n500# a_n29_n500# 0.15fF
C59 a_761_n500# a_129_n500# 0.11fF
C60 a_445_n500# a_129_n500# 0.24fF
C61 a_603_n500# a_n187_n500# 0.09fF
C62 a_761_n500# a_n187_n500# 0.07fF
C63 a_n661_n500# a_919_n500# 0.04fF
C64 a_603_n500# a_n345_n500# 0.07fF
C65 a_603_n500# a_n503_n500# 0.06fF
C66 a_445_n500# a_n187_n500# 0.11fF
C67 a_761_n500# a_n503_n500# 0.05fF
C68 a_761_n500# a_n345_n500# 0.06fF
C69 a_445_n500# a_n345_n500# 0.09fF
C70 a_445_n500# a_n503_n500# 0.07fF
C71 a_n29_n500# a_287_n500# 0.24fF
C72 a_129_n500# a_287_n500# 0.56fF
C73 a_n187_n500# a_287_n500# 0.15fF
C74 a_129_n500# a_n29_n500# 0.56fF
C75 a_n345_n500# a_287_n500# 0.11fF
C76 a_n503_n500# a_287_n500# 0.09fF
C77 a_n661_n500# a_603_n500# 0.05fF
C78 a_n187_n500# a_n29_n500# 0.56fF
C79 a_n661_n500# a_761_n500# 0.05fF
C80 a_n345_n500# a_n29_n500# 0.24fF
C81 a_n29_n500# a_n503_n500# 0.15fF
C82 a_n187_n500# a_129_n500# 0.24fF
C83 a_n661_n500# a_445_n500# 0.06fF
C84 a_129_n500# a_n345_n500# 0.15fF
C85 a_129_n500# a_n503_n500# 0.11fF
C86 a_603_n500# a_n977_n500# 0.04fF
C87 a_n187_n500# a_n345_n500# 0.56fF
C88 a_603_n500# a_n819_n500# 0.05fF
C89 a_445_n500# a_n977_n500# 0.05fF
C90 a_n187_n500# a_n503_n500# 0.24fF
C91 a_761_n500# a_n819_n500# 0.04fF
C92 a_n345_n500# a_n503_n500# 0.56fF
C93 a_445_n500# a_n819_n500# 0.05fF
C94 a_n661_n500# a_287_n500# 0.07fF
C95 a_n661_n500# a_n29_n500# 0.11fF
C96 a_445_n500# a_n1135_n500# 0.04fF
C97 a_287_n500# a_n977_n500# 0.05fF
C98 a_n661_n500# a_129_n500# 0.09fF
C99 a_n819_n500# a_287_n500# 0.06fF
C100 a_n661_n500# a_n187_n500# 0.15fF
C101 a_n29_n500# a_n977_n500# 0.07fF
C102 a_n661_n500# a_n345_n500# 0.24fF
C103 a_n819_n500# a_n29_n500# 0.09fF
C104 a_n661_n500# a_n503_n500# 0.56fF
C105 a_129_n500# a_n977_n500# 0.06fF
C106 a_n1135_n500# a_287_n500# 0.05fF
C107 a_n187_n500# a_n977_n500# 0.09fF
C108 a_129_n500# a_n819_n500# 0.07fF
C109 a_n29_n500# a_n1135_n500# 0.06fF
C110 a_n345_n500# a_n977_n500# 0.11fF
C111 a_n187_n500# a_n819_n500# 0.11fF
C112 a_n503_n500# a_n977_n500# 0.15fF
C113 a_129_n500# a_n1135_n500# 0.05fF
C114 a_287_n500# a_n1293_n500# 0.04fF
C115 a_n345_n500# a_n819_n500# 0.15fF
C116 a_n819_n500# a_n503_n500# 0.24fF
C117 a_n29_n500# a_n1451_n500# 0.05fF
C118 a_n187_n500# a_n1135_n500# 0.07fF
C119 a_n29_n500# a_n1293_n500# 0.05fF
C120 a_n345_n500# a_n1135_n500# 0.09fF
C121 a_129_n500# a_n1451_n500# 0.04fF
C122 a_n29_n500# a_n1609_n500# 0.04fF
C123 a_n1135_n500# a_n503_n500# 0.11fF
C124 a_129_n500# a_n1293_n500# 0.05fF
C125 a_n187_n500# a_n1451_n500# 0.05fF
C126 a_n187_n500# a_n1293_n500# 0.06fF
C127 a_n345_n500# a_n1451_n500# 0.06fF
C128 a_n661_n500# a_n977_n500# 0.24fF
C129 a_n345_n500# a_n1293_n500# 0.07fF
C130 a_n503_n500# a_n1451_n500# 0.07fF
C131 a_n187_n500# a_n1609_n500# 0.05fF
C132 a_n503_n500# a_n1293_n500# 0.09fF
C133 a_n345_n500# a_n1609_n500# 0.05fF
C134 a_n1609_n500# a_n503_n500# 0.06fF
C135 a_n661_n500# a_n819_n500# 0.56fF
C136 a_n661_n500# a_n1135_n500# 0.15fF
C137 a_n819_n500# a_n977_n500# 0.56fF
C138 a_n661_n500# a_n1451_n500# 0.09fF
C139 a_n1135_n500# a_n977_n500# 0.56fF
C140 a_n661_n500# a_n1293_n500# 0.11fF
C141 a_n819_n500# a_n1135_n500# 0.24fF
C142 a_n661_n500# a_n1609_n500# 0.07fF
C143 a_n1451_n500# a_n977_n500# 0.15fF
C144 a_n1293_n500# a_n977_n500# 0.24fF
C145 a_n819_n500# a_n1451_n500# 0.11fF
C146 a_n1609_n500# a_n977_n500# 0.11fF
C147 a_n819_n500# a_n1293_n500# 0.15fF
C148 a_n819_n500# a_n1609_n500# 0.09fF
C149 a_n1135_n500# a_n1451_n500# 0.24fF
C150 a_n1135_n500# a_n1293_n500# 0.56fF
C151 a_n1135_n500# a_n1609_n500# 0.15fF
C152 a_n1293_n500# a_n1451_n500# 0.56fF
C153 a_n1609_n500# a_n1451_n500# 0.56fF
C154 a_n1609_n500# a_n1293_n500# 0.24fF
C155 a_1451_n588# a_1135_n588# 0.04fF
C156 a_1451_n588# a_1293_n588# 0.12fF
C157 a_1451_n588# a_977_n588# 0.02fF
C158 a_1135_n588# a_1293_n588# 0.12fF
C159 a_819_n588# a_1451_n588# 0.02fF
C160 a_1135_n588# a_977_n588# 0.12fF
C161 a_1293_n588# a_977_n588# 0.04fF
C162 a_819_n588# a_1135_n588# 0.04fF
C163 a_819_n588# a_1293_n588# 0.02fF
C164 a_819_n588# a_977_n588# 0.12fF
C165 a_1451_n588# a_503_n588# 0.01fF
C166 a_1451_n588# a_661_n588# 0.01fF
C167 a_1135_n588# a_503_n588# 0.02fF
C168 a_1293_n588# a_503_n588# 0.01fF
C169 a_1135_n588# a_661_n588# 0.02fF
C170 a_661_n588# a_1293_n588# 0.02fF
C171 a_977_n588# a_503_n588# 0.02fF
C172 a_661_n588# a_977_n588# 0.04fF
C173 a_819_n588# a_503_n588# 0.04fF
C174 a_819_n588# a_661_n588# 0.12fF
C175 a_1451_n588# a_345_n588# 0.01fF
C176 a_187_n588# a_1451_n588# 0.01fF
C177 a_1451_n588# a_29_n588# 0.01fF
C178 a_1135_n588# a_345_n588# 0.01fF
C179 a_1451_n588# a_n129_n588# 0.01fF
C180 a_187_n588# a_1135_n588# 0.01fF
C181 a_345_n588# a_1293_n588# 0.01fF
C182 a_187_n588# a_1293_n588# 0.01fF
C183 a_1135_n588# a_29_n588# 0.01fF
C184 a_345_n588# a_977_n588# 0.02fF
C185 a_1293_n588# a_29_n588# 0.01fF
C186 a_661_n588# a_503_n588# 0.12fF
C187 a_187_n588# a_977_n588# 0.01fF
C188 a_29_n588# a_977_n588# 0.01fF
C189 a_n129_n588# a_1135_n588# 0.01fF
C190 a_n129_n588# a_1293_n588# 0.01fF
C191 a_n445_n588# a_1135_n588# 0.01fF
C192 a_819_n588# a_345_n588# 0.02fF
C193 a_n129_n588# a_977_n588# 0.01fF
C194 a_187_n588# a_819_n588# 0.02fF
C195 a_1135_n588# a_n287_n588# 0.01fF
C196 a_1293_n588# a_n287_n588# 0.01fF
C197 a_819_n588# a_29_n588# 0.01fF
C198 a_n445_n588# a_977_n588# 0.01fF
C199 a_n287_n588# a_977_n588# 0.01fF
C200 a_819_n588# a_n129_n588# 0.01fF
C201 a_n603_n588# a_977_n588# 0.01fF
C202 a_819_n588# a_n445_n588# 0.01fF
C203 a_819_n588# a_n287_n588# 0.01fF
C204 a_345_n588# a_503_n588# 0.12fF
C205 a_187_n588# a_503_n588# 0.04fF
C206 a_345_n588# a_661_n588# 0.04fF
C207 a_187_n588# a_661_n588# 0.02fF
C208 a_29_n588# a_503_n588# 0.02fF
C209 a_819_n588# a_n603_n588# 0.01fF
C210 a_661_n588# a_29_n588# 0.02fF
C211 a_n129_n588# a_503_n588# 0.02fF
C212 a_n129_n588# a_661_n588# 0.01fF
C213 a_819_n588# a_n761_n588# 0.01fF
C214 a_n445_n588# a_503_n588# 0.01fF
C215 a_n445_n588# a_661_n588# 0.01fF
C216 a_n287_n588# a_503_n588# 0.01fF
C217 a_661_n588# a_n287_n588# 0.01fF
C218 a_n603_n588# a_503_n588# 0.01fF
C219 a_661_n588# a_n603_n588# 0.01fF
C220 a_187_n588# a_345_n588# 0.12fF
C221 a_503_n588# a_n761_n588# 0.01fF
C222 a_661_n588# a_n761_n588# 0.01fF
C223 a_345_n588# a_29_n588# 0.04fF
C224 a_187_n588# a_29_n588# 0.12fF
C225 a_n919_n588# a_503_n588# 0.01fF
C226 a_661_n588# a_n919_n588# 0.01fF
C227 a_n129_n588# a_345_n588# 0.02fF
C228 a_187_n588# a_n129_n588# 0.04fF
C229 a_n129_n588# a_29_n588# 0.12fF
C230 a_n445_n588# a_345_n588# 0.01fF
C231 a_187_n588# a_n445_n588# 0.02fF
C232 a_n445_n588# a_29_n588# 0.02fF
C233 a_345_n588# a_n287_n588# 0.02fF
C234 a_187_n588# a_n287_n588# 0.02fF
C235 a_29_n588# a_n287_n588# 0.04fF
C236 a_345_n588# a_n603_n588# 0.01fF
C237 a_187_n588# a_n603_n588# 0.01fF
C238 a_n1077_n588# a_503_n588# 0.01fF
C239 a_n603_n588# a_29_n588# 0.02fF
C240 a_n445_n588# a_n129_n588# 0.04fF
C241 a_n129_n588# a_n287_n588# 0.12fF
C242 a_345_n588# a_n761_n588# 0.01fF
C243 a_187_n588# a_n761_n588# 0.01fF
C244 a_n445_n588# a_n287_n588# 0.12fF
C245 a_29_n588# a_n761_n588# 0.01fF
C246 a_n129_n588# a_n603_n588# 0.02fF
C247 a_345_n588# a_n919_n588# 0.01fF
C248 a_187_n588# a_n919_n588# 0.01fF
C249 a_n445_n588# a_n603_n588# 0.12fF
C250 a_n919_n588# a_29_n588# 0.01fF
C251 a_n603_n588# a_n287_n588# 0.04fF
C252 a_n129_n588# a_n761_n588# 0.02fF
C253 a_n445_n588# a_n761_n588# 0.04fF
C254 a_n129_n588# a_n919_n588# 0.01fF
C255 a_n287_n588# a_n761_n588# 0.02fF
C256 a_n445_n588# a_n919_n588# 0.02fF
C257 a_n919_n588# a_n287_n588# 0.02fF
C258 a_345_n588# a_n1077_n588# 0.01fF
C259 a_n603_n588# a_n761_n588# 0.12fF
C260 a_187_n588# a_n1077_n588# 0.01fF
C261 a_n919_n588# a_n603_n588# 0.04fF
C262 a_n1077_n588# a_29_n588# 0.01fF
C263 a_345_n588# a_n1235_n588# 0.01fF
C264 a_187_n588# a_n1235_n588# 0.01fF
C265 a_n129_n588# a_n1077_n588# 0.01fF
C266 a_n919_n588# a_n761_n588# 0.12fF
C267 a_n1235_n588# a_29_n588# 0.01fF
C268 a_n445_n588# a_n1077_n588# 0.02fF
C269 a_n129_n588# a_n1235_n588# 0.01fF
C270 a_n1077_n588# a_n287_n588# 0.01fF
C271 a_187_n588# a_n1393_n588# 0.01fF
C272 a_29_n588# a_n1393_n588# 0.01fF
C273 a_n445_n588# a_n1235_n588# 0.01fF
C274 a_n1077_n588# a_n603_n588# 0.02fF
C275 a_n1551_n588# a_29_n588# 0.01fF
C276 a_n1235_n588# a_n287_n588# 0.01fF
C277 a_n129_n588# a_n1393_n588# 0.01fF
C278 a_n1235_n588# a_n603_n588# 0.02fF
C279 a_n1551_n588# a_n129_n588# 0.01fF
C280 a_n1077_n588# a_n761_n588# 0.04fF
C281 a_n445_n588# a_n1393_n588# 0.01fF
C282 a_n1551_n588# a_n445_n588# 0.01fF
C283 a_n919_n588# a_n1077_n588# 0.12fF
C284 a_n1551_n588# a_n287_n588# 0.01fF
C285 a_n287_n588# a_n1393_n588# 0.01fF
C286 a_n1235_n588# a_n761_n588# 0.02fF
C287 a_n603_n588# a_n1393_n588# 0.01fF
C288 a_n1551_n588# a_n603_n588# 0.01fF
C289 a_n919_n588# a_n1235_n588# 0.04fF
C290 a_n1393_n588# a_n761_n588# 0.02fF
C291 a_n1551_n588# a_n761_n588# 0.01fF
C292 a_n919_n588# a_n1393_n588# 0.02fF
C293 a_n1551_n588# a_n919_n588# 0.02fF
C294 a_n1077_n588# a_n1235_n588# 0.12fF
C295 a_n1077_n588# a_n1393_n588# 0.04fF
C296 a_n1551_n588# a_n1077_n588# 0.02fF
C297 a_n1235_n588# a_n1393_n588# 0.12fF
C298 a_n1551_n588# a_n1235_n588# 0.04fF
C299 a_n1551_n588# a_n1393_n588# 0.12fF
C300 a_1551_n500# a_n1743_n722# 0.30fF
C301 a_1393_n500# a_n1743_n722# 0.13fF
C302 a_1235_n500# a_n1743_n722# 0.09fF
C303 a_1077_n500# a_n1743_n722# 0.07fF
C304 a_919_n500# a_n1743_n722# 0.06fF
C305 a_761_n500# a_n1743_n722# 0.05fF
C306 a_603_n500# a_n1743_n722# 0.05fF
C307 a_445_n500# a_n1743_n722# 0.04fF
C308 a_287_n500# a_n1743_n722# 0.04fF
C309 a_129_n500# a_n1743_n722# 0.04fF
C310 a_n29_n500# a_n1743_n722# 0.02fF
C311 a_n187_n500# a_n1743_n722# 0.04fF
C312 a_n345_n500# a_n1743_n722# 0.04fF
C313 a_n503_n500# a_n1743_n722# 0.04fF
C314 a_n661_n500# a_n1743_n722# 0.05fF
C315 a_n819_n500# a_n1743_n722# 0.05fF
C316 a_n977_n500# a_n1743_n722# 0.06fF
C317 a_n1135_n500# a_n1743_n722# 0.07fF
C318 a_n1293_n500# a_n1743_n722# 0.09fF
C319 a_n1451_n500# a_n1743_n722# 0.13fF
C320 a_n1609_n500# a_n1743_n722# 0.30fF
C321 a_1451_n588# a_n1743_n722# 0.28fF
C322 a_1293_n588# a_n1743_n722# 0.23fF
C323 a_1135_n588# a_n1743_n722# 0.24fF
C324 a_977_n588# a_n1743_n722# 0.25fF
C325 a_819_n588# a_n1743_n722# 0.26fF
C326 a_661_n588# a_n1743_n722# 0.26fF
C327 a_503_n588# a_n1743_n722# 0.27fF
C328 a_345_n588# a_n1743_n722# 0.28fF
C329 a_187_n588# a_n1743_n722# 0.28fF
C330 a_29_n588# a_n1743_n722# 0.28fF
C331 a_n129_n588# a_n1743_n722# 0.28fF
C332 a_n287_n588# a_n1743_n722# 0.28fF
C333 a_n445_n588# a_n1743_n722# 0.28fF
C334 a_n603_n588# a_n1743_n722# 0.28fF
C335 a_n761_n588# a_n1743_n722# 0.28fF
C336 a_n919_n588# a_n1743_n722# 0.28fF
C337 a_n1077_n588# a_n1743_n722# 0.28fF
C338 a_n1235_n588# a_n1743_n722# 0.29fF
C339 a_n1393_n588# a_n1743_n722# 0.29fF
C340 a_n1551_n588# a_n1743_n722# 0.34fF
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CADZ46 a_n345_n500# a_n1609_n500# a_n1135_n500#
+ a_29_n597# a_n977_n500# a_n129_n597# a_187_n597# a_n503_n500# a_129_n500# a_n1293_n500#
+ a_n287_n597# a_819_n597# a_n1077_n597# a_287_n500# a_n661_n500# a_345_n597# a_n919_n597#
+ a_n1451_n500# a_977_n597# a_n445_n597# a_919_n500# a_n1235_n597# a_445_n500# a_503_n597#
+ w_n1809_n797# a_n603_n597# a_1077_n500# a_1135_n597# a_661_n597# a_n1393_n597# a_603_n500#
+ a_1293_n597# a_n761_n597# a_1235_n500# a_n1551_n597# a_761_n500# a_n29_n500# a_1451_n597#
+ a_1393_n500# a_n187_n500# a_1551_n500# a_n819_n500# VSUBS
X0 a_n819_n500# a_n919_n597# a_n977_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n597# a_n819_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n597# a_761_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n597# a_n345_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n597# a_603_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n597# a_129_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n597# a_n1451_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n597# a_1235_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n597# a_n503_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n597# a_n29_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n597# a_287_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n597# a_n1609_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n597# a_1393_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n597# a_n1135_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_1077_n500# a_977_n597# a_919_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X15 a_n503_n500# a_n603_n597# a_n661_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n597# a_n187_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n597# a_445_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n597# a_n1293_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n597# a_1077_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_n1077_n597# a_n445_n597# 0.02fF
C1 a_n1077_n597# a_n603_n597# 0.02fF
C2 w_n1809_n797# a_129_n500# 0.04fF
C3 a_n1077_n597# a_n761_n597# 0.04fF
C4 a_n1077_n597# a_n919_n597# 0.12fF
C5 a_n29_n500# w_n1809_n797# 0.02fF
C6 w_n1809_n797# a_n187_n500# 0.04fF
C7 a_n345_n500# w_n1809_n797# 0.04fF
C8 a_n503_n500# w_n1809_n797# 0.04fF
C9 w_n1809_n797# a_n819_n500# 0.05fF
C10 w_n1809_n797# a_n661_n500# 0.05fF
C11 a_n977_n500# w_n1809_n797# 0.06fF
C12 a_n1135_n500# w_n1809_n797# 0.07fF
C13 a_n1293_n500# w_n1809_n797# 0.09fF
C14 w_n1809_n797# a_n1451_n500# 0.13fF
C15 w_n1809_n797# a_n1609_n500# 0.30fF
C16 a_1451_n597# w_n1809_n797# 0.24fF
C17 a_1293_n597# w_n1809_n797# 0.19fF
C18 a_1135_n597# w_n1809_n797# 0.20fF
C19 a_977_n597# w_n1809_n797# 0.20fF
C20 a_819_n597# w_n1809_n797# 0.21fF
C21 w_n1809_n797# a_661_n597# 0.22fF
C22 w_n1809_n797# a_503_n597# 0.23fF
C23 w_n1809_n797# a_29_n597# 0.24fF
C24 w_n1809_n797# a_187_n597# 0.24fF
C25 a_n129_n597# w_n1809_n797# 0.24fF
C26 a_345_n597# w_n1809_n797# 0.23fF
C27 a_29_n597# a_n1551_n597# 0.01fF
C28 a_n1393_n597# a_29_n597# 0.01fF
C29 a_n1393_n597# a_187_n597# 0.01fF
C30 a_n129_n597# a_n1551_n597# 0.01fF
C31 a_n1393_n597# a_n129_n597# 0.01fF
C32 a_n1235_n597# a_29_n597# 0.01fF
C33 a_n287_n597# w_n1809_n797# 0.24fF
C34 a_n1235_n597# a_187_n597# 0.01fF
C35 a_n129_n597# a_n1235_n597# 0.01fF
C36 a_345_n597# a_n1235_n597# 0.01fF
C37 a_n287_n597# a_n1551_n597# 0.01fF
C38 w_n1809_n797# a_n445_n597# 0.24fF
C39 w_n1809_n797# a_n603_n597# 0.24fF
C40 a_n1393_n597# a_n287_n597# 0.01fF
C41 a_n1235_n597# a_n287_n597# 0.01fF
C42 a_n1551_n597# a_n603_n597# 0.01fF
C43 a_n445_n597# a_n1551_n597# 0.01fF
C44 w_n1809_n797# a_n761_n597# 0.24fF
C45 a_n1393_n597# a_n603_n597# 0.01fF
C46 a_n1393_n597# a_n445_n597# 0.01fF
C47 a_n1235_n597# a_n603_n597# 0.02fF
C48 a_n919_n597# w_n1809_n797# 0.24fF
C49 a_n1235_n597# a_n445_n597# 0.01fF
C50 a_n1551_n597# a_n761_n597# 0.01fF
C51 a_n1393_n597# a_n761_n597# 0.02fF
C52 a_n1235_n597# a_n761_n597# 0.02fF
C53 a_n919_n597# a_n1551_n597# 0.02fF
C54 a_n1393_n597# a_n919_n597# 0.02fF
C55 a_n1077_n597# w_n1809_n797# 0.24fF
C56 a_n1235_n597# a_n919_n597# 0.04fF
C57 a_n1077_n597# a_n1551_n597# 0.02fF
C58 a_n1393_n597# a_n1077_n597# 0.04fF
C59 a_n1077_n597# a_n1235_n597# 0.12fF
C60 a_1393_n500# a_1551_n500# 0.56fF
C61 a_1551_n500# a_1235_n500# 0.24fF
C62 a_1393_n500# a_1235_n500# 0.56fF
C63 a_1551_n500# a_919_n500# 0.11fF
C64 a_1393_n500# a_919_n500# 0.15fF
C65 a_919_n500# a_1235_n500# 0.24fF
C66 a_1551_n500# a_1077_n500# 0.15fF
C67 a_1077_n500# a_1235_n500# 0.56fF
C68 a_1393_n500# a_1077_n500# 0.24fF
C69 a_1077_n500# a_919_n500# 0.56fF
C70 a_1551_n500# a_445_n500# 0.06fF
C71 a_445_n500# a_1235_n500# 0.09fF
C72 a_1393_n500# a_445_n500# 0.07fF
C73 a_1551_n500# a_287_n500# 0.05fF
C74 a_1551_n500# a_603_n500# 0.07fF
C75 a_1393_n500# a_287_n500# 0.06fF
C76 a_287_n500# a_1235_n500# 0.07fF
C77 a_919_n500# a_445_n500# 0.15fF
C78 a_1551_n500# a_761_n500# 0.09fF
C79 a_1077_n500# a_445_n500# 0.11fF
C80 a_1393_n500# a_603_n500# 0.09fF
C81 a_287_n500# a_919_n500# 0.11fF
C82 a_1235_n500# a_603_n500# 0.11fF
C83 a_919_n500# a_603_n500# 0.24fF
C84 a_1393_n500# a_761_n500# 0.11fF
C85 a_287_n500# a_1077_n500# 0.09fF
C86 a_761_n500# a_1235_n500# 0.15fF
C87 a_761_n500# a_919_n500# 0.56fF
C88 a_1077_n500# a_603_n500# 0.15fF
C89 a_287_n500# a_445_n500# 0.56fF
C90 a_761_n500# a_1077_n500# 0.24fF
C91 a_445_n500# a_603_n500# 0.56fF
C92 a_761_n500# a_445_n500# 0.24fF
C93 a_287_n500# a_603_n500# 0.24fF
C94 a_761_n500# a_287_n500# 0.15fF
C95 a_761_n500# a_603_n500# 0.56fF
C96 a_1551_n500# a_129_n500# 0.05fF
C97 a_1393_n500# a_129_n500# 0.05fF
C98 a_129_n500# a_1235_n500# 0.06fF
C99 a_129_n500# a_919_n500# 0.09fF
C100 a_1077_n500# a_129_n500# 0.07fF
C101 a_129_n500# a_445_n500# 0.24fF
C102 a_287_n500# a_129_n500# 0.56fF
C103 a_n29_n500# a_1551_n500# 0.04fF
C104 a_129_n500# a_603_n500# 0.15fF
C105 a_761_n500# a_129_n500# 0.11fF
C106 a_n29_n500# a_1393_n500# 0.05fF
C107 a_n29_n500# a_1235_n500# 0.05fF
C108 a_n29_n500# a_919_n500# 0.07fF
C109 a_n29_n500# a_1077_n500# 0.06fF
C110 a_n187_n500# a_1235_n500# 0.05fF
C111 a_1393_n500# a_n187_n500# 0.04fF
C112 a_n29_n500# a_445_n500# 0.15fF
C113 a_n29_n500# a_287_n500# 0.24fF
C114 a_919_n500# a_n187_n500# 0.06fF
C115 a_n29_n500# a_603_n500# 0.11fF
C116 a_1077_n500# a_n187_n500# 0.05fF
C117 a_n29_n500# a_761_n500# 0.09fF
C118 a_n187_n500# a_445_n500# 0.11fF
C119 w_n1809_n797# a_n1551_n597# 0.30fF
C120 a_n1393_n597# w_n1809_n797# 0.25fF
C121 a_287_n500# a_n187_n500# 0.15fF
C122 a_n187_n500# a_603_n500# 0.09fF
C123 a_761_n500# a_n187_n500# 0.07fF
C124 a_n1235_n597# w_n1809_n797# 0.24fF
C125 a_n1393_n597# a_n1551_n597# 0.12fF
C126 a_n1235_n597# a_n1551_n597# 0.04fF
C127 a_n1393_n597# a_n1235_n597# 0.12fF
C128 a_n345_n500# a_1235_n500# 0.04fF
C129 a_n345_n500# a_919_n500# 0.05fF
C130 a_n29_n500# a_129_n500# 0.56fF
C131 a_n345_n500# a_1077_n500# 0.05fF
C132 a_n503_n500# a_919_n500# 0.05fF
C133 a_n503_n500# a_1077_n500# 0.04fF
C134 a_n345_n500# a_445_n500# 0.09fF
C135 a_919_n500# a_n661_n500# 0.04fF
C136 a_129_n500# a_n187_n500# 0.24fF
C137 a_n345_n500# a_287_n500# 0.11fF
C138 a_n503_n500# a_445_n500# 0.07fF
C139 a_n345_n500# a_603_n500# 0.07fF
C140 a_n503_n500# a_287_n500# 0.09fF
C141 a_445_n500# a_n661_n500# 0.06fF
C142 a_n503_n500# a_603_n500# 0.06fF
C143 a_n819_n500# a_445_n500# 0.05fF
C144 a_761_n500# a_n345_n500# 0.06fF
C145 a_761_n500# a_n503_n500# 0.05fF
C146 a_287_n500# a_n661_n500# 0.07fF
C147 a_287_n500# a_n819_n500# 0.06fF
C148 a_n819_n500# a_603_n500# 0.05fF
C149 a_n661_n500# a_603_n500# 0.05fF
C150 a_n977_n500# a_445_n500# 0.05fF
C151 a_761_n500# a_n819_n500# 0.04fF
C152 a_761_n500# a_n661_n500# 0.05fF
C153 a_n977_n500# a_287_n500# 0.05fF
C154 a_n977_n500# a_603_n500# 0.04fF
C155 a_n29_n500# a_n187_n500# 0.56fF
C156 a_n1135_n500# a_445_n500# 0.04fF
C157 a_n1135_n500# a_287_n500# 0.05fF
C158 a_n345_n500# a_129_n500# 0.15fF
C159 a_n503_n500# a_129_n500# 0.11fF
C160 a_129_n500# a_n819_n500# 0.07fF
C161 a_129_n500# a_n661_n500# 0.09fF
C162 a_n977_n500# a_129_n500# 0.06fF
C163 a_n29_n500# a_n345_n500# 0.24fF
C164 a_n29_n500# a_n503_n500# 0.15fF
C165 a_n1293_n500# a_287_n500# 0.04fF
C166 a_n1135_n500# a_129_n500# 0.05fF
C167 a_n29_n500# a_n819_n500# 0.09fF
C168 a_n29_n500# a_n661_n500# 0.11fF
C169 a_n345_n500# a_n187_n500# 0.56fF
C170 a_n503_n500# a_n187_n500# 0.24fF
C171 a_n29_n500# a_n977_n500# 0.07fF
C172 a_n819_n500# a_n187_n500# 0.11fF
C173 a_n187_n500# a_n661_n500# 0.15fF
C174 a_n29_n500# a_n1135_n500# 0.06fF
C175 a_n977_n500# a_n187_n500# 0.09fF
C176 a_n1135_n500# a_n187_n500# 0.07fF
C177 a_n1293_n500# a_129_n500# 0.05fF
C178 a_n503_n500# a_n345_n500# 0.56fF
C179 a_n345_n500# a_n661_n500# 0.24fF
C180 a_n345_n500# a_n819_n500# 0.15fF
C181 a_n503_n500# a_n819_n500# 0.24fF
C182 a_n503_n500# a_n661_n500# 0.56fF
C183 a_n29_n500# a_n1293_n500# 0.05fF
C184 a_129_n500# a_n1451_n500# 0.04fF
C185 a_n977_n500# a_n345_n500# 0.11fF
C186 a_n819_n500# a_n661_n500# 0.56fF
C187 a_n977_n500# a_n503_n500# 0.15fF
C188 a_n1293_n500# a_n187_n500# 0.06fF
C189 a_n977_n500# a_n819_n500# 0.56fF
C190 a_n977_n500# a_n661_n500# 0.24fF
C191 a_n345_n500# a_n1135_n500# 0.09fF
C192 a_n503_n500# a_n1135_n500# 0.11fF
C193 a_n29_n500# a_n1451_n500# 0.05fF
C194 a_n1135_n500# a_n819_n500# 0.24fF
C195 a_n1135_n500# a_n661_n500# 0.15fF
C196 a_n29_n500# a_n1609_n500# 0.04fF
C197 a_n977_n500# a_n1135_n500# 0.56fF
C198 a_n187_n500# a_n1451_n500# 0.05fF
C199 a_n187_n500# a_n1609_n500# 0.05fF
C200 a_n1293_n500# a_n345_n500# 0.07fF
C201 a_n1293_n500# a_n503_n500# 0.09fF
C202 a_n1293_n500# a_n819_n500# 0.15fF
C203 a_n1293_n500# a_n661_n500# 0.11fF
C204 a_n977_n500# a_n1293_n500# 0.24fF
C205 a_n345_n500# a_n1451_n500# 0.06fF
C206 a_n503_n500# a_n1451_n500# 0.07fF
C207 a_n1293_n500# a_n1135_n500# 0.56fF
C208 a_n819_n500# a_n1451_n500# 0.11fF
C209 a_n661_n500# a_n1451_n500# 0.09fF
C210 a_n345_n500# a_n1609_n500# 0.05fF
C211 a_n503_n500# a_n1609_n500# 0.06fF
C212 a_n977_n500# a_n1451_n500# 0.15fF
C213 a_n819_n500# a_n1609_n500# 0.09fF
C214 a_n1609_n500# a_n661_n500# 0.07fF
C215 a_n977_n500# a_n1609_n500# 0.11fF
C216 a_n1135_n500# a_n1451_n500# 0.24fF
C217 a_n1135_n500# a_n1609_n500# 0.15fF
C218 a_n1293_n500# a_n1451_n500# 0.56fF
C219 a_n1293_n500# a_n1609_n500# 0.24fF
C220 a_n1609_n500# a_n1451_n500# 0.56fF
C221 a_1293_n597# a_1451_n597# 0.12fF
C222 a_977_n597# a_1451_n597# 0.02fF
C223 a_1135_n597# a_1451_n597# 0.04fF
C224 a_819_n597# a_1451_n597# 0.02fF
C225 a_1451_n597# a_661_n597# 0.01fF
C226 a_977_n597# a_1293_n597# 0.04fF
C227 a_1135_n597# a_1293_n597# 0.12fF
C228 a_819_n597# a_1293_n597# 0.02fF
C229 a_1293_n597# a_661_n597# 0.02fF
C230 a_1135_n597# a_977_n597# 0.12fF
C231 a_1451_n597# a_503_n597# 0.01fF
C232 a_819_n597# a_977_n597# 0.12fF
C233 a_819_n597# a_1135_n597# 0.04fF
C234 a_977_n597# a_661_n597# 0.04fF
C235 a_1135_n597# a_661_n597# 0.02fF
C236 a_819_n597# a_661_n597# 0.12fF
C237 a_1451_n597# a_29_n597# 0.01fF
C238 a_1293_n597# a_503_n597# 0.01fF
C239 a_1451_n597# a_187_n597# 0.01fF
C240 a_n129_n597# a_1451_n597# 0.01fF
C241 a_345_n597# a_1451_n597# 0.01fF
C242 a_977_n597# a_503_n597# 0.02fF
C243 a_1135_n597# a_503_n597# 0.02fF
C244 a_1293_n597# a_29_n597# 0.01fF
C245 a_1293_n597# a_187_n597# 0.01fF
C246 a_n129_n597# a_1293_n597# 0.01fF
C247 a_345_n597# a_1293_n597# 0.01fF
C248 a_819_n597# a_503_n597# 0.04fF
C249 a_503_n597# a_661_n597# 0.12fF
C250 a_977_n597# a_29_n597# 0.01fF
C251 a_n129_n597# a_977_n597# 0.01fF
C252 a_1135_n597# a_29_n597# 0.01fF
C253 a_1135_n597# a_187_n597# 0.01fF
C254 a_1293_n597# a_n287_n597# 0.01fF
C255 a_977_n597# a_187_n597# 0.01fF
C256 a_n129_n597# a_1135_n597# 0.01fF
C257 a_345_n597# a_977_n597# 0.02fF
C258 a_345_n597# a_1135_n597# 0.01fF
C259 a_819_n597# a_29_n597# 0.01fF
C260 a_819_n597# a_187_n597# 0.02fF
C261 a_n129_n597# a_819_n597# 0.01fF
C262 a_29_n597# a_661_n597# 0.02fF
C263 a_661_n597# a_187_n597# 0.02fF
C264 a_345_n597# a_819_n597# 0.02fF
C265 a_n129_n597# a_661_n597# 0.01fF
C266 a_1135_n597# a_n287_n597# 0.01fF
C267 a_977_n597# a_n287_n597# 0.01fF
C268 a_345_n597# a_661_n597# 0.04fF
C269 a_819_n597# a_n287_n597# 0.01fF
C270 a_977_n597# a_n603_n597# 0.01fF
C271 a_n287_n597# a_661_n597# 0.01fF
C272 a_1135_n597# a_n445_n597# 0.01fF
C273 a_977_n597# a_n445_n597# 0.01fF
C274 a_819_n597# a_n603_n597# 0.01fF
C275 a_819_n597# a_n445_n597# 0.01fF
C276 a_29_n597# a_503_n597# 0.02fF
C277 a_503_n597# a_187_n597# 0.04fF
C278 a_661_n597# a_n603_n597# 0.01fF
C279 a_n129_n597# a_503_n597# 0.02fF
C280 a_661_n597# a_n445_n597# 0.01fF
C281 a_345_n597# a_503_n597# 0.12fF
C282 a_819_n597# a_n761_n597# 0.01fF
C283 a_661_n597# a_n761_n597# 0.01fF
C284 a_n287_n597# a_503_n597# 0.01fF
C285 a_n919_n597# a_661_n597# 0.01fF
C286 a_29_n597# a_187_n597# 0.12fF
C287 a_n129_n597# a_187_n597# 0.04fF
C288 a_n129_n597# a_29_n597# 0.12fF
C289 a_345_n597# a_29_n597# 0.04fF
C290 a_345_n597# a_187_n597# 0.12fF
C291 a_n129_n597# a_345_n597# 0.02fF
C292 a_503_n597# a_n603_n597# 0.01fF
C293 a_503_n597# a_n445_n597# 0.01fF
C294 a_n287_n597# a_29_n597# 0.04fF
C295 a_n287_n597# a_187_n597# 0.02fF
C296 a_n129_n597# a_n287_n597# 0.12fF
C297 a_503_n597# a_n761_n597# 0.01fF
C298 a_345_n597# a_n287_n597# 0.02fF
C299 a_n919_n597# a_503_n597# 0.01fF
C300 a_29_n597# a_n603_n597# 0.02fF
C301 a_29_n597# a_n445_n597# 0.02fF
C302 a_187_n597# a_n603_n597# 0.01fF
C303 a_n445_n597# a_187_n597# 0.02fF
C304 a_n129_n597# a_n445_n597# 0.04fF
C305 a_n129_n597# a_n603_n597# 0.02fF
C306 a_345_n597# a_n603_n597# 0.01fF
C307 a_345_n597# a_n445_n597# 0.01fF
C308 a_29_n597# a_n761_n597# 0.01fF
C309 a_187_n597# a_n761_n597# 0.01fF
C310 a_n129_n597# a_n761_n597# 0.02fF
C311 a_n1077_n597# a_503_n597# 0.01fF
C312 a_345_n597# a_n761_n597# 0.01fF
C313 a_n287_n597# a_n445_n597# 0.12fF
C314 a_n287_n597# a_n603_n597# 0.04fF
C315 a_n919_n597# a_29_n597# 0.01fF
C316 a_n919_n597# a_187_n597# 0.01fF
C317 a_n129_n597# a_n919_n597# 0.01fF
C318 a_345_n597# a_n919_n597# 0.01fF
C319 a_n287_n597# a_n761_n597# 0.02fF
C320 a_n445_n597# a_n603_n597# 0.12fF
C321 a_1551_n500# w_n1809_n797# 0.30fF
C322 a_n1077_n597# a_29_n597# 0.01fF
C323 a_1393_n500# w_n1809_n797# 0.13fF
C324 w_n1809_n797# a_1235_n500# 0.09fF
C325 a_n287_n597# a_n919_n597# 0.02fF
C326 a_n1077_n597# a_187_n597# 0.01fF
C327 a_n129_n597# a_n1077_n597# 0.01fF
C328 w_n1809_n797# a_919_n500# 0.06fF
C329 a_1077_n500# w_n1809_n797# 0.07fF
C330 a_n761_n597# a_n603_n597# 0.12fF
C331 a_345_n597# a_n1077_n597# 0.01fF
C332 a_n445_n597# a_n761_n597# 0.04fF
C333 w_n1809_n797# a_445_n500# 0.04fF
C334 a_287_n500# w_n1809_n797# 0.04fF
C335 w_n1809_n797# a_603_n500# 0.05fF
C336 a_n919_n597# a_n603_n597# 0.04fF
C337 a_n919_n597# a_n445_n597# 0.02fF
C338 a_761_n500# w_n1809_n797# 0.05fF
C339 a_n1077_n597# a_n287_n597# 0.01fF
C340 a_n919_n597# a_n761_n597# 0.12fF
C341 w_n1809_n797# VSUBS 17.30fF
.ends

.subckt esd_cell esd VDD VSS
Xsky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0 VSS VSS VSS VSS VSS VSS esd VSS VSS VSS esd
+ VSS esd VSS VSS VSS VSS esd VSS esd esd VSS VSS VSS VSS VSS VSS esd VSS VSS VSS
+ VSS esd VSS VSS esd VSS VSS VSS VSS VSS esd sky130_fd_pr__nfet_g5v0d10v5_BRTJC6
Xsky130_fd_pr__pfet_g5v0d10v5_CADZ46_0 VDD VDD esd VDD VDD VDD VDD esd esd VDD VDD
+ VDD VDD VDD VDD VDD VDD esd VDD VDD VDD VDD esd VDD VDD VDD esd VDD VDD VDD VDD
+ VDD VDD VDD VDD esd VDD VDD esd esd VDD esd VSS sky130_fd_pr__pfet_g5v0d10v5_CADZ46
C0 VDD esd 4.35fF
C1 VDD VSS -182.19fF
C2 esd VSS 22.39fF
.ends

