magic
tech sky130A
magscale 1 2
timestamp 1653034865
<< nmos >>
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
<< ndiff >>
rect -652 128 -594 140
rect -652 -128 -640 128
rect -606 -128 -594 128
rect -652 -140 -594 -128
rect -474 128 -416 140
rect -474 -128 -462 128
rect -428 -128 -416 128
rect -474 -140 -416 -128
rect -296 128 -238 140
rect -296 -128 -284 128
rect -250 -128 -238 128
rect -296 -140 -238 -128
rect -118 128 -60 140
rect -118 -128 -106 128
rect -72 -128 -60 128
rect -118 -140 -60 -128
rect 60 128 118 140
rect 60 -128 72 128
rect 106 -128 118 128
rect 60 -140 118 -128
rect 238 128 296 140
rect 238 -128 250 128
rect 284 -128 296 128
rect 238 -140 296 -128
rect 416 128 474 140
rect 416 -128 428 128
rect 462 -128 474 128
rect 416 -140 474 -128
rect 594 128 652 140
rect 594 -128 606 128
rect 640 -128 652 128
rect 594 -140 652 -128
<< ndiffc >>
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
<< poly >>
rect -572 212 -496 228
rect -572 195 -556 212
rect -594 178 -556 195
rect -512 195 -496 212
rect -394 212 -318 228
rect -394 195 -378 212
rect -512 178 -474 195
rect -594 140 -474 178
rect -416 178 -378 195
rect -334 195 -318 212
rect -216 212 -140 228
rect -216 195 -200 212
rect -334 178 -296 195
rect -416 140 -296 178
rect -238 178 -200 195
rect -156 195 -140 212
rect -38 212 38 228
rect -38 195 -22 212
rect -156 178 -118 195
rect -238 140 -118 178
rect -60 178 -22 195
rect 22 195 38 212
rect 140 212 216 228
rect 140 195 156 212
rect 22 178 60 195
rect -60 140 60 178
rect 118 178 156 195
rect 200 195 216 212
rect 318 212 394 228
rect 318 195 334 212
rect 200 178 238 195
rect 118 140 238 178
rect 296 178 334 195
rect 378 195 394 212
rect 496 212 572 228
rect 496 195 512 212
rect 378 178 416 195
rect 296 140 416 178
rect 474 178 512 195
rect 556 195 572 212
rect 556 178 594 195
rect 474 140 594 178
rect -594 -178 -474 -140
rect -594 -195 -556 -178
rect -572 -212 -556 -195
rect -512 -195 -474 -178
rect -416 -178 -296 -140
rect -416 -195 -378 -178
rect -512 -212 -496 -195
rect -572 -228 -496 -212
rect -394 -212 -378 -195
rect -334 -195 -296 -178
rect -238 -178 -118 -140
rect -238 -195 -200 -178
rect -334 -212 -318 -195
rect -394 -228 -318 -212
rect -216 -212 -200 -195
rect -156 -195 -118 -178
rect -60 -178 60 -140
rect -60 -195 -22 -178
rect -156 -212 -140 -195
rect -216 -228 -140 -212
rect -38 -212 -22 -195
rect 22 -195 60 -178
rect 118 -178 238 -140
rect 118 -195 156 -178
rect 22 -212 38 -195
rect -38 -228 38 -212
rect 140 -212 156 -195
rect 200 -195 238 -178
rect 296 -178 416 -140
rect 296 -195 334 -178
rect 200 -212 216 -195
rect 140 -228 216 -212
rect 318 -212 334 -195
rect 378 -195 416 -178
rect 474 -178 594 -140
rect 474 -195 512 -178
rect 378 -212 394 -195
rect 318 -228 394 -212
rect 496 -212 512 -195
rect 556 -195 594 -178
rect 556 -212 572 -195
rect 496 -228 572 -212
<< polycont >>
rect -556 178 -512 212
rect -378 178 -334 212
rect -200 178 -156 212
rect -22 178 22 212
rect 156 178 200 212
rect 334 178 378 212
rect 512 178 556 212
rect -556 -212 -512 -178
rect -378 -212 -334 -178
rect -200 -212 -156 -178
rect -22 -212 22 -178
rect 156 -212 200 -178
rect 334 -212 378 -178
rect 512 -212 556 -178
<< locali >>
rect -572 178 -556 212
rect -512 178 -496 212
rect -394 178 -378 212
rect -334 178 -318 212
rect -216 178 -200 212
rect -156 178 -140 212
rect -38 178 -22 212
rect 22 178 38 212
rect 140 178 156 212
rect 200 178 216 212
rect 318 178 334 212
rect 378 178 394 212
rect 496 178 512 212
rect 556 178 572 212
rect -640 128 -606 144
rect -640 -144 -606 -128
rect -462 128 -428 144
rect -462 -144 -428 -128
rect -284 128 -250 144
rect -284 -144 -250 -128
rect -106 128 -72 144
rect -106 -144 -72 -128
rect 72 128 106 144
rect 72 -144 106 -128
rect 250 128 284 144
rect 250 -144 284 -128
rect 428 128 462 144
rect 428 -144 462 -128
rect 606 128 640 144
rect 606 -144 640 -128
rect -572 -212 -556 -178
rect -512 -212 -496 -178
rect -394 -212 -378 -178
rect -334 -212 -318 -178
rect -216 -212 -200 -178
rect -156 -212 -140 -178
rect -38 -212 -22 -178
rect 22 -212 38 -178
rect 140 -212 156 -178
rect 200 -212 216 -178
rect 318 -212 334 -178
rect 378 -212 394 -178
rect 496 -212 512 -178
rect 556 -212 572 -178
<< viali >>
rect -556 178 -512 212
rect -378 178 -334 212
rect -200 178 -156 212
rect -22 178 22 212
rect 156 178 200 212
rect 334 178 378 212
rect 512 178 556 212
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect -556 -212 -512 -178
rect -378 -212 -334 -178
rect -200 -212 -156 -178
rect -22 -212 22 -178
rect 156 -212 200 -178
rect 334 -212 378 -178
rect 512 -212 556 -178
<< metal1 >>
rect -572 212 -496 228
rect -572 178 -556 212
rect -512 178 -496 212
rect -572 172 -496 178
rect -394 212 -318 228
rect -394 178 -378 212
rect -334 178 -318 212
rect -394 172 -318 178
rect -216 212 -140 228
rect -216 178 -200 212
rect -156 178 -140 212
rect -216 172 -140 178
rect -38 212 38 228
rect -38 178 -22 212
rect 22 178 38 212
rect -38 172 38 178
rect 140 212 216 228
rect 140 178 156 212
rect 200 178 216 212
rect 140 172 216 178
rect 318 212 394 228
rect 318 178 334 212
rect 378 178 394 212
rect 318 172 394 178
rect 496 212 572 228
rect 496 178 512 212
rect 556 178 572 212
rect 496 172 572 178
rect -646 128 -600 140
rect -646 -128 -640 128
rect -606 -128 -600 128
rect -646 -140 -600 -128
rect -468 128 -422 140
rect -468 -128 -462 128
rect -428 -128 -422 128
rect -468 -140 -422 -128
rect -290 128 -244 140
rect -290 -128 -284 128
rect -250 -128 -244 128
rect -290 -140 -244 -128
rect -112 128 -66 140
rect -112 -128 -106 128
rect -72 -128 -66 128
rect -112 -140 -66 -128
rect 66 128 112 140
rect 66 -128 72 128
rect 106 -128 112 128
rect 66 -140 112 -128
rect 244 128 290 140
rect 244 -128 250 128
rect 284 -128 290 128
rect 244 -140 290 -128
rect 422 128 468 140
rect 422 -128 428 128
rect 462 -128 468 128
rect 422 -140 468 -128
rect 600 128 646 140
rect 600 -128 606 128
rect 640 -128 646 128
rect 600 -140 646 -128
rect -572 -178 -496 -172
rect -572 -212 -556 -178
rect -512 -212 -496 -178
rect -572 -228 -496 -212
rect -394 -178 -318 -172
rect -394 -212 -378 -178
rect -334 -212 -318 -178
rect -394 -228 -318 -212
rect -216 -178 -140 -172
rect -216 -212 -200 -178
rect -156 -212 -140 -178
rect -216 -228 -140 -212
rect -38 -178 38 -172
rect -38 -212 -22 -178
rect 22 -212 38 -178
rect -38 -228 38 -212
rect 140 -178 216 -172
rect 140 -212 156 -178
rect 200 -212 216 -178
rect 140 -228 216 -212
rect 318 -178 394 -172
rect 318 -212 334 -178
rect 378 -212 394 -178
rect 318 -228 394 -212
rect 496 -178 572 -172
rect 496 -212 512 -178
rect 556 -212 572 -178
rect 496 -228 572 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 7 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
