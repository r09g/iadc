magic
tech sky130A
timestamp 1655484843
<< metal1 >>
rect -13 13 13 16
rect -13 -16 13 -13
<< via1 >>
rect -13 -13 13 13
<< metal2 >>
rect -16 -13 -13 13
rect 13 -13 16 13
<< properties >>
string GDS_END 505162
string GDS_FILE digital_filter_3a.gds
string GDS_START 504966
<< end >>
