magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< nwell >>
rect -2112 -241 2112 241
<< pmos >>
rect -2018 -140 -1898 140
rect -1840 -140 -1720 140
rect -1662 -140 -1542 140
rect -1484 -140 -1364 140
rect -1306 -140 -1186 140
rect -1128 -140 -1008 140
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
rect 1008 -140 1128 140
rect 1186 -140 1306 140
rect 1364 -140 1484 140
rect 1542 -140 1662 140
rect 1720 -140 1840 140
rect 1898 -140 2018 140
<< pdiff >>
rect -2076 128 -2018 140
rect -2076 -128 -2064 128
rect -2030 -128 -2018 128
rect -2076 -140 -2018 -128
rect -1898 128 -1840 140
rect -1898 -128 -1886 128
rect -1852 -128 -1840 128
rect -1898 -140 -1840 -128
rect -1720 128 -1662 140
rect -1720 -128 -1708 128
rect -1674 -128 -1662 128
rect -1720 -140 -1662 -128
rect -1542 128 -1484 140
rect -1542 -128 -1530 128
rect -1496 -128 -1484 128
rect -1542 -140 -1484 -128
rect -1364 128 -1306 140
rect -1364 -128 -1352 128
rect -1318 -128 -1306 128
rect -1364 -140 -1306 -128
rect -1186 128 -1128 140
rect -1186 -128 -1174 128
rect -1140 -128 -1128 128
rect -1186 -140 -1128 -128
rect -1008 128 -950 140
rect -1008 -128 -996 128
rect -962 -128 -950 128
rect -1008 -140 -950 -128
rect -830 128 -772 140
rect -830 -128 -818 128
rect -784 -128 -772 128
rect -830 -140 -772 -128
rect -652 128 -594 140
rect -652 -128 -640 128
rect -606 -128 -594 128
rect -652 -140 -594 -128
rect -474 128 -416 140
rect -474 -128 -462 128
rect -428 -128 -416 128
rect -474 -140 -416 -128
rect -296 128 -238 140
rect -296 -128 -284 128
rect -250 -128 -238 128
rect -296 -140 -238 -128
rect -118 128 -60 140
rect -118 -128 -106 128
rect -72 -128 -60 128
rect -118 -140 -60 -128
rect 60 128 118 140
rect 60 -128 72 128
rect 106 -128 118 128
rect 60 -140 118 -128
rect 238 128 296 140
rect 238 -128 250 128
rect 284 -128 296 128
rect 238 -140 296 -128
rect 416 128 474 140
rect 416 -128 428 128
rect 462 -128 474 128
rect 416 -140 474 -128
rect 594 128 652 140
rect 594 -128 606 128
rect 640 -128 652 128
rect 594 -140 652 -128
rect 772 128 830 140
rect 772 -128 784 128
rect 818 -128 830 128
rect 772 -140 830 -128
rect 950 128 1008 140
rect 950 -128 962 128
rect 996 -128 1008 128
rect 950 -140 1008 -128
rect 1128 128 1186 140
rect 1128 -128 1140 128
rect 1174 -128 1186 128
rect 1128 -140 1186 -128
rect 1306 128 1364 140
rect 1306 -128 1318 128
rect 1352 -128 1364 128
rect 1306 -140 1364 -128
rect 1484 128 1542 140
rect 1484 -128 1496 128
rect 1530 -128 1542 128
rect 1484 -140 1542 -128
rect 1662 128 1720 140
rect 1662 -128 1674 128
rect 1708 -128 1720 128
rect 1662 -140 1720 -128
rect 1840 128 1898 140
rect 1840 -128 1852 128
rect 1886 -128 1898 128
rect 1840 -140 1898 -128
rect 2018 128 2076 140
rect 2018 -128 2030 128
rect 2064 -128 2076 128
rect 2018 -140 2076 -128
<< pdiffc >>
rect -2064 -128 -2030 128
rect -1886 -128 -1852 128
rect -1708 -128 -1674 128
rect -1530 -128 -1496 128
rect -1352 -128 -1318 128
rect -1174 -128 -1140 128
rect -996 -128 -962 128
rect -818 -128 -784 128
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect 784 -128 818 128
rect 962 -128 996 128
rect 1140 -128 1174 128
rect 1318 -128 1352 128
rect 1496 -128 1530 128
rect 1674 -128 1708 128
rect 1852 -128 1886 128
rect 2030 -128 2064 128
<< poly >>
rect -1996 221 -1920 237
rect -1996 205 -1980 221
rect -2018 187 -1980 205
rect -1936 205 -1920 221
rect -1818 221 -1742 237
rect -1818 205 -1802 221
rect -1936 187 -1898 205
rect -2018 140 -1898 187
rect -1840 187 -1802 205
rect -1758 205 -1742 221
rect -1640 221 -1564 237
rect -1640 205 -1624 221
rect -1758 187 -1720 205
rect -1840 140 -1720 187
rect -1662 187 -1624 205
rect -1580 205 -1564 221
rect -1462 221 -1386 237
rect -1462 205 -1446 221
rect -1580 187 -1542 205
rect -1662 140 -1542 187
rect -1484 187 -1446 205
rect -1402 205 -1386 221
rect -1284 221 -1208 237
rect -1284 205 -1268 221
rect -1402 187 -1364 205
rect -1484 140 -1364 187
rect -1306 187 -1268 205
rect -1224 205 -1208 221
rect -1106 221 -1030 237
rect -1106 205 -1090 221
rect -1224 187 -1186 205
rect -1306 140 -1186 187
rect -1128 187 -1090 205
rect -1046 205 -1030 221
rect -928 221 -852 237
rect -928 205 -912 221
rect -1046 187 -1008 205
rect -1128 140 -1008 187
rect -950 187 -912 205
rect -868 205 -852 221
rect -750 221 -674 237
rect -750 205 -734 221
rect -868 187 -830 205
rect -950 140 -830 187
rect -772 187 -734 205
rect -690 205 -674 221
rect -572 221 -496 237
rect -572 205 -556 221
rect -690 187 -652 205
rect -772 140 -652 187
rect -594 187 -556 205
rect -512 205 -496 221
rect -394 221 -318 237
rect -394 205 -378 221
rect -512 187 -474 205
rect -594 140 -474 187
rect -416 187 -378 205
rect -334 205 -318 221
rect -216 221 -140 237
rect -216 205 -200 221
rect -334 187 -296 205
rect -416 140 -296 187
rect -238 187 -200 205
rect -156 205 -140 221
rect -38 221 38 237
rect -38 205 -22 221
rect -156 187 -118 205
rect -238 140 -118 187
rect -60 187 -22 205
rect 22 205 38 221
rect 140 221 216 237
rect 140 205 156 221
rect 22 187 60 205
rect -60 140 60 187
rect 118 187 156 205
rect 200 205 216 221
rect 318 221 394 237
rect 318 205 334 221
rect 200 187 238 205
rect 118 140 238 187
rect 296 187 334 205
rect 378 205 394 221
rect 496 221 572 237
rect 496 205 512 221
rect 378 187 416 205
rect 296 140 416 187
rect 474 187 512 205
rect 556 205 572 221
rect 674 221 750 237
rect 674 205 690 221
rect 556 187 594 205
rect 474 140 594 187
rect 652 187 690 205
rect 734 205 750 221
rect 852 221 928 237
rect 852 205 868 221
rect 734 187 772 205
rect 652 140 772 187
rect 830 187 868 205
rect 912 205 928 221
rect 1030 221 1106 237
rect 1030 205 1046 221
rect 912 187 950 205
rect 830 140 950 187
rect 1008 187 1046 205
rect 1090 205 1106 221
rect 1208 221 1284 237
rect 1208 205 1224 221
rect 1090 187 1128 205
rect 1008 140 1128 187
rect 1186 187 1224 205
rect 1268 205 1284 221
rect 1386 221 1462 237
rect 1386 205 1402 221
rect 1268 187 1306 205
rect 1186 140 1306 187
rect 1364 187 1402 205
rect 1446 205 1462 221
rect 1564 221 1640 237
rect 1564 205 1580 221
rect 1446 187 1484 205
rect 1364 140 1484 187
rect 1542 187 1580 205
rect 1624 205 1640 221
rect 1742 221 1818 237
rect 1742 205 1758 221
rect 1624 187 1662 205
rect 1542 140 1662 187
rect 1720 187 1758 205
rect 1802 205 1818 221
rect 1920 221 1996 237
rect 1920 205 1936 221
rect 1802 187 1840 205
rect 1720 140 1840 187
rect 1898 187 1936 205
rect 1980 205 1996 221
rect 1980 187 2018 205
rect 1898 140 2018 187
rect -2018 -187 -1898 -140
rect -2018 -205 -1980 -187
rect -1996 -221 -1980 -205
rect -1936 -205 -1898 -187
rect -1840 -187 -1720 -140
rect -1840 -205 -1802 -187
rect -1936 -221 -1920 -205
rect -1996 -237 -1920 -221
rect -1818 -221 -1802 -205
rect -1758 -205 -1720 -187
rect -1662 -187 -1542 -140
rect -1662 -205 -1624 -187
rect -1758 -221 -1742 -205
rect -1818 -237 -1742 -221
rect -1640 -221 -1624 -205
rect -1580 -205 -1542 -187
rect -1484 -187 -1364 -140
rect -1484 -205 -1446 -187
rect -1580 -221 -1564 -205
rect -1640 -237 -1564 -221
rect -1462 -221 -1446 -205
rect -1402 -205 -1364 -187
rect -1306 -187 -1186 -140
rect -1306 -205 -1268 -187
rect -1402 -221 -1386 -205
rect -1462 -237 -1386 -221
rect -1284 -221 -1268 -205
rect -1224 -205 -1186 -187
rect -1128 -187 -1008 -140
rect -1128 -205 -1090 -187
rect -1224 -221 -1208 -205
rect -1284 -237 -1208 -221
rect -1106 -221 -1090 -205
rect -1046 -205 -1008 -187
rect -950 -187 -830 -140
rect -950 -205 -912 -187
rect -1046 -221 -1030 -205
rect -1106 -237 -1030 -221
rect -928 -221 -912 -205
rect -868 -205 -830 -187
rect -772 -187 -652 -140
rect -772 -205 -734 -187
rect -868 -221 -852 -205
rect -928 -237 -852 -221
rect -750 -221 -734 -205
rect -690 -205 -652 -187
rect -594 -187 -474 -140
rect -594 -205 -556 -187
rect -690 -221 -674 -205
rect -750 -237 -674 -221
rect -572 -221 -556 -205
rect -512 -205 -474 -187
rect -416 -187 -296 -140
rect -416 -205 -378 -187
rect -512 -221 -496 -205
rect -572 -237 -496 -221
rect -394 -221 -378 -205
rect -334 -205 -296 -187
rect -238 -187 -118 -140
rect -238 -205 -200 -187
rect -334 -221 -318 -205
rect -394 -237 -318 -221
rect -216 -221 -200 -205
rect -156 -205 -118 -187
rect -60 -187 60 -140
rect -60 -205 -22 -187
rect -156 -221 -140 -205
rect -216 -237 -140 -221
rect -38 -221 -22 -205
rect 22 -205 60 -187
rect 118 -187 238 -140
rect 118 -205 156 -187
rect 22 -221 38 -205
rect -38 -237 38 -221
rect 140 -221 156 -205
rect 200 -205 238 -187
rect 296 -187 416 -140
rect 296 -205 334 -187
rect 200 -221 216 -205
rect 140 -237 216 -221
rect 318 -221 334 -205
rect 378 -205 416 -187
rect 474 -187 594 -140
rect 474 -205 512 -187
rect 378 -221 394 -205
rect 318 -237 394 -221
rect 496 -221 512 -205
rect 556 -205 594 -187
rect 652 -187 772 -140
rect 652 -205 690 -187
rect 556 -221 572 -205
rect 496 -237 572 -221
rect 674 -221 690 -205
rect 734 -205 772 -187
rect 830 -187 950 -140
rect 830 -205 868 -187
rect 734 -221 750 -205
rect 674 -237 750 -221
rect 852 -221 868 -205
rect 912 -205 950 -187
rect 1008 -187 1128 -140
rect 1008 -205 1046 -187
rect 912 -221 928 -205
rect 852 -237 928 -221
rect 1030 -221 1046 -205
rect 1090 -205 1128 -187
rect 1186 -187 1306 -140
rect 1186 -205 1224 -187
rect 1090 -221 1106 -205
rect 1030 -237 1106 -221
rect 1208 -221 1224 -205
rect 1268 -205 1306 -187
rect 1364 -187 1484 -140
rect 1364 -205 1402 -187
rect 1268 -221 1284 -205
rect 1208 -237 1284 -221
rect 1386 -221 1402 -205
rect 1446 -205 1484 -187
rect 1542 -187 1662 -140
rect 1542 -205 1580 -187
rect 1446 -221 1462 -205
rect 1386 -237 1462 -221
rect 1564 -221 1580 -205
rect 1624 -205 1662 -187
rect 1720 -187 1840 -140
rect 1720 -205 1758 -187
rect 1624 -221 1640 -205
rect 1564 -237 1640 -221
rect 1742 -221 1758 -205
rect 1802 -205 1840 -187
rect 1898 -187 2018 -140
rect 1898 -205 1936 -187
rect 1802 -221 1818 -205
rect 1742 -237 1818 -221
rect 1920 -221 1936 -205
rect 1980 -205 2018 -187
rect 1980 -221 1996 -205
rect 1920 -237 1996 -221
<< polycont >>
rect -1980 187 -1936 221
rect -1802 187 -1758 221
rect -1624 187 -1580 221
rect -1446 187 -1402 221
rect -1268 187 -1224 221
rect -1090 187 -1046 221
rect -912 187 -868 221
rect -734 187 -690 221
rect -556 187 -512 221
rect -378 187 -334 221
rect -200 187 -156 221
rect -22 187 22 221
rect 156 187 200 221
rect 334 187 378 221
rect 512 187 556 221
rect 690 187 734 221
rect 868 187 912 221
rect 1046 187 1090 221
rect 1224 187 1268 221
rect 1402 187 1446 221
rect 1580 187 1624 221
rect 1758 187 1802 221
rect 1936 187 1980 221
rect -1980 -221 -1936 -187
rect -1802 -221 -1758 -187
rect -1624 -221 -1580 -187
rect -1446 -221 -1402 -187
rect -1268 -221 -1224 -187
rect -1090 -221 -1046 -187
rect -912 -221 -868 -187
rect -734 -221 -690 -187
rect -556 -221 -512 -187
rect -378 -221 -334 -187
rect -200 -221 -156 -187
rect -22 -221 22 -187
rect 156 -221 200 -187
rect 334 -221 378 -187
rect 512 -221 556 -187
rect 690 -221 734 -187
rect 868 -221 912 -187
rect 1046 -221 1090 -187
rect 1224 -221 1268 -187
rect 1402 -221 1446 -187
rect 1580 -221 1624 -187
rect 1758 -221 1802 -187
rect 1936 -221 1980 -187
<< locali >>
rect -1996 187 -1980 221
rect -1936 187 -1920 221
rect -1818 187 -1802 221
rect -1758 187 -1742 221
rect -1640 187 -1624 221
rect -1580 187 -1564 221
rect -1462 187 -1446 221
rect -1402 187 -1386 221
rect -1284 187 -1268 221
rect -1224 187 -1208 221
rect -1106 187 -1090 221
rect -1046 187 -1030 221
rect -928 187 -912 221
rect -868 187 -852 221
rect -750 187 -734 221
rect -690 187 -674 221
rect -572 187 -556 221
rect -512 187 -496 221
rect -394 187 -378 221
rect -334 187 -318 221
rect -216 187 -200 221
rect -156 187 -140 221
rect -38 187 -22 221
rect 22 187 38 221
rect 140 187 156 221
rect 200 187 216 221
rect 318 187 334 221
rect 378 187 394 221
rect 496 187 512 221
rect 556 187 572 221
rect 674 187 690 221
rect 734 187 750 221
rect 852 187 868 221
rect 912 187 928 221
rect 1030 187 1046 221
rect 1090 187 1106 221
rect 1208 187 1224 221
rect 1268 187 1284 221
rect 1386 187 1402 221
rect 1446 187 1462 221
rect 1564 187 1580 221
rect 1624 187 1640 221
rect 1742 187 1758 221
rect 1802 187 1818 221
rect 1920 187 1936 221
rect 1980 187 1996 221
rect -2064 128 -2030 144
rect -2064 -144 -2030 -128
rect -1886 128 -1852 144
rect -1886 -144 -1852 -128
rect -1708 128 -1674 144
rect -1708 -144 -1674 -128
rect -1530 128 -1496 144
rect -1530 -144 -1496 -128
rect -1352 128 -1318 144
rect -1352 -144 -1318 -128
rect -1174 128 -1140 144
rect -1174 -144 -1140 -128
rect -996 128 -962 144
rect -996 -144 -962 -128
rect -818 128 -784 144
rect -818 -144 -784 -128
rect -640 128 -606 144
rect -640 -144 -606 -128
rect -462 128 -428 144
rect -462 -144 -428 -128
rect -284 128 -250 144
rect -284 -144 -250 -128
rect -106 128 -72 144
rect -106 -144 -72 -128
rect 72 128 106 144
rect 72 -144 106 -128
rect 250 128 284 144
rect 250 -144 284 -128
rect 428 128 462 144
rect 428 -144 462 -128
rect 606 128 640 144
rect 606 -144 640 -128
rect 784 128 818 144
rect 784 -144 818 -128
rect 962 128 996 144
rect 962 -144 996 -128
rect 1140 128 1174 144
rect 1140 -144 1174 -128
rect 1318 128 1352 144
rect 1318 -144 1352 -128
rect 1496 128 1530 144
rect 1496 -144 1530 -128
rect 1674 128 1708 144
rect 1674 -144 1708 -128
rect 1852 128 1886 144
rect 1852 -144 1886 -128
rect 2030 128 2064 144
rect 2030 -144 2064 -128
rect -1996 -221 -1980 -187
rect -1936 -221 -1920 -187
rect -1818 -221 -1802 -187
rect -1758 -221 -1742 -187
rect -1640 -221 -1624 -187
rect -1580 -221 -1564 -187
rect -1462 -221 -1446 -187
rect -1402 -221 -1386 -187
rect -1284 -221 -1268 -187
rect -1224 -221 -1208 -187
rect -1106 -221 -1090 -187
rect -1046 -221 -1030 -187
rect -928 -221 -912 -187
rect -868 -221 -852 -187
rect -750 -221 -734 -187
rect -690 -221 -674 -187
rect -572 -221 -556 -187
rect -512 -221 -496 -187
rect -394 -221 -378 -187
rect -334 -221 -318 -187
rect -216 -221 -200 -187
rect -156 -221 -140 -187
rect -38 -221 -22 -187
rect 22 -221 38 -187
rect 140 -221 156 -187
rect 200 -221 216 -187
rect 318 -221 334 -187
rect 378 -221 394 -187
rect 496 -221 512 -187
rect 556 -221 572 -187
rect 674 -221 690 -187
rect 734 -221 750 -187
rect 852 -221 868 -187
rect 912 -221 928 -187
rect 1030 -221 1046 -187
rect 1090 -221 1106 -187
rect 1208 -221 1224 -187
rect 1268 -221 1284 -187
rect 1386 -221 1402 -187
rect 1446 -221 1462 -187
rect 1564 -221 1580 -187
rect 1624 -221 1640 -187
rect 1742 -221 1758 -187
rect 1802 -221 1818 -187
rect 1920 -221 1936 -187
rect 1980 -221 1996 -187
<< viali >>
rect -1980 187 -1936 221
rect -1802 187 -1758 221
rect -1624 187 -1580 221
rect -1446 187 -1402 221
rect -1268 187 -1224 221
rect -1090 187 -1046 221
rect -912 187 -868 221
rect -734 187 -690 221
rect -556 187 -512 221
rect -378 187 -334 221
rect -200 187 -156 221
rect -22 187 22 221
rect 156 187 200 221
rect 334 187 378 221
rect 512 187 556 221
rect 690 187 734 221
rect 868 187 912 221
rect 1046 187 1090 221
rect 1224 187 1268 221
rect 1402 187 1446 221
rect 1580 187 1624 221
rect 1758 187 1802 221
rect 1936 187 1980 221
rect -2064 -128 -2030 128
rect -1886 -128 -1852 128
rect -1708 -128 -1674 128
rect -1530 -128 -1496 128
rect -1352 -128 -1318 128
rect -1174 -128 -1140 128
rect -996 -128 -962 128
rect -818 -128 -784 128
rect -640 -128 -606 128
rect -462 -128 -428 128
rect -284 -128 -250 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 250 -128 284 128
rect 428 -128 462 128
rect 606 -128 640 128
rect 784 -128 818 128
rect 962 -128 996 128
rect 1140 -128 1174 128
rect 1318 -128 1352 128
rect 1496 -128 1530 128
rect 1674 -128 1708 128
rect 1852 -128 1886 128
rect 2030 -128 2064 128
rect -1980 -221 -1936 -187
rect -1802 -221 -1758 -187
rect -1624 -221 -1580 -187
rect -1446 -221 -1402 -187
rect -1268 -221 -1224 -187
rect -1090 -221 -1046 -187
rect -912 -221 -868 -187
rect -734 -221 -690 -187
rect -556 -221 -512 -187
rect -378 -221 -334 -187
rect -200 -221 -156 -187
rect -22 -221 22 -187
rect 156 -221 200 -187
rect 334 -221 378 -187
rect 512 -221 556 -187
rect 690 -221 734 -187
rect 868 -221 912 -187
rect 1046 -221 1090 -187
rect 1224 -221 1268 -187
rect 1402 -221 1446 -187
rect 1580 -221 1624 -187
rect 1758 -221 1802 -187
rect 1936 -221 1980 -187
<< metal1 >>
rect -1996 221 -1920 237
rect -1996 187 -1980 221
rect -1936 187 -1920 221
rect -1996 181 -1920 187
rect -1818 221 -1742 237
rect -1818 187 -1802 221
rect -1758 187 -1742 221
rect -1818 181 -1742 187
rect -1640 221 -1564 237
rect -1640 187 -1624 221
rect -1580 187 -1564 221
rect -1640 181 -1564 187
rect -1462 221 -1386 237
rect -1462 187 -1446 221
rect -1402 187 -1386 221
rect -1462 181 -1386 187
rect -1284 221 -1208 237
rect -1284 187 -1268 221
rect -1224 187 -1208 221
rect -1284 181 -1208 187
rect -1106 221 -1030 237
rect -1106 187 -1090 221
rect -1046 187 -1030 221
rect -1106 181 -1030 187
rect -928 221 -852 237
rect -928 187 -912 221
rect -868 187 -852 221
rect -928 181 -852 187
rect -750 221 -674 237
rect -750 187 -734 221
rect -690 187 -674 221
rect -750 181 -674 187
rect -572 221 -496 237
rect -572 187 -556 221
rect -512 187 -496 221
rect -572 181 -496 187
rect -394 221 -318 237
rect -394 187 -378 221
rect -334 187 -318 221
rect -394 181 -318 187
rect -216 221 -140 237
rect -216 187 -200 221
rect -156 187 -140 221
rect -216 181 -140 187
rect -38 221 38 237
rect -38 187 -22 221
rect 22 187 38 221
rect -38 181 38 187
rect 140 221 216 237
rect 140 187 156 221
rect 200 187 216 221
rect 140 181 216 187
rect 318 221 394 237
rect 318 187 334 221
rect 378 187 394 221
rect 318 181 394 187
rect 496 221 572 237
rect 496 187 512 221
rect 556 187 572 221
rect 496 181 572 187
rect 674 221 750 237
rect 674 187 690 221
rect 734 187 750 221
rect 674 181 750 187
rect 852 221 928 237
rect 852 187 868 221
rect 912 187 928 221
rect 852 181 928 187
rect 1030 221 1106 237
rect 1030 187 1046 221
rect 1090 187 1106 221
rect 1030 181 1106 187
rect 1208 221 1284 237
rect 1208 187 1224 221
rect 1268 187 1284 221
rect 1208 181 1284 187
rect 1386 221 1462 237
rect 1386 187 1402 221
rect 1446 187 1462 221
rect 1386 181 1462 187
rect 1564 221 1640 237
rect 1564 187 1580 221
rect 1624 187 1640 221
rect 1564 181 1640 187
rect 1742 221 1818 237
rect 1742 187 1758 221
rect 1802 187 1818 221
rect 1742 181 1818 187
rect 1920 221 1996 237
rect 1920 187 1936 221
rect 1980 187 1996 221
rect 1920 181 1996 187
rect -2070 128 -2024 140
rect -2070 -128 -2064 128
rect -2030 -128 -2024 128
rect -2070 -140 -2024 -128
rect -1892 128 -1846 140
rect -1892 -128 -1886 128
rect -1852 -128 -1846 128
rect -1892 -140 -1846 -128
rect -1714 128 -1668 140
rect -1714 -128 -1708 128
rect -1674 -128 -1668 128
rect -1714 -140 -1668 -128
rect -1536 128 -1490 140
rect -1536 -128 -1530 128
rect -1496 -128 -1490 128
rect -1536 -140 -1490 -128
rect -1358 128 -1312 140
rect -1358 -128 -1352 128
rect -1318 -128 -1312 128
rect -1358 -140 -1312 -128
rect -1180 128 -1134 140
rect -1180 -128 -1174 128
rect -1140 -128 -1134 128
rect -1180 -140 -1134 -128
rect -1002 128 -956 140
rect -1002 -128 -996 128
rect -962 -128 -956 128
rect -1002 -140 -956 -128
rect -824 128 -778 140
rect -824 -128 -818 128
rect -784 -128 -778 128
rect -824 -140 -778 -128
rect -646 128 -600 140
rect -646 -128 -640 128
rect -606 -128 -600 128
rect -646 -140 -600 -128
rect -468 128 -422 140
rect -468 -128 -462 128
rect -428 -128 -422 128
rect -468 -140 -422 -128
rect -290 128 -244 140
rect -290 -128 -284 128
rect -250 -128 -244 128
rect -290 -140 -244 -128
rect -112 128 -66 140
rect -112 -128 -106 128
rect -72 -128 -66 128
rect -112 -140 -66 -128
rect 66 128 112 140
rect 66 -128 72 128
rect 106 -128 112 128
rect 66 -140 112 -128
rect 244 128 290 140
rect 244 -128 250 128
rect 284 -128 290 128
rect 244 -140 290 -128
rect 422 128 468 140
rect 422 -128 428 128
rect 462 -128 468 128
rect 422 -140 468 -128
rect 600 128 646 140
rect 600 -128 606 128
rect 640 -128 646 128
rect 600 -140 646 -128
rect 778 128 824 140
rect 778 -128 784 128
rect 818 -128 824 128
rect 778 -140 824 -128
rect 956 128 1002 140
rect 956 -128 962 128
rect 996 -128 1002 128
rect 956 -140 1002 -128
rect 1134 128 1180 140
rect 1134 -128 1140 128
rect 1174 -128 1180 128
rect 1134 -140 1180 -128
rect 1312 128 1358 140
rect 1312 -128 1318 128
rect 1352 -128 1358 128
rect 1312 -140 1358 -128
rect 1490 128 1536 140
rect 1490 -128 1496 128
rect 1530 -128 1536 128
rect 1490 -140 1536 -128
rect 1668 128 1714 140
rect 1668 -128 1674 128
rect 1708 -128 1714 128
rect 1668 -140 1714 -128
rect 1846 128 1892 140
rect 1846 -128 1852 128
rect 1886 -128 1892 128
rect 1846 -140 1892 -128
rect 2024 128 2070 140
rect 2024 -128 2030 128
rect 2064 -128 2070 128
rect 2024 -140 2070 -128
rect -1996 -187 -1920 -181
rect -1996 -221 -1980 -187
rect -1936 -221 -1920 -187
rect -1996 -237 -1920 -221
rect -1818 -187 -1742 -181
rect -1818 -221 -1802 -187
rect -1758 -221 -1742 -187
rect -1818 -237 -1742 -221
rect -1640 -187 -1564 -181
rect -1640 -221 -1624 -187
rect -1580 -221 -1564 -187
rect -1640 -237 -1564 -221
rect -1462 -187 -1386 -181
rect -1462 -221 -1446 -187
rect -1402 -221 -1386 -187
rect -1462 -237 -1386 -221
rect -1284 -187 -1208 -181
rect -1284 -221 -1268 -187
rect -1224 -221 -1208 -187
rect -1284 -237 -1208 -221
rect -1106 -187 -1030 -181
rect -1106 -221 -1090 -187
rect -1046 -221 -1030 -187
rect -1106 -237 -1030 -221
rect -928 -187 -852 -181
rect -928 -221 -912 -187
rect -868 -221 -852 -187
rect -928 -237 -852 -221
rect -750 -187 -674 -181
rect -750 -221 -734 -187
rect -690 -221 -674 -187
rect -750 -237 -674 -221
rect -572 -187 -496 -181
rect -572 -221 -556 -187
rect -512 -221 -496 -187
rect -572 -237 -496 -221
rect -394 -187 -318 -181
rect -394 -221 -378 -187
rect -334 -221 -318 -187
rect -394 -237 -318 -221
rect -216 -187 -140 -181
rect -216 -221 -200 -187
rect -156 -221 -140 -187
rect -216 -237 -140 -221
rect -38 -187 38 -181
rect -38 -221 -22 -187
rect 22 -221 38 -187
rect -38 -237 38 -221
rect 140 -187 216 -181
rect 140 -221 156 -187
rect 200 -221 216 -187
rect 140 -237 216 -221
rect 318 -187 394 -181
rect 318 -221 334 -187
rect 378 -221 394 -187
rect 318 -237 394 -221
rect 496 -187 572 -181
rect 496 -221 512 -187
rect 556 -221 572 -187
rect 496 -237 572 -221
rect 674 -187 750 -181
rect 674 -221 690 -187
rect 734 -221 750 -187
rect 674 -237 750 -221
rect 852 -187 928 -181
rect 852 -221 868 -187
rect 912 -221 928 -187
rect 852 -237 928 -221
rect 1030 -187 1106 -181
rect 1030 -221 1046 -187
rect 1090 -221 1106 -187
rect 1030 -237 1106 -221
rect 1208 -187 1284 -181
rect 1208 -221 1224 -187
rect 1268 -221 1284 -187
rect 1208 -237 1284 -221
rect 1386 -187 1462 -181
rect 1386 -221 1402 -187
rect 1446 -221 1462 -187
rect 1386 -237 1462 -221
rect 1564 -187 1640 -181
rect 1564 -221 1580 -187
rect 1624 -221 1640 -187
rect 1564 -237 1640 -221
rect 1742 -187 1818 -181
rect 1742 -221 1758 -187
rect 1802 -221 1818 -187
rect 1742 -237 1818 -221
rect 1920 -187 1996 -181
rect 1920 -221 1936 -187
rect 1980 -221 1996 -187
rect 1920 -237 1996 -221
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 23 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
