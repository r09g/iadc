magic
tech sky130A
timestamp 1654711401
<< error_p >>
rect -734 86 -705 89
rect -638 86 -609 89
rect -542 86 -513 89
rect -446 86 -417 89
rect -350 86 -321 89
rect -254 86 -225 89
rect -158 86 -129 89
rect -62 86 -33 89
rect 33 86 62 89
rect 129 86 158 89
rect 225 86 254 89
rect 321 86 350 89
rect 417 86 446 89
rect 513 86 542 89
rect 609 86 638 89
rect 705 86 734 89
rect -734 69 -728 86
rect -638 69 -632 86
rect -542 69 -536 86
rect -446 69 -440 86
rect -350 69 -344 86
rect -254 69 -248 86
rect -158 69 -152 86
rect -62 69 -56 86
rect 33 69 39 86
rect 129 69 135 86
rect 225 69 231 86
rect 321 69 327 86
rect 417 69 423 86
rect 513 69 519 86
rect 609 69 615 86
rect 705 69 711 86
rect -734 66 -705 69
rect -638 66 -609 69
rect -542 66 -513 69
rect -446 66 -417 69
rect -350 66 -321 69
rect -254 66 -225 69
rect -158 66 -129 69
rect -62 66 -33 69
rect 33 66 62 69
rect 129 66 158 69
rect 225 66 254 69
rect 321 66 350 69
rect 417 66 446 69
rect 513 66 542 69
rect 609 66 638 69
rect 705 66 734 69
<< pwell >>
rect -899 -155 899 155
<< nmos >>
rect -799 -50 -784 50
rect -751 -50 -736 50
rect -703 -50 -688 50
rect -655 -50 -640 50
rect -607 -50 -592 50
rect -559 -50 -544 50
rect -511 -50 -496 50
rect -463 -50 -448 50
rect -415 -50 -400 50
rect -367 -50 -352 50
rect -319 -50 -304 50
rect -271 -50 -256 50
rect -223 -50 -208 50
rect -175 -50 -160 50
rect -127 -50 -112 50
rect -79 -50 -64 50
rect -31 -50 -16 50
rect 16 -50 31 50
rect 64 -50 79 50
rect 112 -50 127 50
rect 160 -50 175 50
rect 208 -50 223 50
rect 256 -50 271 50
rect 304 -50 319 50
rect 352 -50 367 50
rect 400 -50 415 50
rect 448 -50 463 50
rect 496 -50 511 50
rect 544 -50 559 50
rect 592 -50 607 50
rect 640 -50 655 50
rect 688 -50 703 50
rect 736 -50 751 50
rect 784 -50 799 50
<< ndiff >>
rect -830 44 -799 50
rect -830 -44 -824 44
rect -807 -44 -799 44
rect -830 -50 -799 -44
rect -784 44 -751 50
rect -784 -44 -776 44
rect -759 -44 -751 44
rect -784 -50 -751 -44
rect -736 44 -703 50
rect -736 -44 -728 44
rect -711 -44 -703 44
rect -736 -50 -703 -44
rect -688 44 -655 50
rect -688 -44 -680 44
rect -663 -44 -655 44
rect -688 -50 -655 -44
rect -640 44 -607 50
rect -640 -44 -632 44
rect -615 -44 -607 44
rect -640 -50 -607 -44
rect -592 44 -559 50
rect -592 -44 -584 44
rect -567 -44 -559 44
rect -592 -50 -559 -44
rect -544 44 -511 50
rect -544 -44 -536 44
rect -519 -44 -511 44
rect -544 -50 -511 -44
rect -496 44 -463 50
rect -496 -44 -488 44
rect -471 -44 -463 44
rect -496 -50 -463 -44
rect -448 44 -415 50
rect -448 -44 -440 44
rect -423 -44 -415 44
rect -448 -50 -415 -44
rect -400 44 -367 50
rect -400 -44 -392 44
rect -375 -44 -367 44
rect -400 -50 -367 -44
rect -352 44 -319 50
rect -352 -44 -344 44
rect -327 -44 -319 44
rect -352 -50 -319 -44
rect -304 44 -271 50
rect -304 -44 -296 44
rect -279 -44 -271 44
rect -304 -50 -271 -44
rect -256 44 -223 50
rect -256 -44 -248 44
rect -231 -44 -223 44
rect -256 -50 -223 -44
rect -208 44 -175 50
rect -208 -44 -200 44
rect -183 -44 -175 44
rect -208 -50 -175 -44
rect -160 44 -127 50
rect -160 -44 -152 44
rect -135 -44 -127 44
rect -160 -50 -127 -44
rect -112 44 -79 50
rect -112 -44 -104 44
rect -87 -44 -79 44
rect -112 -50 -79 -44
rect -64 44 -31 50
rect -64 -44 -56 44
rect -39 -44 -31 44
rect -64 -50 -31 -44
rect -16 44 16 50
rect -16 -44 -8 44
rect 8 -44 16 44
rect -16 -50 16 -44
rect 31 44 64 50
rect 31 -44 39 44
rect 56 -44 64 44
rect 31 -50 64 -44
rect 79 44 112 50
rect 79 -44 87 44
rect 104 -44 112 44
rect 79 -50 112 -44
rect 127 44 160 50
rect 127 -44 135 44
rect 152 -44 160 44
rect 127 -50 160 -44
rect 175 44 208 50
rect 175 -44 183 44
rect 200 -44 208 44
rect 175 -50 208 -44
rect 223 44 256 50
rect 223 -44 231 44
rect 248 -44 256 44
rect 223 -50 256 -44
rect 271 44 304 50
rect 271 -44 279 44
rect 296 -44 304 44
rect 271 -50 304 -44
rect 319 44 352 50
rect 319 -44 327 44
rect 344 -44 352 44
rect 319 -50 352 -44
rect 367 44 400 50
rect 367 -44 375 44
rect 392 -44 400 44
rect 367 -50 400 -44
rect 415 44 448 50
rect 415 -44 423 44
rect 440 -44 448 44
rect 415 -50 448 -44
rect 463 44 496 50
rect 463 -44 471 44
rect 488 -44 496 44
rect 463 -50 496 -44
rect 511 44 544 50
rect 511 -44 519 44
rect 536 -44 544 44
rect 511 -50 544 -44
rect 559 44 592 50
rect 559 -44 567 44
rect 584 -44 592 44
rect 559 -50 592 -44
rect 607 44 640 50
rect 607 -44 615 44
rect 632 -44 640 44
rect 607 -50 640 -44
rect 655 44 688 50
rect 655 -44 663 44
rect 680 -44 688 44
rect 655 -50 688 -44
rect 703 44 736 50
rect 703 -44 711 44
rect 728 -44 736 44
rect 703 -50 736 -44
rect 751 44 784 50
rect 751 -44 759 44
rect 776 -44 784 44
rect 751 -50 784 -44
rect 799 44 830 50
rect 799 -44 807 44
rect 824 -44 830 44
rect 799 -50 830 -44
<< ndiffc >>
rect -824 -44 -807 44
rect -776 -44 -759 44
rect -728 -44 -711 44
rect -680 -44 -663 44
rect -632 -44 -615 44
rect -584 -44 -567 44
rect -536 -44 -519 44
rect -488 -44 -471 44
rect -440 -44 -423 44
rect -392 -44 -375 44
rect -344 -44 -327 44
rect -296 -44 -279 44
rect -248 -44 -231 44
rect -200 -44 -183 44
rect -152 -44 -135 44
rect -104 -44 -87 44
rect -56 -44 -39 44
rect -8 -44 8 44
rect 39 -44 56 44
rect 87 -44 104 44
rect 135 -44 152 44
rect 183 -44 200 44
rect 231 -44 248 44
rect 279 -44 296 44
rect 327 -44 344 44
rect 375 -44 392 44
rect 423 -44 440 44
rect 471 -44 488 44
rect 519 -44 536 44
rect 567 -44 584 44
rect 615 -44 632 44
rect 663 -44 680 44
rect 711 -44 728 44
rect 759 -44 776 44
rect 807 -44 824 44
<< psubdiff >>
rect -881 120 -833 137
rect 833 120 881 137
rect -881 89 -864 120
rect 864 89 881 120
rect -881 -120 -864 -89
rect 864 -120 881 -89
rect -881 -137 -833 -120
rect 833 -137 881 -120
<< psubdiffcont >>
rect -833 120 833 137
rect -881 -89 -864 89
rect 864 -89 881 89
rect -833 -137 833 -120
<< poly >>
rect -760 86 760 94
rect -760 69 -728 86
rect -711 69 -632 86
rect -615 69 -536 86
rect -519 69 -440 86
rect -423 69 -344 86
rect -327 69 -248 86
rect -231 69 -152 86
rect -135 69 -56 86
rect -39 69 39 86
rect 56 69 135 86
rect 152 69 231 86
rect 248 69 327 86
rect 344 69 423 86
rect 440 69 519 86
rect 536 69 615 86
rect 632 69 711 86
rect 728 69 760 86
rect -799 50 -784 63
rect -760 61 760 69
rect -751 50 -736 61
rect -703 50 -688 61
rect -655 50 -640 61
rect -607 50 -592 61
rect -559 50 -544 61
rect -511 50 -496 61
rect -463 50 -448 61
rect -415 50 -400 61
rect -367 50 -352 61
rect -319 50 -304 61
rect -271 50 -256 61
rect -223 50 -208 61
rect -175 50 -160 61
rect -127 50 -112 61
rect -79 50 -64 61
rect -31 50 -16 61
rect 16 50 31 61
rect 64 50 79 61
rect 112 50 127 61
rect 160 50 175 61
rect 208 50 223 61
rect 256 50 271 61
rect 304 50 319 61
rect 352 50 367 61
rect 400 50 415 61
rect 448 50 463 61
rect 496 50 511 61
rect 544 50 559 61
rect 592 50 607 61
rect 640 50 655 61
rect 688 50 703 61
rect 736 50 751 61
rect 784 50 799 63
rect -799 -61 -784 -50
rect -808 -69 -775 -61
rect -751 -63 -736 -50
rect -703 -63 -688 -50
rect -655 -63 -640 -50
rect -607 -63 -592 -50
rect -559 -63 -544 -50
rect -511 -63 -496 -50
rect -463 -63 -448 -50
rect -415 -63 -400 -50
rect -367 -63 -352 -50
rect -319 -63 -304 -50
rect -271 -63 -256 -50
rect -223 -63 -208 -50
rect -175 -63 -160 -50
rect -127 -63 -112 -50
rect -79 -63 -64 -50
rect -31 -63 -16 -50
rect 16 -63 31 -50
rect 64 -63 79 -50
rect 112 -63 127 -50
rect 160 -63 175 -50
rect 208 -63 223 -50
rect 256 -63 271 -50
rect 304 -63 319 -50
rect 352 -63 367 -50
rect 400 -63 415 -50
rect 448 -63 463 -50
rect 496 -63 511 -50
rect 544 -63 559 -50
rect 592 -63 607 -50
rect 640 -63 655 -50
rect 688 -63 703 -50
rect 736 -63 751 -50
rect 784 -63 799 -50
rect -808 -86 -800 -69
rect -783 -86 -775 -69
rect -808 -94 -775 -86
rect 775 -71 808 -63
rect 775 -88 783 -71
rect 800 -88 808 -71
rect 775 -96 808 -88
<< polycont >>
rect -728 69 -711 86
rect -632 69 -615 86
rect -536 69 -519 86
rect -440 69 -423 86
rect -344 69 -327 86
rect -248 69 -231 86
rect -152 69 -135 86
rect -56 69 -39 86
rect 39 69 56 86
rect 135 69 152 86
rect 231 69 248 86
rect 327 69 344 86
rect 423 69 440 86
rect 519 69 536 86
rect 615 69 632 86
rect 711 69 728 86
rect -800 -86 -783 -69
rect 783 -88 800 -71
<< locali >>
rect -881 120 -833 137
rect 833 120 881 137
rect -881 89 -864 120
rect 864 89 881 120
rect -736 69 -728 86
rect -711 69 -703 86
rect -640 69 -632 86
rect -615 69 -607 86
rect -544 69 -536 86
rect -519 69 -511 86
rect -448 69 -440 86
rect -423 69 -415 86
rect -352 69 -344 86
rect -327 69 -319 86
rect -256 69 -248 86
rect -231 69 -223 86
rect -160 69 -152 86
rect -135 69 -127 86
rect -64 69 -56 86
rect -39 69 -31 86
rect 31 69 39 86
rect 56 69 64 86
rect 127 69 135 86
rect 152 69 160 86
rect 223 69 231 86
rect 248 69 256 86
rect 319 69 327 86
rect 344 69 352 86
rect 415 69 423 86
rect 440 69 448 86
rect 511 69 519 86
rect 536 69 544 86
rect 607 69 615 86
rect 632 69 640 86
rect 703 69 711 86
rect 728 69 736 86
rect -881 -120 -864 -89
rect -824 44 -807 52
rect -824 -69 -807 -44
rect -776 44 -759 52
rect -776 -52 -759 -44
rect -728 44 -711 52
rect -728 -52 -711 -44
rect -680 44 -663 52
rect -680 -52 -663 -44
rect -632 44 -615 52
rect -632 -52 -615 -44
rect -584 44 -567 52
rect -584 -52 -567 -44
rect -536 44 -519 52
rect -536 -52 -519 -44
rect -488 44 -471 52
rect -488 -52 -471 -44
rect -440 44 -423 52
rect -440 -52 -423 -44
rect -392 44 -375 52
rect -392 -52 -375 -44
rect -344 44 -327 52
rect -344 -52 -327 -44
rect -296 44 -279 52
rect -296 -52 -279 -44
rect -248 44 -231 52
rect -248 -52 -231 -44
rect -200 44 -183 52
rect -200 -52 -183 -44
rect -152 44 -135 52
rect -152 -52 -135 -44
rect -104 44 -87 52
rect -104 -52 -87 -44
rect -56 44 -39 52
rect -56 -52 -39 -44
rect -8 44 8 52
rect -8 -52 8 -44
rect 39 44 56 52
rect 39 -52 56 -44
rect 87 44 104 52
rect 87 -52 104 -44
rect 135 44 152 52
rect 135 -52 152 -44
rect 183 44 200 52
rect 183 -52 200 -44
rect 231 44 248 52
rect 231 -52 248 -44
rect 279 44 296 52
rect 279 -52 296 -44
rect 327 44 344 52
rect 327 -52 344 -44
rect 375 44 392 52
rect 375 -52 392 -44
rect 423 44 440 52
rect 423 -52 440 -44
rect 471 44 488 52
rect 471 -52 488 -44
rect 519 44 536 52
rect 519 -52 536 -44
rect 567 44 584 52
rect 567 -52 584 -44
rect 615 44 632 52
rect 615 -52 632 -44
rect 663 44 680 52
rect 663 -52 680 -44
rect 711 44 728 52
rect 711 -52 728 -44
rect 759 44 776 52
rect 759 -52 776 -44
rect 807 44 824 52
rect -824 -86 -800 -69
rect -783 -86 -775 -69
rect 807 -71 824 -44
rect -824 -120 -807 -86
rect 775 -88 783 -71
rect 800 -88 824 -71
rect 807 -120 824 -88
rect 864 -120 881 -89
rect -881 -137 -833 -120
rect 833 -137 881 -120
<< viali >>
rect -728 69 -711 86
rect -632 69 -615 86
rect -536 69 -519 86
rect -440 69 -423 86
rect -344 69 -327 86
rect -248 69 -231 86
rect -152 69 -135 86
rect -56 69 -39 86
rect 39 69 56 86
rect 135 69 152 86
rect 231 69 248 86
rect 327 69 344 86
rect 423 69 440 86
rect 519 69 536 86
rect 615 69 632 86
rect 711 69 728 86
<< metal1 >>
rect -734 86 -705 89
rect -734 69 -728 86
rect -711 69 -705 86
rect -734 66 -705 69
rect -638 86 -609 89
rect -638 69 -632 86
rect -615 69 -609 86
rect -638 66 -609 69
rect -542 86 -513 89
rect -542 69 -536 86
rect -519 69 -513 86
rect -542 66 -513 69
rect -446 86 -417 89
rect -446 69 -440 86
rect -423 69 -417 86
rect -446 66 -417 69
rect -350 86 -321 89
rect -350 69 -344 86
rect -327 69 -321 86
rect -350 66 -321 69
rect -254 86 -225 89
rect -254 69 -248 86
rect -231 69 -225 86
rect -254 66 -225 69
rect -158 86 -129 89
rect -158 69 -152 86
rect -135 69 -129 86
rect -158 66 -129 69
rect -62 86 -33 89
rect -62 69 -56 86
rect -39 69 -33 86
rect -62 66 -33 69
rect 33 86 62 89
rect 33 69 39 86
rect 56 69 62 86
rect 33 66 62 69
rect 129 86 158 89
rect 129 69 135 86
rect 152 69 158 86
rect 129 66 158 69
rect 225 86 254 89
rect 225 69 231 86
rect 248 69 254 86
rect 225 66 254 69
rect 321 86 350 89
rect 321 69 327 86
rect 344 69 350 86
rect 321 66 350 69
rect 417 86 446 89
rect 417 69 423 86
rect 440 69 446 86
rect 417 66 446 69
rect 513 86 542 89
rect 513 69 519 86
rect 536 69 542 86
rect 513 66 542 69
rect 609 86 638 89
rect 609 69 615 86
rect 632 69 638 86
rect 609 66 638 69
rect 705 86 734 89
rect 705 69 711 86
rect 728 69 734 86
rect 705 66 734 69
<< properties >>
string FIXED_BBOX -873 -128 873 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 34 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
