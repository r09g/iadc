magic
tech sky130A
magscale 1 2
timestamp 1655495960
<< nwell >>
rect -3377 -295 -2714 26
rect -3377 -1383 -2469 -817
rect -3377 -2471 -2469 -1905
rect -3377 -3559 -2469 -2993
rect -3377 -4647 -2469 -4081
rect -3377 -5735 -2469 -5169
rect -3377 -6823 -2223 -6257
rect -3377 -7911 -2469 -7345
rect -3377 -8999 -2469 -8433
rect -3377 -10087 -2469 -9521
rect -3377 -11175 -2469 -10609
rect -3377 -12263 -2469 -11697
rect -3377 -13351 -2469 -12785
rect -3377 -14194 -2714 -13873
<< pwell >>
rect -3034 -535 17037 -361
rect -3034 -751 17037 -577
rect -3034 -1623 17037 -1449
rect -3034 -1839 17037 -1665
rect -3034 -2711 17037 -2537
rect -3034 -2927 17037 -2753
rect -3034 -3799 17037 -3625
rect -3034 -4015 17037 -3841
rect -3034 -4887 17037 -4713
rect -3034 -5103 17037 -4929
rect -948 -5793 -896 -5780
rect -3034 -5975 17037 -5801
rect -3034 -6191 17037 -6017
rect -3034 -7063 17037 -6889
rect -3034 -7279 17037 -7105
rect -3035 -8124 17044 -7976
rect -3034 -8151 17037 -8124
rect -3034 -8220 17037 -8193
rect -3034 -8368 17044 -8220
rect -3035 -9212 17044 -9064
rect -3034 -9239 17037 -9212
rect -3034 -9308 17037 -9281
rect -3034 -9456 17044 -9308
rect -3035 -10300 17044 -10152
rect -3034 -10327 17037 -10300
rect -3034 -10396 17037 -10369
rect -3034 -10544 17044 -10396
rect -3035 -11388 17044 -11240
rect -3034 -11415 17037 -11388
rect -3034 -11484 17037 -11457
rect -3034 -11632 17044 -11484
rect -3035 -12476 17044 -12328
rect -3034 -12503 17037 -12476
rect -3034 -12572 17037 -12545
rect -3034 -12720 17044 -12572
rect -3035 -13564 17044 -13416
rect -3034 -13591 17037 -13564
rect -3034 -13660 17037 -13633
rect -3034 -13808 17044 -13660
<< psubdiff >>
rect 16908 -402 16972 -378
rect 16908 -490 16972 -466
rect 16908 -646 16972 -622
rect 16908 -734 16972 -710
rect 16908 -1490 16972 -1466
rect 16908 -1578 16972 -1554
rect 16908 -1734 16972 -1710
rect 16908 -1822 16972 -1798
rect 16908 -2578 16972 -2554
rect 16908 -2666 16972 -2642
rect 16908 -2822 16972 -2798
rect 16908 -2910 16972 -2886
rect 16908 -3666 16972 -3642
rect 16908 -3754 16972 -3730
rect 16908 -3910 16972 -3886
rect 16908 -3998 16972 -3974
rect 16908 -4754 16972 -4730
rect 16908 -4842 16972 -4818
rect 16908 -4998 16972 -4974
rect 16908 -5086 16972 -5062
rect 16908 -5842 16972 -5818
rect 16908 -5930 16972 -5906
rect 16908 -6086 16972 -6062
rect 16908 -6174 16972 -6150
rect 16908 -6930 16972 -6906
rect 16908 -7018 16972 -6994
rect 16908 -7174 16972 -7150
rect 16908 -7262 16972 -7238
rect 16908 -8018 16972 -7994
rect 16908 -8106 16972 -8082
rect 16908 -8262 16972 -8238
rect 16908 -8350 16972 -8326
rect 16908 -9106 16972 -9082
rect 16908 -9194 16972 -9170
rect 16908 -9350 16972 -9326
rect 16908 -9438 16972 -9414
rect 16908 -10194 16972 -10170
rect 16908 -10282 16972 -10258
rect 16908 -10438 16972 -10414
rect 16908 -10526 16972 -10502
rect 16908 -11282 16972 -11258
rect 16908 -11370 16972 -11346
rect 16908 -11526 16972 -11502
rect 16908 -11614 16972 -11590
rect 16908 -12370 16972 -12346
rect 16908 -12458 16972 -12434
rect 16908 -12614 16972 -12590
rect 16908 -12702 16972 -12678
rect 16908 -13458 16972 -13434
rect 16908 -13546 16972 -13522
rect 16908 -13702 16972 -13678
rect 16908 -13790 16972 -13766
<< nsubdiff >>
rect -3279 -104 -3215 -80
rect -3279 -192 -3215 -168
rect -3279 -947 -3215 -923
rect -3279 -1035 -3215 -1011
rect -3279 -1192 -3215 -1168
rect -3279 -1280 -3215 -1256
rect -3279 -2035 -3215 -2011
rect -3279 -2123 -3215 -2099
rect -3279 -2280 -3215 -2256
rect -3279 -2368 -3215 -2344
rect -3279 -3123 -3215 -3099
rect -3279 -3211 -3215 -3187
rect -3279 -3368 -3215 -3344
rect -3279 -3456 -3215 -3432
rect -3279 -4211 -3215 -4187
rect -3279 -4299 -3215 -4275
rect -3279 -4456 -3215 -4432
rect -3279 -4544 -3215 -4520
rect -3279 -5299 -3215 -5275
rect -3279 -5387 -3215 -5363
rect -3279 -5544 -3215 -5520
rect -3279 -5632 -3215 -5608
rect -3279 -6387 -3215 -6363
rect -3279 -6475 -3215 -6451
rect -3279 -6632 -3215 -6608
rect -3279 -6720 -3215 -6696
rect -3279 -7475 -3215 -7451
rect -3279 -7563 -3215 -7539
rect -3279 -7720 -3215 -7696
rect -3279 -7808 -3215 -7784
rect -3279 -8563 -3215 -8539
rect -3279 -8651 -3215 -8627
rect -3279 -8808 -3215 -8784
rect -3279 -8896 -3215 -8872
rect -3279 -9651 -3215 -9627
rect -3279 -9739 -3215 -9715
rect -3279 -9896 -3215 -9872
rect -3279 -9984 -3215 -9960
rect -3279 -10739 -3215 -10715
rect -3279 -10827 -3215 -10803
rect -3279 -10984 -3215 -10960
rect -3279 -11072 -3215 -11048
rect -3279 -11827 -3215 -11803
rect -3279 -11915 -3215 -11891
rect -3279 -12072 -3215 -12048
rect -3279 -12160 -3215 -12136
rect -3279 -12915 -3215 -12891
rect -3279 -13003 -3215 -12979
rect -3279 -13160 -3215 -13136
rect -3279 -13248 -3215 -13224
rect -3279 -14003 -3215 -13979
rect -3279 -14091 -3215 -14067
<< psubdiffcont >>
rect 16908 -466 16972 -402
rect 16908 -710 16972 -646
rect 16908 -1554 16972 -1490
rect 16908 -1798 16972 -1734
rect 16908 -2642 16972 -2578
rect 16908 -2886 16972 -2822
rect 16908 -3730 16972 -3666
rect 16908 -3974 16972 -3910
rect 16908 -4818 16972 -4754
rect 16908 -5062 16972 -4998
rect 16908 -5906 16972 -5842
rect 16908 -6150 16972 -6086
rect 16908 -6994 16972 -6930
rect 16908 -7238 16972 -7174
rect 16908 -8082 16972 -8018
rect 16908 -8326 16972 -8262
rect 16908 -9170 16972 -9106
rect 16908 -9414 16972 -9350
rect 16908 -10258 16972 -10194
rect 16908 -10502 16972 -10438
rect 16908 -11346 16972 -11282
rect 16908 -11590 16972 -11526
rect 16908 -12434 16972 -12370
rect 16908 -12678 16972 -12614
rect 16908 -13522 16972 -13458
rect 16908 -13766 16972 -13702
<< nsubdiffcont >>
rect -3279 -168 -3215 -104
rect -3279 -1011 -3215 -947
rect -3279 -1256 -3215 -1192
rect -3279 -2099 -3215 -2035
rect -3279 -2344 -3215 -2280
rect -3279 -3187 -3215 -3123
rect -3279 -3432 -3215 -3368
rect -3279 -4275 -3215 -4211
rect -3279 -4520 -3215 -4456
rect -3279 -5363 -3215 -5299
rect -3279 -5608 -3215 -5544
rect -3279 -6451 -3215 -6387
rect -3279 -6696 -3215 -6632
rect -3279 -7539 -3215 -7475
rect -3279 -7784 -3215 -7720
rect -3279 -8627 -3215 -8563
rect -3279 -8872 -3215 -8808
rect -3279 -9715 -3215 -9651
rect -3279 -9960 -3215 -9896
rect -3279 -10803 -3215 -10739
rect -3279 -11048 -3215 -10984
rect -3279 -11891 -3215 -11827
rect -3279 -12136 -3215 -12072
rect -3279 -12979 -3215 -12915
rect -3279 -13224 -3215 -13160
rect -3279 -14067 -3215 -14003
<< locali >>
rect -3311 -29 -2971 5
rect -3311 -104 -3183 -29
rect -3311 -168 -3279 -104
rect -3215 -168 -3183 -104
rect -3311 -947 -3183 -168
rect 434 -294 468 -260
rect 16878 -402 17006 5
rect 16878 -466 16908 -402
rect 16972 -466 17006 -402
rect 16878 -539 17006 -466
rect 16662 -573 17006 -539
rect 16878 -646 17006 -573
rect 16878 -710 16908 -646
rect 16972 -710 17006 -646
rect -3311 -1011 -3279 -947
rect -3215 -1011 -3183 -947
rect -3311 -1083 -3183 -1011
rect -3311 -1117 -2992 -1083
rect -3311 -1192 -3183 -1117
rect -3311 -1256 -3279 -1192
rect -3215 -1256 -3183 -1192
rect -3311 -2035 -3183 -1256
rect 16878 -1490 17006 -710
rect 16878 -1554 16908 -1490
rect 16972 -1554 17006 -1490
rect 16878 -1627 17006 -1554
rect 16662 -1661 17006 -1627
rect 16878 -1734 17006 -1661
rect 16878 -1798 16908 -1734
rect 16972 -1798 17006 -1734
rect -857 -1934 -856 -1900
rect -3311 -2099 -3279 -2035
rect -3215 -2099 -3183 -2035
rect -3311 -2171 -3183 -2099
rect -3311 -2205 -2968 -2171
rect -3311 -2280 -3183 -2205
rect -3311 -2344 -3279 -2280
rect -3215 -2344 -3183 -2280
rect -3311 -3123 -3183 -2344
rect 16878 -2578 17006 -1798
rect 16878 -2642 16908 -2578
rect 16972 -2642 17006 -2578
rect 16878 -2715 17006 -2642
rect 16662 -2749 17006 -2715
rect 16878 -2822 17006 -2749
rect 16878 -2886 16908 -2822
rect 16972 -2886 17006 -2822
rect -3311 -3187 -3279 -3123
rect -3215 -3187 -3183 -3123
rect -3311 -3259 -3183 -3187
rect -3311 -3293 -2968 -3259
rect -3311 -3368 -3183 -3293
rect -3311 -3432 -3279 -3368
rect -3215 -3432 -3183 -3368
rect -3311 -4211 -3183 -3432
rect 16878 -3666 17006 -2886
rect 16878 -3730 16908 -3666
rect 16972 -3730 17006 -3666
rect 16878 -3803 17006 -3730
rect 16662 -3837 17006 -3803
rect 16878 -3910 17006 -3837
rect 16878 -3974 16908 -3910
rect 16972 -3974 17006 -3910
rect -3311 -4275 -3279 -4211
rect -3215 -4275 -3183 -4211
rect -3311 -4347 -3183 -4275
rect -3311 -4381 -2968 -4347
rect -3311 -4456 -3183 -4381
rect -3311 -4520 -3279 -4456
rect -3215 -4520 -3183 -4456
rect -3311 -5299 -3183 -4520
rect 16878 -4754 17006 -3974
rect 16878 -4818 16908 -4754
rect 16972 -4818 17006 -4754
rect 16878 -4891 17006 -4818
rect 16662 -4925 17006 -4891
rect 16878 -4998 17006 -4925
rect 16878 -5062 16908 -4998
rect 16972 -5062 17006 -4998
rect -3311 -5363 -3279 -5299
rect -3215 -5363 -3183 -5299
rect -3311 -5435 -3183 -5363
rect -3311 -5469 -2968 -5435
rect -3311 -5544 -3183 -5469
rect -3311 -5608 -3279 -5544
rect -3215 -5608 -3183 -5544
rect -3311 -6387 -3183 -5608
rect 16878 -5842 17006 -5062
rect 16878 -5906 16908 -5842
rect 16972 -5906 17006 -5842
rect 16878 -5979 17006 -5906
rect 16662 -6013 17006 -5979
rect 16878 -6086 17006 -6013
rect 16878 -6150 16908 -6086
rect 16972 -6150 17006 -6086
rect 434 -6292 468 -6258
rect -3311 -6451 -3279 -6387
rect -3215 -6451 -3183 -6387
rect -3311 -6523 -3183 -6451
rect -3311 -6557 -2968 -6523
rect -3311 -6632 -3183 -6557
rect -3311 -6696 -3279 -6632
rect -3215 -6696 -3183 -6632
rect -3311 -7475 -3183 -6696
rect 16878 -6930 17006 -6150
rect 16878 -6994 16908 -6930
rect 16972 -6994 17006 -6930
rect 16878 -7067 17006 -6994
rect 16662 -7101 17006 -7067
rect 16878 -7174 17006 -7101
rect 16878 -7238 16908 -7174
rect 16972 -7238 17006 -7174
rect -3311 -7539 -3279 -7475
rect -3215 -7539 -3183 -7475
rect -3311 -7611 -3183 -7539
rect -3311 -7645 -2968 -7611
rect -3311 -7720 -3183 -7645
rect -3311 -7784 -3279 -7720
rect -3215 -7784 -3183 -7720
rect -3311 -8563 -3183 -7784
rect 434 -7910 468 -7876
rect 16878 -8018 17006 -7238
rect 16878 -8082 16908 -8018
rect 16972 -8082 17006 -8018
rect 16878 -8155 17006 -8082
rect 16662 -8189 17006 -8155
rect 16878 -8262 17006 -8189
rect 16878 -8326 16908 -8262
rect 16972 -8326 17006 -8262
rect -3311 -8627 -3279 -8563
rect -3215 -8627 -3183 -8563
rect -3311 -8699 -3183 -8627
rect -3311 -8733 -2968 -8699
rect -3311 -8808 -3183 -8733
rect -3311 -8872 -3279 -8808
rect -3215 -8872 -3183 -8808
rect -3311 -9651 -3183 -8872
rect 16878 -9106 17006 -8326
rect 16878 -9170 16908 -9106
rect 16972 -9170 17006 -9106
rect 16878 -9243 17006 -9170
rect 16662 -9277 17006 -9243
rect 16878 -9350 17006 -9277
rect 16878 -9414 16908 -9350
rect 16972 -9414 17006 -9350
rect -857 -9550 -856 -9516
rect -3311 -9715 -3279 -9651
rect -3215 -9715 -3183 -9651
rect -3311 -9787 -3183 -9715
rect -3311 -9821 -2968 -9787
rect -3311 -9896 -3183 -9821
rect -3311 -9960 -3279 -9896
rect -3215 -9960 -3183 -9896
rect -3311 -10739 -3183 -9960
rect 16878 -10194 17006 -9414
rect 16878 -10258 16908 -10194
rect 16972 -10258 17006 -10194
rect 16878 -10331 17006 -10258
rect 16662 -10365 17006 -10331
rect 16878 -10438 17006 -10365
rect 16878 -10502 16908 -10438
rect 16972 -10502 17006 -10438
rect -3311 -10803 -3279 -10739
rect -3215 -10803 -3183 -10739
rect -3311 -10875 -3183 -10803
rect -3311 -10909 -2968 -10875
rect -3311 -10984 -3183 -10909
rect -3311 -11048 -3279 -10984
rect -3215 -11048 -3183 -10984
rect -3311 -11827 -3183 -11048
rect 16878 -11282 17006 -10502
rect 16878 -11346 16908 -11282
rect 16972 -11346 17006 -11282
rect 16878 -11419 17006 -11346
rect 16662 -11453 17006 -11419
rect 16878 -11526 17006 -11453
rect 16878 -11590 16908 -11526
rect 16972 -11590 17006 -11526
rect -3311 -11891 -3279 -11827
rect -3215 -11891 -3183 -11827
rect -3311 -11963 -3183 -11891
rect -3311 -11997 -2968 -11963
rect -3311 -12072 -3183 -11997
rect -3311 -12136 -3279 -12072
rect -3215 -12136 -3183 -12072
rect -3311 -12915 -3183 -12136
rect 16878 -12370 17006 -11590
rect 16878 -12434 16908 -12370
rect 16972 -12434 17006 -12370
rect 16878 -12507 17006 -12434
rect 16662 -12541 17006 -12507
rect 16878 -12614 17006 -12541
rect 16878 -12678 16908 -12614
rect 16972 -12678 17006 -12614
rect -3311 -12979 -3279 -12915
rect -3215 -12979 -3183 -12915
rect -3311 -13051 -3183 -12979
rect -3311 -13085 -2968 -13051
rect -3311 -13160 -3183 -13085
rect -3311 -13224 -3279 -13160
rect -3215 -13224 -3183 -13160
rect -3311 -14003 -3183 -13224
rect 16878 -13458 17006 -12678
rect 16878 -13522 16908 -13458
rect 16972 -13522 17006 -13458
rect 16878 -13595 17006 -13522
rect 16663 -13629 17006 -13595
rect 16878 -13702 17006 -13629
rect 16878 -13766 16908 -13702
rect 16972 -13766 17006 -13702
rect 434 -13908 468 -13874
rect -850 -13960 -816 -13926
rect -3311 -14067 -3279 -14003
rect -3215 -14067 -3183 -14003
rect -3311 -14139 -3183 -14067
rect -3311 -14173 -2968 -14139
rect 16878 -14173 17006 -13766
<< viali >>
rect -943 -335 -909 -301
rect -762 -335 -728 -301
rect -30 -341 4 -307
rect 106 -341 140 -307
rect 242 -341 276 -307
rect 434 -379 468 -345
rect 1076 -346 1110 -312
rect 1171 -340 1205 -306
rect 1263 -340 1297 -306
rect 2369 -335 2403 -301
rect 3015 -336 3049 -302
rect 6876 -336 6910 -302
rect 7522 -336 7556 -302
rect 8164 -337 8198 -303
rect 8811 -335 8845 -301
rect 9453 -335 9487 -301
rect 10099 -334 10133 -300
rect 10741 -335 10775 -301
rect 10832 -335 10866 -301
rect 11129 -302 11163 -268
rect 10925 -336 10959 -302
rect 11017 -336 11051 -302
rect 11250 -333 11284 -299
rect 11344 -333 11378 -299
rect -848 -446 -814 -412
rect -769 -446 -735 -412
rect 1076 -419 1110 -385
rect 1052 -809 1086 -775
rect 3012 -809 3046 -775
rect 3626 -809 3660 -775
rect 5586 -809 5620 -775
rect 6200 -809 6234 -775
rect 8160 -809 8194 -775
rect 8774 -809 8808 -775
rect 10737 -811 10771 -777
rect 11369 -812 11403 -778
rect 13685 -780 13719 -746
rect 15248 -762 15282 -728
rect 15340 -763 15374 -729
rect 433 -846 467 -812
rect 15248 -858 15282 -824
rect 15341 -858 15375 -824
rect 11387 -1389 11421 -1355
rect 15248 -1372 15282 -1338
rect 15340 -1373 15374 -1339
rect 432 -1426 466 -1392
rect 1082 -1423 1116 -1389
rect 3042 -1423 3076 -1389
rect 3656 -1423 3690 -1389
rect 5616 -1423 5650 -1389
rect 6230 -1423 6264 -1389
rect 8190 -1423 8224 -1389
rect 8804 -1423 8838 -1389
rect 10764 -1423 10798 -1389
rect 12558 -1426 12592 -1392
rect 12642 -1426 12676 -1392
rect 12739 -1426 12773 -1392
rect 12836 -1426 12870 -1392
rect 12942 -1426 12976 -1392
rect 13038 -1419 13072 -1385
rect 13684 -1456 13718 -1422
rect 13038 -1491 13072 -1457
rect 15248 -1468 15282 -1434
rect 15341 -1468 15375 -1434
rect -210 -1899 -176 -1865
rect 1054 -1900 1088 -1866
rect 3014 -1900 3048 -1866
rect 3628 -1900 3662 -1866
rect 5588 -1900 5622 -1866
rect 6202 -1900 6236 -1866
rect 8162 -1900 8196 -1866
rect 8776 -1900 8810 -1866
rect 10736 -1900 10770 -1866
rect 11386 -1897 11420 -1863
rect 13685 -1866 13719 -1832
rect 15248 -1850 15282 -1816
rect 15340 -1851 15374 -1817
rect -856 -1934 -822 -1900
rect 432 -1934 466 -1900
rect 15248 -1946 15282 -1912
rect 15341 -1946 15375 -1912
rect 12480 -2441 12514 -2407
rect 436 -2514 470 -2480
rect 1081 -2512 1115 -2478
rect 3041 -2512 3075 -2478
rect 3655 -2512 3689 -2478
rect 5615 -2512 5649 -2478
rect 6229 -2512 6263 -2478
rect 8189 -2512 8223 -2478
rect 8806 -2512 8840 -2478
rect 10763 -2512 10797 -2478
rect 11386 -2479 11420 -2445
rect 15248 -2460 15282 -2426
rect 15340 -2460 15374 -2426
rect 12480 -2515 12514 -2481
rect 12568 -2513 12602 -2479
rect 12659 -2513 12693 -2479
rect 12765 -2513 12799 -2479
rect 12858 -2511 12892 -2477
rect 12942 -2511 12976 -2477
rect 13039 -2500 13073 -2466
rect 12480 -2587 12514 -2553
rect 13042 -2577 13076 -2543
rect 13685 -2544 13719 -2510
rect 15248 -2556 15282 -2522
rect 15341 -2556 15375 -2522
rect -1783 -2949 -1749 -2915
rect -1960 -2986 -1926 -2952
rect 1072 -2986 1106 -2952
rect 3016 -2987 3050 -2953
rect 3630 -2987 3664 -2953
rect 5590 -2987 5624 -2953
rect 6204 -2987 6238 -2953
rect 8164 -2987 8198 -2953
rect 8778 -2987 8812 -2953
rect 429 -3021 463 -2987
rect 10738 -2988 10772 -2954
rect 11384 -2986 11418 -2952
rect 432 -3565 466 -3531
rect 1070 -3602 1104 -3568
rect 3016 -3599 3050 -3565
rect 3630 -3599 3664 -3565
rect 5590 -3599 5624 -3565
rect 6204 -3599 6238 -3565
rect 8164 -3599 8198 -3565
rect 8778 -3599 8812 -3565
rect 10735 -3602 10769 -3568
rect 11383 -3601 11417 -3567
rect 12480 -3999 12514 -3965
rect 13042 -4009 13076 -3975
rect 436 -4074 470 -4040
rect 1081 -4074 1115 -4040
rect 3041 -4074 3075 -4040
rect 3655 -4074 3689 -4040
rect 5615 -4074 5649 -4040
rect 6229 -4074 6263 -4040
rect 8189 -4074 8223 -4040
rect 8806 -4074 8840 -4040
rect 10763 -4074 10797 -4040
rect 12480 -4071 12514 -4037
rect 12568 -4073 12602 -4039
rect 12659 -4073 12693 -4039
rect 12765 -4073 12799 -4039
rect 12858 -4075 12892 -4041
rect 12942 -4075 12976 -4041
rect 13685 -4042 13719 -4008
rect 15248 -4030 15282 -3996
rect 15341 -4030 15375 -3996
rect 11386 -4111 11420 -4077
rect 13039 -4086 13073 -4052
rect 12480 -4145 12514 -4111
rect 15248 -4126 15282 -4092
rect 15340 -4126 15374 -4092
rect -855 -4653 -821 -4619
rect 433 -4653 467 -4619
rect 15248 -4640 15282 -4606
rect 15341 -4640 15375 -4606
rect -210 -4690 -176 -4656
rect 1054 -4686 1088 -4652
rect 3014 -4686 3048 -4652
rect 3628 -4686 3662 -4652
rect 5588 -4686 5622 -4652
rect 6202 -4686 6236 -4652
rect 8162 -4686 8196 -4652
rect 8776 -4686 8810 -4652
rect 10736 -4686 10770 -4652
rect 11384 -4691 11418 -4657
rect 13685 -4720 13719 -4686
rect 15248 -4736 15282 -4702
rect 15340 -4735 15374 -4701
rect 13038 -5095 13072 -5061
rect 436 -5162 470 -5128
rect 1082 -5163 1116 -5129
rect 3042 -5163 3076 -5129
rect 3656 -5163 3690 -5129
rect 5616 -5163 5650 -5129
rect 6230 -5163 6264 -5129
rect 8190 -5163 8224 -5129
rect 8804 -5163 8838 -5129
rect 10764 -5163 10798 -5129
rect 12558 -5160 12592 -5126
rect 12642 -5160 12676 -5126
rect 12739 -5160 12773 -5126
rect 12836 -5160 12870 -5126
rect 12942 -5160 12976 -5126
rect 13684 -5130 13718 -5096
rect 15248 -5118 15282 -5084
rect 15341 -5118 15375 -5084
rect 11389 -5196 11423 -5162
rect 13038 -5167 13072 -5133
rect 15248 -5214 15282 -5180
rect 15340 -5213 15374 -5179
rect 432 -5742 466 -5708
rect 15248 -5728 15282 -5694
rect 15341 -5728 15375 -5694
rect 1052 -5777 1086 -5743
rect 3012 -5777 3046 -5743
rect 3626 -5777 3660 -5743
rect 5586 -5777 5620 -5743
rect 6200 -5777 6234 -5743
rect 8160 -5777 8194 -5743
rect 8774 -5777 8808 -5743
rect 10737 -5775 10771 -5741
rect 11369 -5774 11403 -5740
rect 13685 -5806 13719 -5772
rect 15248 -5824 15282 -5790
rect 15340 -5823 15374 -5789
rect -848 -6140 -814 -6106
rect -769 -6140 -735 -6106
rect 1076 -6167 1110 -6133
rect 434 -6207 468 -6173
rect -932 -6252 -898 -6218
rect -760 -6251 -726 -6217
rect -30 -6245 4 -6211
rect 106 -6245 140 -6211
rect 242 -6245 276 -6211
rect 1076 -6240 1110 -6206
rect 1171 -6246 1205 -6212
rect 1263 -6246 1297 -6212
rect 2369 -6251 2403 -6217
rect 3015 -6250 3049 -6216
rect 6876 -6250 6910 -6216
rect 7522 -6250 7556 -6216
rect 8164 -6249 8198 -6215
rect 8811 -6251 8845 -6217
rect 9453 -6251 9487 -6217
rect 10099 -6252 10133 -6218
rect 10741 -6251 10775 -6217
rect 10832 -6251 10866 -6217
rect 10925 -6250 10959 -6216
rect 11017 -6250 11051 -6216
rect 11129 -6284 11163 -6250
rect 11250 -6253 11284 -6219
rect 11344 -6253 11378 -6219
rect -2599 -6864 -2565 -6830
rect -2343 -6916 -2309 -6882
rect -940 -6914 -906 -6880
rect -1233 -6994 -1199 -6960
rect 3111 -7225 3145 -7191
rect 3852 -7222 3886 -7188
rect 4955 -7238 4989 -7204
rect 6245 -7214 6279 -7180
rect 2934 -7304 2968 -7270
rect 7356 -7298 7390 -7264
rect 3747 -7338 3781 -7304
rect 3928 -7339 3962 -7305
rect 4565 -7338 4599 -7304
rect 5036 -7340 5070 -7306
rect 7604 -7324 7638 -7290
rect 5171 -7407 5205 -7373
rect 7605 -7398 7639 -7364
rect -937 -7952 -903 -7918
rect -762 -7951 -728 -7917
rect -30 -7957 4 -7923
rect 106 -7957 140 -7923
rect 242 -7957 276 -7923
rect 434 -7995 468 -7961
rect 1076 -7962 1110 -7928
rect 1171 -7956 1205 -7922
rect 1263 -7956 1297 -7922
rect 2369 -7951 2403 -7917
rect 3015 -7952 3049 -7918
rect 6876 -7952 6910 -7918
rect 7522 -7952 7556 -7918
rect 8164 -7953 8198 -7919
rect 8811 -7951 8845 -7917
rect 9453 -7951 9487 -7917
rect 10099 -7950 10133 -7916
rect 10741 -7951 10775 -7917
rect 10832 -7951 10866 -7917
rect 11129 -7918 11163 -7884
rect 10925 -7952 10959 -7918
rect 11017 -7952 11051 -7918
rect 11250 -7949 11284 -7915
rect 11344 -7949 11378 -7915
rect -848 -8062 -814 -8028
rect -769 -8062 -735 -8028
rect 1076 -8035 1110 -8001
rect 1052 -8425 1086 -8391
rect 3012 -8425 3046 -8391
rect 3626 -8425 3660 -8391
rect 5586 -8425 5620 -8391
rect 6200 -8425 6234 -8391
rect 8160 -8425 8194 -8391
rect 8774 -8425 8808 -8391
rect 10737 -8427 10771 -8393
rect 11369 -8428 11403 -8394
rect 13685 -8396 13719 -8362
rect 15248 -8378 15282 -8344
rect 15340 -8379 15374 -8345
rect 433 -8462 467 -8428
rect 15248 -8474 15282 -8440
rect 15341 -8474 15375 -8440
rect 11387 -9005 11421 -8971
rect 15248 -8988 15282 -8954
rect 15340 -8989 15374 -8955
rect 432 -9042 466 -9008
rect 1082 -9039 1116 -9005
rect 3042 -9039 3076 -9005
rect 3656 -9039 3690 -9005
rect 5616 -9039 5650 -9005
rect 6230 -9039 6264 -9005
rect 8190 -9039 8224 -9005
rect 8804 -9039 8838 -9005
rect 10764 -9039 10798 -9005
rect 12558 -9042 12592 -9008
rect 12642 -9042 12676 -9008
rect 12739 -9042 12773 -9008
rect 12836 -9042 12870 -9008
rect 12942 -9042 12976 -9008
rect 13038 -9035 13072 -9001
rect 13684 -9072 13718 -9038
rect 13038 -9107 13072 -9073
rect 15248 -9084 15282 -9050
rect 15341 -9084 15375 -9050
rect -210 -9515 -176 -9481
rect 1054 -9516 1088 -9482
rect 3014 -9516 3048 -9482
rect 3628 -9516 3662 -9482
rect 5588 -9516 5622 -9482
rect 6202 -9516 6236 -9482
rect 8162 -9516 8196 -9482
rect 8776 -9516 8810 -9482
rect 10736 -9516 10770 -9482
rect 11386 -9513 11420 -9479
rect 13685 -9482 13719 -9448
rect 15248 -9466 15282 -9432
rect 15340 -9467 15374 -9433
rect -856 -9550 -822 -9516
rect 432 -9550 466 -9516
rect 15248 -9562 15282 -9528
rect 15341 -9562 15375 -9528
rect 12480 -10057 12514 -10023
rect 436 -10130 470 -10096
rect 1081 -10128 1115 -10094
rect 3041 -10128 3075 -10094
rect 3655 -10128 3689 -10094
rect 5615 -10128 5649 -10094
rect 6229 -10128 6263 -10094
rect 8189 -10128 8223 -10094
rect 8806 -10128 8840 -10094
rect 10763 -10128 10797 -10094
rect 11386 -10095 11420 -10061
rect 15248 -10076 15282 -10042
rect 15340 -10076 15374 -10042
rect 12480 -10131 12514 -10097
rect 12568 -10129 12602 -10095
rect 12659 -10129 12693 -10095
rect 12765 -10129 12799 -10095
rect 12858 -10127 12892 -10093
rect 12942 -10127 12976 -10093
rect 13039 -10116 13073 -10082
rect 12480 -10203 12514 -10169
rect 13042 -10193 13076 -10159
rect 13685 -10160 13719 -10126
rect 15248 -10172 15282 -10138
rect 15341 -10172 15375 -10138
rect -1961 -10533 -1927 -10499
rect -1813 -10568 -1779 -10534
rect 1072 -10602 1106 -10568
rect 3016 -10603 3050 -10569
rect 3630 -10603 3664 -10569
rect 5590 -10603 5624 -10569
rect 6204 -10603 6238 -10569
rect 8164 -10603 8198 -10569
rect 8778 -10603 8812 -10569
rect 429 -10637 463 -10603
rect 10738 -10604 10772 -10570
rect 11384 -10602 11418 -10568
rect 432 -11181 466 -11147
rect 1070 -11218 1104 -11184
rect 3016 -11215 3050 -11181
rect 3630 -11215 3664 -11181
rect 5590 -11215 5624 -11181
rect 6204 -11215 6238 -11181
rect 8164 -11215 8198 -11181
rect 8778 -11215 8812 -11181
rect 10735 -11218 10769 -11184
rect 11383 -11217 11417 -11183
rect 12480 -11615 12514 -11581
rect 13042 -11625 13076 -11591
rect 436 -11690 470 -11656
rect 1081 -11690 1115 -11656
rect 3041 -11690 3075 -11656
rect 3655 -11690 3689 -11656
rect 5615 -11690 5649 -11656
rect 6229 -11690 6263 -11656
rect 8189 -11690 8223 -11656
rect 8806 -11690 8840 -11656
rect 10763 -11690 10797 -11656
rect 12480 -11687 12514 -11653
rect 12568 -11689 12602 -11655
rect 12659 -11689 12693 -11655
rect 12765 -11689 12799 -11655
rect 12858 -11691 12892 -11657
rect 12942 -11691 12976 -11657
rect 13685 -11658 13719 -11624
rect 15248 -11646 15282 -11612
rect 15341 -11646 15375 -11612
rect 11386 -11727 11420 -11693
rect 13039 -11702 13073 -11668
rect 12480 -11761 12514 -11727
rect 15248 -11742 15282 -11708
rect 15340 -11742 15374 -11708
rect -855 -12269 -821 -12235
rect 433 -12269 467 -12235
rect 15248 -12256 15282 -12222
rect 15341 -12256 15375 -12222
rect -210 -12306 -176 -12272
rect 1054 -12302 1088 -12268
rect 3014 -12302 3048 -12268
rect 3628 -12302 3662 -12268
rect 5588 -12302 5622 -12268
rect 6202 -12302 6236 -12268
rect 8162 -12302 8196 -12268
rect 8776 -12302 8810 -12268
rect 10736 -12302 10770 -12268
rect 11384 -12307 11418 -12273
rect 13685 -12336 13719 -12302
rect 15248 -12352 15282 -12318
rect 15340 -12351 15374 -12317
rect 13038 -12711 13072 -12677
rect 436 -12778 470 -12744
rect 1082 -12779 1116 -12745
rect 3042 -12779 3076 -12745
rect 3656 -12779 3690 -12745
rect 5616 -12779 5650 -12745
rect 6230 -12779 6264 -12745
rect 8190 -12779 8224 -12745
rect 8804 -12779 8838 -12745
rect 10764 -12779 10798 -12745
rect 12558 -12776 12592 -12742
rect 12642 -12776 12676 -12742
rect 12739 -12776 12773 -12742
rect 12836 -12776 12870 -12742
rect 12942 -12776 12976 -12742
rect 13684 -12746 13718 -12712
rect 15248 -12734 15282 -12700
rect 15341 -12734 15375 -12700
rect 11389 -12812 11423 -12778
rect 13038 -12783 13072 -12749
rect 15248 -12830 15282 -12796
rect 15340 -12829 15374 -12795
rect 432 -13358 466 -13324
rect 15248 -13344 15282 -13310
rect 15341 -13344 15375 -13310
rect 1052 -13393 1086 -13359
rect 3012 -13393 3046 -13359
rect 3626 -13393 3660 -13359
rect 5586 -13393 5620 -13359
rect 6200 -13393 6234 -13359
rect 8160 -13393 8194 -13359
rect 8774 -13393 8808 -13359
rect 10737 -13391 10771 -13357
rect 11369 -13390 11403 -13356
rect 13685 -13422 13719 -13388
rect 15248 -13440 15282 -13406
rect 15340 -13439 15374 -13405
rect -848 -13756 -814 -13722
rect -769 -13756 -735 -13722
rect 1076 -13783 1110 -13749
rect 434 -13823 468 -13789
rect -932 -13868 -898 -13834
rect -764 -13869 -730 -13835
rect -30 -13861 4 -13827
rect 106 -13861 140 -13827
rect 242 -13861 276 -13827
rect 1076 -13856 1110 -13822
rect 1171 -13862 1205 -13828
rect 1263 -13862 1297 -13828
rect 2369 -13867 2403 -13833
rect 3015 -13866 3049 -13832
rect 6876 -13866 6910 -13832
rect 7522 -13866 7556 -13832
rect 8164 -13865 8198 -13831
rect 8811 -13867 8845 -13833
rect 9453 -13867 9487 -13833
rect 10099 -13868 10133 -13834
rect 10741 -13867 10775 -13833
rect 10832 -13867 10866 -13833
rect 10925 -13866 10959 -13832
rect 11017 -13866 11051 -13832
rect 11129 -13900 11163 -13866
rect 11250 -13869 11284 -13835
rect 11344 -13869 11378 -13835
<< metal1 >>
rect 308 -212 11419 -127
rect -1802 -343 -1792 -291
rect -1740 -294 -1730 -291
rect -1740 -301 -896 -294
rect -1740 -335 -943 -301
rect -909 -335 -896 -301
rect -1740 -342 -896 -335
rect -781 -342 -771 -290
rect -719 -342 -709 -290
rect 308 -298 387 -212
rect 1153 -284 1310 -283
rect -57 -307 389 -298
rect -57 -341 -30 -307
rect 4 -341 106 -307
rect 140 -341 242 -307
rect 276 -341 389 -307
rect -1740 -343 -1730 -342
rect -57 -346 389 -341
rect -57 -347 16 -346
rect 94 -347 152 -346
rect 227 -347 389 -346
rect 418 -312 1122 -294
rect 418 -325 1076 -312
rect 418 -345 982 -325
rect -57 -403 12 -347
rect 418 -379 434 -345
rect 468 -377 982 -345
rect 1034 -346 1076 -325
rect 1110 -346 1122 -312
rect 1034 -377 1122 -346
rect 468 -379 1122 -377
rect 418 -385 1122 -379
rect -862 -412 13 -403
rect 418 -405 1076 -385
rect 418 -409 485 -405
rect -862 -446 -848 -412
rect -814 -446 -769 -412
rect -735 -446 13 -412
rect -862 -452 13 -446
rect 1064 -419 1076 -405
rect 1110 -419 1122 -385
rect 1153 -301 2449 -284
rect 1153 -306 2369 -301
rect 1153 -340 1171 -306
rect 1205 -340 1263 -306
rect 1297 -335 2369 -306
rect 2403 -335 2449 -301
rect 1297 -340 2449 -335
rect 1153 -346 2449 -340
rect 2994 -302 6963 -282
rect 2994 -336 3015 -302
rect 3049 -336 6876 -302
rect 6910 -336 6963 -302
rect 1153 -406 1310 -346
rect 2994 -353 6963 -336
rect 7509 -302 8255 -281
rect 7509 -336 7522 -302
rect 7556 -303 8255 -302
rect 7556 -336 8164 -303
rect 7509 -337 8164 -336
rect 8198 -337 8255 -303
rect 7509 -355 8255 -337
rect 8799 -301 9545 -283
rect 8799 -335 8811 -301
rect 8845 -335 9453 -301
rect 9487 -335 9545 -301
rect 8799 -354 9545 -335
rect 10086 -296 11058 -278
rect 10086 -300 11063 -296
rect 10086 -334 10099 -300
rect 10133 -301 11063 -300
rect 10133 -334 10741 -301
rect 10086 -335 10741 -334
rect 10775 -335 10832 -301
rect 10866 -302 11063 -301
rect 10866 -335 10925 -302
rect 10086 -336 10925 -335
rect 10959 -336 11017 -302
rect 11051 -336 11063 -302
rect 11110 -311 11120 -259
rect 11172 -311 11182 -259
rect 11233 -299 11418 -212
rect 10086 -342 11063 -336
rect 11233 -333 11250 -299
rect 11284 -333 11344 -299
rect 11378 -333 11418 -299
rect 11233 -341 11418 -333
rect 10086 -348 11058 -342
rect 1064 -474 1122 -419
rect 1070 -478 1116 -474
rect 13669 -681 13738 -679
rect 966 -733 982 -681
rect 1034 -682 13738 -681
rect 1034 -733 12753 -682
rect 966 -734 12753 -733
rect 12805 -734 13738 -682
rect 966 -736 13738 -734
rect 13669 -746 13738 -736
rect 1040 -770 1098 -769
rect 3000 -770 3058 -769
rect 1040 -775 3058 -770
rect 413 -854 423 -802
rect 475 -854 485 -802
rect 1040 -809 1052 -775
rect 1086 -809 3012 -775
rect 3046 -809 3058 -775
rect 1040 -814 3058 -809
rect 1040 -815 1098 -814
rect 3000 -815 3058 -814
rect 3614 -770 3672 -769
rect 5574 -770 5632 -769
rect 3614 -775 5632 -770
rect 3614 -809 3626 -775
rect 3660 -809 5586 -775
rect 5620 -809 5632 -775
rect 3614 -814 5632 -809
rect 3614 -815 3672 -814
rect 5574 -815 5632 -814
rect 6188 -770 6246 -769
rect 8148 -770 8206 -769
rect 6188 -775 8206 -770
rect 6188 -809 6200 -775
rect 6234 -809 8160 -775
rect 8194 -809 8206 -775
rect 6188 -814 8206 -809
rect 6188 -815 6246 -814
rect 8148 -815 8206 -814
rect 8762 -770 8820 -769
rect 8762 -771 10131 -770
rect 8762 -775 10783 -771
rect 8762 -809 8774 -775
rect 8808 -777 10783 -775
rect 8808 -809 10737 -777
rect 8762 -811 10737 -809
rect 10771 -811 10783 -777
rect 8762 -814 10783 -811
rect 8762 -815 8820 -814
rect 10129 -815 10783 -814
rect 10725 -817 10783 -815
rect 11338 -778 11430 -771
rect 11338 -812 11369 -778
rect 11403 -812 11430 -778
rect 11338 -828 11430 -812
rect 13669 -780 13685 -746
rect 13719 -780 13738 -746
rect 13669 -823 13738 -780
rect 15236 -728 15294 -722
rect 15328 -728 15386 -723
rect 15236 -762 15248 -728
rect 15282 -729 15394 -728
rect 15282 -762 15340 -729
rect 15236 -763 15340 -762
rect 15374 -763 15394 -729
rect 15236 -808 15394 -763
rect 15236 -824 16946 -808
rect 11338 -883 12463 -828
rect 11339 -887 12463 -883
rect 12522 -887 12532 -828
rect 15236 -858 15248 -824
rect 15282 -858 15341 -824
rect 15375 -848 16946 -824
rect 15375 -858 15394 -848
rect 15236 -864 15294 -858
rect 15329 -864 15387 -858
rect 7161 -1232 11181 -1231
rect 7161 -1235 11118 -1232
rect 7155 -1287 7165 -1235
rect 7217 -1284 11118 -1235
rect 11170 -1284 11181 -1232
rect 7217 -1287 11181 -1284
rect 7161 -1293 11181 -1287
rect 15236 -1338 15294 -1332
rect 15328 -1338 15386 -1333
rect 413 -1435 423 -1383
rect 475 -1435 485 -1383
rect 1070 -1384 1128 -1383
rect 3030 -1384 3088 -1383
rect 1070 -1389 3088 -1384
rect 1070 -1423 1082 -1389
rect 1116 -1423 3042 -1389
rect 3076 -1423 3088 -1389
rect 1070 -1428 3088 -1423
rect 1070 -1429 1128 -1428
rect 3030 -1429 3088 -1428
rect 3644 -1384 3702 -1383
rect 5604 -1384 5662 -1383
rect 3644 -1389 5662 -1384
rect 3644 -1423 3656 -1389
rect 3690 -1423 5616 -1389
rect 5650 -1423 5662 -1389
rect 3644 -1428 5662 -1423
rect 3644 -1429 3702 -1428
rect 5604 -1429 5662 -1428
rect 6218 -1384 6276 -1383
rect 8178 -1384 8236 -1383
rect 6218 -1389 8236 -1384
rect 6218 -1423 6230 -1389
rect 6264 -1423 8190 -1389
rect 8224 -1423 8236 -1389
rect 6218 -1428 8236 -1423
rect 6218 -1429 6276 -1428
rect 8178 -1429 8236 -1428
rect 8792 -1384 8850 -1383
rect 10752 -1384 10810 -1383
rect 8792 -1389 10810 -1384
rect 8792 -1423 8804 -1389
rect 8838 -1423 10764 -1389
rect 10798 -1423 10810 -1389
rect 11368 -1397 11378 -1345
rect 11430 -1397 11440 -1345
rect 15236 -1372 15248 -1338
rect 15282 -1339 15394 -1338
rect 15282 -1372 15340 -1339
rect 15236 -1373 15340 -1372
rect 15374 -1352 15394 -1339
rect 15374 -1373 16946 -1352
rect 13026 -1380 13084 -1379
rect 12548 -1386 12752 -1382
rect 12546 -1392 12752 -1386
rect 12804 -1392 12992 -1382
rect 8792 -1428 10810 -1423
rect 8792 -1429 8850 -1428
rect 10752 -1429 10810 -1428
rect 12546 -1426 12558 -1392
rect 12592 -1426 12642 -1392
rect 12676 -1426 12739 -1392
rect 12804 -1426 12836 -1392
rect 12870 -1426 12942 -1392
rect 12976 -1426 12992 -1392
rect 12546 -1432 12752 -1426
rect 12548 -1434 12752 -1432
rect 12804 -1434 12992 -1426
rect 12548 -1435 12992 -1434
rect 13026 -1385 13737 -1380
rect 13026 -1419 13038 -1385
rect 13072 -1419 13737 -1385
rect 13026 -1422 13737 -1419
rect 13026 -1456 13684 -1422
rect 13718 -1456 13737 -1422
rect 13026 -1457 13737 -1456
rect 13026 -1491 13038 -1457
rect 13072 -1490 13737 -1457
rect 15236 -1392 16946 -1373
rect 15236 -1434 15394 -1392
rect 15236 -1468 15248 -1434
rect 15282 -1468 15341 -1434
rect 15375 -1468 15394 -1434
rect 15236 -1474 15294 -1468
rect 15329 -1474 15387 -1468
rect 13072 -1491 13084 -1490
rect 13026 -1498 13084 -1491
rect 13671 -1762 13735 -1761
rect 7153 -1763 13735 -1762
rect 7153 -1815 7163 -1763
rect 7215 -1766 13735 -1763
rect 7215 -1815 12756 -1766
rect 7153 -1816 12756 -1815
rect 12746 -1818 12756 -1816
rect 12808 -1816 13735 -1766
rect 12808 -1818 12818 -1816
rect 13671 -1832 13735 -1816
rect -952 -1943 -942 -1891
rect -890 -1893 -880 -1891
rect -890 -1900 -809 -1893
rect -890 -1934 -856 -1900
rect -822 -1934 -809 -1900
rect -227 -1906 -217 -1854
rect -165 -1906 -155 -1854
rect 1042 -1861 1100 -1860
rect 3002 -1861 3060 -1860
rect 1042 -1866 3060 -1861
rect -890 -1941 -809 -1934
rect -890 -1943 -880 -1941
rect 413 -1942 423 -1890
rect 475 -1942 485 -1890
rect 1042 -1900 1054 -1866
rect 1088 -1900 3014 -1866
rect 3048 -1900 3060 -1866
rect 1042 -1905 3060 -1900
rect 1042 -1906 1100 -1905
rect 3002 -1906 3060 -1905
rect 3616 -1861 3674 -1860
rect 5576 -1861 5634 -1860
rect 3616 -1866 5634 -1861
rect 3616 -1900 3628 -1866
rect 3662 -1900 5588 -1866
rect 5622 -1900 5634 -1866
rect 3616 -1905 5634 -1900
rect 3616 -1906 3674 -1905
rect 5576 -1906 5634 -1905
rect 6190 -1861 6248 -1860
rect 8150 -1861 8208 -1860
rect 6190 -1866 8208 -1861
rect 6190 -1900 6202 -1866
rect 6236 -1900 8162 -1866
rect 8196 -1900 8208 -1866
rect 6190 -1905 8208 -1900
rect 6190 -1906 6248 -1905
rect 8150 -1906 8208 -1905
rect 8764 -1861 8822 -1860
rect 10724 -1861 10782 -1860
rect 8764 -1866 10782 -1861
rect 8764 -1900 8776 -1866
rect 8810 -1900 10736 -1866
rect 10770 -1900 10782 -1866
rect 8764 -1905 10782 -1900
rect 8764 -1906 8822 -1905
rect 10724 -1906 10782 -1905
rect 11365 -1908 11375 -1856
rect 11427 -1908 11437 -1856
rect 13671 -1866 13685 -1832
rect 13719 -1866 13735 -1832
rect 13671 -1910 13735 -1866
rect 15236 -1816 15294 -1810
rect 15328 -1816 15386 -1811
rect 15236 -1850 15248 -1816
rect 15282 -1817 15394 -1816
rect 15282 -1850 15340 -1817
rect 15236 -1851 15340 -1850
rect 15374 -1851 15394 -1817
rect 15236 -1896 15394 -1851
rect 15236 -1912 16946 -1896
rect 15236 -1946 15248 -1912
rect 15282 -1946 15341 -1912
rect 15375 -1936 16946 -1912
rect 15375 -1946 15394 -1936
rect 15236 -1952 15294 -1946
rect 15329 -1952 15387 -1946
rect 12467 -2407 12520 -2375
rect 12467 -2414 12480 -2407
rect 12514 -2414 12520 -2407
rect 418 -2521 428 -2469
rect 480 -2521 490 -2469
rect 1069 -2473 1127 -2472
rect 3029 -2473 3087 -2472
rect 1069 -2478 3087 -2473
rect 1069 -2512 1081 -2478
rect 1115 -2512 3041 -2478
rect 3075 -2512 3087 -2478
rect 1069 -2517 3087 -2512
rect 1069 -2518 1127 -2517
rect 3029 -2518 3087 -2517
rect 3643 -2473 3701 -2472
rect 5603 -2473 5661 -2472
rect 3643 -2478 5661 -2473
rect 3643 -2512 3655 -2478
rect 3689 -2512 5615 -2478
rect 5649 -2512 5661 -2478
rect 3643 -2517 5661 -2512
rect 3643 -2518 3701 -2517
rect 5603 -2518 5661 -2517
rect 6217 -2473 6275 -2472
rect 8177 -2473 8235 -2472
rect 6217 -2478 8235 -2473
rect 6217 -2512 6229 -2478
rect 6263 -2512 8189 -2478
rect 8223 -2512 8235 -2478
rect 6217 -2517 8235 -2512
rect 6217 -2518 6275 -2517
rect 8177 -2518 8235 -2517
rect 8791 -2473 8849 -2472
rect 10751 -2473 10809 -2472
rect 8791 -2478 10809 -2473
rect 8791 -2512 8806 -2478
rect 8840 -2512 10763 -2478
rect 10797 -2512 10809 -2478
rect 11368 -2488 11378 -2436
rect 11430 -2488 11440 -2436
rect 12456 -2466 12466 -2414
rect 12518 -2466 12520 -2414
rect 15236 -2426 15294 -2420
rect 15328 -2426 15386 -2420
rect 13027 -2461 13085 -2460
rect 12467 -2481 12520 -2466
rect 13023 -2466 13738 -2461
rect 12846 -2472 12991 -2471
rect 8791 -2517 10809 -2512
rect 8791 -2518 8849 -2517
rect 10751 -2518 10809 -2517
rect 12467 -2515 12480 -2481
rect 12514 -2515 12520 -2481
rect 12467 -2528 12520 -2515
rect 12548 -2479 12755 -2472
rect 12807 -2477 12993 -2472
rect 12548 -2513 12568 -2479
rect 12602 -2513 12659 -2479
rect 12693 -2513 12755 -2479
rect 12807 -2511 12858 -2477
rect 12892 -2511 12942 -2477
rect 12976 -2511 12993 -2477
rect 12548 -2521 12755 -2513
rect 12745 -2524 12755 -2521
rect 12807 -2521 12993 -2511
rect 13023 -2500 13039 -2466
rect 13073 -2500 13738 -2466
rect 13916 -2485 13926 -2433
rect 13978 -2440 13988 -2433
rect 15236 -2440 15248 -2426
rect 13978 -2460 15248 -2440
rect 15282 -2460 15340 -2426
rect 15374 -2440 15394 -2426
rect 15374 -2460 16946 -2440
rect 13978 -2480 16946 -2460
rect 13978 -2485 13988 -2480
rect 13023 -2510 13738 -2500
rect 12807 -2524 12817 -2521
rect 12456 -2580 12466 -2528
rect 12518 -2580 12520 -2528
rect 12467 -2587 12480 -2580
rect 12514 -2587 12520 -2580
rect 13023 -2543 13685 -2510
rect 13023 -2577 13042 -2543
rect 13076 -2544 13685 -2543
rect 13719 -2544 13738 -2510
rect 13076 -2577 13738 -2544
rect 15236 -2522 15394 -2480
rect 15236 -2556 15248 -2522
rect 15282 -2556 15341 -2522
rect 15375 -2556 15394 -2522
rect 15236 -2562 15294 -2556
rect 15329 -2562 15387 -2556
rect 13023 -2584 13738 -2577
rect 12467 -2612 12520 -2587
rect -1978 -2996 -1968 -2944
rect -1916 -2996 -1906 -2944
rect -1802 -2958 -1792 -2906
rect -1740 -2958 -1730 -2906
rect 1035 -2952 3062 -2946
rect -225 -2981 479 -2979
rect -231 -3033 -221 -2981
rect -169 -2987 479 -2981
rect -169 -3021 429 -2987
rect 463 -3021 479 -2987
rect 1035 -2986 1072 -2952
rect 1106 -2953 3062 -2952
rect 1106 -2986 3016 -2953
rect 1035 -2987 3016 -2986
rect 3050 -2987 3062 -2953
rect 1035 -2993 3062 -2987
rect 3618 -2948 3676 -2947
rect 5578 -2948 5636 -2947
rect 3618 -2953 5636 -2948
rect 3618 -2987 3630 -2953
rect 3664 -2987 5590 -2953
rect 5624 -2987 5636 -2953
rect 3618 -2992 5636 -2987
rect 3618 -2993 3676 -2992
rect 5578 -2993 5636 -2992
rect 6192 -2948 6250 -2947
rect 8152 -2948 8210 -2947
rect 6192 -2953 8210 -2948
rect 6192 -2987 6204 -2953
rect 6238 -2987 8164 -2953
rect 8198 -2987 8210 -2953
rect 6192 -2992 8210 -2987
rect 6192 -2993 6250 -2992
rect 8152 -2993 8210 -2992
rect 8766 -2948 8824 -2947
rect 8766 -2953 10784 -2948
rect 8766 -2987 8778 -2953
rect 8812 -2954 10784 -2953
rect 8812 -2987 10738 -2954
rect 8766 -2988 10738 -2987
rect 10772 -2988 10784 -2954
rect 8766 -2994 10784 -2988
rect 11366 -2995 11376 -2943
rect 11428 -2995 11438 -2943
rect -169 -3033 479 -3021
rect -1968 -3059 -1201 -3058
rect -1968 -3062 -1272 -3059
rect -1978 -3114 -1968 -3062
rect -1916 -3114 -1272 -3062
rect -1968 -3118 -1272 -3114
rect -1213 -3118 -1201 -3059
rect -1968 -3119 -1201 -3118
rect 105 -3573 115 -3521
rect 167 -3523 177 -3521
rect 167 -3531 481 -3523
rect 167 -3565 432 -3531
rect 466 -3565 481 -3531
rect 167 -3572 481 -3565
rect 1033 -3565 3062 -3559
rect 1033 -3568 3016 -3565
rect 167 -3573 177 -3572
rect 1033 -3602 1070 -3568
rect 1104 -3599 3016 -3568
rect 3050 -3599 3062 -3565
rect 1104 -3602 3062 -3599
rect 1033 -3610 3062 -3602
rect 3618 -3560 3676 -3559
rect 5578 -3560 5636 -3559
rect 3618 -3565 5636 -3560
rect 3618 -3599 3630 -3565
rect 3664 -3599 5590 -3565
rect 5624 -3599 5636 -3565
rect 3618 -3604 5636 -3599
rect 3618 -3605 3676 -3604
rect 5578 -3605 5636 -3604
rect 6192 -3560 6250 -3559
rect 8152 -3560 8210 -3559
rect 6192 -3565 8210 -3560
rect 6192 -3599 6204 -3565
rect 6238 -3599 8164 -3565
rect 8198 -3599 8210 -3565
rect 6192 -3604 8210 -3599
rect 6192 -3605 6250 -3604
rect 8152 -3605 8210 -3604
rect 8766 -3565 10783 -3557
rect 8766 -3599 8778 -3565
rect 8812 -3568 10783 -3565
rect 8812 -3599 10735 -3568
rect 8766 -3602 10735 -3599
rect 10769 -3602 10783 -3568
rect 8766 -3607 10783 -3602
rect 10723 -3608 10781 -3607
rect 11363 -3609 11373 -3557
rect 11425 -3609 11435 -3557
rect 12467 -3965 12520 -3940
rect 12467 -3972 12480 -3965
rect 12514 -3972 12520 -3965
rect 12456 -4024 12466 -3972
rect 12518 -4024 12520 -3972
rect 417 -4083 427 -4031
rect 479 -4083 489 -4031
rect 1069 -4035 1127 -4034
rect 3029 -4035 3087 -4034
rect 1069 -4040 3087 -4035
rect 1069 -4074 1081 -4040
rect 1115 -4074 3041 -4040
rect 3075 -4074 3087 -4040
rect 1069 -4079 3087 -4074
rect 1069 -4080 1127 -4079
rect 3029 -4080 3087 -4079
rect 3643 -4035 3701 -4034
rect 5603 -4035 5661 -4034
rect 3643 -4040 5661 -4035
rect 3643 -4074 3655 -4040
rect 3689 -4074 5615 -4040
rect 5649 -4074 5661 -4040
rect 3643 -4079 5661 -4074
rect 3643 -4080 3701 -4079
rect 5603 -4080 5661 -4079
rect 6217 -4035 6275 -4034
rect 8177 -4035 8235 -4034
rect 6217 -4040 8235 -4035
rect 6217 -4074 6229 -4040
rect 6263 -4074 8189 -4040
rect 8223 -4074 8235 -4040
rect 6217 -4079 8235 -4074
rect 6217 -4080 6275 -4079
rect 8177 -4080 8235 -4079
rect 8791 -4035 8849 -4034
rect 10751 -4035 10809 -4034
rect 8791 -4040 10809 -4035
rect 8791 -4074 8806 -4040
rect 8840 -4074 10763 -4040
rect 10797 -4074 10809 -4040
rect 12467 -4037 12520 -4024
rect 13023 -3975 13738 -3968
rect 13023 -4009 13042 -3975
rect 13076 -4008 13738 -3975
rect 13076 -4009 13685 -4008
rect 12745 -4031 12755 -4028
rect 8791 -4079 10809 -4074
rect 8791 -4080 8849 -4079
rect 10751 -4080 10809 -4079
rect 11367 -4119 11377 -4067
rect 11429 -4119 11439 -4067
rect 12467 -4071 12480 -4037
rect 12514 -4071 12520 -4037
rect 12467 -4086 12520 -4071
rect 12548 -4039 12755 -4031
rect 12807 -4031 12817 -4028
rect 12548 -4073 12568 -4039
rect 12602 -4073 12659 -4039
rect 12693 -4073 12755 -4039
rect 12807 -4041 12993 -4031
rect 12548 -4080 12755 -4073
rect 12807 -4075 12858 -4041
rect 12892 -4075 12942 -4041
rect 12976 -4075 12993 -4041
rect 12807 -4080 12993 -4075
rect 13023 -4042 13685 -4009
rect 13719 -4042 13738 -4008
rect 13023 -4052 13738 -4042
rect 12846 -4081 12991 -4080
rect 12456 -4138 12466 -4086
rect 12518 -4138 12520 -4086
rect 13023 -4086 13039 -4052
rect 13073 -4086 13738 -4052
rect 15236 -3996 15294 -3990
rect 15329 -3996 15387 -3990
rect 15236 -4030 15248 -3996
rect 15282 -4030 15341 -3996
rect 15375 -4030 15394 -3996
rect 13023 -4091 13738 -4086
rect 13027 -4092 13085 -4091
rect 14618 -4118 14628 -4064
rect 14682 -4072 14692 -4064
rect 15236 -4072 15394 -4030
rect 14682 -4092 16946 -4072
rect 14682 -4112 15248 -4092
rect 14682 -4118 14692 -4112
rect 15236 -4126 15248 -4112
rect 15282 -4126 15340 -4092
rect 15374 -4112 16946 -4092
rect 15374 -4126 15394 -4112
rect 15236 -4132 15294 -4126
rect 15328 -4132 15386 -4126
rect 12467 -4145 12480 -4138
rect 12514 -4145 12520 -4138
rect 12467 -4177 12520 -4145
rect 15236 -4606 15294 -4600
rect 15329 -4606 15387 -4600
rect -866 -4613 -771 -4608
rect -867 -4619 -771 -4613
rect -867 -4653 -855 -4619
rect -821 -4653 -771 -4619
rect -867 -4659 -771 -4653
rect -866 -4663 -771 -4659
rect -716 -4663 -706 -4608
rect 105 -4647 115 -4643
rect -866 -4666 -706 -4663
rect -253 -4656 115 -4647
rect -253 -4690 -210 -4656
rect -176 -4690 115 -4656
rect -253 -4693 115 -4690
rect -222 -4696 -164 -4693
rect 105 -4695 115 -4693
rect 167 -4695 177 -4643
rect 414 -4662 424 -4610
rect 476 -4662 486 -4610
rect 15236 -4640 15248 -4606
rect 15282 -4640 15341 -4606
rect 15375 -4616 15394 -4606
rect 15375 -4640 16946 -4616
rect 1042 -4647 1100 -4646
rect 3002 -4647 3060 -4646
rect 1042 -4652 3060 -4647
rect 1042 -4686 1054 -4652
rect 1088 -4686 3014 -4652
rect 3048 -4686 3060 -4652
rect 1042 -4691 3060 -4686
rect 1042 -4692 1100 -4691
rect 3002 -4692 3060 -4691
rect 3616 -4647 3674 -4646
rect 5576 -4647 5634 -4646
rect 3616 -4652 5634 -4647
rect 3616 -4686 3628 -4652
rect 3662 -4686 5588 -4652
rect 5622 -4686 5634 -4652
rect 3616 -4691 5634 -4686
rect 3616 -4692 3674 -4691
rect 5576 -4692 5634 -4691
rect 6190 -4647 6248 -4646
rect 8150 -4647 8208 -4646
rect 6190 -4652 8208 -4647
rect 6190 -4686 6202 -4652
rect 6236 -4686 8162 -4652
rect 8196 -4686 8208 -4652
rect 6190 -4691 8208 -4686
rect 6190 -4692 6248 -4691
rect 8150 -4692 8208 -4691
rect 8764 -4647 8822 -4646
rect 10724 -4647 10782 -4646
rect 8764 -4652 10782 -4647
rect 8764 -4686 8776 -4652
rect 8810 -4686 10736 -4652
rect 10770 -4686 10782 -4652
rect 8764 -4691 10782 -4686
rect 8764 -4692 8822 -4691
rect 10724 -4692 10782 -4691
rect 11365 -4697 11375 -4645
rect 11427 -4697 11437 -4645
rect 13671 -4686 13735 -4642
rect 13671 -4720 13685 -4686
rect 13719 -4720 13735 -4686
rect 12746 -4736 12756 -4734
rect 7153 -4737 12756 -4736
rect 7153 -4789 7163 -4737
rect 7215 -4786 12756 -4737
rect 12808 -4736 12818 -4734
rect 13671 -4736 13735 -4720
rect 12808 -4786 13735 -4736
rect 15236 -4656 16946 -4640
rect 15236 -4701 15394 -4656
rect 15236 -4702 15340 -4701
rect 15236 -4736 15248 -4702
rect 15282 -4735 15340 -4702
rect 15374 -4735 15394 -4701
rect 15282 -4736 15394 -4735
rect 15236 -4742 15294 -4736
rect 15328 -4741 15386 -4736
rect 7215 -4789 13735 -4786
rect 7153 -4790 13735 -4789
rect 13671 -4791 13735 -4790
rect 13026 -5061 13084 -5054
rect 13026 -5095 13038 -5061
rect 13072 -5062 13084 -5061
rect 13072 -5095 13737 -5062
rect 13026 -5096 13737 -5095
rect 12548 -5118 12992 -5117
rect 12548 -5120 12752 -5118
rect 417 -5172 427 -5120
rect 479 -5172 489 -5120
rect 1070 -5124 1128 -5123
rect 3030 -5124 3088 -5123
rect 1070 -5129 3088 -5124
rect 1070 -5163 1082 -5129
rect 1116 -5163 3042 -5129
rect 3076 -5163 3088 -5129
rect 1070 -5168 3088 -5163
rect 1070 -5169 1128 -5168
rect 3030 -5169 3088 -5168
rect 3644 -5124 3702 -5123
rect 5604 -5124 5662 -5123
rect 3644 -5129 5662 -5124
rect 3644 -5163 3656 -5129
rect 3690 -5163 5616 -5129
rect 5650 -5163 5662 -5129
rect 3644 -5168 5662 -5163
rect 3644 -5169 3702 -5168
rect 5604 -5169 5662 -5168
rect 6218 -5124 6276 -5123
rect 8178 -5124 8236 -5123
rect 6218 -5129 8236 -5124
rect 6218 -5163 6230 -5129
rect 6264 -5163 8190 -5129
rect 8224 -5163 8236 -5129
rect 6218 -5168 8236 -5163
rect 6218 -5169 6276 -5168
rect 8178 -5169 8236 -5168
rect 8792 -5124 8850 -5123
rect 10752 -5124 10810 -5123
rect 8792 -5129 10810 -5124
rect 8792 -5163 8804 -5129
rect 8838 -5163 10764 -5129
rect 10798 -5163 10810 -5129
rect 12546 -5126 12752 -5120
rect 12804 -5126 12992 -5118
rect 8792 -5168 10810 -5163
rect 8792 -5169 8850 -5168
rect 10752 -5169 10810 -5168
rect 11370 -5204 11380 -5152
rect 11432 -5204 11442 -5152
rect 12546 -5160 12558 -5126
rect 12592 -5160 12642 -5126
rect 12676 -5160 12739 -5126
rect 12804 -5160 12836 -5126
rect 12870 -5160 12942 -5126
rect 12976 -5160 12992 -5126
rect 12546 -5166 12752 -5160
rect 12548 -5170 12752 -5166
rect 12804 -5170 12992 -5160
rect 13026 -5130 13684 -5096
rect 13718 -5130 13737 -5096
rect 13026 -5133 13737 -5130
rect 13026 -5167 13038 -5133
rect 13072 -5167 13737 -5133
rect 13026 -5172 13737 -5167
rect 15236 -5084 15294 -5078
rect 15329 -5084 15387 -5078
rect 15236 -5118 15248 -5084
rect 15282 -5118 15341 -5084
rect 15375 -5118 15394 -5084
rect 15236 -5160 15394 -5118
rect 13026 -5173 13084 -5172
rect 15236 -5179 16946 -5160
rect 15236 -5180 15340 -5179
rect 15236 -5214 15248 -5180
rect 15282 -5213 15340 -5180
rect 15374 -5200 16946 -5179
rect 15374 -5213 15394 -5200
rect 15282 -5214 15394 -5213
rect 15236 -5220 15294 -5214
rect 15328 -5219 15386 -5214
rect 7161 -5265 11181 -5259
rect 7155 -5317 7165 -5265
rect 7217 -5268 11181 -5265
rect 7217 -5317 11118 -5268
rect 7161 -5320 11118 -5317
rect 11170 -5320 11181 -5268
rect 7161 -5321 11181 -5320
rect 11339 -5669 12463 -5665
rect 11338 -5699 12463 -5669
rect 412 -5751 422 -5699
rect 474 -5751 484 -5699
rect 11338 -5724 11586 -5699
rect 12030 -5724 12463 -5699
rect 12522 -5724 12532 -5665
rect 15236 -5694 15294 -5688
rect 15329 -5694 15387 -5688
rect 10725 -5737 10783 -5735
rect 1040 -5738 1098 -5737
rect 3000 -5738 3058 -5737
rect 1040 -5743 3058 -5738
rect 1040 -5777 1052 -5743
rect 1086 -5777 3012 -5743
rect 3046 -5777 3058 -5743
rect 1040 -5782 3058 -5777
rect 1040 -5783 1098 -5782
rect 3000 -5783 3058 -5782
rect 3614 -5738 3672 -5737
rect 5574 -5738 5632 -5737
rect 3614 -5743 5632 -5738
rect 3614 -5777 3626 -5743
rect 3660 -5777 5586 -5743
rect 5620 -5777 5632 -5743
rect 3614 -5782 5632 -5777
rect 3614 -5783 3672 -5782
rect 5574 -5783 5632 -5782
rect 6188 -5738 6246 -5737
rect 8148 -5738 8206 -5737
rect 6188 -5743 8206 -5738
rect 6188 -5777 6200 -5743
rect 6234 -5777 8160 -5743
rect 8194 -5777 8206 -5743
rect 6188 -5782 8206 -5777
rect 6188 -5783 6246 -5782
rect 8148 -5783 8206 -5782
rect 8762 -5738 8820 -5737
rect 10133 -5738 10783 -5737
rect 8762 -5741 10783 -5738
rect 8762 -5743 10737 -5741
rect 8762 -5777 8774 -5743
rect 8808 -5775 10737 -5743
rect 10771 -5775 10783 -5741
rect 8808 -5777 10783 -5775
rect 8762 -5781 10783 -5777
rect 11338 -5740 11430 -5724
rect 15236 -5728 15248 -5694
rect 15282 -5728 15341 -5694
rect 15375 -5704 15394 -5694
rect 15375 -5728 16946 -5704
rect 11338 -5774 11369 -5740
rect 11403 -5774 11430 -5740
rect 11338 -5781 11430 -5774
rect 13669 -5772 13738 -5729
rect 8762 -5782 10231 -5781
rect 8762 -5783 8820 -5782
rect 13669 -5806 13685 -5772
rect 13719 -5806 13738 -5772
rect 13669 -5816 13738 -5806
rect 966 -5818 13738 -5816
rect 966 -5819 12753 -5818
rect 966 -5871 982 -5819
rect 1034 -5870 12753 -5819
rect 12805 -5870 13738 -5818
rect 15236 -5744 16946 -5728
rect 15236 -5789 15394 -5744
rect 15236 -5790 15340 -5789
rect 15236 -5824 15248 -5790
rect 15282 -5823 15340 -5790
rect 15374 -5823 15394 -5789
rect 15282 -5824 15394 -5823
rect 15236 -5830 15294 -5824
rect 15328 -5829 15386 -5824
rect 1034 -5871 13738 -5870
rect 13669 -5873 13738 -5871
rect 1070 -6078 1116 -6074
rect -862 -6106 13 -6100
rect -862 -6140 -848 -6106
rect -814 -6140 -769 -6106
rect -735 -6140 13 -6106
rect -862 -6149 13 -6140
rect 1064 -6133 1122 -6078
rect 418 -6147 485 -6143
rect 1064 -6147 1076 -6133
rect -57 -6205 12 -6149
rect 418 -6167 1076 -6147
rect 1110 -6167 1122 -6133
rect 418 -6173 1122 -6167
rect -57 -6206 16 -6205
rect 94 -6206 152 -6205
rect 227 -6206 389 -6205
rect -954 -6263 -944 -6207
rect -886 -6263 -876 -6207
rect -782 -6263 -772 -6207
rect -714 -6263 -704 -6207
rect -57 -6211 389 -6206
rect -57 -6245 -30 -6211
rect 4 -6245 106 -6211
rect 140 -6245 242 -6211
rect 276 -6245 389 -6211
rect -57 -6254 389 -6245
rect 418 -6207 434 -6173
rect 468 -6175 1122 -6173
rect 468 -6207 982 -6175
rect 418 -6227 982 -6207
rect 1034 -6206 1122 -6175
rect 1034 -6227 1076 -6206
rect 418 -6240 1076 -6227
rect 1110 -6240 1122 -6206
rect 308 -6340 387 -6254
rect 418 -6258 1122 -6240
rect 1153 -6206 1310 -6146
rect 1153 -6212 2449 -6206
rect 1153 -6246 1171 -6212
rect 1205 -6246 1263 -6212
rect 1297 -6217 2449 -6212
rect 1297 -6246 2369 -6217
rect 1153 -6251 2369 -6246
rect 2403 -6251 2449 -6217
rect 1153 -6268 2449 -6251
rect 2994 -6216 6963 -6199
rect 2994 -6250 3015 -6216
rect 3049 -6250 6876 -6216
rect 6910 -6250 6963 -6216
rect 1153 -6269 1310 -6268
rect 2994 -6270 6963 -6250
rect 7509 -6215 8255 -6197
rect 7509 -6216 8164 -6215
rect 7509 -6250 7522 -6216
rect 7556 -6249 8164 -6216
rect 8198 -6249 8255 -6215
rect 7556 -6250 8255 -6249
rect 7509 -6271 8255 -6250
rect 8799 -6217 9545 -6198
rect 8799 -6251 8811 -6217
rect 8845 -6251 9453 -6217
rect 9487 -6251 9545 -6217
rect 8799 -6269 9545 -6251
rect 10086 -6210 11058 -6204
rect 10086 -6216 11063 -6210
rect 10086 -6217 10925 -6216
rect 10086 -6218 10741 -6217
rect 10086 -6252 10099 -6218
rect 10133 -6251 10741 -6218
rect 10775 -6251 10832 -6217
rect 10866 -6250 10925 -6217
rect 10959 -6250 11017 -6216
rect 11051 -6250 11063 -6216
rect 11233 -6219 11418 -6211
rect 10866 -6251 11063 -6250
rect 10133 -6252 11063 -6251
rect 10086 -6256 11063 -6252
rect 10086 -6274 11058 -6256
rect 11110 -6293 11120 -6241
rect 11172 -6293 11182 -6241
rect 11233 -6253 11250 -6219
rect 11284 -6253 11344 -6219
rect 11378 -6253 11418 -6219
rect 11233 -6340 11418 -6253
rect 14617 -6274 14627 -6219
rect 14682 -6226 14692 -6219
rect 15824 -6226 15834 -6219
rect 14682 -6266 15834 -6226
rect 14682 -6274 14692 -6266
rect 15824 -6274 15834 -6266
rect 15889 -6274 15899 -6219
rect -1281 -6409 -1271 -6353
rect -1213 -6356 -1203 -6353
rect -1213 -6409 -768 -6356
rect -715 -6409 -705 -6356
rect -1267 -6410 -705 -6409
rect 308 -6425 11419 -6340
rect -787 -6671 7349 -6670
rect -787 -6727 -772 -6671
rect -714 -6726 7349 -6671
rect 7407 -6726 7417 -6670
rect -714 -6727 7403 -6726
rect -787 -6728 7403 -6727
rect -2617 -6824 -2607 -6821
rect -3193 -6870 -2607 -6824
rect -2617 -6873 -2607 -6870
rect -2554 -6873 -2544 -6821
rect 5018 -6840 5028 -6786
rect 5082 -6840 13925 -6786
rect 13979 -6840 13989 -6786
rect -2356 -6875 -2299 -6868
rect -952 -6875 -894 -6874
rect -2356 -6880 -894 -6875
rect -2356 -6882 -940 -6880
rect -2356 -6916 -2343 -6882
rect -2309 -6914 -940 -6882
rect -906 -6914 -894 -6880
rect -2309 -6916 -894 -6914
rect -2356 -6917 -894 -6916
rect -2356 -6923 -2299 -6917
rect -952 -6920 -894 -6917
rect -1978 -7003 -1968 -6951
rect -1915 -6954 -1908 -6951
rect -1915 -6960 -1183 -6954
rect -415 -6958 -405 -6899
rect -346 -6958 3736 -6899
rect 3795 -6958 3805 -6899
rect -1915 -6994 -1233 -6960
rect -1199 -6994 -1183 -6960
rect 4934 -6977 4945 -6923
rect 4999 -6977 15832 -6923
rect 15886 -6977 15896 -6923
rect -1915 -7000 -1183 -6994
rect -1915 -7003 -1908 -7000
rect 5736 -7180 6293 -7173
rect 3840 -7185 3898 -7182
rect 3099 -7188 3898 -7185
rect 3099 -7191 3852 -7188
rect 3099 -7225 3111 -7191
rect 3145 -7222 3852 -7191
rect 3886 -7222 3898 -7188
rect 3145 -7225 3898 -7222
rect 3099 -7228 3898 -7225
rect 3099 -7230 3872 -7228
rect 3099 -7231 3157 -7230
rect 4935 -7249 4945 -7195
rect 4999 -7249 5009 -7195
rect 5736 -7214 6245 -7180
rect 6279 -7214 6293 -7180
rect 5736 -7220 6293 -7214
rect 2724 -7317 2736 -7258
rect 2795 -7270 2991 -7258
rect 2795 -7304 2934 -7270
rect 2968 -7304 2991 -7270
rect 2795 -7317 2991 -7304
rect 2724 -7318 2991 -7317
rect 3726 -7351 3736 -7292
rect 3795 -7351 3805 -7292
rect 4553 -7299 4611 -7298
rect 3906 -7304 4611 -7299
rect 3906 -7305 4565 -7304
rect 3906 -7339 3928 -7305
rect 3962 -7338 4565 -7305
rect 4599 -7338 4611 -7304
rect 3962 -7339 4611 -7338
rect 3906 -7344 4611 -7339
rect 5028 -7299 5082 -7290
rect 3906 -7348 4599 -7344
rect 5028 -7372 5082 -7353
rect 5736 -7367 5783 -7220
rect 7339 -7310 7349 -7254
rect 7407 -7310 7417 -7254
rect 7582 -7267 16044 -7265
rect 7582 -7290 15971 -7267
rect 5131 -7373 5783 -7367
rect 5131 -7407 5171 -7373
rect 5205 -7407 5783 -7373
rect 5131 -7414 5783 -7407
rect 7582 -7324 7604 -7290
rect 7638 -7324 15971 -7290
rect 7582 -7326 15971 -7324
rect 16030 -7326 16044 -7267
rect 7582 -7330 16044 -7326
rect 7582 -7364 7661 -7330
rect 7582 -7398 7605 -7364
rect 7639 -7398 7661 -7364
rect 7582 -7408 7661 -7398
rect -631 -7498 -620 -7439
rect -561 -7498 2736 -7439
rect 2795 -7498 2805 -7439
rect 308 -7828 11419 -7743
rect -629 -7906 -619 -7902
rect -1978 -7960 -1968 -7908
rect -1915 -7911 -1905 -7908
rect -1915 -7918 -889 -7911
rect -1915 -7952 -937 -7918
rect -903 -7952 -889 -7918
rect -1915 -7958 -889 -7952
rect -781 -7917 -619 -7906
rect -781 -7951 -762 -7917
rect -728 -7951 -619 -7917
rect -781 -7957 -619 -7951
rect -781 -7958 -709 -7957
rect -1915 -7960 -1905 -7958
rect -629 -7961 -619 -7957
rect -560 -7961 -550 -7902
rect 308 -7914 387 -7828
rect 1153 -7900 1310 -7899
rect -57 -7923 389 -7914
rect -57 -7957 -30 -7923
rect 4 -7957 106 -7923
rect 140 -7957 242 -7923
rect 276 -7957 389 -7923
rect -57 -7962 389 -7957
rect -57 -7963 16 -7962
rect 94 -7963 152 -7962
rect 227 -7963 389 -7962
rect 418 -7928 1122 -7910
rect 418 -7941 1076 -7928
rect 418 -7961 982 -7941
rect -57 -8019 12 -7963
rect 418 -7995 434 -7961
rect 468 -7993 982 -7961
rect 1034 -7962 1076 -7941
rect 1110 -7962 1122 -7928
rect 1034 -7993 1122 -7962
rect 468 -7995 1122 -7993
rect 418 -8001 1122 -7995
rect -862 -8028 13 -8019
rect 418 -8021 1076 -8001
rect 418 -8025 485 -8021
rect -862 -8062 -848 -8028
rect -814 -8062 -769 -8028
rect -735 -8062 13 -8028
rect -862 -8068 13 -8062
rect 1064 -8035 1076 -8021
rect 1110 -8035 1122 -8001
rect 1153 -7917 2449 -7900
rect 1153 -7922 2369 -7917
rect 1153 -7956 1171 -7922
rect 1205 -7956 1263 -7922
rect 1297 -7951 2369 -7922
rect 2403 -7951 2449 -7917
rect 1297 -7956 2449 -7951
rect 1153 -7962 2449 -7956
rect 2994 -7918 6963 -7898
rect 2994 -7952 3015 -7918
rect 3049 -7952 6876 -7918
rect 6910 -7952 6963 -7918
rect 1153 -8022 1310 -7962
rect 2994 -7969 6963 -7952
rect 7509 -7918 8255 -7897
rect 7509 -7952 7522 -7918
rect 7556 -7919 8255 -7918
rect 7556 -7952 8164 -7919
rect 7509 -7953 8164 -7952
rect 8198 -7953 8255 -7919
rect 7509 -7971 8255 -7953
rect 8799 -7917 9545 -7899
rect 8799 -7951 8811 -7917
rect 8845 -7951 9453 -7917
rect 9487 -7951 9545 -7917
rect 8799 -7970 9545 -7951
rect 10086 -7912 11058 -7894
rect 10086 -7916 11063 -7912
rect 10086 -7950 10099 -7916
rect 10133 -7917 11063 -7916
rect 10133 -7950 10741 -7917
rect 10086 -7951 10741 -7950
rect 10775 -7951 10832 -7917
rect 10866 -7918 11063 -7917
rect 10866 -7951 10925 -7918
rect 10086 -7952 10925 -7951
rect 10959 -7952 11017 -7918
rect 11051 -7952 11063 -7918
rect 11110 -7927 11120 -7875
rect 11172 -7927 11182 -7875
rect 11233 -7915 11418 -7828
rect 10086 -7958 11063 -7952
rect 11233 -7949 11250 -7915
rect 11284 -7949 11344 -7915
rect 11378 -7949 11418 -7915
rect 11233 -7957 11418 -7949
rect 10086 -7964 11058 -7958
rect 1064 -8090 1122 -8035
rect 1070 -8094 1116 -8090
rect 16662 -8220 16946 -8124
rect 13669 -8297 13738 -8295
rect 966 -8349 982 -8297
rect 1034 -8298 13738 -8297
rect 1034 -8349 12753 -8298
rect 966 -8350 12753 -8349
rect 12805 -8350 13738 -8298
rect 966 -8352 13738 -8350
rect 13669 -8362 13738 -8352
rect 1040 -8386 1098 -8385
rect 3000 -8386 3058 -8385
rect 1040 -8391 3058 -8386
rect 413 -8470 423 -8418
rect 475 -8470 485 -8418
rect 1040 -8425 1052 -8391
rect 1086 -8425 3012 -8391
rect 3046 -8425 3058 -8391
rect 1040 -8430 3058 -8425
rect 1040 -8431 1098 -8430
rect 3000 -8431 3058 -8430
rect 3614 -8386 3672 -8385
rect 5574 -8386 5632 -8385
rect 3614 -8391 5632 -8386
rect 3614 -8425 3626 -8391
rect 3660 -8425 5586 -8391
rect 5620 -8425 5632 -8391
rect 3614 -8430 5632 -8425
rect 3614 -8431 3672 -8430
rect 5574 -8431 5632 -8430
rect 6188 -8386 6246 -8385
rect 8148 -8386 8206 -8385
rect 6188 -8391 8206 -8386
rect 6188 -8425 6200 -8391
rect 6234 -8425 8160 -8391
rect 8194 -8425 8206 -8391
rect 6188 -8430 8206 -8425
rect 6188 -8431 6246 -8430
rect 8148 -8431 8206 -8430
rect 8762 -8386 8820 -8385
rect 8762 -8387 10320 -8386
rect 8762 -8391 10783 -8387
rect 8762 -8425 8774 -8391
rect 8808 -8393 10783 -8391
rect 8808 -8425 10737 -8393
rect 8762 -8427 10737 -8425
rect 10771 -8427 10783 -8393
rect 8762 -8430 10783 -8427
rect 8762 -8431 8820 -8430
rect 10131 -8431 10783 -8430
rect 10725 -8433 10783 -8431
rect 11338 -8394 11430 -8387
rect 11338 -8428 11369 -8394
rect 11403 -8428 11430 -8394
rect 11338 -8444 11430 -8428
rect 13669 -8396 13685 -8362
rect 13719 -8396 13738 -8362
rect 13669 -8439 13738 -8396
rect 15236 -8344 15294 -8338
rect 15328 -8344 15386 -8339
rect 15236 -8378 15248 -8344
rect 15282 -8345 15394 -8344
rect 15282 -8378 15340 -8345
rect 15236 -8379 15340 -8378
rect 15374 -8379 15394 -8345
rect 15236 -8424 15394 -8379
rect 15962 -8424 15972 -8416
rect 15236 -8440 15972 -8424
rect 11338 -8499 12463 -8444
rect 11339 -8503 12463 -8499
rect 12522 -8503 12532 -8444
rect 15236 -8474 15248 -8440
rect 15282 -8474 15341 -8440
rect 15375 -8464 15972 -8440
rect 15375 -8474 15394 -8464
rect 15236 -8480 15294 -8474
rect 15329 -8480 15387 -8474
rect 15962 -8475 15972 -8464
rect 16031 -8424 16041 -8416
rect 16031 -8464 16946 -8424
rect 16031 -8475 16041 -8464
rect 7161 -8848 11181 -8847
rect 7161 -8851 11118 -8848
rect 7155 -8903 7165 -8851
rect 7217 -8900 11118 -8851
rect 11170 -8900 11181 -8848
rect 7217 -8903 11181 -8900
rect 7161 -8909 11181 -8903
rect 15236 -8954 15294 -8948
rect 15328 -8954 15386 -8949
rect 413 -9051 423 -8999
rect 475 -9051 485 -8999
rect 1070 -9000 1128 -8999
rect 3030 -9000 3088 -8999
rect 1070 -9005 3088 -9000
rect 1070 -9039 1082 -9005
rect 1116 -9039 3042 -9005
rect 3076 -9039 3088 -9005
rect 1070 -9044 3088 -9039
rect 1070 -9045 1128 -9044
rect 3030 -9045 3088 -9044
rect 3644 -9000 3702 -8999
rect 5604 -9000 5662 -8999
rect 3644 -9005 5662 -9000
rect 3644 -9039 3656 -9005
rect 3690 -9039 5616 -9005
rect 5650 -9039 5662 -9005
rect 3644 -9044 5662 -9039
rect 3644 -9045 3702 -9044
rect 5604 -9045 5662 -9044
rect 6218 -9000 6276 -8999
rect 8178 -9000 8236 -8999
rect 6218 -9005 8236 -9000
rect 6218 -9039 6230 -9005
rect 6264 -9039 8190 -9005
rect 8224 -9039 8236 -9005
rect 6218 -9044 8236 -9039
rect 6218 -9045 6276 -9044
rect 8178 -9045 8236 -9044
rect 8792 -9000 8850 -8999
rect 10752 -9000 10810 -8999
rect 8792 -9005 10810 -9000
rect 8792 -9039 8804 -9005
rect 8838 -9039 10764 -9005
rect 10798 -9039 10810 -9005
rect 11368 -9013 11378 -8961
rect 11430 -9013 11440 -8961
rect 15236 -8988 15248 -8954
rect 15282 -8955 15394 -8954
rect 15282 -8988 15340 -8955
rect 15236 -8989 15340 -8988
rect 15374 -8968 15394 -8955
rect 15374 -8989 16946 -8968
rect 13026 -8996 13084 -8995
rect 12548 -9002 12752 -8998
rect 12546 -9008 12752 -9002
rect 12804 -9008 12992 -8998
rect 8792 -9044 10810 -9039
rect 8792 -9045 8850 -9044
rect 10752 -9045 10810 -9044
rect 12546 -9042 12558 -9008
rect 12592 -9042 12642 -9008
rect 12676 -9042 12739 -9008
rect 12804 -9042 12836 -9008
rect 12870 -9042 12942 -9008
rect 12976 -9042 12992 -9008
rect 12546 -9048 12752 -9042
rect 12548 -9050 12752 -9048
rect 12804 -9050 12992 -9042
rect 12548 -9051 12992 -9050
rect 13026 -9001 13737 -8996
rect 13026 -9035 13038 -9001
rect 13072 -9035 13737 -9001
rect 13026 -9038 13737 -9035
rect 13026 -9072 13684 -9038
rect 13718 -9072 13737 -9038
rect 13026 -9073 13737 -9072
rect 13026 -9107 13038 -9073
rect 13072 -9106 13737 -9073
rect 15236 -9008 16946 -8989
rect 15236 -9050 15394 -9008
rect 15236 -9084 15248 -9050
rect 15282 -9084 15341 -9050
rect 15375 -9084 15394 -9050
rect 15236 -9090 15294 -9084
rect 15329 -9090 15387 -9084
rect 13072 -9107 13084 -9106
rect 13026 -9114 13084 -9107
rect 13671 -9378 13735 -9377
rect 7153 -9379 13735 -9378
rect 7153 -9431 7163 -9379
rect 7215 -9382 13735 -9379
rect 7215 -9431 12756 -9382
rect 7153 -9432 12756 -9431
rect 12746 -9434 12756 -9432
rect 12808 -9432 13735 -9382
rect 12808 -9434 12818 -9432
rect 13671 -9448 13735 -9432
rect -952 -9559 -942 -9507
rect -890 -9509 -880 -9507
rect -890 -9516 -809 -9509
rect -890 -9550 -856 -9516
rect -822 -9550 -809 -9516
rect -227 -9522 -217 -9470
rect -165 -9522 -155 -9470
rect 1042 -9477 1100 -9476
rect 3002 -9477 3060 -9476
rect 1042 -9482 3060 -9477
rect -890 -9557 -809 -9550
rect -890 -9559 -880 -9557
rect 413 -9558 423 -9506
rect 475 -9558 485 -9506
rect 1042 -9516 1054 -9482
rect 1088 -9516 3014 -9482
rect 3048 -9516 3060 -9482
rect 1042 -9521 3060 -9516
rect 1042 -9522 1100 -9521
rect 3002 -9522 3060 -9521
rect 3616 -9477 3674 -9476
rect 5576 -9477 5634 -9476
rect 3616 -9482 5634 -9477
rect 3616 -9516 3628 -9482
rect 3662 -9516 5588 -9482
rect 5622 -9516 5634 -9482
rect 3616 -9521 5634 -9516
rect 3616 -9522 3674 -9521
rect 5576 -9522 5634 -9521
rect 6190 -9477 6248 -9476
rect 8150 -9477 8208 -9476
rect 6190 -9482 8208 -9477
rect 6190 -9516 6202 -9482
rect 6236 -9516 8162 -9482
rect 8196 -9516 8208 -9482
rect 6190 -9521 8208 -9516
rect 6190 -9522 6248 -9521
rect 8150 -9522 8208 -9521
rect 8764 -9477 8822 -9476
rect 10724 -9477 10782 -9476
rect 8764 -9482 10782 -9477
rect 8764 -9516 8776 -9482
rect 8810 -9516 10736 -9482
rect 10770 -9516 10782 -9482
rect 8764 -9521 10782 -9516
rect 8764 -9522 8822 -9521
rect 10724 -9522 10782 -9521
rect 11365 -9524 11375 -9472
rect 11427 -9524 11437 -9472
rect 13671 -9482 13685 -9448
rect 13719 -9482 13735 -9448
rect 13671 -9526 13735 -9482
rect 15236 -9432 15294 -9426
rect 15328 -9432 15386 -9427
rect 15236 -9466 15248 -9432
rect 15282 -9433 15394 -9432
rect 15282 -9466 15340 -9433
rect 15236 -9467 15340 -9466
rect 15374 -9467 15394 -9433
rect 15236 -9512 15394 -9467
rect 15236 -9528 16946 -9512
rect 15236 -9562 15248 -9528
rect 15282 -9562 15341 -9528
rect 15375 -9552 16946 -9528
rect 15375 -9562 15394 -9552
rect 15236 -9568 15294 -9562
rect 15329 -9568 15387 -9562
rect 12467 -10023 12520 -9991
rect 12467 -10030 12480 -10023
rect 12514 -10030 12520 -10023
rect 418 -10137 428 -10085
rect 480 -10137 490 -10085
rect 1069 -10089 1127 -10088
rect 3029 -10089 3087 -10088
rect 1069 -10094 3087 -10089
rect 1069 -10128 1081 -10094
rect 1115 -10128 3041 -10094
rect 3075 -10128 3087 -10094
rect 1069 -10133 3087 -10128
rect 1069 -10134 1127 -10133
rect 3029 -10134 3087 -10133
rect 3643 -10089 3701 -10088
rect 5603 -10089 5661 -10088
rect 3643 -10094 5661 -10089
rect 3643 -10128 3655 -10094
rect 3689 -10128 5615 -10094
rect 5649 -10128 5661 -10094
rect 3643 -10133 5661 -10128
rect 3643 -10134 3701 -10133
rect 5603 -10134 5661 -10133
rect 6217 -10089 6275 -10088
rect 8177 -10089 8235 -10088
rect 6217 -10094 8235 -10089
rect 6217 -10128 6229 -10094
rect 6263 -10128 8189 -10094
rect 8223 -10128 8235 -10094
rect 6217 -10133 8235 -10128
rect 6217 -10134 6275 -10133
rect 8177 -10134 8235 -10133
rect 8791 -10089 8849 -10088
rect 10751 -10089 10809 -10088
rect 8791 -10094 10809 -10089
rect 8791 -10128 8806 -10094
rect 8840 -10128 10763 -10094
rect 10797 -10128 10809 -10094
rect 11368 -10104 11378 -10052
rect 11430 -10104 11440 -10052
rect 12456 -10082 12466 -10030
rect 12518 -10082 12520 -10030
rect 15236 -10042 15294 -10036
rect 15328 -10042 15386 -10036
rect 15236 -10076 15248 -10042
rect 15282 -10076 15340 -10042
rect 15374 -10056 15394 -10042
rect 15374 -10076 16946 -10056
rect 13027 -10077 13085 -10076
rect 12467 -10097 12520 -10082
rect 13023 -10082 13738 -10077
rect 12846 -10088 12991 -10087
rect 8791 -10133 10809 -10128
rect 8791 -10134 8849 -10133
rect 10751 -10134 10809 -10133
rect 12467 -10131 12480 -10097
rect 12514 -10131 12520 -10097
rect 12467 -10144 12520 -10131
rect 12548 -10095 12755 -10088
rect 12807 -10093 12993 -10088
rect 12548 -10129 12568 -10095
rect 12602 -10129 12659 -10095
rect 12693 -10129 12755 -10095
rect 12807 -10127 12858 -10093
rect 12892 -10127 12942 -10093
rect 12976 -10127 12993 -10093
rect 12548 -10137 12755 -10129
rect 12745 -10140 12755 -10137
rect 12807 -10137 12993 -10127
rect 13023 -10116 13039 -10082
rect 13073 -10116 13738 -10082
rect 13023 -10126 13738 -10116
rect 12807 -10140 12817 -10137
rect 12456 -10196 12466 -10144
rect 12518 -10196 12520 -10144
rect 12467 -10203 12480 -10196
rect 12514 -10203 12520 -10196
rect 13023 -10159 13685 -10126
rect 13023 -10193 13042 -10159
rect 13076 -10160 13685 -10159
rect 13719 -10160 13738 -10126
rect 13076 -10193 13738 -10160
rect 15236 -10096 16946 -10076
rect 15236 -10138 15394 -10096
rect 15236 -10172 15248 -10138
rect 15282 -10172 15341 -10138
rect 15375 -10172 15394 -10138
rect 15236 -10178 15294 -10172
rect 15329 -10178 15387 -10172
rect 13023 -10200 13738 -10193
rect 12467 -10228 12520 -10203
rect -2617 -10490 -1969 -10489
rect -2617 -10543 -2607 -10490
rect -2554 -10543 -1969 -10490
rect -1915 -10543 -1905 -10489
rect -1833 -10579 -1823 -10525
rect -1769 -10579 -1759 -10525
rect 1035 -10564 2469 -10562
rect 3004 -10564 3062 -10563
rect 1035 -10568 3062 -10564
rect -225 -10597 479 -10595
rect -231 -10649 -221 -10597
rect -169 -10603 479 -10597
rect -169 -10637 429 -10603
rect 463 -10637 479 -10603
rect 1035 -10602 1072 -10568
rect 1106 -10569 3062 -10568
rect 1106 -10602 3016 -10569
rect 1035 -10603 3016 -10602
rect 3050 -10603 3062 -10569
rect 1035 -10608 3062 -10603
rect 1035 -10609 2469 -10608
rect 3004 -10609 3062 -10608
rect 3618 -10564 3676 -10563
rect 5578 -10564 5636 -10563
rect 3618 -10569 5636 -10564
rect 3618 -10603 3630 -10569
rect 3664 -10603 5590 -10569
rect 5624 -10603 5636 -10569
rect 3618 -10608 5636 -10603
rect 3618 -10609 3676 -10608
rect 5578 -10609 5636 -10608
rect 6192 -10564 6250 -10563
rect 8152 -10564 8210 -10563
rect 6192 -10569 8210 -10564
rect 6192 -10603 6204 -10569
rect 6238 -10603 8164 -10569
rect 8198 -10603 8210 -10569
rect 6192 -10608 8210 -10603
rect 6192 -10609 6250 -10608
rect 8152 -10609 8210 -10608
rect 8766 -10564 8824 -10563
rect 10145 -10564 10783 -10562
rect 8766 -10569 10784 -10564
rect 8766 -10603 8778 -10569
rect 8812 -10570 10784 -10569
rect 8812 -10603 10738 -10570
rect 8766 -10604 10738 -10603
rect 10772 -10604 10784 -10570
rect 8766 -10608 10784 -10604
rect 8766 -10609 8824 -10608
rect 10145 -10610 10784 -10608
rect 10145 -10614 10783 -10610
rect 11366 -10611 11376 -10559
rect 11428 -10611 11438 -10559
rect -169 -10649 479 -10637
rect 105 -11189 115 -11137
rect 167 -11139 177 -11137
rect 167 -11147 481 -11139
rect 167 -11181 432 -11147
rect 466 -11181 481 -11147
rect 3004 -11176 3062 -11175
rect 2409 -11177 3062 -11176
rect 167 -11188 481 -11181
rect 1033 -11181 3062 -11177
rect 1033 -11184 3016 -11181
rect 167 -11189 177 -11188
rect 1033 -11218 1070 -11184
rect 1104 -11215 3016 -11184
rect 3050 -11215 3062 -11181
rect 1104 -11218 3062 -11215
rect 1033 -11220 3062 -11218
rect 1033 -11226 2499 -11220
rect 3004 -11221 3062 -11220
rect 3618 -11176 3676 -11175
rect 5578 -11176 5636 -11175
rect 3618 -11181 5636 -11176
rect 3618 -11215 3630 -11181
rect 3664 -11215 5590 -11181
rect 5624 -11215 5636 -11181
rect 3618 -11220 5636 -11215
rect 3618 -11221 3676 -11220
rect 5578 -11221 5636 -11220
rect 6192 -11176 6250 -11175
rect 8152 -11176 8210 -11175
rect 6192 -11181 8210 -11176
rect 6192 -11215 6204 -11181
rect 6238 -11215 8164 -11181
rect 8198 -11215 8210 -11181
rect 6192 -11220 8210 -11215
rect 6192 -11221 6250 -11220
rect 8152 -11221 8210 -11220
rect 8766 -11176 8824 -11175
rect 10147 -11176 10783 -11173
rect 8766 -11181 10783 -11176
rect 8766 -11215 8778 -11181
rect 8812 -11184 10783 -11181
rect 8812 -11215 10735 -11184
rect 8766 -11218 10735 -11215
rect 10769 -11218 10783 -11184
rect 8766 -11220 10783 -11218
rect 8766 -11221 8824 -11220
rect 10147 -11223 10783 -11220
rect 10723 -11224 10781 -11223
rect 11363 -11225 11373 -11173
rect 11425 -11225 11435 -11173
rect 12467 -11581 12520 -11556
rect 12467 -11588 12480 -11581
rect 12514 -11588 12520 -11581
rect 12456 -11640 12466 -11588
rect 12518 -11640 12520 -11588
rect 417 -11699 427 -11647
rect 479 -11699 489 -11647
rect 1069 -11651 1127 -11650
rect 3029 -11651 3087 -11650
rect 1069 -11656 3087 -11651
rect 1069 -11690 1081 -11656
rect 1115 -11690 3041 -11656
rect 3075 -11690 3087 -11656
rect 1069 -11695 3087 -11690
rect 1069 -11696 1127 -11695
rect 3029 -11696 3087 -11695
rect 3643 -11651 3701 -11650
rect 5603 -11651 5661 -11650
rect 3643 -11656 5661 -11651
rect 3643 -11690 3655 -11656
rect 3689 -11690 5615 -11656
rect 5649 -11690 5661 -11656
rect 3643 -11695 5661 -11690
rect 3643 -11696 3701 -11695
rect 5603 -11696 5661 -11695
rect 6217 -11651 6275 -11650
rect 8177 -11651 8235 -11650
rect 6217 -11656 8235 -11651
rect 6217 -11690 6229 -11656
rect 6263 -11690 8189 -11656
rect 8223 -11690 8235 -11656
rect 6217 -11695 8235 -11690
rect 6217 -11696 6275 -11695
rect 8177 -11696 8235 -11695
rect 8791 -11651 8849 -11650
rect 10751 -11651 10809 -11650
rect 8791 -11656 10809 -11651
rect 8791 -11690 8806 -11656
rect 8840 -11690 10763 -11656
rect 10797 -11690 10809 -11656
rect 12467 -11653 12520 -11640
rect 13023 -11591 13738 -11584
rect 13023 -11625 13042 -11591
rect 13076 -11624 13738 -11591
rect 13076 -11625 13685 -11624
rect 12745 -11647 12755 -11644
rect 8791 -11695 10809 -11690
rect 8791 -11696 8849 -11695
rect 10751 -11696 10809 -11695
rect 11367 -11735 11377 -11683
rect 11429 -11735 11439 -11683
rect 12467 -11687 12480 -11653
rect 12514 -11687 12520 -11653
rect 12467 -11702 12520 -11687
rect 12548 -11655 12755 -11647
rect 12807 -11647 12817 -11644
rect 12548 -11689 12568 -11655
rect 12602 -11689 12659 -11655
rect 12693 -11689 12755 -11655
rect 12807 -11657 12993 -11647
rect 12548 -11696 12755 -11689
rect 12807 -11691 12858 -11657
rect 12892 -11691 12942 -11657
rect 12976 -11691 12993 -11657
rect 12807 -11696 12993 -11691
rect 13023 -11658 13685 -11625
rect 13719 -11658 13738 -11624
rect 13023 -11668 13738 -11658
rect 12846 -11697 12991 -11696
rect 12456 -11754 12466 -11702
rect 12518 -11754 12520 -11702
rect 13023 -11702 13039 -11668
rect 13073 -11702 13738 -11668
rect 13023 -11707 13738 -11702
rect 15236 -11612 15294 -11606
rect 15329 -11612 15387 -11606
rect 15236 -11646 15248 -11612
rect 15282 -11646 15341 -11612
rect 15375 -11646 15394 -11612
rect 15236 -11688 15394 -11646
rect 13027 -11708 13085 -11707
rect 15236 -11708 16946 -11688
rect 15236 -11742 15248 -11708
rect 15282 -11742 15340 -11708
rect 15374 -11728 16946 -11708
rect 15374 -11742 15394 -11728
rect 15236 -11748 15294 -11742
rect 15328 -11748 15386 -11742
rect 12467 -11761 12480 -11754
rect 12514 -11761 12520 -11754
rect 12467 -11793 12520 -11761
rect 15236 -12222 15294 -12216
rect 15329 -12222 15387 -12216
rect -866 -12229 -404 -12224
rect -867 -12235 -404 -12229
rect -867 -12269 -855 -12235
rect -821 -12269 -404 -12235
rect -867 -12275 -404 -12269
rect -866 -12282 -404 -12275
rect -346 -12282 -336 -12224
rect 105 -12263 115 -12259
rect -253 -12272 115 -12263
rect -253 -12306 -210 -12272
rect -176 -12306 115 -12272
rect -253 -12309 115 -12306
rect -222 -12312 -164 -12309
rect 105 -12311 115 -12309
rect 167 -12311 177 -12259
rect 414 -12278 424 -12226
rect 476 -12278 486 -12226
rect 15236 -12256 15248 -12222
rect 15282 -12256 15341 -12222
rect 15375 -12232 15394 -12222
rect 15375 -12256 16946 -12232
rect 1042 -12263 1100 -12262
rect 3002 -12263 3060 -12262
rect 1042 -12268 3060 -12263
rect 1042 -12302 1054 -12268
rect 1088 -12302 3014 -12268
rect 3048 -12302 3060 -12268
rect 1042 -12307 3060 -12302
rect 1042 -12308 1100 -12307
rect 3002 -12308 3060 -12307
rect 3616 -12263 3674 -12262
rect 5576 -12263 5634 -12262
rect 3616 -12268 5634 -12263
rect 3616 -12302 3628 -12268
rect 3662 -12302 5588 -12268
rect 5622 -12302 5634 -12268
rect 3616 -12307 5634 -12302
rect 3616 -12308 3674 -12307
rect 5576 -12308 5634 -12307
rect 6190 -12263 6248 -12262
rect 8150 -12263 8208 -12262
rect 6190 -12268 8208 -12263
rect 6190 -12302 6202 -12268
rect 6236 -12302 8162 -12268
rect 8196 -12302 8208 -12268
rect 6190 -12307 8208 -12302
rect 6190 -12308 6248 -12307
rect 8150 -12308 8208 -12307
rect 8764 -12263 8822 -12262
rect 10724 -12263 10782 -12262
rect 8764 -12268 10782 -12263
rect 8764 -12302 8776 -12268
rect 8810 -12302 10736 -12268
rect 10770 -12302 10782 -12268
rect 8764 -12307 10782 -12302
rect 8764 -12308 8822 -12307
rect 10724 -12308 10782 -12307
rect 11365 -12313 11375 -12261
rect 11427 -12313 11437 -12261
rect 13671 -12302 13735 -12258
rect 13671 -12336 13685 -12302
rect 13719 -12336 13735 -12302
rect 12746 -12352 12756 -12350
rect 7153 -12353 12756 -12352
rect 7153 -12405 7163 -12353
rect 7215 -12402 12756 -12353
rect 12808 -12352 12818 -12350
rect 13671 -12352 13735 -12336
rect 12808 -12402 13735 -12352
rect 15236 -12272 16946 -12256
rect 15236 -12317 15394 -12272
rect 15236 -12318 15340 -12317
rect 15236 -12352 15248 -12318
rect 15282 -12351 15340 -12318
rect 15374 -12351 15394 -12317
rect 15282 -12352 15394 -12351
rect 15236 -12358 15294 -12352
rect 15328 -12357 15386 -12352
rect 7215 -12405 13735 -12402
rect 7153 -12406 13735 -12405
rect 13671 -12407 13735 -12406
rect 13026 -12677 13084 -12670
rect 13026 -12711 13038 -12677
rect 13072 -12678 13084 -12677
rect 13072 -12711 13737 -12678
rect 13026 -12712 13737 -12711
rect 12548 -12734 12992 -12733
rect 12548 -12736 12752 -12734
rect 417 -12788 427 -12736
rect 479 -12788 489 -12736
rect 1070 -12740 1128 -12739
rect 3030 -12740 3088 -12739
rect 1070 -12745 3088 -12740
rect 1070 -12779 1082 -12745
rect 1116 -12779 3042 -12745
rect 3076 -12779 3088 -12745
rect 1070 -12784 3088 -12779
rect 1070 -12785 1128 -12784
rect 3030 -12785 3088 -12784
rect 3644 -12740 3702 -12739
rect 5604 -12740 5662 -12739
rect 3644 -12745 5662 -12740
rect 3644 -12779 3656 -12745
rect 3690 -12779 5616 -12745
rect 5650 -12779 5662 -12745
rect 3644 -12784 5662 -12779
rect 3644 -12785 3702 -12784
rect 5604 -12785 5662 -12784
rect 6218 -12740 6276 -12739
rect 8178 -12740 8236 -12739
rect 6218 -12745 8236 -12740
rect 6218 -12779 6230 -12745
rect 6264 -12779 8190 -12745
rect 8224 -12779 8236 -12745
rect 6218 -12784 8236 -12779
rect 6218 -12785 6276 -12784
rect 8178 -12785 8236 -12784
rect 8792 -12740 8850 -12739
rect 10752 -12740 10810 -12739
rect 8792 -12745 10810 -12740
rect 8792 -12779 8804 -12745
rect 8838 -12779 10764 -12745
rect 10798 -12779 10810 -12745
rect 12546 -12742 12752 -12736
rect 12804 -12742 12992 -12734
rect 8792 -12784 10810 -12779
rect 8792 -12785 8850 -12784
rect 10752 -12785 10810 -12784
rect 11370 -12820 11380 -12768
rect 11432 -12820 11442 -12768
rect 12546 -12776 12558 -12742
rect 12592 -12776 12642 -12742
rect 12676 -12776 12739 -12742
rect 12804 -12776 12836 -12742
rect 12870 -12776 12942 -12742
rect 12976 -12776 12992 -12742
rect 12546 -12782 12752 -12776
rect 12548 -12786 12752 -12782
rect 12804 -12786 12992 -12776
rect 13026 -12746 13684 -12712
rect 13718 -12746 13737 -12712
rect 13026 -12749 13737 -12746
rect 13026 -12783 13038 -12749
rect 13072 -12783 13737 -12749
rect 13026 -12788 13737 -12783
rect 15236 -12700 15294 -12694
rect 15329 -12700 15387 -12694
rect 15236 -12734 15248 -12700
rect 15282 -12734 15341 -12700
rect 15375 -12734 15394 -12700
rect 15236 -12776 15394 -12734
rect 13026 -12789 13084 -12788
rect 15236 -12795 16946 -12776
rect 15236 -12796 15340 -12795
rect 15236 -12830 15248 -12796
rect 15282 -12829 15340 -12796
rect 15374 -12816 16946 -12795
rect 15374 -12829 15394 -12816
rect 15282 -12830 15394 -12829
rect 15236 -12836 15294 -12830
rect 15328 -12835 15386 -12830
rect 7161 -12881 11181 -12875
rect 7155 -12933 7165 -12881
rect 7217 -12884 11181 -12881
rect 7217 -12933 11118 -12884
rect 7161 -12936 11118 -12933
rect 11170 -12936 11181 -12884
rect 7161 -12937 11181 -12936
rect 11339 -13285 12463 -13281
rect 412 -13367 422 -13315
rect 474 -13367 484 -13315
rect 11338 -13340 12463 -13285
rect 12522 -13340 12532 -13281
rect 15236 -13310 15294 -13304
rect 15329 -13310 15387 -13304
rect 10725 -13353 10783 -13351
rect 1040 -13354 1098 -13353
rect 3000 -13354 3058 -13353
rect 1040 -13359 3058 -13354
rect 1040 -13393 1052 -13359
rect 1086 -13393 3012 -13359
rect 3046 -13393 3058 -13359
rect 1040 -13398 3058 -13393
rect 1040 -13399 1098 -13398
rect 3000 -13399 3058 -13398
rect 3614 -13354 3672 -13353
rect 5574 -13354 5632 -13353
rect 3614 -13359 5632 -13354
rect 3614 -13393 3626 -13359
rect 3660 -13393 5586 -13359
rect 5620 -13393 5632 -13359
rect 3614 -13398 5632 -13393
rect 3614 -13399 3672 -13398
rect 5574 -13399 5632 -13398
rect 6188 -13354 6246 -13353
rect 8148 -13354 8206 -13353
rect 6188 -13359 8206 -13354
rect 6188 -13393 6200 -13359
rect 6234 -13393 8160 -13359
rect 8194 -13393 8206 -13359
rect 6188 -13398 8206 -13393
rect 6188 -13399 6246 -13398
rect 8148 -13399 8206 -13398
rect 8762 -13354 8820 -13353
rect 10139 -13354 10783 -13353
rect 8762 -13357 10783 -13354
rect 8762 -13359 10737 -13357
rect 8762 -13393 8774 -13359
rect 8808 -13391 10737 -13359
rect 10771 -13391 10783 -13357
rect 8808 -13393 10783 -13391
rect 8762 -13397 10783 -13393
rect 11338 -13356 11430 -13340
rect 15236 -13344 15248 -13310
rect 15282 -13344 15341 -13310
rect 15375 -13320 15394 -13310
rect 15375 -13344 16946 -13320
rect 11338 -13390 11369 -13356
rect 11403 -13390 11430 -13356
rect 11338 -13397 11430 -13390
rect 13669 -13388 13738 -13345
rect 8762 -13398 10273 -13397
rect 8762 -13399 8820 -13398
rect 13669 -13422 13685 -13388
rect 13719 -13422 13738 -13388
rect 13669 -13432 13738 -13422
rect 966 -13434 13738 -13432
rect 966 -13435 12753 -13434
rect 966 -13487 982 -13435
rect 1034 -13486 12753 -13435
rect 12805 -13486 13738 -13434
rect 15236 -13360 16946 -13344
rect 15236 -13405 15394 -13360
rect 15236 -13406 15340 -13405
rect 15236 -13440 15248 -13406
rect 15282 -13439 15340 -13406
rect 15374 -13439 15394 -13405
rect 15282 -13440 15394 -13439
rect 15236 -13446 15294 -13440
rect 15328 -13445 15386 -13440
rect 1034 -13487 13738 -13486
rect 13669 -13489 13738 -13487
rect 1070 -13694 1116 -13690
rect -862 -13722 13 -13716
rect -862 -13756 -848 -13722
rect -814 -13756 -769 -13722
rect -735 -13756 13 -13722
rect -862 -13765 13 -13756
rect 1064 -13749 1122 -13694
rect 418 -13763 485 -13759
rect 1064 -13763 1076 -13749
rect -57 -13821 12 -13765
rect 418 -13783 1076 -13763
rect 1110 -13783 1122 -13749
rect 418 -13789 1122 -13783
rect -57 -13822 16 -13821
rect 94 -13822 152 -13821
rect 227 -13822 389 -13821
rect -954 -13879 -944 -13823
rect -886 -13879 -876 -13823
rect -778 -13829 -723 -13826
rect -57 -13827 389 -13822
rect -778 -13835 -718 -13829
rect -778 -13869 -764 -13835
rect -730 -13869 -718 -13835
rect -778 -13875 -718 -13869
rect -57 -13861 -30 -13827
rect 4 -13861 106 -13827
rect 140 -13861 242 -13827
rect 276 -13861 389 -13827
rect -57 -13870 389 -13861
rect 418 -13823 434 -13789
rect 468 -13791 1122 -13789
rect 468 -13823 982 -13791
rect 418 -13843 982 -13823
rect 1034 -13822 1122 -13791
rect 1034 -13843 1076 -13822
rect 418 -13856 1076 -13843
rect 1110 -13856 1122 -13822
rect -778 -13916 -723 -13875
rect -1834 -13971 -1824 -13916
rect -1769 -13971 -723 -13916
rect 308 -13956 387 -13870
rect 418 -13874 1122 -13856
rect 1153 -13822 1310 -13762
rect 1153 -13828 2449 -13822
rect 1153 -13862 1171 -13828
rect 1205 -13862 1263 -13828
rect 1297 -13833 2449 -13828
rect 1297 -13862 2369 -13833
rect 1153 -13867 2369 -13862
rect 2403 -13867 2449 -13833
rect 1153 -13884 2449 -13867
rect 2994 -13832 6963 -13815
rect 2994 -13866 3015 -13832
rect 3049 -13866 6876 -13832
rect 6910 -13866 6963 -13832
rect 1153 -13885 1310 -13884
rect 2994 -13886 6963 -13866
rect 7509 -13831 8255 -13813
rect 7509 -13832 8164 -13831
rect 7509 -13866 7522 -13832
rect 7556 -13865 8164 -13832
rect 8198 -13865 8255 -13831
rect 7556 -13866 8255 -13865
rect 7509 -13887 8255 -13866
rect 8799 -13833 9545 -13814
rect 8799 -13867 8811 -13833
rect 8845 -13867 9453 -13833
rect 9487 -13867 9545 -13833
rect 8799 -13885 9545 -13867
rect 10086 -13826 11058 -13820
rect 10086 -13832 11063 -13826
rect 10086 -13833 10925 -13832
rect 10086 -13834 10741 -13833
rect 10086 -13868 10099 -13834
rect 10133 -13867 10741 -13834
rect 10775 -13867 10832 -13833
rect 10866 -13866 10925 -13833
rect 10959 -13866 11017 -13832
rect 11051 -13866 11063 -13832
rect 11233 -13835 11418 -13827
rect 10866 -13867 11063 -13866
rect 10133 -13868 11063 -13867
rect 10086 -13872 11063 -13868
rect 10086 -13890 11058 -13872
rect 11110 -13909 11120 -13857
rect 11172 -13909 11182 -13857
rect 11233 -13869 11250 -13835
rect 11284 -13869 11344 -13835
rect 11378 -13869 11418 -13835
rect 11233 -13956 11418 -13869
rect 308 -13992 11419 -13956
<< via1 >>
rect -1792 -343 -1740 -291
rect -771 -301 -719 -290
rect -771 -335 -762 -301
rect -762 -335 -728 -301
rect -728 -335 -719 -301
rect -771 -342 -719 -335
rect 982 -377 1034 -325
rect 11120 -268 11172 -259
rect 11120 -302 11129 -268
rect 11129 -302 11163 -268
rect 11163 -302 11172 -268
rect 11120 -311 11172 -302
rect 982 -733 1034 -681
rect 12753 -734 12805 -682
rect 423 -812 475 -802
rect 423 -846 433 -812
rect 433 -846 467 -812
rect 467 -846 475 -812
rect 423 -854 475 -846
rect 12463 -887 12522 -828
rect 7165 -1287 7217 -1235
rect 11118 -1284 11170 -1232
rect 423 -1392 475 -1383
rect 423 -1426 432 -1392
rect 432 -1426 466 -1392
rect 466 -1426 475 -1392
rect 423 -1435 475 -1426
rect 11378 -1355 11430 -1345
rect 11378 -1389 11387 -1355
rect 11387 -1389 11421 -1355
rect 11421 -1389 11430 -1355
rect 11378 -1397 11430 -1389
rect 12752 -1392 12804 -1382
rect 12752 -1426 12773 -1392
rect 12773 -1426 12804 -1392
rect 12752 -1434 12804 -1426
rect 7163 -1815 7215 -1763
rect 12756 -1818 12808 -1766
rect -942 -1943 -890 -1891
rect -217 -1865 -165 -1854
rect -217 -1899 -210 -1865
rect -210 -1899 -176 -1865
rect -176 -1899 -165 -1865
rect -217 -1906 -165 -1899
rect 423 -1900 475 -1890
rect 423 -1934 432 -1900
rect 432 -1934 466 -1900
rect 466 -1934 475 -1900
rect 423 -1942 475 -1934
rect 11375 -1863 11427 -1856
rect 11375 -1897 11386 -1863
rect 11386 -1897 11420 -1863
rect 11420 -1897 11427 -1863
rect 11375 -1908 11427 -1897
rect 428 -2480 480 -2469
rect 428 -2514 436 -2480
rect 436 -2514 470 -2480
rect 470 -2514 480 -2480
rect 428 -2521 480 -2514
rect 11378 -2445 11430 -2436
rect 11378 -2479 11386 -2445
rect 11386 -2479 11420 -2445
rect 11420 -2479 11430 -2445
rect 11378 -2488 11430 -2479
rect 12466 -2441 12480 -2414
rect 12480 -2441 12514 -2414
rect 12514 -2441 12518 -2414
rect 12466 -2466 12518 -2441
rect 12755 -2479 12807 -2472
rect 12755 -2513 12765 -2479
rect 12765 -2513 12799 -2479
rect 12799 -2513 12807 -2479
rect 12755 -2524 12807 -2513
rect 13926 -2485 13978 -2433
rect 12466 -2553 12518 -2528
rect 12466 -2580 12480 -2553
rect 12480 -2580 12514 -2553
rect 12514 -2580 12518 -2553
rect -1968 -2952 -1916 -2944
rect -1968 -2986 -1960 -2952
rect -1960 -2986 -1926 -2952
rect -1926 -2986 -1916 -2952
rect -1968 -2996 -1916 -2986
rect -1792 -2915 -1740 -2906
rect -1792 -2949 -1783 -2915
rect -1783 -2949 -1749 -2915
rect -1749 -2949 -1740 -2915
rect -1792 -2958 -1740 -2949
rect -221 -3033 -169 -2981
rect 11376 -2952 11428 -2943
rect 11376 -2986 11384 -2952
rect 11384 -2986 11418 -2952
rect 11418 -2986 11428 -2952
rect 11376 -2995 11428 -2986
rect -1968 -3114 -1916 -3062
rect -1272 -3118 -1213 -3059
rect 115 -3573 167 -3521
rect 11373 -3567 11425 -3557
rect 11373 -3601 11383 -3567
rect 11383 -3601 11417 -3567
rect 11417 -3601 11425 -3567
rect 11373 -3609 11425 -3601
rect 12466 -3999 12480 -3972
rect 12480 -3999 12514 -3972
rect 12514 -3999 12518 -3972
rect 12466 -4024 12518 -3999
rect 427 -4040 479 -4031
rect 427 -4074 436 -4040
rect 436 -4074 470 -4040
rect 470 -4074 479 -4040
rect 427 -4083 479 -4074
rect 11377 -4077 11429 -4067
rect 11377 -4111 11386 -4077
rect 11386 -4111 11420 -4077
rect 11420 -4111 11429 -4077
rect 11377 -4119 11429 -4111
rect 12755 -4039 12807 -4028
rect 12755 -4073 12765 -4039
rect 12765 -4073 12799 -4039
rect 12799 -4073 12807 -4039
rect 12755 -4080 12807 -4073
rect 12466 -4111 12518 -4086
rect 12466 -4138 12480 -4111
rect 12480 -4138 12514 -4111
rect 12514 -4138 12518 -4111
rect 14628 -4118 14682 -4064
rect -771 -4663 -716 -4608
rect 115 -4695 167 -4643
rect 424 -4619 476 -4610
rect 424 -4653 433 -4619
rect 433 -4653 467 -4619
rect 467 -4653 476 -4619
rect 424 -4662 476 -4653
rect 11375 -4657 11427 -4645
rect 11375 -4691 11384 -4657
rect 11384 -4691 11418 -4657
rect 11418 -4691 11427 -4657
rect 11375 -4697 11427 -4691
rect 7163 -4789 7215 -4737
rect 12756 -4786 12808 -4734
rect 427 -5128 479 -5120
rect 427 -5162 436 -5128
rect 436 -5162 470 -5128
rect 470 -5162 479 -5128
rect 427 -5172 479 -5162
rect 12752 -5126 12804 -5118
rect 11380 -5162 11432 -5152
rect 11380 -5196 11389 -5162
rect 11389 -5196 11423 -5162
rect 11423 -5196 11432 -5162
rect 11380 -5204 11432 -5196
rect 12752 -5160 12773 -5126
rect 12773 -5160 12804 -5126
rect 12752 -5170 12804 -5160
rect 7165 -5317 7217 -5265
rect 11118 -5320 11170 -5268
rect 422 -5708 474 -5699
rect 422 -5742 432 -5708
rect 432 -5742 466 -5708
rect 466 -5742 474 -5708
rect 422 -5751 474 -5742
rect 12463 -5724 12522 -5665
rect 982 -5871 1034 -5819
rect 12753 -5870 12805 -5818
rect -944 -6218 -886 -6207
rect -944 -6252 -932 -6218
rect -932 -6252 -898 -6218
rect -898 -6252 -886 -6218
rect -944 -6263 -886 -6252
rect -772 -6217 -714 -6207
rect -772 -6251 -760 -6217
rect -760 -6251 -726 -6217
rect -726 -6251 -714 -6217
rect -772 -6263 -714 -6251
rect 982 -6227 1034 -6175
rect 11120 -6250 11172 -6241
rect 11120 -6284 11129 -6250
rect 11129 -6284 11163 -6250
rect 11163 -6284 11172 -6250
rect 11120 -6293 11172 -6284
rect 14627 -6274 14682 -6219
rect 15834 -6274 15889 -6219
rect -1271 -6409 -1213 -6353
rect -768 -6409 -715 -6356
rect -772 -6727 -714 -6671
rect 7349 -6726 7407 -6670
rect -2607 -6830 -2554 -6821
rect -2607 -6864 -2599 -6830
rect -2599 -6864 -2565 -6830
rect -2565 -6864 -2554 -6830
rect -2607 -6873 -2554 -6864
rect 5028 -6840 5082 -6786
rect 13925 -6840 13979 -6786
rect -1968 -7003 -1915 -6951
rect -405 -6958 -346 -6899
rect 3736 -6958 3795 -6899
rect 4945 -6977 4999 -6923
rect 15832 -6977 15886 -6923
rect 4945 -7204 4999 -7195
rect 4945 -7238 4955 -7204
rect 4955 -7238 4989 -7204
rect 4989 -7238 4999 -7204
rect 4945 -7249 4999 -7238
rect 2736 -7317 2795 -7258
rect 3736 -7304 3795 -7292
rect 3736 -7338 3747 -7304
rect 3747 -7338 3781 -7304
rect 3781 -7338 3795 -7304
rect 3736 -7351 3795 -7338
rect 5028 -7306 5082 -7299
rect 5028 -7340 5036 -7306
rect 5036 -7340 5070 -7306
rect 5070 -7340 5082 -7306
rect 5028 -7353 5082 -7340
rect 7349 -7264 7407 -7254
rect 7349 -7298 7356 -7264
rect 7356 -7298 7390 -7264
rect 7390 -7298 7407 -7264
rect 7349 -7310 7407 -7298
rect 15971 -7326 16030 -7267
rect -620 -7498 -561 -7439
rect 2736 -7498 2795 -7439
rect -1968 -7960 -1915 -7908
rect -619 -7961 -560 -7902
rect 982 -7993 1034 -7941
rect 11120 -7884 11172 -7875
rect 11120 -7918 11129 -7884
rect 11129 -7918 11163 -7884
rect 11163 -7918 11172 -7884
rect 11120 -7927 11172 -7918
rect 982 -8349 1034 -8297
rect 12753 -8350 12805 -8298
rect 423 -8428 475 -8418
rect 423 -8462 433 -8428
rect 433 -8462 467 -8428
rect 467 -8462 475 -8428
rect 423 -8470 475 -8462
rect 12463 -8503 12522 -8444
rect 15972 -8475 16031 -8416
rect 7165 -8903 7217 -8851
rect 11118 -8900 11170 -8848
rect 423 -9008 475 -8999
rect 423 -9042 432 -9008
rect 432 -9042 466 -9008
rect 466 -9042 475 -9008
rect 423 -9051 475 -9042
rect 11378 -8971 11430 -8961
rect 11378 -9005 11387 -8971
rect 11387 -9005 11421 -8971
rect 11421 -9005 11430 -8971
rect 11378 -9013 11430 -9005
rect 12752 -9008 12804 -8998
rect 12752 -9042 12773 -9008
rect 12773 -9042 12804 -9008
rect 12752 -9050 12804 -9042
rect 7163 -9431 7215 -9379
rect 12756 -9434 12808 -9382
rect -942 -9559 -890 -9507
rect -217 -9481 -165 -9470
rect -217 -9515 -210 -9481
rect -210 -9515 -176 -9481
rect -176 -9515 -165 -9481
rect -217 -9522 -165 -9515
rect 423 -9516 475 -9506
rect 423 -9550 432 -9516
rect 432 -9550 466 -9516
rect 466 -9550 475 -9516
rect 423 -9558 475 -9550
rect 11375 -9479 11427 -9472
rect 11375 -9513 11386 -9479
rect 11386 -9513 11420 -9479
rect 11420 -9513 11427 -9479
rect 11375 -9524 11427 -9513
rect 428 -10096 480 -10085
rect 428 -10130 436 -10096
rect 436 -10130 470 -10096
rect 470 -10130 480 -10096
rect 428 -10137 480 -10130
rect 11378 -10061 11430 -10052
rect 11378 -10095 11386 -10061
rect 11386 -10095 11420 -10061
rect 11420 -10095 11430 -10061
rect 11378 -10104 11430 -10095
rect 12466 -10057 12480 -10030
rect 12480 -10057 12514 -10030
rect 12514 -10057 12518 -10030
rect 12466 -10082 12518 -10057
rect 12755 -10095 12807 -10088
rect 12755 -10129 12765 -10095
rect 12765 -10129 12799 -10095
rect 12799 -10129 12807 -10095
rect 12755 -10140 12807 -10129
rect 12466 -10169 12518 -10144
rect 12466 -10196 12480 -10169
rect 12480 -10196 12514 -10169
rect 12514 -10196 12518 -10169
rect -2607 -10543 -2554 -10490
rect -1969 -10499 -1915 -10489
rect -1969 -10533 -1961 -10499
rect -1961 -10533 -1927 -10499
rect -1927 -10533 -1915 -10499
rect -1969 -10543 -1915 -10533
rect -1823 -10534 -1769 -10525
rect -1823 -10568 -1813 -10534
rect -1813 -10568 -1779 -10534
rect -1779 -10568 -1769 -10534
rect -1823 -10579 -1769 -10568
rect -221 -10649 -169 -10597
rect 11376 -10568 11428 -10559
rect 11376 -10602 11384 -10568
rect 11384 -10602 11418 -10568
rect 11418 -10602 11428 -10568
rect 11376 -10611 11428 -10602
rect 115 -11189 167 -11137
rect 11373 -11183 11425 -11173
rect 11373 -11217 11383 -11183
rect 11383 -11217 11417 -11183
rect 11417 -11217 11425 -11183
rect 11373 -11225 11425 -11217
rect 12466 -11615 12480 -11588
rect 12480 -11615 12514 -11588
rect 12514 -11615 12518 -11588
rect 12466 -11640 12518 -11615
rect 427 -11656 479 -11647
rect 427 -11690 436 -11656
rect 436 -11690 470 -11656
rect 470 -11690 479 -11656
rect 427 -11699 479 -11690
rect 11377 -11693 11429 -11683
rect 11377 -11727 11386 -11693
rect 11386 -11727 11420 -11693
rect 11420 -11727 11429 -11693
rect 11377 -11735 11429 -11727
rect 12755 -11655 12807 -11644
rect 12755 -11689 12765 -11655
rect 12765 -11689 12799 -11655
rect 12799 -11689 12807 -11655
rect 12755 -11696 12807 -11689
rect 12466 -11727 12518 -11702
rect 12466 -11754 12480 -11727
rect 12480 -11754 12514 -11727
rect 12514 -11754 12518 -11727
rect -404 -12282 -346 -12224
rect 115 -12311 167 -12259
rect 424 -12235 476 -12226
rect 424 -12269 433 -12235
rect 433 -12269 467 -12235
rect 467 -12269 476 -12235
rect 424 -12278 476 -12269
rect 11375 -12273 11427 -12261
rect 11375 -12307 11384 -12273
rect 11384 -12307 11418 -12273
rect 11418 -12307 11427 -12273
rect 11375 -12313 11427 -12307
rect 7163 -12405 7215 -12353
rect 12756 -12402 12808 -12350
rect 427 -12744 479 -12736
rect 427 -12778 436 -12744
rect 436 -12778 470 -12744
rect 470 -12778 479 -12744
rect 427 -12788 479 -12778
rect 12752 -12742 12804 -12734
rect 11380 -12778 11432 -12768
rect 11380 -12812 11389 -12778
rect 11389 -12812 11423 -12778
rect 11423 -12812 11432 -12778
rect 11380 -12820 11432 -12812
rect 12752 -12776 12773 -12742
rect 12773 -12776 12804 -12742
rect 12752 -12786 12804 -12776
rect 7165 -12933 7217 -12881
rect 11118 -12936 11170 -12884
rect 422 -13324 474 -13315
rect 422 -13358 432 -13324
rect 432 -13358 466 -13324
rect 466 -13358 474 -13324
rect 422 -13367 474 -13358
rect 12463 -13340 12522 -13281
rect 982 -13487 1034 -13435
rect 12753 -13486 12805 -13434
rect -944 -13834 -886 -13823
rect -944 -13868 -932 -13834
rect -932 -13868 -898 -13834
rect -898 -13868 -886 -13834
rect -944 -13879 -886 -13868
rect 982 -13843 1034 -13791
rect -1824 -13971 -1769 -13916
rect 11120 -13866 11172 -13857
rect 11120 -13900 11129 -13866
rect 11129 -13900 11163 -13866
rect 11163 -13900 11172 -13866
rect 11120 -13909 11172 -13900
<< metal2 >>
rect 11110 -259 11178 -243
rect -1792 -291 -1740 -280
rect -1792 -2906 -1740 -343
rect -771 -290 -716 -279
rect -719 -342 -716 -290
rect 11110 -311 11120 -259
rect 11172 -311 11178 -259
rect -1968 -2944 -1915 -2933
rect -1916 -2996 -1915 -2944
rect -1792 -2988 -1740 -2958
rect -944 -1891 -886 -1879
rect -944 -1943 -942 -1891
rect -890 -1943 -886 -1891
rect -1968 -3062 -1915 -2996
rect -1916 -3114 -1915 -3062
rect -2607 -6821 -2554 -6811
rect -2607 -10490 -2554 -6873
rect -1968 -6951 -1915 -3114
rect -1272 -3059 -1213 -3049
rect -1272 -6353 -1213 -3118
rect -944 -6207 -886 -1943
rect -771 -4608 -716 -342
rect 979 -325 1039 -314
rect 979 -377 982 -325
rect 1034 -377 1039 -325
rect 979 -681 1039 -377
rect 979 -733 982 -681
rect 1034 -733 1039 -681
rect 979 -743 1039 -733
rect 423 -802 475 -792
rect 423 -1383 475 -854
rect 423 -1445 475 -1435
rect 7154 -1235 7223 -1225
rect 7154 -1287 7165 -1235
rect 7217 -1287 7223 -1235
rect 7154 -1763 7223 -1287
rect 11110 -1232 11178 -311
rect 12751 -682 12806 -671
rect 12751 -734 12753 -682
rect 12805 -734 12806 -682
rect 11110 -1284 11118 -1232
rect 11170 -1284 11178 -1232
rect 11110 -1294 11178 -1284
rect 12463 -828 12522 -818
rect 7154 -1815 7163 -1763
rect 7215 -1815 7223 -1763
rect 7154 -1821 7223 -1815
rect 11372 -1345 11434 -1332
rect 11372 -1397 11378 -1345
rect 11430 -1397 11434 -1345
rect 7163 -1825 7215 -1821
rect -217 -1854 -165 -1844
rect -227 -1906 -217 -1860
rect 11372 -1856 11434 -1397
rect -165 -1906 -164 -1860
rect 427 -1880 476 -1879
rect -227 -2981 -164 -1906
rect 423 -1890 476 -1880
rect 475 -1942 476 -1890
rect 11372 -1908 11375 -1856
rect 11427 -1908 11434 -1856
rect 11372 -1921 11434 -1908
rect 423 -1952 476 -1942
rect 427 -2459 476 -1952
rect 12463 -2414 12522 -887
rect 12751 -1382 12806 -734
rect 12751 -1434 12752 -1382
rect 12804 -1434 12806 -1382
rect 12751 -1435 12806 -1434
rect 12752 -1444 12804 -1435
rect 11374 -2436 11433 -2423
rect 427 -2469 480 -2459
rect 427 -2521 428 -2469
rect 427 -2531 480 -2521
rect 11374 -2488 11378 -2436
rect 11430 -2488 11433 -2436
rect 427 -2533 476 -2531
rect -227 -3033 -221 -2981
rect -169 -3033 -164 -2981
rect 11374 -2943 11433 -2488
rect 12463 -2466 12466 -2414
rect 12518 -2466 12522 -2414
rect 12463 -2528 12522 -2466
rect 12463 -2580 12466 -2528
rect 12518 -2580 12522 -2528
rect 12753 -1766 12812 -1753
rect 12753 -1818 12756 -1766
rect 12808 -1818 12812 -1766
rect 12753 -2472 12812 -1818
rect 12753 -2524 12755 -2472
rect 12807 -2524 12812 -2472
rect 12753 -2538 12812 -2524
rect 13925 -2433 13979 -2422
rect 13925 -2485 13926 -2433
rect 13978 -2485 13979 -2433
rect 12463 -2593 12522 -2580
rect 11374 -2995 11376 -2943
rect 11428 -2995 11433 -2943
rect 11374 -3008 11433 -2995
rect -227 -3048 -164 -3033
rect -771 -4673 -716 -4663
rect 113 -3521 170 -3507
rect 113 -3573 115 -3521
rect 167 -3573 170 -3521
rect 11375 -3547 11426 -3545
rect 113 -4643 170 -3573
rect 11373 -3557 11426 -3547
rect 11425 -3609 11426 -3557
rect 11373 -3619 11426 -3609
rect 425 -4031 480 -4018
rect 425 -4083 427 -4031
rect 479 -4083 480 -4031
rect 425 -4600 480 -4083
rect 11375 -4057 11426 -3619
rect 12463 -3972 12522 -3959
rect 12463 -4024 12466 -3972
rect 12518 -4024 12522 -3972
rect 11375 -4067 11429 -4057
rect 11375 -4119 11377 -4067
rect 11375 -4129 11429 -4119
rect 12463 -4086 12522 -4024
rect 11375 -4132 11426 -4129
rect 113 -4695 115 -4643
rect 167 -4695 170 -4643
rect 424 -4610 480 -4600
rect 476 -4662 480 -4610
rect 12463 -4138 12466 -4086
rect 12518 -4138 12522 -4086
rect 424 -4672 480 -4662
rect 425 -4675 480 -4672
rect 11373 -4645 11435 -4633
rect 113 -4701 170 -4695
rect 11373 -4697 11375 -4645
rect 11427 -4697 11435 -4645
rect 115 -4705 167 -4701
rect 7163 -4731 7215 -4727
rect 7154 -4737 7223 -4731
rect 7154 -4789 7163 -4737
rect 7215 -4789 7223 -4737
rect 424 -5110 476 -5107
rect 424 -5120 479 -5110
rect 424 -5172 427 -5120
rect 424 -5182 479 -5172
rect 424 -5689 476 -5182
rect 7154 -5265 7223 -4789
rect 11373 -5152 11435 -4697
rect 11373 -5204 11380 -5152
rect 11432 -5204 11435 -5152
rect 11373 -5217 11435 -5204
rect 7154 -5317 7165 -5265
rect 7217 -5317 7223 -5265
rect 7154 -5327 7223 -5317
rect 11110 -5268 11178 -5258
rect 11110 -5320 11118 -5268
rect 11170 -5320 11178 -5268
rect 422 -5699 476 -5689
rect 474 -5751 476 -5699
rect 422 -5761 476 -5751
rect 424 -5764 476 -5761
rect 979 -5819 1039 -5809
rect 979 -5871 982 -5819
rect 1034 -5871 1039 -5819
rect 979 -6175 1039 -5871
rect -944 -6273 -886 -6263
rect -773 -6207 -712 -6194
rect -773 -6263 -772 -6207
rect -714 -6263 -712 -6207
rect 979 -6227 982 -6175
rect 1034 -6227 1039 -6175
rect 979 -6238 1039 -6227
rect -1272 -6409 -1271 -6353
rect -1272 -6420 -1213 -6409
rect -773 -6356 -712 -6263
rect 11110 -6241 11178 -5320
rect 12463 -5665 12522 -4138
rect 12753 -4028 12812 -4014
rect 12753 -4080 12755 -4028
rect 12807 -4080 12812 -4028
rect 12753 -4734 12812 -4080
rect 12753 -4786 12756 -4734
rect 12808 -4786 12812 -4734
rect 12753 -4799 12812 -4786
rect 12752 -5117 12804 -5108
rect 12463 -5734 12522 -5724
rect 12751 -5118 12806 -5117
rect 12751 -5170 12752 -5118
rect 12804 -5170 12806 -5118
rect 12751 -5818 12806 -5170
rect 12751 -5870 12753 -5818
rect 12805 -5870 12806 -5818
rect 12751 -5881 12806 -5870
rect 11110 -6293 11120 -6241
rect 11172 -6293 11178 -6241
rect 11110 -6309 11178 -6293
rect -773 -6409 -768 -6356
rect -715 -6409 -712 -6356
rect -773 -6671 -712 -6409
rect -773 -6709 -772 -6671
rect -714 -6709 -712 -6671
rect 7345 -6670 7409 -6658
rect -772 -6737 -714 -6727
rect 7345 -6726 7349 -6670
rect 7407 -6726 7409 -6670
rect 5028 -6786 5082 -6776
rect -1968 -7010 -1915 -7003
rect -405 -6899 -346 -6889
rect -620 -7439 -561 -7429
rect -561 -7498 -559 -7460
rect -2607 -10553 -2554 -10543
rect -1969 -7908 -1915 -7898
rect -1969 -7960 -1968 -7908
rect -1969 -10489 -1915 -7960
rect -620 -7902 -559 -7498
rect -620 -7961 -619 -7902
rect -560 -7961 -559 -7902
rect -620 -7973 -559 -7961
rect -944 -9507 -886 -9495
rect -944 -9559 -942 -9507
rect -890 -9559 -886 -9507
rect -1969 -10556 -1915 -10543
rect -1824 -10525 -1769 -10514
rect -1824 -10579 -1823 -10525
rect -1824 -13916 -1769 -10579
rect -944 -13823 -886 -9559
rect -405 -12224 -346 -6958
rect 3736 -6899 3795 -6889
rect 2736 -7255 2795 -7248
rect 2735 -7258 2796 -7255
rect 2735 -7317 2736 -7258
rect 2795 -7317 2796 -7258
rect 2735 -7439 2796 -7317
rect 3736 -7292 3795 -6958
rect 4945 -6923 4999 -6905
rect 4945 -7195 4999 -6977
rect 4945 -7259 4999 -7249
rect 3736 -7361 3795 -7351
rect 5028 -7299 5082 -6840
rect 7345 -7254 7409 -6726
rect 13925 -6786 13979 -2485
rect 14627 -4064 14682 -4053
rect 14627 -4118 14628 -4064
rect 14627 -6219 14682 -4118
rect 14627 -6284 14682 -6274
rect 15829 -6219 15892 -6206
rect 15829 -6274 15834 -6219
rect 15889 -6274 15892 -6219
rect 13925 -6850 13979 -6840
rect 15829 -6923 15892 -6274
rect 15829 -6977 15832 -6923
rect 15886 -6977 15892 -6923
rect 15829 -6991 15892 -6977
rect 7345 -7310 7349 -7254
rect 7407 -7310 7409 -7254
rect 15971 -7262 16030 -7257
rect 7345 -7339 7409 -7310
rect 15968 -7267 16033 -7262
rect 15968 -7326 15971 -7267
rect 16030 -7326 16033 -7267
rect 5028 -7363 5082 -7353
rect 2735 -7498 2736 -7439
rect 2795 -7498 2796 -7439
rect 2735 -7508 2796 -7498
rect 11110 -7875 11178 -7859
rect 11110 -7927 11120 -7875
rect 11172 -7927 11178 -7875
rect 979 -7941 1039 -7930
rect 979 -7993 982 -7941
rect 1034 -7993 1039 -7941
rect 979 -8297 1039 -7993
rect 979 -8349 982 -8297
rect 1034 -8349 1039 -8297
rect 979 -8359 1039 -8349
rect 423 -8418 475 -8408
rect 423 -8999 475 -8470
rect 423 -9061 475 -9051
rect 7154 -8851 7223 -8841
rect 7154 -8903 7165 -8851
rect 7217 -8903 7223 -8851
rect 7154 -9379 7223 -8903
rect 11110 -8848 11178 -7927
rect 12751 -8298 12806 -8287
rect 12751 -8350 12753 -8298
rect 12805 -8350 12806 -8298
rect 11110 -8900 11118 -8848
rect 11170 -8900 11178 -8848
rect 11110 -8910 11178 -8900
rect 12463 -8444 12522 -8434
rect 7154 -9431 7163 -9379
rect 7215 -9431 7223 -9379
rect 7154 -9437 7223 -9431
rect 11372 -8961 11434 -8948
rect 11372 -9013 11378 -8961
rect 11430 -9013 11434 -8961
rect 7163 -9441 7215 -9437
rect -217 -9470 -165 -9460
rect -227 -9522 -217 -9476
rect 11372 -9472 11434 -9013
rect -165 -9522 -164 -9476
rect 427 -9496 476 -9495
rect -227 -10597 -164 -9522
rect 423 -9506 476 -9496
rect 475 -9558 476 -9506
rect 11372 -9524 11375 -9472
rect 11427 -9524 11434 -9472
rect 11372 -9537 11434 -9524
rect 423 -9568 476 -9558
rect 427 -10075 476 -9568
rect 12463 -10030 12522 -8503
rect 12751 -8998 12806 -8350
rect 15968 -8416 16033 -7326
rect 15968 -8475 15972 -8416
rect 16031 -8475 16033 -8416
rect 15968 -8489 16033 -8475
rect 12751 -9050 12752 -8998
rect 12804 -9050 12806 -8998
rect 12751 -9051 12806 -9050
rect 12752 -9060 12804 -9051
rect 11374 -10052 11433 -10039
rect 427 -10085 480 -10075
rect 427 -10137 428 -10085
rect 427 -10147 480 -10137
rect 11374 -10104 11378 -10052
rect 11430 -10104 11433 -10052
rect 427 -10149 476 -10147
rect -227 -10649 -221 -10597
rect -169 -10649 -164 -10597
rect 11374 -10559 11433 -10104
rect 12463 -10082 12466 -10030
rect 12518 -10082 12522 -10030
rect 12463 -10144 12522 -10082
rect 12463 -10196 12466 -10144
rect 12518 -10196 12522 -10144
rect 12753 -9382 12812 -9369
rect 12753 -9434 12756 -9382
rect 12808 -9434 12812 -9382
rect 12753 -10088 12812 -9434
rect 12753 -10140 12755 -10088
rect 12807 -10140 12812 -10088
rect 12753 -10154 12812 -10140
rect 12463 -10209 12522 -10196
rect 11374 -10611 11376 -10559
rect 11428 -10611 11433 -10559
rect 11374 -10624 11433 -10611
rect -227 -10664 -164 -10649
rect -405 -12282 -404 -12224
rect -405 -12293 -346 -12282
rect 113 -11137 170 -11123
rect 113 -11189 115 -11137
rect 167 -11189 170 -11137
rect 11375 -11163 11426 -11161
rect 113 -12259 170 -11189
rect 11373 -11173 11426 -11163
rect 11425 -11225 11426 -11173
rect 11373 -11235 11426 -11225
rect 425 -11647 480 -11634
rect 425 -11699 427 -11647
rect 479 -11699 480 -11647
rect 425 -12216 480 -11699
rect 11375 -11673 11426 -11235
rect 12463 -11588 12522 -11575
rect 12463 -11640 12466 -11588
rect 12518 -11640 12522 -11588
rect 11375 -11683 11429 -11673
rect 11375 -11735 11377 -11683
rect 11375 -11745 11429 -11735
rect 12463 -11702 12522 -11640
rect 11375 -11748 11426 -11745
rect 113 -12311 115 -12259
rect 167 -12311 170 -12259
rect 424 -12226 480 -12216
rect 476 -12278 480 -12226
rect 12463 -11754 12466 -11702
rect 12518 -11754 12522 -11702
rect 424 -12288 480 -12278
rect 425 -12291 480 -12288
rect 11373 -12261 11435 -12249
rect 113 -12317 170 -12311
rect 11373 -12313 11375 -12261
rect 11427 -12313 11435 -12261
rect 115 -12321 167 -12317
rect 7163 -12347 7215 -12343
rect 7154 -12353 7223 -12347
rect 7154 -12405 7163 -12353
rect 7215 -12405 7223 -12353
rect 424 -12726 476 -12723
rect 424 -12736 479 -12726
rect 424 -12788 427 -12736
rect 424 -12798 479 -12788
rect 424 -13305 476 -12798
rect 7154 -12881 7223 -12405
rect 11373 -12768 11435 -12313
rect 11373 -12820 11380 -12768
rect 11432 -12820 11435 -12768
rect 11373 -12833 11435 -12820
rect 7154 -12933 7165 -12881
rect 7217 -12933 7223 -12881
rect 7154 -12943 7223 -12933
rect 11110 -12884 11178 -12874
rect 11110 -12936 11118 -12884
rect 11170 -12936 11178 -12884
rect 422 -13315 476 -13305
rect 474 -13367 476 -13315
rect 422 -13377 476 -13367
rect 424 -13380 476 -13377
rect 979 -13435 1039 -13425
rect 979 -13487 982 -13435
rect 1034 -13487 1039 -13435
rect 979 -13791 1039 -13487
rect 979 -13843 982 -13791
rect 1034 -13843 1039 -13791
rect 979 -13854 1039 -13843
rect -944 -13889 -886 -13879
rect 11110 -13857 11178 -12936
rect 12463 -13281 12522 -11754
rect 12753 -11644 12812 -11630
rect 12753 -11696 12755 -11644
rect 12807 -11696 12812 -11644
rect 12753 -12350 12812 -11696
rect 12753 -12402 12756 -12350
rect 12808 -12402 12812 -12350
rect 12753 -12415 12812 -12402
rect 12752 -12733 12804 -12724
rect 12463 -13350 12522 -13340
rect 12751 -12734 12806 -12733
rect 12751 -12786 12752 -12734
rect 12804 -12786 12806 -12734
rect 12751 -13434 12806 -12786
rect 12751 -13486 12753 -13434
rect 12805 -13486 12806 -13434
rect 12751 -13497 12806 -13486
rect 11110 -13909 11120 -13857
rect 11172 -13909 11178 -13857
rect 11110 -13925 11178 -13909
rect -1824 -13981 -1769 -13971
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 13655 0 -1 -556
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_1
timestamp 1655495960
transform 1 0 13655 0 -1 -1644
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_2
timestamp 1655495960
transform 1 0 13655 0 1 -1644
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_3
timestamp 1655495960
transform 1 0 13655 0 1 -2732
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_4
timestamp 1655495960
transform 1 0 13655 0 -1 -3820
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_5
timestamp 1655495960
transform 1 0 13655 0 1 -4908
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_6
timestamp 1655495960
transform 1 0 13655 0 -1 -4908
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_7
timestamp 1655495960
transform 1 0 13655 0 1 -5996
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_8
timestamp 1655495960
transform 1 0 13655 0 1 -13612
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_9
timestamp 1655495960
transform 1 0 13655 0 -1 -12524
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_10
timestamp 1655495960
transform 1 0 13655 0 1 -12524
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_11
timestamp 1655495960
transform 1 0 13655 0 -1 -11436
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_12
timestamp 1655495960
transform 1 0 13655 0 1 -10348
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_13
timestamp 1655495960
transform 1 0 13655 0 -1 -9260
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_14
timestamp 1655495960
transform 1 0 13655 0 1 -9260
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_15
timestamp 1655495960
transform 1 0 13655 0 -1 -8172
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 2339 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_1
timestamp 1655495960
transform 1 0 6847 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_2
timestamp 1655495960
transform 1 0 8135 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_3
timestamp 1655495960
transform 1 0 9423 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_5
timestamp 1655495960
transform -1 0 11447 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_6
timestamp 1655495960
transform -1 0 8871 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_8
timestamp 1655495960
transform -1 0 6295 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_10
timestamp 1655495960
transform -1 0 3719 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_11
timestamp 1655495960
transform -1 0 3719 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_13
timestamp 1655495960
transform -1 0 6295 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_15
timestamp 1655495960
transform -1 0 8871 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_17
timestamp 1655495960
transform -1 0 11447 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_18
timestamp 1655495960
transform 1 0 2983 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_20
timestamp 1655495960
transform 1 0 5559 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_22
timestamp 1655495960
transform 1 0 8135 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_24
timestamp 1655495960
transform 1 0 10711 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_25
timestamp 1655495960
transform 1 0 2983 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_27
timestamp 1655495960
transform 1 0 5559 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_29
timestamp 1655495960
transform 1 0 8135 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_31
timestamp 1655495960
transform 1 0 10711 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_32
timestamp 1655495960
transform -1 0 3719 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_34
timestamp 1655495960
transform -1 0 6295 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_36
timestamp 1655495960
transform -1 0 8871 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_38
timestamp 1655495960
transform -1 0 11447 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_39
timestamp 1655495960
transform -1 0 1143 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_42
timestamp 1655495960
transform -1 0 1143 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_44
timestamp 1655495960
transform 1 0 407 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_47
timestamp 1655495960
transform 1 0 407 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_48
timestamp 1655495960
transform -1 0 1143 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_49
timestamp 1655495960
transform -1 0 -145 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_50
timestamp 1655495960
transform -1 0 1143 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_52
timestamp 1655495960
transform -1 0 3719 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_54
timestamp 1655495960
transform -1 0 6295 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_56
timestamp 1655495960
transform -1 0 8871 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_58
timestamp 1655495960
transform -1 0 11447 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_59
timestamp 1655495960
transform 1 0 407 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_61
timestamp 1655495960
transform 1 0 2983 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_63
timestamp 1655495960
transform 1 0 5559 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_65
timestamp 1655495960
transform 1 0 8135 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_67
timestamp 1655495960
transform 1 0 10711 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_68
timestamp 1655495960
transform -1 0 -145 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_69
timestamp 1655495960
transform -1 0 1143 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_71
timestamp 1655495960
transform -1 0 3719 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_73
timestamp 1655495960
transform -1 0 6295 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_75
timestamp 1655495960
transform -1 0 8871 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_77
timestamp 1655495960
transform -1 0 11447 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_78
timestamp 1655495960
transform 1 0 407 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_80
timestamp 1655495960
transform 1 0 2983 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_82
timestamp 1655495960
transform 1 0 5559 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_84
timestamp 1655495960
transform 1 0 8135 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_86
timestamp 1655495960
transform 1 0 10711 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_87
timestamp 1655495960
transform -1 0 1143 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_89
timestamp 1655495960
transform 1 0 2339 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_90
timestamp 1655495960
transform -1 0 3719 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_92
timestamp 1655495960
transform -1 0 6295 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_93
timestamp 1655495960
transform 1 0 6847 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_95
timestamp 1655495960
transform 1 0 8135 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_96
timestamp 1655495960
transform -1 0 8871 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_97
timestamp 1655495960
transform 1 0 9423 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_99
timestamp 1655495960
transform -1 0 11447 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_100
timestamp 1655495960
transform 1 0 2339 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_101
timestamp 1655495960
transform 1 0 6847 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_102
timestamp 1655495960
transform 1 0 8135 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_103
timestamp 1655495960
transform 1 0 9423 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_104
timestamp 1655495960
transform -1 0 1143 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_107
timestamp 1655495960
transform -1 0 3719 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_108
timestamp 1655495960
transform -1 0 6295 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_109
timestamp 1655495960
transform -1 0 8871 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_112
timestamp 1655495960
transform -1 0 11447 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_113
timestamp 1655495960
transform 1 0 407 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_116
timestamp 1655495960
transform 1 0 2983 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_117
timestamp 1655495960
transform 1 0 5559 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_118
timestamp 1655495960
transform 1 0 8135 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_121
timestamp 1655495960
transform 1 0 10711 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_122
timestamp 1655495960
transform -1 0 -145 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_123
timestamp 1655495960
transform -1 0 1143 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_125
timestamp 1655495960
transform -1 0 3719 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_127
timestamp 1655495960
transform -1 0 6295 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_129
timestamp 1655495960
transform -1 0 8871 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_131
timestamp 1655495960
transform -1 0 11447 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_132
timestamp 1655495960
transform 1 0 407 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_134
timestamp 1655495960
transform 1 0 2983 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_136
timestamp 1655495960
transform 1 0 5559 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_138
timestamp 1655495960
transform 1 0 8135 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_140
timestamp 1655495960
transform 1 0 10711 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_141
timestamp 1655495960
transform -1 0 1143 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_142
timestamp 1655495960
transform -1 0 1143 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_146
timestamp 1655495960
transform -1 0 3719 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_147
timestamp 1655495960
transform -1 0 3719 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_149
timestamp 1655495960
transform -1 0 6295 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_150
timestamp 1655495960
transform -1 0 6295 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_152
timestamp 1655495960
transform -1 0 8871 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_154
timestamp 1655495960
transform -1 0 8871 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_157
timestamp 1655495960
transform -1 0 11447 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_158
timestamp 1655495960
transform -1 0 11447 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_159
timestamp 1655495960
transform 1 0 407 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_162
timestamp 1655495960
transform 1 0 2983 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_163
timestamp 1655495960
transform 1 0 5559 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_164
timestamp 1655495960
transform 1 0 8135 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_167
timestamp 1655495960
transform 1 0 10711 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_168
timestamp 1655495960
transform -1 0 1143 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_169
timestamp 1655495960
transform -1 0 -145 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_172
timestamp 1655495960
transform -1 0 3719 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_173
timestamp 1655495960
transform -1 0 6295 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_174
timestamp 1655495960
transform -1 0 8871 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_177
timestamp 1655495960
transform -1 0 11447 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_178
timestamp 1655495960
transform 1 0 407 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_180
timestamp 1655495960
transform 1 0 2983 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_182
timestamp 1655495960
transform 1 0 5559 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_184
timestamp 1655495960
transform 1 0 8135 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_186
timestamp 1655495960
transform 1 0 10711 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_187
timestamp 1655495960
transform -1 0 1143 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_190
timestamp 1655495960
transform -1 0 3719 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_191
timestamp 1655495960
transform -1 0 6295 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_193
timestamp 1655495960
transform -1 0 8871 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_195
timestamp 1655495960
transform -1 0 11447 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_196
timestamp 1655495960
transform 1 0 2339 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_197
timestamp 1655495960
transform 1 0 6847 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_198
timestamp 1655495960
transform 1 0 8135 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  sky130_fd_sc_hd__clkdlybuf4s50_1_199
timestamp 1655495960
transform 1 0 9423 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 1051 0 1 -556
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_1
timestamp 1655495960
transform 1 0 1051 0 -1 -5996
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_2
timestamp 1655495960
transform 1 0 1051 0 -1 -13612
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_3
timestamp 1655495960
transform 1 0 1051 0 1 -8172
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_4
timestamp 1655495960
transform -1 0 3167 0 -1 -7084
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_5
timestamp 1655495960
transform 1 0 -1985 0 -1 -2732
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  sky130_fd_sc_hd__clkinv_1_6
timestamp 1655495960
transform 1 0 -1985 0 -1 -10348
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 -145 0 1 -556
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1655495960
transform 1 0 12459 0 1 -1644
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1655495960
transform 1 0 12459 0 1 -2732
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1655495960
transform 1 0 12459 0 -1 -3820
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_4
timestamp 1655495960
transform 1 0 12459 0 -1 -4908
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_5
timestamp 1655495960
transform 1 0 -145 0 -1 -5996
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_6
timestamp 1655495960
transform 1 0 -145 0 -1 -13612
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_7
timestamp 1655495960
transform 1 0 12459 0 -1 -12524
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_8
timestamp 1655495960
transform 1 0 12459 0 -1 -11436
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_9
timestamp 1655495960
transform 1 0 12459 0 1 -10348
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_10
timestamp 1655495960
transform 1 0 12459 0 1 -9260
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_11
timestamp 1655495960
transform 1 0 -145 0 1 -8172
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 -2997 0 1 -7084
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 -1433 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1655495960
transform 1 0 591 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1655495960
transform 1 0 1419 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1655495960
transform 1 0 1879 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1655495960
transform 1 0 6387 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1655495960
transform 1 0 7675 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1655495960
transform 1 0 8963 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_7
timestamp 1655495960
transform 1 0 10251 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_8
timestamp 1655495960
transform 1 0 -605 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_9
timestamp 1655495960
transform 1 0 11631 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_10
timestamp 1655495960
transform -1 0 11999 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_11
timestamp 1655495960
transform -1 0 10711 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_12
timestamp 1655495960
transform -1 0 9331 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_13
timestamp 1655495960
transform -1 0 8043 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_14
timestamp 1655495960
transform -1 0 6755 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_15
timestamp 1655495960
transform -1 0 5467 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_16
timestamp 1655495960
transform -1 0 4179 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_17
timestamp 1655495960
transform -1 0 2891 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_18
timestamp 1655495960
transform -1 0 2891 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_19
timestamp 1655495960
transform -1 0 4179 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_20
timestamp 1655495960
transform -1 0 5467 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_21
timestamp 1655495960
transform -1 0 6755 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_22
timestamp 1655495960
transform -1 0 8043 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_23
timestamp 1655495960
transform -1 0 9331 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_24
timestamp 1655495960
transform -1 0 10711 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_25
timestamp 1655495960
transform -1 0 11999 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_26
timestamp 1655495960
transform -1 0 2891 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_27
timestamp 1655495960
transform -1 0 4179 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_28
timestamp 1655495960
transform -1 0 5467 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_29
timestamp 1655495960
transform -1 0 6755 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_30
timestamp 1655495960
transform -1 0 8043 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_31
timestamp 1655495960
transform -1 0 9331 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_32
timestamp 1655495960
transform -1 0 10711 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_33
timestamp 1655495960
transform -1 0 11999 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_34
timestamp 1655495960
transform -1 0 2891 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_35
timestamp 1655495960
transform -1 0 4179 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_36
timestamp 1655495960
transform -1 0 5467 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_37
timestamp 1655495960
transform -1 0 6755 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_38
timestamp 1655495960
transform -1 0 8043 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_39
timestamp 1655495960
transform -1 0 9331 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_40
timestamp 1655495960
transform -1 0 10711 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_41
timestamp 1655495960
transform -1 0 11999 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_42
timestamp 1655495960
transform -1 0 2891 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_43
timestamp 1655495960
transform -1 0 4179 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_44
timestamp 1655495960
transform -1 0 5467 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_45
timestamp 1655495960
transform -1 0 6755 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_46
timestamp 1655495960
transform -1 0 8043 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_47
timestamp 1655495960
transform -1 0 9331 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_48
timestamp 1655495960
transform -1 0 10711 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_49
timestamp 1655495960
transform -1 0 11999 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_50
timestamp 1655495960
transform -1 0 315 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_51
timestamp 1655495960
transform -1 0 1603 0 -1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_52
timestamp 1655495960
transform -1 0 1603 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_53
timestamp 1655495960
transform -1 0 315 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_54
timestamp 1655495960
transform -1 0 1603 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_55
timestamp 1655495960
transform -1 0 315 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_56
timestamp 1655495960
transform -1 0 1603 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_57
timestamp 1655495960
transform -1 0 1603 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_58
timestamp 1655495960
transform -1 0 315 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_59
timestamp 1655495960
transform -1 0 315 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_60
timestamp 1655495960
transform 1 0 3167 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_61
timestamp 1655495960
transform -1 0 315 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_62
timestamp 1655495960
transform 1 0 13195 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_63
timestamp 1655495960
transform 1 0 13195 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_64
timestamp 1655495960
transform -1 0 1603 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_65
timestamp 1655495960
transform -1 0 2891 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_66
timestamp 1655495960
transform -1 0 4179 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_67
timestamp 1655495960
transform -1 0 5467 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_68
timestamp 1655495960
transform -1 0 6755 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_69
timestamp 1655495960
transform -1 0 8043 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_70
timestamp 1655495960
transform -1 0 9331 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_71
timestamp 1655495960
transform -1 0 10711 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_72
timestamp 1655495960
transform -1 0 11999 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_73
timestamp 1655495960
transform -1 0 315 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_74
timestamp 1655495960
transform -1 0 1603 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_75
timestamp 1655495960
transform -1 0 2891 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_76
timestamp 1655495960
transform -1 0 4179 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_77
timestamp 1655495960
transform -1 0 5467 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_78
timestamp 1655495960
transform -1 0 6755 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_79
timestamp 1655495960
transform -1 0 8043 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_80
timestamp 1655495960
transform -1 0 9331 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_81
timestamp 1655495960
transform -1 0 10711 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_82
timestamp 1655495960
transform -1 0 11999 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_83
timestamp 1655495960
transform 1 0 13195 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_84
timestamp 1655495960
transform -1 0 315 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_85
timestamp 1655495960
transform -1 0 1603 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_86
timestamp 1655495960
transform -1 0 2891 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_87
timestamp 1655495960
transform -1 0 4179 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_88
timestamp 1655495960
transform -1 0 5467 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_89
timestamp 1655495960
transform -1 0 6755 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_90
timestamp 1655495960
transform -1 0 8043 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_91
timestamp 1655495960
transform -1 0 9331 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_92
timestamp 1655495960
transform -1 0 10711 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_93
timestamp 1655495960
transform -1 0 11999 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_94
timestamp 1655495960
transform -1 0 315 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_95
timestamp 1655495960
transform -1 0 1603 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_96
timestamp 1655495960
transform -1 0 2891 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_97
timestamp 1655495960
transform -1 0 4179 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_98
timestamp 1655495960
transform -1 0 5467 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_99
timestamp 1655495960
transform -1 0 6755 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_100
timestamp 1655495960
transform -1 0 8043 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_101
timestamp 1655495960
transform -1 0 9331 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_102
timestamp 1655495960
transform -1 0 10711 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_103
timestamp 1655495960
transform -1 0 11999 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_104
timestamp 1655495960
transform 1 0 13195 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_105
timestamp 1655495960
transform 1 0 -1433 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_106
timestamp 1655495960
transform 1 0 -605 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_107
timestamp 1655495960
transform -1 0 315 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_108
timestamp 1655495960
transform 1 0 591 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_109
timestamp 1655495960
transform 1 0 1419 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_110
timestamp 1655495960
transform -1 0 1603 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_111
timestamp 1655495960
transform 1 0 1879 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_112
timestamp 1655495960
transform -1 0 2891 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_113
timestamp 1655495960
transform 1 0 3167 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_114
timestamp 1655495960
transform -1 0 4179 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_115
timestamp 1655495960
transform -1 0 5467 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_116
timestamp 1655495960
transform 1 0 6387 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_117
timestamp 1655495960
transform -1 0 6755 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_118
timestamp 1655495960
transform 1 0 7675 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_119
timestamp 1655495960
transform -1 0 8043 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_120
timestamp 1655495960
transform 1 0 8963 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_121
timestamp 1655495960
transform -1 0 9331 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_122
timestamp 1655495960
transform 1 0 10251 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_123
timestamp 1655495960
transform -1 0 10711 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_124
timestamp 1655495960
transform 1 0 11631 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_125
timestamp 1655495960
transform -1 0 11999 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_126
timestamp 1655495960
transform 1 0 -1433 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_127
timestamp 1655495960
transform 1 0 591 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_128
timestamp 1655495960
transform 1 0 -605 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_129
timestamp 1655495960
transform 1 0 1419 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_130
timestamp 1655495960
transform 1 0 1879 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_131
timestamp 1655495960
transform 1 0 3167 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_132
timestamp 1655495960
transform 1 0 6387 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_133
timestamp 1655495960
transform 1 0 7675 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_134
timestamp 1655495960
transform 1 0 8963 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_135
timestamp 1655495960
transform 1 0 10251 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_136
timestamp 1655495960
transform 1 0 11631 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_137
timestamp 1655495960
transform -1 0 315 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_138
timestamp 1655495960
transform -1 0 2891 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_139
timestamp 1655495960
transform -1 0 1603 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_140
timestamp 1655495960
transform -1 0 4179 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_141
timestamp 1655495960
transform -1 0 6755 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_142
timestamp 1655495960
transform -1 0 5467 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_143
timestamp 1655495960
transform -1 0 8043 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_144
timestamp 1655495960
transform -1 0 9331 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_145
timestamp 1655495960
transform -1 0 11999 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_146
timestamp 1655495960
transform -1 0 10711 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_147
timestamp 1655495960
transform -1 0 315 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_148
timestamp 1655495960
transform -1 0 2891 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_149
timestamp 1655495960
transform -1 0 1603 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_150
timestamp 1655495960
transform -1 0 4179 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_151
timestamp 1655495960
transform -1 0 6755 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_152
timestamp 1655495960
transform -1 0 5467 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_153
timestamp 1655495960
transform -1 0 8043 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_154
timestamp 1655495960
transform -1 0 9331 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_155
timestamp 1655495960
transform -1 0 11999 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_156
timestamp 1655495960
transform -1 0 10711 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_157
timestamp 1655495960
transform 1 0 13195 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_158
timestamp 1655495960
transform -1 0 315 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_159
timestamp 1655495960
transform -1 0 1603 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_160
timestamp 1655495960
transform -1 0 2891 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_161
timestamp 1655495960
transform -1 0 4179 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_162
timestamp 1655495960
transform -1 0 5467 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_163
timestamp 1655495960
transform -1 0 6755 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_164
timestamp 1655495960
transform -1 0 8043 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_165
timestamp 1655495960
transform -1 0 9331 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_166
timestamp 1655495960
transform -1 0 10711 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_167
timestamp 1655495960
transform -1 0 11999 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_168
timestamp 1655495960
transform -1 0 315 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_169
timestamp 1655495960
transform -1 0 1603 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_170
timestamp 1655495960
transform -1 0 2891 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_171
timestamp 1655495960
transform -1 0 4179 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_172
timestamp 1655495960
transform -1 0 5467 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_173
timestamp 1655495960
transform -1 0 6755 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_174
timestamp 1655495960
transform -1 0 8043 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_175
timestamp 1655495960
transform -1 0 9331 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_176
timestamp 1655495960
transform -1 0 10711 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_177
timestamp 1655495960
transform -1 0 11999 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_178
timestamp 1655495960
transform 1 0 13195 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_179
timestamp 1655495960
transform -1 0 315 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_180
timestamp 1655495960
transform -1 0 315 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_181
timestamp 1655495960
transform -1 0 1603 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_182
timestamp 1655495960
transform -1 0 2891 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_183
timestamp 1655495960
transform -1 0 1603 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_184
timestamp 1655495960
transform -1 0 2891 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_185
timestamp 1655495960
transform -1 0 4179 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_186
timestamp 1655495960
transform -1 0 4179 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_187
timestamp 1655495960
transform -1 0 6755 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_188
timestamp 1655495960
transform -1 0 5467 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_189
timestamp 1655495960
transform -1 0 5467 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_190
timestamp 1655495960
transform -1 0 6755 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_191
timestamp 1655495960
transform -1 0 8043 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_192
timestamp 1655495960
transform -1 0 8043 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_193
timestamp 1655495960
transform -1 0 9331 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_194
timestamp 1655495960
transform -1 0 9331 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_195
timestamp 1655495960
transform -1 0 11999 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_196
timestamp 1655495960
transform -1 0 10711 0 -1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_197
timestamp 1655495960
transform -1 0 10711 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_198
timestamp 1655495960
transform -1 0 11999 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_199
timestamp 1655495960
transform -1 0 315 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_200
timestamp 1655495960
transform -1 0 2891 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_201
timestamp 1655495960
transform -1 0 1603 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_202
timestamp 1655495960
transform -1 0 4179 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_203
timestamp 1655495960
transform -1 0 6755 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_204
timestamp 1655495960
transform -1 0 5467 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_205
timestamp 1655495960
transform -1 0 8043 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_206
timestamp 1655495960
transform -1 0 9331 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_207
timestamp 1655495960
transform -1 0 11999 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_208
timestamp 1655495960
transform -1 0 10711 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_209
timestamp 1655495960
transform 1 0 13195 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_210
timestamp 1655495960
transform -1 0 315 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_211
timestamp 1655495960
transform -1 0 2891 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_212
timestamp 1655495960
transform -1 0 1603 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_213
timestamp 1655495960
transform -1 0 4179 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_214
timestamp 1655495960
transform -1 0 6755 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_215
timestamp 1655495960
transform -1 0 5467 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_216
timestamp 1655495960
transform -1 0 8043 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_217
timestamp 1655495960
transform -1 0 9331 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_218
timestamp 1655495960
transform -1 0 11999 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_219
timestamp 1655495960
transform -1 0 10711 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_220
timestamp 1655495960
transform -1 0 315 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_221
timestamp 1655495960
transform -1 0 1603 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_222
timestamp 1655495960
transform -1 0 2891 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_223
timestamp 1655495960
transform -1 0 4179 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_224
timestamp 1655495960
transform -1 0 5467 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_225
timestamp 1655495960
transform -1 0 6755 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_226
timestamp 1655495960
transform -1 0 8043 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_227
timestamp 1655495960
transform -1 0 9331 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_228
timestamp 1655495960
transform -1 0 10711 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_229
timestamp 1655495960
transform -1 0 11999 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_230
timestamp 1655495960
transform 1 0 13195 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_231
timestamp 1655495960
transform -1 0 315 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_232
timestamp 1655495960
transform -1 0 1603 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_233
timestamp 1655495960
transform -1 0 2891 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_234
timestamp 1655495960
transform -1 0 4179 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_235
timestamp 1655495960
transform -1 0 6755 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_236
timestamp 1655495960
transform -1 0 5467 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_237
timestamp 1655495960
transform -1 0 8043 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_238
timestamp 1655495960
transform -1 0 9331 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_239
timestamp 1655495960
transform -1 0 11999 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_240
timestamp 1655495960
transform -1 0 10711 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_241
timestamp 1655495960
transform 1 0 -1433 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_242
timestamp 1655495960
transform 1 0 591 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_243
timestamp 1655495960
transform 1 0 -605 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_244
timestamp 1655495960
transform 1 0 1419 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_245
timestamp 1655495960
transform 1 0 1879 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_246
timestamp 1655495960
transform 1 0 3167 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_247
timestamp 1655495960
transform 1 0 6387 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_248
timestamp 1655495960
transform 1 0 7675 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_249
timestamp 1655495960
transform 1 0 8963 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_250
timestamp 1655495960
transform 1 0 10251 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_251
timestamp 1655495960
transform 1 0 11631 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_252
timestamp 1655495960
transform -1 0 3627 0 -1 -7084
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_253
timestamp 1655495960
transform -1 0 4455 0 -1 -7084
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_254
timestamp 1655495960
transform -1 0 5835 0 -1 -7084
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_255
timestamp 1655495960
transform -1 0 2615 0 -1 -7084
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform -1 0 -145 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1655495960
transform -1 0 -881 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1655495960
transform 1 0 -1617 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1655495960
transform 1 0 -881 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1655495960
transform -1 0 -881 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1655495960
transform 1 0 -1617 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1655495960
transform 1 0 -881 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1655495960
transform -1 0 -881 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1655495960
transform -1 0 -145 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1655495960
transform 1 0 15955 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1655495960
transform -1 0 16691 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_11
timestamp 1655495960
transform -1 0 -881 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_12
timestamp 1655495960
transform -1 0 -145 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_13
timestamp 1655495960
transform -1 0 16691 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_14
timestamp 1655495960
transform 1 0 -1617 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_15
timestamp 1655495960
transform 1 0 -881 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_16
timestamp 1655495960
transform -1 0 -881 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_17
timestamp 1655495960
transform 1 0 -1617 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_18
timestamp 1655495960
transform 1 0 -881 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_19
timestamp 1655495960
transform -1 0 -881 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_20
timestamp 1655495960
transform -1 0 -145 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_21
timestamp 1655495960
transform 1 0 15955 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_22
timestamp 1655495960
transform 1 0 15955 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_23
timestamp 1655495960
transform -1 0 -881 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_24
timestamp 1655495960
transform -1 0 -145 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_25
timestamp 1655495960
transform 1 0 -1617 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_26
timestamp 1655495960
transform 1 0 -881 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_27
timestamp 1655495960
transform -1 0 -881 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_28
timestamp 1655495960
transform 1 0 -1617 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_29
timestamp 1655495960
transform 1 0 -881 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_30
timestamp 1655495960
transform -1 0 -881 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_31
timestamp 1655495960
transform -1 0 -881 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_32
timestamp 1655495960
transform -1 0 -145 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_33
timestamp 1655495960
transform -1 0 -145 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_34
timestamp 1655495960
transform -1 0 16691 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_35
timestamp 1655495960
transform -1 0 16691 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_36
timestamp 1655495960
transform 1 0 -1617 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_37
timestamp 1655495960
transform 1 0 -881 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_38
timestamp 1655495960
transform -1 0 -881 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_39
timestamp 1655495960
transform 1 0 -1617 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_40
timestamp 1655495960
transform 1 0 -881 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_41
timestamp 1655495960
transform -1 0 -881 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_42
timestamp 1655495960
transform -1 0 -145 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_43
timestamp 1655495960
transform 1 0 15955 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_44
timestamp 1655495960
transform 1 0 -1617 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_45
timestamp 1655495960
transform 1 0 -881 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_46
timestamp 1655495960
transform 1 0 -2997 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_47
timestamp 1655495960
transform -1 0 -145 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_48
timestamp 1655495960
transform 1 0 -53 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_49
timestamp 1655495960
transform 1 0 683 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_50
timestamp 1655495960
transform -1 0 683 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_51
timestamp 1655495960
transform -1 0 1419 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_52
timestamp 1655495960
transform 1 0 7767 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_53
timestamp 1655495960
transform 1 0 1511 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_54
timestamp 1655495960
transform 1 0 8503 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_55
timestamp 1655495960
transform -1 0 2247 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_56
timestamp 1655495960
transform -1 0 2983 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_57
timestamp 1655495960
transform -1 0 4547 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_58
timestamp 1655495960
transform -1 0 3811 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_59
timestamp 1655495960
transform -1 0 6111 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_60
timestamp 1655495960
transform -1 0 5375 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_61
timestamp 1655495960
transform -1 0 6939 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_62
timestamp 1655495960
transform -1 0 7675 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_63
timestamp 1655495960
transform -1 0 8503 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_64
timestamp 1655495960
transform 1 0 15955 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_65
timestamp 1655495960
transform -1 0 9239 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_66
timestamp 1655495960
transform -1 0 16691 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_67
timestamp 1655495960
transform -1 0 -2261 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_68
timestamp 1655495960
transform 1 0 -2997 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_69
timestamp 1655495960
transform -1 0 -2261 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_70
timestamp 1655495960
transform 1 0 -2997 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_71
timestamp 1655495960
transform -1 0 -2261 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_72
timestamp 1655495960
transform 1 0 -2997 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_73
timestamp 1655495960
transform -1 0 -2261 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_74
timestamp 1655495960
transform -1 0 -2261 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_75
timestamp 1655495960
transform 1 0 -2997 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_76
timestamp 1655495960
transform -1 0 -2261 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_77
timestamp 1655495960
transform 1 0 -2997 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_78
timestamp 1655495960
transform -1 0 -2261 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_79
timestamp 1655495960
transform 1 0 -2997 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_80
timestamp 1655495960
transform -1 0 -2261 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_81
timestamp 1655495960
transform 1 0 -2997 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_82
timestamp 1655495960
transform -1 0 -2261 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_83
timestamp 1655495960
transform 1 0 -2997 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_84
timestamp 1655495960
transform -1 0 -2261 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_85
timestamp 1655495960
transform 1 0 -2997 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_86
timestamp 1655495960
transform -1 0 -2261 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_87
timestamp 1655495960
transform 1 0 -2997 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_88
timestamp 1655495960
transform -1 0 -2261 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_89
timestamp 1655495960
transform -1 0 -2261 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_90
timestamp 1655495960
transform 1 0 -2997 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_91
timestamp 1655495960
transform -1 0 2431 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_92
timestamp 1655495960
transform 1 0 1695 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_93
timestamp 1655495960
transform -1 0 2431 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_94
timestamp 1655495960
transform 1 0 1695 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_95
timestamp 1655495960
transform -1 0 2431 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_96
timestamp 1655495960
transform 1 0 1695 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_97
timestamp 1655495960
transform -1 0 2431 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_98
timestamp 1655495960
transform 1 0 1695 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_99
timestamp 1655495960
transform -1 0 2431 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_100
timestamp 1655495960
transform 1 0 1695 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_101
timestamp 1655495960
transform 1 0 4271 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_102
timestamp 1655495960
transform 1 0 4271 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_103
timestamp 1655495960
transform -1 0 5007 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_104
timestamp 1655495960
transform 1 0 4271 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_105
timestamp 1655495960
transform -1 0 5007 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_106
timestamp 1655495960
transform -1 0 5007 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_107
timestamp 1655495960
transform 1 0 4271 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_108
timestamp 1655495960
transform -1 0 5007 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_109
timestamp 1655495960
transform 1 0 4271 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_110
timestamp 1655495960
transform -1 0 5007 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_111
timestamp 1655495960
transform -1 0 7583 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_112
timestamp 1655495960
transform 1 0 6847 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_113
timestamp 1655495960
transform -1 0 7583 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_114
timestamp 1655495960
transform 1 0 6847 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_115
timestamp 1655495960
transform -1 0 7583 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_116
timestamp 1655495960
transform 1 0 6847 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_117
timestamp 1655495960
transform -1 0 7583 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_118
timestamp 1655495960
transform 1 0 6847 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_119
timestamp 1655495960
transform -1 0 7583 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_120
timestamp 1655495960
transform 1 0 6847 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_121
timestamp 1655495960
transform -1 0 10159 0 -1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_122
timestamp 1655495960
transform 1 0 9423 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_123
timestamp 1655495960
transform -1 0 10159 0 -1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_124
timestamp 1655495960
transform 1 0 9423 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_125
timestamp 1655495960
transform -1 0 10159 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_126
timestamp 1655495960
transform 1 0 9423 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_127
timestamp 1655495960
transform -1 0 10159 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_128
timestamp 1655495960
transform 1 0 9423 0 1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_129
timestamp 1655495960
transform -1 0 10159 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_130
timestamp 1655495960
transform 1 0 9423 0 1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_131
timestamp 1655495960
transform -1 0 2431 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_132
timestamp 1655495960
transform 1 0 1695 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_133
timestamp 1655495960
transform -1 0 2431 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_134
timestamp 1655495960
transform 1 0 1695 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_135
timestamp 1655495960
transform -1 0 2431 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_136
timestamp 1655495960
transform 1 0 1695 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_137
timestamp 1655495960
transform -1 0 2431 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_138
timestamp 1655495960
transform 1 0 1695 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_139
timestamp 1655495960
transform -1 0 2431 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_140
timestamp 1655495960
transform 1 0 1695 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_141
timestamp 1655495960
transform -1 0 5007 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_142
timestamp 1655495960
transform 1 0 4271 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_143
timestamp 1655495960
transform -1 0 5007 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_144
timestamp 1655495960
transform 1 0 4271 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_145
timestamp 1655495960
transform -1 0 5007 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_146
timestamp 1655495960
transform 1 0 4271 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_147
timestamp 1655495960
transform -1 0 5007 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_148
timestamp 1655495960
transform 1 0 4271 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_149
timestamp 1655495960
transform -1 0 5007 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_150
timestamp 1655495960
transform 1 0 4271 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_151
timestamp 1655495960
transform -1 0 7583 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_152
timestamp 1655495960
transform 1 0 6847 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_153
timestamp 1655495960
transform -1 0 7583 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_154
timestamp 1655495960
transform 1 0 6847 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_155
timestamp 1655495960
transform -1 0 7583 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_156
timestamp 1655495960
transform 1 0 6847 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_157
timestamp 1655495960
transform -1 0 7583 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_158
timestamp 1655495960
transform 1 0 6847 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_159
timestamp 1655495960
transform 1 0 6847 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_160
timestamp 1655495960
transform -1 0 7583 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_161
timestamp 1655495960
transform 1 0 9423 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_162
timestamp 1655495960
transform -1 0 10159 0 -1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_163
timestamp 1655495960
transform 1 0 9423 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_164
timestamp 1655495960
transform -1 0 10159 0 -1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_165
timestamp 1655495960
transform 1 0 9423 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_166
timestamp 1655495960
transform -1 0 10159 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_167
timestamp 1655495960
transform 1 0 9423 0 1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_168
timestamp 1655495960
transform -1 0 10159 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_169
timestamp 1655495960
transform 1 0 9423 0 1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_170
timestamp 1655495960
transform -1 0 10159 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 4363 0 1 -556
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_1
timestamp 1655495960
transform 1 0 13563 0 1 -556
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_2
timestamp 1655495960
transform 1 0 14759 0 1 -556
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_3
timestamp 1655495960
transform 1 0 15587 0 1 -1644
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_4
timestamp 1655495960
transform -1 0 16691 0 -1 -556
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_5
timestamp 1655495960
transform -1 0 16691 0 -1 -1644
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_6
timestamp 1655495960
transform 1 0 15587 0 1 -2732
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_7
timestamp 1655495960
transform -1 0 14667 0 -1 -2732
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_8
timestamp 1655495960
transform -1 0 15863 0 -1 -2732
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_9
timestamp 1655495960
transform -1 0 14667 0 1 -3820
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_10
timestamp 1655495960
transform -1 0 15863 0 1 -3820
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_11
timestamp 1655495960
transform 1 0 15587 0 -1 -3820
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_12
timestamp 1655495960
transform -1 0 16691 0 1 -4908
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_13
timestamp 1655495960
transform 1 0 15587 0 -1 -4908
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_14
timestamp 1655495960
transform 1 0 4363 0 -1 -5996
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_15
timestamp 1655495960
transform 1 0 13563 0 -1 -5996
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_16
timestamp 1655495960
transform 1 0 14759 0 -1 -5996
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_17
timestamp 1655495960
transform -1 0 16691 0 1 -5996
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_18
timestamp 1655495960
transform 1 0 4363 0 -1 -13612
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_19
timestamp 1655495960
transform 1 0 13563 0 -1 -13612
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_20
timestamp 1655495960
transform 1 0 14759 0 -1 -13612
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_21
timestamp 1655495960
transform -1 0 16691 0 1 -13612
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_22
timestamp 1655495960
transform 1 0 15587 0 -1 -12524
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_23
timestamp 1655495960
transform -1 0 16691 0 1 -12524
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_24
timestamp 1655495960
transform 1 0 15587 0 -1 -11436
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_25
timestamp 1655495960
transform -1 0 14667 0 -1 -10348
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_26
timestamp 1655495960
transform -1 0 14667 0 1 -11436
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_27
timestamp 1655495960
transform -1 0 15863 0 -1 -10348
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_28
timestamp 1655495960
transform -1 0 15863 0 1 -11436
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_29
timestamp 1655495960
transform 1 0 15587 0 1 -10348
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_30
timestamp 1655495960
transform -1 0 16691 0 -1 -9260
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_31
timestamp 1655495960
transform 1 0 15587 0 1 -9260
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_32
timestamp 1655495960
transform -1 0 16691 0 -1 -8172
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_33
timestamp 1655495960
transform 1 0 4363 0 1 -8172
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_34
timestamp 1655495960
transform 1 0 13563 0 1 -8172
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_35
timestamp 1655495960
transform 1 0 14759 0 1 -8172
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform -1 0 7675 0 -1 -7084
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1655495960
transform 1 0 -2629 0 1 -7084
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform -1 0 11631 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1655495960
transform -1 0 10711 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1655495960
transform -1 0 10343 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1655495960
transform -1 0 10343 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1655495960
transform -1 0 10711 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1655495960
transform -1 0 11631 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1655495960
transform -1 0 10343 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1655495960
transform -1 0 10711 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1655495960
transform -1 0 11631 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1655495960
transform -1 0 10343 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1655495960
transform -1 0 10711 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1655495960
transform -1 0 11631 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1655495960
transform -1 0 10343 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1655495960
transform -1 0 10711 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1655495960
transform -1 0 11631 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1655495960
transform -1 0 13563 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1655495960
transform 1 0 5835 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1655495960
transform -1 0 13563 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1655495960
transform -1 0 10343 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1655495960
transform -1 0 10711 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1655495960
transform -1 0 11631 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1655495960
transform -1 0 10343 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1655495960
transform -1 0 10711 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1655495960
transform -1 0 11631 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1655495960
transform -1 0 10343 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1655495960
transform -1 0 10711 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1655495960
transform -1 0 11631 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1655495960
transform -1 0 13563 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1655495960
transform -1 0 10343 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1655495960
transform -1 0 10711 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1655495960
transform -1 0 11631 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1655495960
transform 1 0 5835 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1655495960
transform -1 0 10343 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1655495960
transform -1 0 10711 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1655495960
transform -1 0 11631 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1655495960
transform -1 0 13563 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1655495960
transform 1 0 5835 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_37
timestamp 1655495960
transform -1 0 10343 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_38
timestamp 1655495960
transform -1 0 11631 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_39
timestamp 1655495960
transform -1 0 10711 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_40
timestamp 1655495960
transform -1 0 13563 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_41
timestamp 1655495960
transform -1 0 10343 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_42
timestamp 1655495960
transform -1 0 11631 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_43
timestamp 1655495960
transform -1 0 10711 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_44
timestamp 1655495960
transform -1 0 10343 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_45
timestamp 1655495960
transform -1 0 10711 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_46
timestamp 1655495960
transform -1 0 11631 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_47
timestamp 1655495960
transform -1 0 13563 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_48
timestamp 1655495960
transform -1 0 10343 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_49
timestamp 1655495960
transform -1 0 10711 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_50
timestamp 1655495960
transform -1 0 11631 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_51
timestamp 1655495960
transform -1 0 10343 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_52
timestamp 1655495960
transform -1 0 10343 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_53
timestamp 1655495960
transform -1 0 11631 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_54
timestamp 1655495960
transform -1 0 10711 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_55
timestamp 1655495960
transform -1 0 10711 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_56
timestamp 1655495960
transform -1 0 11631 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_57
timestamp 1655495960
transform -1 0 10343 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_58
timestamp 1655495960
transform -1 0 11631 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_59
timestamp 1655495960
transform -1 0 10711 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_60
timestamp 1655495960
transform -1 0 10343 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_61
timestamp 1655495960
transform -1 0 11631 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_62
timestamp 1655495960
transform -1 0 10711 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_63
timestamp 1655495960
transform -1 0 13563 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_64
timestamp 1655495960
transform -1 0 10343 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_65
timestamp 1655495960
transform -1 0 10711 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_66
timestamp 1655495960
transform -1 0 11631 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_67
timestamp 1655495960
transform -1 0 10343 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_68
timestamp 1655495960
transform -1 0 11631 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_69
timestamp 1655495960
transform -1 0 10711 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_70
timestamp 1655495960
transform -1 0 13563 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_71
timestamp 1655495960
transform 1 0 5835 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform -1 0 -1617 0 -1 -556
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_1
timestamp 1655495960
transform 1 0 -1617 0 -1 -5996
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_2
timestamp 1655495960
transform 1 0 -1617 0 -1 -13612
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_3
timestamp 1655495960
transform 1 0 -1617 0 1 -8172
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_4
timestamp 1655495960
transform -1 0 2799 0 -1 -7084
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_5
timestamp 1655495960
transform 1 0 -1801 0 1 -1644
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_6
timestamp 1655495960
transform 1 0 -1801 0 1 -2732
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_7
timestamp 1655495960
transform -1 0 -1617 0 -1 -1644
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_8
timestamp 1655495960
transform -1 0 -1985 0 -1 -2732
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_9
timestamp 1655495960
transform 1 0 -1801 0 1 -3820
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_10
timestamp 1655495960
transform -1 0 -1617 0 -1 -3820
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_11
timestamp 1655495960
transform -1 0 -1617 0 -1 -4908
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_12
timestamp 1655495960
transform 1 0 -1801 0 1 -4908
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_13
timestamp 1655495960
transform -1 0 -1617 0 -1 -5996
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_14
timestamp 1655495960
transform 1 0 -1801 0 1 -5996
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_15
timestamp 1655495960
transform 1 0 -1617 0 1 -556
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_16
timestamp 1655495960
transform -1 0 -1617 0 1 -556
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_17
timestamp 1655495960
transform -1 0 -1617 0 -1 -7084
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_18
timestamp 1655495960
transform 1 0 -1801 0 1 -8172
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_19
timestamp 1655495960
transform -1 0 -1617 0 -1 -8172
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_20
timestamp 1655495960
transform 1 0 -1801 0 1 -9260
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_21
timestamp 1655495960
transform -1 0 -1617 0 -1 -9260
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_22
timestamp 1655495960
transform 1 0 -1801 0 1 -10348
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_23
timestamp 1655495960
transform -1 0 -1985 0 -1 -10348
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_24
timestamp 1655495960
transform 1 0 -1801 0 1 -11436
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_25
timestamp 1655495960
transform -1 0 -1617 0 -1 -11436
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_26
timestamp 1655495960
transform 1 0 -1801 0 1 -12524
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_27
timestamp 1655495960
transform -1 0 -1617 0 -1 -12524
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_28
timestamp 1655495960
transform -1 0 -1617 0 -1 -13612
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  sky130_fd_sc_hd__fill_2_29
timestamp 1655495960
transform 1 0 -1801 0 1 -13612
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 5927 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_1
timestamp 1655495960
transform 1 0 5467 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_2
timestamp 1655495960
transform 1 0 11999 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_3
timestamp 1655495960
transform 1 0 11999 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_4
timestamp 1655495960
transform 1 0 11999 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_5
timestamp 1655495960
transform 1 0 11999 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_6
timestamp 1655495960
transform 1 0 5927 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_7
timestamp 1655495960
transform 1 0 5467 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_8
timestamp 1655495960
transform 1 0 5467 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_9
timestamp 1655495960
transform 1 0 5927 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_10
timestamp 1655495960
transform 1 0 11999 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_11
timestamp 1655495960
transform 1 0 11999 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_12
timestamp 1655495960
transform 1 0 11999 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_13
timestamp 1655495960
transform 1 0 11999 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_14
timestamp 1655495960
transform 1 0 5927 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_15
timestamp 1655495960
transform 1 0 5467 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_16
timestamp 1655495960
transform 1 0 -2169 0 1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_17
timestamp 1655495960
transform -1 0 -1801 0 -1 -7084
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_18
timestamp 1655495960
transform -1 0 -1801 0 -1 -556
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_19
timestamp 1655495960
transform 1 0 -2169 0 1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_20
timestamp 1655495960
transform -1 0 -1801 0 -1 -1644
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_21
timestamp 1655495960
transform 1 0 -2169 0 1 -2732
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_22
timestamp 1655495960
transform 1 0 -2169 0 1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_23
timestamp 1655495960
transform -1 0 -1801 0 -1 -3820
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_24
timestamp 1655495960
transform -1 0 -1801 0 -1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_25
timestamp 1655495960
transform 1 0 -2169 0 1 -4908
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_26
timestamp 1655495960
transform -1 0 -1801 0 -1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_27
timestamp 1655495960
transform 1 0 -2169 0 1 -5996
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_28
timestamp 1655495960
transform 1 0 -2169 0 1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_29
timestamp 1655495960
transform -1 0 -1801 0 -1 -8172
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_30
timestamp 1655495960
transform 1 0 -2169 0 1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_31
timestamp 1655495960
transform -1 0 -1801 0 -1 -9260
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_32
timestamp 1655495960
transform 1 0 -2169 0 1 -10348
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_33
timestamp 1655495960
transform 1 0 -2169 0 1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_34
timestamp 1655495960
transform -1 0 -1801 0 -1 -11436
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_35
timestamp 1655495960
transform -1 0 -1801 0 -1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_36
timestamp 1655495960
transform 1 0 -2169 0 1 -12524
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_37
timestamp 1655495960
transform -1 0 -1801 0 -1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  sky130_fd_sc_hd__fill_4_38
timestamp 1655495960
transform 1 0 -2169 0 1 -13612
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform -1 0 12735 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1655495960
transform -1 0 13471 0 -1 -1644
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1655495960
transform 1 0 3627 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1655495960
transform -1 0 12735 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1655495960
transform -1 0 13471 0 -1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1655495960
transform 1 0 11999 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_6
timestamp 1655495960
transform 1 0 12735 0 1 -556
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_7
timestamp 1655495960
transform -1 0 13471 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_8
timestamp 1655495960
transform -1 0 12735 0 -1 -2732
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_9
timestamp 1655495960
transform -1 0 12735 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_10
timestamp 1655495960
transform -1 0 13471 0 1 -3820
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_11
timestamp 1655495960
transform -1 0 12735 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_12
timestamp 1655495960
transform -1 0 13471 0 1 -4908
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_13
timestamp 1655495960
transform 1 0 3627 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_14
timestamp 1655495960
transform 1 0 11999 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_15
timestamp 1655495960
transform -1 0 12735 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_16
timestamp 1655495960
transform -1 0 13471 0 1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_17
timestamp 1655495960
transform 1 0 12735 0 -1 -5996
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_18
timestamp 1655495960
transform 1 0 3627 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_19
timestamp 1655495960
transform 1 0 11999 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_20
timestamp 1655495960
transform 1 0 12735 0 -1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_21
timestamp 1655495960
transform -1 0 12735 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_22
timestamp 1655495960
transform -1 0 13471 0 1 -13612
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_23
timestamp 1655495960
transform -1 0 12735 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_24
timestamp 1655495960
transform -1 0 13471 0 1 -12524
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_25
timestamp 1655495960
transform -1 0 12735 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_26
timestamp 1655495960
transform -1 0 12735 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_27
timestamp 1655495960
transform -1 0 13471 0 -1 -10348
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_28
timestamp 1655495960
transform -1 0 13471 0 1 -11436
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_29
timestamp 1655495960
transform -1 0 12735 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_30
timestamp 1655495960
transform -1 0 13471 0 -1 -9260
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_31
timestamp 1655495960
transform -1 0 12735 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_32
timestamp 1655495960
transform -1 0 13471 0 -1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_33
timestamp 1655495960
transform 1 0 3627 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_34
timestamp 1655495960
transform 1 0 11999 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_35
timestamp 1655495960
transform 1 0 12735 0 1 -8172
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_36
timestamp 1655495960
transform 1 0 9331 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_37
timestamp 1655495960
transform -1 0 10067 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_38
timestamp 1655495960
transform -1 0 10803 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_39
timestamp 1655495960
transform 1 0 10067 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_40
timestamp 1655495960
transform -1 0 11539 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_41
timestamp 1655495960
transform -1 0 12275 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_42
timestamp 1655495960
transform 1 0 10803 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_43
timestamp 1655495960
transform 1 0 11539 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_44
timestamp 1655495960
transform -1 0 13011 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_45
timestamp 1655495960
transform -1 0 13747 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_46
timestamp 1655495960
transform 1 0 12275 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_47
timestamp 1655495960
transform 1 0 13011 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_48
timestamp 1655495960
transform -1 0 14483 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_49
timestamp 1655495960
transform -1 0 15219 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_50
timestamp 1655495960
transform 1 0 13747 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_51
timestamp 1655495960
transform 1 0 14483 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_52
timestamp 1655495960
transform 1 0 15219 0 1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_53
timestamp 1655495960
transform -1 0 15955 0 -1 -7084
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  sky130_fd_sc_hd__mux2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 4547 0 -1 -7084
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 -973 0 1 -556
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1655495960
transform 1 0 -973 0 -1 -5996
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_2
timestamp 1655495960
transform 1 0 -973 0 -1 -13612
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_3
timestamp 1655495960
transform 1 0 -973 0 1 -8172
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_4
timestamp 1655495960
transform 1 0 3719 0 -1 -7084
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 10711 0 1 -556
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_1
timestamp 1655495960
transform 1 0 10711 0 -1 -5996
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_2
timestamp 1655495960
transform 1 0 10711 0 -1 -13612
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  sky130_fd_sc_hd__nand2_4_3
timestamp 1655495960
transform 1 0 10711 0 1 -8172
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1655495960
transform 1 0 -1065 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1655495960
transform 1 0 -697 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1655495960
transform 1 0 -237 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1655495960
transform 1 0 3535 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1655495960
transform 1 0 499 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1655495960
transform 1 0 959 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1655495960
transform 1 0 1327 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1655495960
transform 1 0 1787 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1655495960
transform 1 0 2247 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1655495960
transform 1 0 6295 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1655495960
transform 1 0 6755 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1655495960
transform 1 0 7583 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1655495960
transform 1 0 8043 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1655495960
transform 1 0 8871 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1655495960
transform 1 0 9331 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1655495960
transform 1 0 10159 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1655495960
transform 1 0 10619 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1655495960
transform 1 0 11539 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1655495960
transform -1 0 11539 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1655495960
transform -1 0 10251 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1655495960
transform -1 0 9423 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1655495960
transform -1 0 8963 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1655495960
transform -1 0 8135 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1655495960
transform -1 0 7675 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1655495960
transform -1 0 6847 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1655495960
transform -1 0 6387 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1655495960
transform -1 0 5559 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1655495960
transform -1 0 5099 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1655495960
transform -1 0 4271 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1655495960
transform -1 0 3811 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1655495960
transform -1 0 2983 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1655495960
transform -1 0 2523 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1655495960
transform -1 0 2523 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1655495960
transform -1 0 2983 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1655495960
transform -1 0 3811 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1655495960
transform -1 0 4271 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1655495960
transform -1 0 5099 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1655495960
transform -1 0 5559 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1655495960
transform -1 0 6387 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1655495960
transform -1 0 6847 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1655495960
transform -1 0 7675 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1655495960
transform -1 0 8135 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1655495960
transform -1 0 8963 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1655495960
transform -1 0 9423 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1655495960
transform -1 0 10251 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1655495960
transform -1 0 11539 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1655495960
transform -1 0 2523 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1655495960
transform -1 0 2983 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1655495960
transform -1 0 3811 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1655495960
transform -1 0 4271 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1655495960
transform -1 0 5559 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1655495960
transform -1 0 5099 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1655495960
transform -1 0 6387 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1655495960
transform -1 0 6847 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1655495960
transform -1 0 7675 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1655495960
transform -1 0 8135 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1655495960
transform -1 0 8963 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1655495960
transform -1 0 9423 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1655495960
transform -1 0 10251 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1655495960
transform -1 0 11539 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1655495960
transform -1 0 2523 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1655495960
transform -1 0 2983 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1655495960
transform -1 0 3811 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1655495960
transform -1 0 4271 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1655495960
transform -1 0 5099 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1655495960
transform -1 0 5559 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1655495960
transform -1 0 6387 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1655495960
transform -1 0 6847 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1655495960
transform -1 0 7675 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1655495960
transform -1 0 8135 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1655495960
transform -1 0 8963 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1655495960
transform -1 0 9423 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1655495960
transform -1 0 10251 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1655495960
transform -1 0 11539 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1655495960
transform -1 0 2523 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1655495960
transform -1 0 2983 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1655495960
transform -1 0 3811 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1655495960
transform -1 0 4271 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1655495960
transform -1 0 5559 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1655495960
transform -1 0 5099 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1655495960
transform -1 0 6387 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1655495960
transform -1 0 6847 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1655495960
transform -1 0 7675 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_83
timestamp 1655495960
transform -1 0 8135 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1655495960
transform -1 0 8963 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1655495960
transform -1 0 9423 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1655495960
transform -1 0 10251 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1655495960
transform -1 0 11539 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1655495960
transform -1 0 1235 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1655495960
transform -1 0 407 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_90
timestamp 1655495960
transform -1 0 -53 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_91
timestamp 1655495960
transform -1 0 1695 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_92
timestamp 1655495960
transform -1 0 1235 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_93
timestamp 1655495960
transform -1 0 1695 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_94
timestamp 1655495960
transform -1 0 407 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_95
timestamp 1655495960
transform -1 0 -53 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_96
timestamp 1655495960
transform -1 0 1235 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_97
timestamp 1655495960
transform -1 0 1695 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_98
timestamp 1655495960
transform -1 0 407 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_99
timestamp 1655495960
transform -1 0 -53 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_100
timestamp 1655495960
transform -1 0 1235 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_101
timestamp 1655495960
transform -1 0 1695 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_102
timestamp 1655495960
transform -1 0 1235 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_103
timestamp 1655495960
transform -1 0 1695 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_104
timestamp 1655495960
transform -1 0 407 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_105
timestamp 1655495960
transform -1 0 407 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_106
timestamp 1655495960
transform -1 0 -53 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_107
timestamp 1655495960
transform -1 0 -53 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_108
timestamp 1655495960
transform 1 0 3075 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_109
timestamp 1655495960
transform -1 0 -53 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_110
timestamp 1655495960
transform -1 0 407 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_111
timestamp 1655495960
transform 1 0 13103 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_112
timestamp 1655495960
transform 1 0 13563 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_113
timestamp 1655495960
transform 1 0 12367 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_114
timestamp 1655495960
transform 1 0 12367 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_115
timestamp 1655495960
transform 1 0 13103 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_116
timestamp 1655495960
transform 1 0 13563 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_117
timestamp 1655495960
transform -1 0 13655 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_118
timestamp 1655495960
transform -1 0 13655 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_119
timestamp 1655495960
transform 1 0 13471 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_120
timestamp 1655495960
transform 1 0 14667 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_121
timestamp 1655495960
transform 1 0 15863 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_122
timestamp 1655495960
transform -1 0 1235 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_123
timestamp 1655495960
transform 1 0 15495 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_124
timestamp 1655495960
transform -1 0 1695 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_125
timestamp 1655495960
transform -1 0 15587 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_126
timestamp 1655495960
transform -1 0 2523 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_127
timestamp 1655495960
transform -1 0 2983 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_128
timestamp 1655495960
transform -1 0 15587 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_129
timestamp 1655495960
transform -1 0 3811 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_130
timestamp 1655495960
transform 1 0 15495 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_131
timestamp 1655495960
transform -1 0 13563 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_132
timestamp 1655495960
transform -1 0 14759 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_133
timestamp 1655495960
transform -1 0 15955 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_134
timestamp 1655495960
transform -1 0 4271 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_135
timestamp 1655495960
transform -1 0 5099 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_136
timestamp 1655495960
transform -1 0 5559 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_137
timestamp 1655495960
transform -1 0 6387 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_138
timestamp 1655495960
transform -1 0 6847 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_139
timestamp 1655495960
transform -1 0 7675 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_140
timestamp 1655495960
transform -1 0 8135 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_141
timestamp 1655495960
transform -1 0 9423 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_142
timestamp 1655495960
transform -1 0 8963 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_143
timestamp 1655495960
transform -1 0 10251 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_144
timestamp 1655495960
transform -1 0 11539 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_145
timestamp 1655495960
transform -1 0 13563 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_146
timestamp 1655495960
transform -1 0 14759 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_147
timestamp 1655495960
transform -1 0 15955 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_148
timestamp 1655495960
transform -1 0 -53 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_149
timestamp 1655495960
transform -1 0 407 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_150
timestamp 1655495960
transform -1 0 1235 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_151
timestamp 1655495960
transform -1 0 1695 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_152
timestamp 1655495960
transform -1 0 2523 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_153
timestamp 1655495960
transform -1 0 2983 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_154
timestamp 1655495960
transform -1 0 3811 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_155
timestamp 1655495960
transform -1 0 4271 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_156
timestamp 1655495960
transform -1 0 5099 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_157
timestamp 1655495960
transform -1 0 5559 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_158
timestamp 1655495960
transform -1 0 6387 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_159
timestamp 1655495960
transform -1 0 6847 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_160
timestamp 1655495960
transform -1 0 7675 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_161
timestamp 1655495960
transform -1 0 8135 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_162
timestamp 1655495960
transform -1 0 9423 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_163
timestamp 1655495960
transform -1 0 8963 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_164
timestamp 1655495960
transform -1 0 10251 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_165
timestamp 1655495960
transform -1 0 11539 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_166
timestamp 1655495960
transform 1 0 12367 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_167
timestamp 1655495960
transform 1 0 13563 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_168
timestamp 1655495960
transform 1 0 13103 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_169
timestamp 1655495960
transform 1 0 15495 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_170
timestamp 1655495960
transform -1 0 -53 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_171
timestamp 1655495960
transform -1 0 407 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_172
timestamp 1655495960
transform -1 0 1235 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_173
timestamp 1655495960
transform -1 0 1695 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_174
timestamp 1655495960
transform -1 0 2523 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_175
timestamp 1655495960
transform -1 0 2983 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_176
timestamp 1655495960
transform -1 0 3811 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_177
timestamp 1655495960
transform -1 0 4271 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_178
timestamp 1655495960
transform -1 0 5099 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_179
timestamp 1655495960
transform -1 0 5559 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_180
timestamp 1655495960
transform -1 0 6387 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_181
timestamp 1655495960
transform -1 0 6847 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_182
timestamp 1655495960
transform -1 0 7675 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_183
timestamp 1655495960
transform -1 0 8135 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_184
timestamp 1655495960
transform -1 0 9423 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_185
timestamp 1655495960
transform -1 0 8963 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_186
timestamp 1655495960
transform -1 0 10251 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_187
timestamp 1655495960
transform -1 0 11539 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_188
timestamp 1655495960
transform -1 0 13655 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_189
timestamp 1655495960
transform -1 0 15587 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_190
timestamp 1655495960
transform -1 0 -53 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_191
timestamp 1655495960
transform -1 0 407 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_192
timestamp 1655495960
transform -1 0 1235 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_193
timestamp 1655495960
transform -1 0 1695 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_194
timestamp 1655495960
transform -1 0 2523 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_195
timestamp 1655495960
transform -1 0 3811 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_196
timestamp 1655495960
transform -1 0 2983 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_197
timestamp 1655495960
transform -1 0 4271 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_198
timestamp 1655495960
transform -1 0 5099 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_199
timestamp 1655495960
transform -1 0 5559 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_200
timestamp 1655495960
transform -1 0 6387 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_201
timestamp 1655495960
transform -1 0 6847 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_202
timestamp 1655495960
transform -1 0 7675 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_203
timestamp 1655495960
transform -1 0 8135 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_204
timestamp 1655495960
transform -1 0 9423 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_205
timestamp 1655495960
transform -1 0 8963 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_206
timestamp 1655495960
transform -1 0 10251 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_207
timestamp 1655495960
transform -1 0 11539 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_208
timestamp 1655495960
transform 1 0 12367 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_209
timestamp 1655495960
transform 1 0 13563 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_210
timestamp 1655495960
transform 1 0 13103 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_211
timestamp 1655495960
transform 1 0 15495 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_212
timestamp 1655495960
transform 1 0 -1065 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_213
timestamp 1655495960
transform 1 0 -697 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_214
timestamp 1655495960
transform -1 0 -53 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_215
timestamp 1655495960
transform -1 0 407 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_216
timestamp 1655495960
transform 1 0 -237 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_217
timestamp 1655495960
transform 1 0 499 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_218
timestamp 1655495960
transform 1 0 1327 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_219
timestamp 1655495960
transform 1 0 959 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_220
timestamp 1655495960
transform -1 0 1235 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_221
timestamp 1655495960
transform 1 0 2247 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_222
timestamp 1655495960
transform 1 0 1787 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_223
timestamp 1655495960
transform -1 0 1695 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_224
timestamp 1655495960
transform -1 0 2523 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_225
timestamp 1655495960
transform 1 0 3075 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_226
timestamp 1655495960
transform 1 0 3535 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_227
timestamp 1655495960
transform -1 0 2983 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_228
timestamp 1655495960
transform -1 0 4271 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_229
timestamp 1655495960
transform -1 0 3811 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_230
timestamp 1655495960
transform -1 0 5099 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_231
timestamp 1655495960
transform -1 0 5559 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_232
timestamp 1655495960
transform 1 0 6295 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_233
timestamp 1655495960
transform -1 0 6387 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_234
timestamp 1655495960
transform 1 0 6755 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_235
timestamp 1655495960
transform -1 0 6847 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_236
timestamp 1655495960
transform 1 0 8043 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_237
timestamp 1655495960
transform 1 0 7583 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_238
timestamp 1655495960
transform -1 0 8135 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_239
timestamp 1655495960
transform -1 0 7675 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_240
timestamp 1655495960
transform 1 0 8871 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_241
timestamp 1655495960
transform -1 0 8963 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_242
timestamp 1655495960
transform 1 0 9331 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_243
timestamp 1655495960
transform -1 0 9423 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_244
timestamp 1655495960
transform 1 0 10159 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_245
timestamp 1655495960
transform -1 0 10251 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_246
timestamp 1655495960
transform 1 0 10619 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_247
timestamp 1655495960
transform 1 0 11539 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_248
timestamp 1655495960
transform -1 0 11539 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_249
timestamp 1655495960
transform -1 0 13655 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_250
timestamp 1655495960
transform 1 0 13471 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_251
timestamp 1655495960
transform 1 0 14667 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_252
timestamp 1655495960
transform -1 0 15587 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_253
timestamp 1655495960
transform 1 0 15863 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_254
timestamp 1655495960
transform 1 0 -237 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_255
timestamp 1655495960
transform 1 0 499 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_256
timestamp 1655495960
transform 1 0 -697 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_257
timestamp 1655495960
transform 1 0 -1065 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_258
timestamp 1655495960
transform 1 0 959 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_259
timestamp 1655495960
transform 1 0 1327 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_260
timestamp 1655495960
transform 1 0 1787 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_261
timestamp 1655495960
transform 1 0 2247 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_262
timestamp 1655495960
transform 1 0 3535 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_263
timestamp 1655495960
transform 1 0 3075 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_264
timestamp 1655495960
transform 1 0 6295 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_265
timestamp 1655495960
transform 1 0 6755 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_266
timestamp 1655495960
transform 1 0 8043 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_267
timestamp 1655495960
transform 1 0 7583 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_268
timestamp 1655495960
transform 1 0 8871 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_269
timestamp 1655495960
transform 1 0 9331 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_270
timestamp 1655495960
transform 1 0 10159 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_271
timestamp 1655495960
transform 1 0 11539 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_272
timestamp 1655495960
transform 1 0 10619 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_273
timestamp 1655495960
transform 1 0 13471 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_274
timestamp 1655495960
transform 1 0 14667 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_275
timestamp 1655495960
transform 1 0 15863 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_276
timestamp 1655495960
transform -1 0 407 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_277
timestamp 1655495960
transform -1 0 -53 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_278
timestamp 1655495960
transform -1 0 2523 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_279
timestamp 1655495960
transform -1 0 1695 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_280
timestamp 1655495960
transform -1 0 1235 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_281
timestamp 1655495960
transform -1 0 3811 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_282
timestamp 1655495960
transform -1 0 4271 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_283
timestamp 1655495960
transform -1 0 2983 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_284
timestamp 1655495960
transform -1 0 6387 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_285
timestamp 1655495960
transform -1 0 5559 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_286
timestamp 1655495960
transform -1 0 5099 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_287
timestamp 1655495960
transform -1 0 7675 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_288
timestamp 1655495960
transform -1 0 8135 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_289
timestamp 1655495960
transform -1 0 6847 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_290
timestamp 1655495960
transform -1 0 10251 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_291
timestamp 1655495960
transform -1 0 9423 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_292
timestamp 1655495960
transform -1 0 8963 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_293
timestamp 1655495960
transform -1 0 11539 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_294
timestamp 1655495960
transform -1 0 13655 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_295
timestamp 1655495960
transform -1 0 15587 0 1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_296
timestamp 1655495960
transform -1 0 407 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_297
timestamp 1655495960
transform -1 0 -53 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_298
timestamp 1655495960
transform -1 0 2523 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_299
timestamp 1655495960
transform -1 0 1695 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_300
timestamp 1655495960
transform -1 0 1235 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_301
timestamp 1655495960
transform -1 0 3811 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_302
timestamp 1655495960
transform -1 0 4271 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_303
timestamp 1655495960
transform -1 0 2983 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_304
timestamp 1655495960
transform -1 0 6387 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_305
timestamp 1655495960
transform -1 0 5559 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_306
timestamp 1655495960
transform -1 0 5099 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_307
timestamp 1655495960
transform -1 0 7675 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_308
timestamp 1655495960
transform -1 0 8135 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_309
timestamp 1655495960
transform -1 0 6847 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_310
timestamp 1655495960
transform -1 0 10251 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_311
timestamp 1655495960
transform -1 0 9423 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_312
timestamp 1655495960
transform -1 0 8963 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_313
timestamp 1655495960
transform -1 0 11539 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_314
timestamp 1655495960
transform 1 0 13563 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_315
timestamp 1655495960
transform 1 0 13103 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_316
timestamp 1655495960
transform 1 0 12367 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_317
timestamp 1655495960
transform 1 0 15495 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_318
timestamp 1655495960
transform -1 0 -53 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_319
timestamp 1655495960
transform -1 0 407 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_320
timestamp 1655495960
transform -1 0 1235 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_321
timestamp 1655495960
transform -1 0 1695 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_322
timestamp 1655495960
transform -1 0 2523 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_323
timestamp 1655495960
transform -1 0 2983 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_324
timestamp 1655495960
transform -1 0 4271 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_325
timestamp 1655495960
transform -1 0 3811 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_326
timestamp 1655495960
transform -1 0 5099 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_327
timestamp 1655495960
transform -1 0 5559 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_328
timestamp 1655495960
transform -1 0 6387 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_329
timestamp 1655495960
transform -1 0 6847 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_330
timestamp 1655495960
transform -1 0 8135 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_331
timestamp 1655495960
transform -1 0 7675 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_332
timestamp 1655495960
transform -1 0 8963 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_333
timestamp 1655495960
transform -1 0 9423 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_334
timestamp 1655495960
transform -1 0 10251 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_335
timestamp 1655495960
transform -1 0 11539 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_336
timestamp 1655495960
transform -1 0 13655 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_337
timestamp 1655495960
transform -1 0 15587 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_338
timestamp 1655495960
transform -1 0 407 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_339
timestamp 1655495960
transform -1 0 -53 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_340
timestamp 1655495960
transform -1 0 1235 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_341
timestamp 1655495960
transform -1 0 1695 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_342
timestamp 1655495960
transform -1 0 2523 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_343
timestamp 1655495960
transform -1 0 2983 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_344
timestamp 1655495960
transform -1 0 3811 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_345
timestamp 1655495960
transform -1 0 4271 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_346
timestamp 1655495960
transform -1 0 5099 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_347
timestamp 1655495960
transform -1 0 5559 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_348
timestamp 1655495960
transform -1 0 6387 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_349
timestamp 1655495960
transform -1 0 6847 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_350
timestamp 1655495960
transform -1 0 7675 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_351
timestamp 1655495960
transform -1 0 8135 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_352
timestamp 1655495960
transform -1 0 8963 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_353
timestamp 1655495960
transform -1 0 9423 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_354
timestamp 1655495960
transform -1 0 10251 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_355
timestamp 1655495960
transform -1 0 11539 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_356
timestamp 1655495960
transform 1 0 12367 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_357
timestamp 1655495960
transform 1 0 13563 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_358
timestamp 1655495960
transform 1 0 13103 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_359
timestamp 1655495960
transform 1 0 15495 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_360
timestamp 1655495960
transform -1 0 407 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_361
timestamp 1655495960
transform -1 0 -53 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_362
timestamp 1655495960
transform -1 0 407 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_363
timestamp 1655495960
transform -1 0 -53 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_364
timestamp 1655495960
transform -1 0 1695 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_365
timestamp 1655495960
transform -1 0 1235 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_366
timestamp 1655495960
transform -1 0 2523 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_367
timestamp 1655495960
transform -1 0 1235 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_368
timestamp 1655495960
transform -1 0 1695 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_369
timestamp 1655495960
transform -1 0 2523 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_370
timestamp 1655495960
transform -1 0 4271 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_371
timestamp 1655495960
transform -1 0 3811 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_372
timestamp 1655495960
transform -1 0 2983 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_373
timestamp 1655495960
transform -1 0 2983 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_374
timestamp 1655495960
transform -1 0 3811 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_375
timestamp 1655495960
transform -1 0 4271 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_376
timestamp 1655495960
transform -1 0 6387 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_377
timestamp 1655495960
transform -1 0 5559 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_378
timestamp 1655495960
transform -1 0 5099 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_379
timestamp 1655495960
transform -1 0 5099 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_380
timestamp 1655495960
transform -1 0 5559 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_381
timestamp 1655495960
transform -1 0 6387 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_382
timestamp 1655495960
transform -1 0 6847 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_383
timestamp 1655495960
transform -1 0 8135 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_384
timestamp 1655495960
transform -1 0 7675 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_385
timestamp 1655495960
transform -1 0 6847 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_386
timestamp 1655495960
transform -1 0 7675 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_387
timestamp 1655495960
transform -1 0 8135 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_388
timestamp 1655495960
transform -1 0 8963 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_389
timestamp 1655495960
transform -1 0 9423 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_390
timestamp 1655495960
transform -1 0 10251 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_391
timestamp 1655495960
transform -1 0 8963 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_392
timestamp 1655495960
transform -1 0 9423 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_393
timestamp 1655495960
transform -1 0 10251 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_394
timestamp 1655495960
transform -1 0 11539 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_395
timestamp 1655495960
transform -1 0 11539 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_396
timestamp 1655495960
transform -1 0 13563 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_397
timestamp 1655495960
transform -1 0 13563 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_398
timestamp 1655495960
transform -1 0 14759 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_399
timestamp 1655495960
transform -1 0 15955 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_400
timestamp 1655495960
transform -1 0 14759 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_401
timestamp 1655495960
transform -1 0 15955 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_402
timestamp 1655495960
transform -1 0 -53 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_403
timestamp 1655495960
transform -1 0 407 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_404
timestamp 1655495960
transform -1 0 2523 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_405
timestamp 1655495960
transform -1 0 1695 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_406
timestamp 1655495960
transform -1 0 1235 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_407
timestamp 1655495960
transform -1 0 3811 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_408
timestamp 1655495960
transform -1 0 4271 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_409
timestamp 1655495960
transform -1 0 2983 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_410
timestamp 1655495960
transform -1 0 6387 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_411
timestamp 1655495960
transform -1 0 5559 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_412
timestamp 1655495960
transform -1 0 5099 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_413
timestamp 1655495960
transform -1 0 7675 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_414
timestamp 1655495960
transform -1 0 8135 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_415
timestamp 1655495960
transform -1 0 6847 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_416
timestamp 1655495960
transform -1 0 10251 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_417
timestamp 1655495960
transform -1 0 9423 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_418
timestamp 1655495960
transform -1 0 8963 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_419
timestamp 1655495960
transform -1 0 11539 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_420
timestamp 1655495960
transform 1 0 13563 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_421
timestamp 1655495960
transform 1 0 13103 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_422
timestamp 1655495960
transform 1 0 12367 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_423
timestamp 1655495960
transform 1 0 15495 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_424
timestamp 1655495960
transform -1 0 -53 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_425
timestamp 1655495960
transform -1 0 407 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_426
timestamp 1655495960
transform -1 0 2523 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_427
timestamp 1655495960
transform -1 0 1695 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_428
timestamp 1655495960
transform -1 0 1235 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_429
timestamp 1655495960
transform -1 0 3811 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_430
timestamp 1655495960
transform -1 0 4271 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_431
timestamp 1655495960
transform -1 0 2983 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_432
timestamp 1655495960
transform -1 0 6387 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_433
timestamp 1655495960
transform -1 0 5559 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_434
timestamp 1655495960
transform -1 0 5099 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_435
timestamp 1655495960
transform -1 0 7675 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_436
timestamp 1655495960
transform -1 0 8135 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_437
timestamp 1655495960
transform -1 0 6847 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_438
timestamp 1655495960
transform -1 0 10251 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_439
timestamp 1655495960
transform -1 0 9423 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_440
timestamp 1655495960
transform -1 0 8963 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_441
timestamp 1655495960
transform -1 0 11539 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_442
timestamp 1655495960
transform -1 0 13655 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_443
timestamp 1655495960
transform -1 0 15587 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_444
timestamp 1655495960
transform -1 0 407 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_445
timestamp 1655495960
transform -1 0 -53 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_446
timestamp 1655495960
transform -1 0 1235 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_447
timestamp 1655495960
transform -1 0 1695 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_448
timestamp 1655495960
transform -1 0 2523 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_449
timestamp 1655495960
transform -1 0 2983 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_450
timestamp 1655495960
transform -1 0 4271 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_451
timestamp 1655495960
transform -1 0 3811 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_452
timestamp 1655495960
transform -1 0 5099 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_453
timestamp 1655495960
transform -1 0 5559 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_454
timestamp 1655495960
transform -1 0 6387 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_455
timestamp 1655495960
transform -1 0 6847 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_456
timestamp 1655495960
transform -1 0 8135 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_457
timestamp 1655495960
transform -1 0 7675 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_458
timestamp 1655495960
transform -1 0 8963 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_459
timestamp 1655495960
transform -1 0 9423 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_460
timestamp 1655495960
transform -1 0 10251 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_461
timestamp 1655495960
transform -1 0 11539 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_462
timestamp 1655495960
transform 1 0 12367 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_463
timestamp 1655495960
transform 1 0 13103 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_464
timestamp 1655495960
transform 1 0 13563 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_465
timestamp 1655495960
transform 1 0 15495 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_466
timestamp 1655495960
transform -1 0 407 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_467
timestamp 1655495960
transform -1 0 -53 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_468
timestamp 1655495960
transform -1 0 1695 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_469
timestamp 1655495960
transform -1 0 1235 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_470
timestamp 1655495960
transform -1 0 2523 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_471
timestamp 1655495960
transform -1 0 4271 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_472
timestamp 1655495960
transform -1 0 2983 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_473
timestamp 1655495960
transform -1 0 3811 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_474
timestamp 1655495960
transform -1 0 6387 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_475
timestamp 1655495960
transform -1 0 5559 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_476
timestamp 1655495960
transform -1 0 5099 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_477
timestamp 1655495960
transform -1 0 6847 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_478
timestamp 1655495960
transform -1 0 8135 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_479
timestamp 1655495960
transform -1 0 7675 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_480
timestamp 1655495960
transform -1 0 8963 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_481
timestamp 1655495960
transform -1 0 9423 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_482
timestamp 1655495960
transform -1 0 10251 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_483
timestamp 1655495960
transform -1 0 11539 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_484
timestamp 1655495960
transform -1 0 13655 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_485
timestamp 1655495960
transform -1 0 15587 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_486
timestamp 1655495960
transform 1 0 499 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_487
timestamp 1655495960
transform 1 0 -237 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_488
timestamp 1655495960
transform 1 0 -697 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_489
timestamp 1655495960
transform 1 0 -1065 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_490
timestamp 1655495960
transform 1 0 1327 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_491
timestamp 1655495960
transform 1 0 959 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_492
timestamp 1655495960
transform 1 0 2247 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_493
timestamp 1655495960
transform 1 0 1787 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_494
timestamp 1655495960
transform 1 0 3075 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_495
timestamp 1655495960
transform 1 0 3535 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_496
timestamp 1655495960
transform 1 0 6295 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_497
timestamp 1655495960
transform 1 0 6755 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_498
timestamp 1655495960
transform 1 0 8043 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_499
timestamp 1655495960
transform 1 0 7583 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_500
timestamp 1655495960
transform 1 0 8871 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_501
timestamp 1655495960
transform 1 0 9331 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_502
timestamp 1655495960
transform 1 0 10159 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_503
timestamp 1655495960
transform 1 0 11539 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_504
timestamp 1655495960
transform 1 0 10619 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_505
timestamp 1655495960
transform 1 0 13471 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_506
timestamp 1655495960
transform 1 0 14667 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_507
timestamp 1655495960
transform 1 0 15863 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_508
timestamp 1655495960
transform 1 0 3167 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_509
timestamp 1655495960
transform 1 0 3627 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_510
timestamp 1655495960
transform 1 0 3995 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_511
timestamp 1655495960
transform 1 0 4455 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_512
timestamp 1655495960
transform 1 0 5375 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_513
timestamp 1655495960
transform 1 0 5835 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_514
timestamp 1655495960
transform 1 0 -145 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_515
timestamp 1655495960
transform -1 0 -53 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_516
timestamp 1655495960
transform 1 0 1419 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_517
timestamp 1655495960
transform -1 0 1511 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_518
timestamp 1655495960
transform 1 0 7675 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_519
timestamp 1655495960
transform -1 0 2891 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_520
timestamp 1655495960
transform 1 0 9239 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_521
timestamp 1655495960
transform -1 0 15955 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_522
timestamp 1655495960
transform -1 0 -1617 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_523
timestamp 1655495960
transform -1 0 -2629 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_524
timestamp 1655495960
transform 1 0 15863 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_525
timestamp 1655495960
transform -1 0 -1617 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_526
timestamp 1655495960
transform -1 0 3075 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_527
timestamp 1655495960
transform -1 0 4639 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_528
timestamp 1655495960
transform -1 0 6203 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_529
timestamp 1655495960
transform -1 0 7767 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_530
timestamp 1655495960
transform -1 0 9331 0 1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_531
timestamp 1655495960
transform 1 0 -2261 0 1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_532
timestamp 1655495960
transform -1 0 -2169 0 -1 -556
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_533
timestamp 1655495960
transform 1 0 -2261 0 1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_534
timestamp 1655495960
transform -1 0 -2169 0 -1 -1644
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_535
timestamp 1655495960
transform 1 0 -2261 0 1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_536
timestamp 1655495960
transform -1 0 -2169 0 -1 -2732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_537
timestamp 1655495960
transform 1 0 -2261 0 1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_538
timestamp 1655495960
transform -1 0 -2169 0 -1 -3820
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_539
timestamp 1655495960
transform -1 0 -2169 0 -1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_540
timestamp 1655495960
transform 1 0 -2261 0 1 -4908
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_541
timestamp 1655495960
transform -1 0 -2169 0 -1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_542
timestamp 1655495960
transform 1 0 -2261 0 1 -5996
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_543
timestamp 1655495960
transform -1 0 -2169 0 -1 -7084
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_544
timestamp 1655495960
transform 1 0 -2261 0 1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_545
timestamp 1655495960
transform -1 0 -2169 0 -1 -8172
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_546
timestamp 1655495960
transform 1 0 -2261 0 1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_547
timestamp 1655495960
transform -1 0 -2169 0 -1 -9260
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_548
timestamp 1655495960
transform 1 0 -2261 0 1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_549
timestamp 1655495960
transform -1 0 -2169 0 -1 -10348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_550
timestamp 1655495960
transform 1 0 -2261 0 1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_551
timestamp 1655495960
transform -1 0 -2169 0 -1 -11436
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_552
timestamp 1655495960
transform 1 0 -2261 0 1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_553
timestamp 1655495960
transform -1 0 -2169 0 -1 -12524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_554
timestamp 1655495960
transform -1 0 -2169 0 -1 -13612
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_555
timestamp 1655495960
transform 1 0 -2261 0 1 -13612
box -38 -48 130 592
<< labels >>
flabel metal1 -3181 -6847 -3181 -6847 1 FreeSans 400 0 0 0 clk
port 1 n
flabel metal1 16932 -828 16932 -828 1 FreeSans 400 0 0 0 B
port 17 n
flabel metal1 16932 -1372 16932 -1372 1 FreeSans 400 0 0 0 B_b
port 16 n
flabel metal1 16932 -1916 16932 -1916 1 FreeSans 400 0 0 0 Bd
port 15 n
flabel metal1 16932 -2460 16932 -2460 1 FreeSans 400 0 0 0 Bd_b
port 14 n
flabel metal1 16932 -4092 16932 -4092 1 FreeSans 400 0 0 0 Ad_b
port 10 n
flabel metal1 16932 -4636 16932 -4636 1 FreeSans 400 0 0 0 Ad
port 11 n
flabel metal1 16932 -5180 16932 -5180 1 FreeSans 400 0 0 0 A_b
port 12 n
flabel metal1 16932 -5724 16932 -5724 1 FreeSans 400 0 0 0 A
port 13 n
flabel metal1 16932 -8444 16932 -8444 1 FreeSans 400 0 0 0 p2
port 5 n
flabel metal1 16932 -8988 16932 -8988 1 FreeSans 400 0 0 0 p2_b
port 4 n
flabel metal1 16932 -9532 16932 -9532 1 FreeSans 400 0 0 0 p2d
port 3 n
flabel metal1 16932 -10076 16932 -10076 1 FreeSans 400 0 0 0 p2d_b
port 2 n
flabel metal1 16932 -11708 16932 -11708 1 FreeSans 400 0 0 0 p1d_b
port 6 n
flabel metal1 16932 -12252 16932 -12252 1 FreeSans 400 0 0 0 p1d
port 7 n
flabel metal1 16932 -12796 16932 -12796 1 FreeSans 400 0 0 0 p1_b
port 8 n
flabel metal1 16932 -13340 16932 -13340 1 FreeSans 400 0 0 0 p1
port 9 n
flabel locali -3248 -12 -3248 -12 1 FreeSans 400 0 0 0 VDD
port 18 n power bidirectional
flabel locali 16943 -11 16943 -11 1 FreeSans 400 0 0 0 VSS
port 19 n power bidirectional
<< end >>
