magic
tech sky130A
magscale 1 2
timestamp 1655495960
<< error_s >>
rect 257 359 315 365
rect 677 359 735 365
rect 1097 359 1155 365
rect 1517 359 1575 365
rect 1937 359 1995 365
rect 2357 359 2415 365
rect 2777 359 2835 365
rect 3197 359 3255 365
rect 3617 359 3675 365
rect 4037 359 4095 365
rect 4457 359 4515 365
rect 4877 359 4935 365
rect 5297 359 5355 365
rect 5717 359 5775 365
rect 6137 359 6195 365
rect 6557 359 6615 365
rect 6977 359 7035 365
rect 7397 359 7455 365
rect 7817 359 7875 365
rect 8237 359 8295 365
rect 257 325 269 359
rect 677 325 689 359
rect 1097 325 1109 359
rect 1517 325 1529 359
rect 1937 325 1949 359
rect 2357 325 2369 359
rect 2777 325 2789 359
rect 3197 325 3209 359
rect 3617 325 3629 359
rect 4037 325 4049 359
rect 4457 325 4469 359
rect 4877 325 4889 359
rect 5297 325 5309 359
rect 5717 325 5729 359
rect 6137 325 6149 359
rect 6557 325 6569 359
rect 6977 325 6989 359
rect 7397 325 7409 359
rect 7817 325 7829 359
rect 8237 325 8249 359
rect 257 319 315 325
rect 677 319 735 325
rect 1097 319 1155 325
rect 1517 319 1575 325
rect 1937 319 1995 325
rect 2357 319 2415 325
rect 2777 319 2835 325
rect 3197 319 3255 325
rect 3617 319 3675 325
rect 4037 319 4095 325
rect 4457 319 4515 325
rect 4877 319 4935 325
rect 5297 319 5355 325
rect 5717 319 5775 325
rect 6137 319 6195 325
rect 6557 319 6615 325
rect 6977 319 7035 325
rect 7397 319 7455 325
rect 7817 319 7875 325
rect 8237 319 8295 325
rect -1 87 61 287
rect 91 87 153 287
rect 209 87 271 287
rect 301 87 363 287
rect 419 87 481 287
rect 511 87 573 287
rect 629 87 691 287
rect 721 87 783 287
rect 839 87 901 287
rect 931 87 993 287
rect 1049 87 1111 287
rect 1141 87 1203 287
rect 1259 87 1321 287
rect 1351 87 1413 287
rect 1469 87 1531 287
rect 1561 87 1623 287
rect 1679 87 1741 287
rect 1771 87 1833 287
rect 1889 87 1951 287
rect 1981 87 2043 287
rect 2099 87 2161 287
rect 2191 87 2253 287
rect 2309 87 2371 287
rect 2401 87 2463 287
rect 2519 87 2581 287
rect 2611 87 2673 287
rect 2729 87 2791 287
rect 2821 87 2883 287
rect 2939 87 3001 287
rect 3031 87 3093 287
rect 3149 87 3211 287
rect 3241 87 3303 287
rect 3359 87 3421 287
rect 3451 87 3513 287
rect 3569 87 3631 287
rect 3661 87 3723 287
rect 3779 87 3841 287
rect 3871 87 3933 287
rect 3989 87 4051 287
rect 4081 87 4143 287
rect 4199 87 4261 287
rect 4291 87 4353 287
rect 4409 87 4471 287
rect 4501 87 4563 287
rect 4619 87 4681 287
rect 4711 87 4773 287
rect 4829 87 4891 287
rect 4921 87 4983 287
rect 5039 87 5101 287
rect 5131 87 5193 287
rect 5249 87 5311 287
rect 5341 87 5403 287
rect 5459 87 5521 287
rect 5551 87 5613 287
rect 5669 87 5731 287
rect 5761 87 5823 287
rect 5879 87 5941 287
rect 5971 87 6033 287
rect 6089 87 6151 287
rect 6181 87 6243 287
rect 6299 87 6361 287
rect 6391 87 6453 287
rect 6509 87 6571 287
rect 6601 87 6663 287
rect 6719 87 6781 287
rect 6811 87 6873 287
rect 6929 87 6991 287
rect 7021 87 7083 287
rect 7139 87 7201 287
rect 7231 87 7293 287
rect 7349 87 7411 287
rect 7441 87 7503 287
rect 7559 87 7621 287
rect 7651 87 7713 287
rect 7769 87 7831 287
rect 7861 87 7923 287
rect 7979 87 8041 287
rect 8071 87 8133 287
rect 8189 87 8251 287
rect 8281 87 8343 287
rect 8399 87 8461 287
rect 8491 87 8553 287
rect 8609 87 8671 287
rect 8701 87 8763 287
rect 467 49 525 55
rect 887 49 945 55
rect 1307 49 1365 55
rect 1727 49 1785 55
rect 2147 49 2205 55
rect 2567 49 2625 55
rect 2987 49 3045 55
rect 3407 49 3465 55
rect 3827 49 3885 55
rect 4247 49 4305 55
rect 4667 49 4725 55
rect 5087 49 5145 55
rect 5507 49 5565 55
rect 5927 49 5985 55
rect 6347 49 6405 55
rect 6767 49 6825 55
rect 7187 49 7245 55
rect 7607 49 7665 55
rect 8027 49 8085 55
rect 8447 49 8505 55
rect 467 15 479 49
rect 887 15 899 49
rect 1307 15 1319 49
rect 1727 15 1739 49
rect 2147 15 2159 49
rect 2567 15 2579 49
rect 2987 15 2999 49
rect 3407 15 3419 49
rect 3827 15 3839 49
rect 4247 15 4259 49
rect 4667 15 4679 49
rect 5087 15 5099 49
rect 5507 15 5519 49
rect 5927 15 5939 49
rect 6347 15 6359 49
rect 6767 15 6779 49
rect 7187 15 7199 49
rect 7607 15 7619 49
rect 8027 15 8039 49
rect 8447 15 8459 49
rect 467 9 525 15
rect 887 9 945 15
rect 1307 9 1365 15
rect 1727 9 1785 15
rect 2147 9 2205 15
rect 2567 9 2625 15
rect 2987 9 3045 15
rect 3407 9 3465 15
rect 3827 9 3885 15
rect 4247 9 4305 15
rect 4667 9 4725 15
rect 5087 9 5145 15
rect 5507 9 5565 15
rect 5927 9 5985 15
rect 6347 9 6405 15
rect 6767 9 6825 15
rect 7187 9 7245 15
rect 7607 9 7665 15
rect 8027 9 8085 15
rect 8447 9 8505 15
rect 257 -81 315 -75
rect 677 -81 735 -75
rect 1097 -81 1155 -75
rect 1517 -81 1575 -75
rect 1937 -81 1995 -75
rect 2357 -81 2415 -75
rect 2777 -81 2835 -75
rect 3197 -81 3255 -75
rect 3617 -81 3675 -75
rect 4037 -81 4095 -75
rect 4457 -81 4515 -75
rect 4877 -81 4935 -75
rect 5297 -81 5355 -75
rect 5717 -81 5775 -75
rect 6137 -81 6195 -75
rect 6557 -81 6615 -75
rect 6977 -81 7035 -75
rect 7397 -81 7455 -75
rect 7817 -81 7875 -75
rect 8237 -81 8295 -75
rect 257 -115 269 -81
rect 677 -115 689 -81
rect 1097 -115 1109 -81
rect 1517 -115 1529 -81
rect 1937 -115 1949 -81
rect 2357 -115 2369 -81
rect 2777 -115 2789 -81
rect 3197 -115 3209 -81
rect 3617 -115 3629 -81
rect 4037 -115 4049 -81
rect 4457 -115 4469 -81
rect 4877 -115 4889 -81
rect 5297 -115 5309 -81
rect 5717 -115 5729 -81
rect 6137 -115 6149 -81
rect 6557 -115 6569 -81
rect 6977 -115 6989 -81
rect 7397 -115 7409 -81
rect 7817 -115 7829 -81
rect 8237 -115 8249 -81
rect 257 -121 315 -115
rect 677 -121 735 -115
rect 1097 -121 1155 -115
rect 1517 -121 1575 -115
rect 1937 -121 1995 -115
rect 2357 -121 2415 -115
rect 2777 -121 2835 -115
rect 3197 -121 3255 -115
rect 3617 -121 3675 -115
rect 4037 -121 4095 -115
rect 4457 -121 4515 -115
rect 4877 -121 4935 -115
rect 5297 -121 5355 -115
rect 5717 -121 5775 -115
rect 6137 -121 6195 -115
rect 6557 -121 6615 -115
rect 6977 -121 7035 -115
rect 7397 -121 7455 -115
rect 7817 -121 7875 -115
rect 8237 -121 8295 -115
rect -1 -353 61 -153
rect 91 -353 153 -153
rect 209 -353 271 -153
rect 301 -353 363 -153
rect 419 -353 481 -153
rect 511 -353 573 -153
rect 629 -353 691 -153
rect 721 -353 783 -153
rect 839 -353 901 -153
rect 931 -353 993 -153
rect 1049 -353 1111 -153
rect 1141 -353 1203 -153
rect 1259 -353 1321 -153
rect 1351 -353 1413 -153
rect 1469 -353 1531 -153
rect 1561 -353 1623 -153
rect 1679 -353 1741 -153
rect 1771 -353 1833 -153
rect 1889 -353 1951 -153
rect 1981 -353 2043 -153
rect 2099 -353 2161 -153
rect 2191 -353 2253 -153
rect 2309 -353 2371 -153
rect 2401 -353 2463 -153
rect 2519 -353 2581 -153
rect 2611 -353 2673 -153
rect 2729 -353 2791 -153
rect 2821 -353 2883 -153
rect 2939 -353 3001 -153
rect 3031 -353 3093 -153
rect 3149 -353 3211 -153
rect 3241 -353 3303 -153
rect 3359 -353 3421 -153
rect 3451 -353 3513 -153
rect 3569 -353 3631 -153
rect 3661 -353 3723 -153
rect 3779 -353 3841 -153
rect 3871 -353 3933 -153
rect 3989 -353 4051 -153
rect 4081 -353 4143 -153
rect 4199 -353 4261 -153
rect 4291 -353 4353 -153
rect 4409 -353 4471 -153
rect 4501 -353 4563 -153
rect 4619 -353 4681 -153
rect 4711 -353 4773 -153
rect 4829 -353 4891 -153
rect 4921 -353 4983 -153
rect 5039 -353 5101 -153
rect 5131 -353 5193 -153
rect 5249 -353 5311 -153
rect 5341 -353 5403 -153
rect 5459 -353 5521 -153
rect 5551 -353 5613 -153
rect 5669 -353 5731 -153
rect 5761 -353 5823 -153
rect 5879 -353 5941 -153
rect 5971 -353 6033 -153
rect 6089 -353 6151 -153
rect 6181 -353 6243 -153
rect 6299 -353 6361 -153
rect 6391 -353 6453 -153
rect 6509 -353 6571 -153
rect 6601 -353 6663 -153
rect 6719 -353 6781 -153
rect 6811 -353 6873 -153
rect 6929 -353 6991 -153
rect 7021 -353 7083 -153
rect 7139 -353 7201 -153
rect 7231 -353 7293 -153
rect 7349 -353 7411 -153
rect 7441 -353 7503 -153
rect 7559 -353 7621 -153
rect 7651 -353 7713 -153
rect 7769 -353 7831 -153
rect 7861 -353 7923 -153
rect 7979 -353 8041 -153
rect 8071 -353 8133 -153
rect 8189 -353 8251 -153
rect 8281 -353 8343 -153
rect 8399 -353 8461 -153
rect 8491 -353 8553 -153
rect 8609 -353 8671 -153
rect 8701 -353 8763 -153
rect 467 -391 525 -385
rect 887 -391 945 -385
rect 1307 -391 1365 -385
rect 1727 -391 1785 -385
rect 2147 -391 2205 -385
rect 2567 -391 2625 -385
rect 2987 -391 3045 -385
rect 3407 -391 3465 -385
rect 3827 -391 3885 -385
rect 4247 -391 4305 -385
rect 4667 -391 4725 -385
rect 5087 -391 5145 -385
rect 5507 -391 5565 -385
rect 5927 -391 5985 -385
rect 6347 -391 6405 -385
rect 6767 -391 6825 -385
rect 7187 -391 7245 -385
rect 7607 -391 7665 -385
rect 8027 -391 8085 -385
rect 8447 -391 8505 -385
rect 467 -425 479 -391
rect 887 -425 899 -391
rect 1307 -425 1319 -391
rect 1727 -425 1739 -391
rect 2147 -425 2159 -391
rect 2567 -425 2579 -391
rect 2987 -425 2999 -391
rect 3407 -425 3419 -391
rect 3827 -425 3839 -391
rect 4247 -425 4259 -391
rect 4667 -425 4679 -391
rect 5087 -425 5099 -391
rect 5507 -425 5519 -391
rect 5927 -425 5939 -391
rect 6347 -425 6359 -391
rect 6767 -425 6779 -391
rect 7187 -425 7199 -391
rect 7607 -425 7619 -391
rect 8027 -425 8039 -391
rect 8447 -425 8459 -391
rect 467 -431 525 -425
rect 887 -431 945 -425
rect 1307 -431 1365 -425
rect 1727 -431 1785 -425
rect 2147 -431 2205 -425
rect 2567 -431 2625 -425
rect 2987 -431 3045 -425
rect 3407 -431 3465 -425
rect 3827 -431 3885 -425
rect 4247 -431 4305 -425
rect 4667 -431 4725 -425
rect 5087 -431 5145 -425
rect 5507 -431 5565 -425
rect 5927 -431 5985 -425
rect 6347 -431 6405 -425
rect 6767 -431 6825 -425
rect 7187 -431 7245 -425
rect 7607 -431 7665 -425
rect 8027 -431 8085 -425
rect 8447 -431 8505 -425
rect 257 -521 315 -515
rect 677 -521 735 -515
rect 1097 -521 1155 -515
rect 1517 -521 1575 -515
rect 1937 -521 1995 -515
rect 2357 -521 2415 -515
rect 2777 -521 2835 -515
rect 3197 -521 3255 -515
rect 3617 -521 3675 -515
rect 4037 -521 4095 -515
rect 4457 -521 4515 -515
rect 4877 -521 4935 -515
rect 5297 -521 5355 -515
rect 5717 -521 5775 -515
rect 6137 -521 6195 -515
rect 6557 -521 6615 -515
rect 6977 -521 7035 -515
rect 7397 -521 7455 -515
rect 7817 -521 7875 -515
rect 8237 -521 8295 -515
rect 257 -555 269 -521
rect 677 -555 689 -521
rect 1097 -555 1109 -521
rect 1517 -555 1529 -521
rect 1937 -555 1949 -521
rect 2357 -555 2369 -521
rect 2777 -555 2789 -521
rect 3197 -555 3209 -521
rect 3617 -555 3629 -521
rect 4037 -555 4049 -521
rect 4457 -555 4469 -521
rect 4877 -555 4889 -521
rect 5297 -555 5309 -521
rect 5717 -555 5729 -521
rect 6137 -555 6149 -521
rect 6557 -555 6569 -521
rect 6977 -555 6989 -521
rect 7397 -555 7409 -521
rect 7817 -555 7829 -521
rect 8237 -555 8249 -521
rect 257 -561 315 -555
rect 677 -561 735 -555
rect 1097 -561 1155 -555
rect 1517 -561 1575 -555
rect 1937 -561 1995 -555
rect 2357 -561 2415 -555
rect 2777 -561 2835 -555
rect 3197 -561 3255 -555
rect 3617 -561 3675 -555
rect 4037 -561 4095 -555
rect 4457 -561 4515 -555
rect 4877 -561 4935 -555
rect 5297 -561 5355 -555
rect 5717 -561 5775 -555
rect 6137 -561 6195 -555
rect 6557 -561 6615 -555
rect 6977 -561 7035 -555
rect 7397 -561 7455 -555
rect 7817 -561 7875 -555
rect 8237 -561 8295 -555
rect -1 -793 61 -593
rect 91 -793 153 -593
rect 209 -793 271 -593
rect 301 -793 363 -593
rect 419 -793 481 -593
rect 511 -793 573 -593
rect 629 -793 691 -593
rect 721 -793 783 -593
rect 839 -793 901 -593
rect 931 -793 993 -593
rect 1049 -793 1111 -593
rect 1141 -793 1203 -593
rect 1259 -793 1321 -593
rect 1351 -793 1413 -593
rect 1469 -793 1531 -593
rect 1561 -793 1623 -593
rect 1679 -793 1741 -593
rect 1771 -793 1833 -593
rect 1889 -793 1951 -593
rect 1981 -793 2043 -593
rect 2099 -793 2161 -593
rect 2191 -793 2253 -593
rect 2309 -793 2371 -593
rect 2401 -793 2463 -593
rect 2519 -793 2581 -593
rect 2611 -793 2673 -593
rect 2729 -793 2791 -593
rect 2821 -793 2883 -593
rect 2939 -793 3001 -593
rect 3031 -793 3093 -593
rect 3149 -793 3211 -593
rect 3241 -793 3303 -593
rect 3359 -793 3421 -593
rect 3451 -793 3513 -593
rect 3569 -793 3631 -593
rect 3661 -793 3723 -593
rect 3779 -793 3841 -593
rect 3871 -793 3933 -593
rect 3989 -793 4051 -593
rect 4081 -793 4143 -593
rect 4199 -793 4261 -593
rect 4291 -793 4353 -593
rect 4409 -793 4471 -593
rect 4501 -793 4563 -593
rect 4619 -793 4681 -593
rect 4711 -793 4773 -593
rect 4829 -793 4891 -593
rect 4921 -793 4983 -593
rect 5039 -793 5101 -593
rect 5131 -793 5193 -593
rect 5249 -793 5311 -593
rect 5341 -793 5403 -593
rect 5459 -793 5521 -593
rect 5551 -793 5613 -593
rect 5669 -793 5731 -593
rect 5761 -793 5823 -593
rect 5879 -793 5941 -593
rect 5971 -793 6033 -593
rect 6089 -793 6151 -593
rect 6181 -793 6243 -593
rect 6299 -793 6361 -593
rect 6391 -793 6453 -593
rect 6509 -793 6571 -593
rect 6601 -793 6663 -593
rect 6719 -793 6781 -593
rect 6811 -793 6873 -593
rect 6929 -793 6991 -593
rect 7021 -793 7083 -593
rect 7139 -793 7201 -593
rect 7231 -793 7293 -593
rect 7349 -793 7411 -593
rect 7441 -793 7503 -593
rect 7559 -793 7621 -593
rect 7651 -793 7713 -593
rect 7769 -793 7831 -593
rect 7861 -793 7923 -593
rect 7979 -793 8041 -593
rect 8071 -793 8133 -593
rect 8189 -793 8251 -593
rect 8281 -793 8343 -593
rect 8399 -793 8461 -593
rect 8491 -793 8553 -593
rect 8609 -793 8671 -593
rect 8701 -793 8763 -593
rect 467 -831 525 -825
rect 887 -831 945 -825
rect 1307 -831 1365 -825
rect 1727 -831 1785 -825
rect 2147 -831 2205 -825
rect 2567 -831 2625 -825
rect 2987 -831 3045 -825
rect 3407 -831 3465 -825
rect 3827 -831 3885 -825
rect 4247 -831 4305 -825
rect 4667 -831 4725 -825
rect 5087 -831 5145 -825
rect 5507 -831 5565 -825
rect 5927 -831 5985 -825
rect 6347 -831 6405 -825
rect 6767 -831 6825 -825
rect 7187 -831 7245 -825
rect 7607 -831 7665 -825
rect 8027 -831 8085 -825
rect 8447 -831 8505 -825
rect 467 -865 479 -831
rect 887 -865 899 -831
rect 1307 -865 1319 -831
rect 1727 -865 1739 -831
rect 2147 -865 2159 -831
rect 2567 -865 2579 -831
rect 2987 -865 2999 -831
rect 3407 -865 3419 -831
rect 3827 -865 3839 -831
rect 4247 -865 4259 -831
rect 4667 -865 4679 -831
rect 5087 -865 5099 -831
rect 5507 -865 5519 -831
rect 5927 -865 5939 -831
rect 6347 -865 6359 -831
rect 6767 -865 6779 -831
rect 7187 -865 7199 -831
rect 7607 -865 7619 -831
rect 8027 -865 8039 -831
rect 8447 -865 8459 -831
rect 467 -871 525 -865
rect 887 -871 945 -865
rect 1307 -871 1365 -865
rect 1727 -871 1785 -865
rect 2147 -871 2205 -865
rect 2567 -871 2625 -865
rect 2987 -871 3045 -865
rect 3407 -871 3465 -865
rect 3827 -871 3885 -865
rect 4247 -871 4305 -865
rect 4667 -871 4725 -865
rect 5087 -871 5145 -865
rect 5507 -871 5565 -865
rect 5927 -871 5985 -865
rect 6347 -871 6405 -865
rect 6767 -871 6825 -865
rect 7187 -871 7245 -865
rect 7607 -871 7665 -865
rect 8027 -871 8085 -865
rect 8447 -871 8505 -865
rect 257 -961 315 -955
rect 677 -961 735 -955
rect 1097 -961 1155 -955
rect 1517 -961 1575 -955
rect 1937 -961 1995 -955
rect 2357 -961 2415 -955
rect 2777 -961 2835 -955
rect 3197 -961 3255 -955
rect 3617 -961 3675 -955
rect 4037 -961 4095 -955
rect 4457 -961 4515 -955
rect 4877 -961 4935 -955
rect 5297 -961 5355 -955
rect 5717 -961 5775 -955
rect 6137 -961 6195 -955
rect 6557 -961 6615 -955
rect 6977 -961 7035 -955
rect 7397 -961 7455 -955
rect 7817 -961 7875 -955
rect 8237 -961 8295 -955
rect 257 -995 269 -961
rect 677 -995 689 -961
rect 1097 -995 1109 -961
rect 1517 -995 1529 -961
rect 1937 -995 1949 -961
rect 2357 -995 2369 -961
rect 2777 -995 2789 -961
rect 3197 -995 3209 -961
rect 3617 -995 3629 -961
rect 4037 -995 4049 -961
rect 4457 -995 4469 -961
rect 4877 -995 4889 -961
rect 5297 -995 5309 -961
rect 5717 -995 5729 -961
rect 6137 -995 6149 -961
rect 6557 -995 6569 -961
rect 6977 -995 6989 -961
rect 7397 -995 7409 -961
rect 7817 -995 7829 -961
rect 8237 -995 8249 -961
rect 257 -1001 315 -995
rect 677 -1001 735 -995
rect 1097 -1001 1155 -995
rect 1517 -1001 1575 -995
rect 1937 -1001 1995 -995
rect 2357 -1001 2415 -995
rect 2777 -1001 2835 -995
rect 3197 -1001 3255 -995
rect 3617 -1001 3675 -995
rect 4037 -1001 4095 -995
rect 4457 -1001 4515 -995
rect 4877 -1001 4935 -995
rect 5297 -1001 5355 -995
rect 5717 -1001 5775 -995
rect 6137 -1001 6195 -995
rect 6557 -1001 6615 -995
rect 6977 -1001 7035 -995
rect 7397 -1001 7455 -995
rect 7817 -1001 7875 -995
rect 8237 -1001 8295 -995
rect -1 -1233 61 -1033
rect 91 -1233 153 -1033
rect 209 -1233 271 -1033
rect 301 -1233 363 -1033
rect 419 -1233 481 -1033
rect 511 -1233 573 -1033
rect 629 -1233 691 -1033
rect 721 -1233 783 -1033
rect 839 -1233 901 -1033
rect 931 -1233 993 -1033
rect 1049 -1233 1111 -1033
rect 1141 -1233 1203 -1033
rect 1259 -1233 1321 -1033
rect 1351 -1233 1413 -1033
rect 1469 -1233 1531 -1033
rect 1561 -1233 1623 -1033
rect 1679 -1233 1741 -1033
rect 1771 -1233 1833 -1033
rect 1889 -1233 1951 -1033
rect 1981 -1233 2043 -1033
rect 2099 -1233 2161 -1033
rect 2191 -1233 2253 -1033
rect 2309 -1233 2371 -1033
rect 2401 -1233 2463 -1033
rect 2519 -1233 2581 -1033
rect 2611 -1233 2673 -1033
rect 2729 -1233 2791 -1033
rect 2821 -1233 2883 -1033
rect 2939 -1233 3001 -1033
rect 3031 -1233 3093 -1033
rect 3149 -1233 3211 -1033
rect 3241 -1233 3303 -1033
rect 3359 -1233 3421 -1033
rect 3451 -1233 3513 -1033
rect 3569 -1233 3631 -1033
rect 3661 -1233 3723 -1033
rect 3779 -1233 3841 -1033
rect 3871 -1233 3933 -1033
rect 3989 -1233 4051 -1033
rect 4081 -1233 4143 -1033
rect 4199 -1233 4261 -1033
rect 4291 -1233 4353 -1033
rect 4409 -1233 4471 -1033
rect 4501 -1233 4563 -1033
rect 4619 -1233 4681 -1033
rect 4711 -1233 4773 -1033
rect 4829 -1233 4891 -1033
rect 4921 -1233 4983 -1033
rect 5039 -1233 5101 -1033
rect 5131 -1233 5193 -1033
rect 5249 -1233 5311 -1033
rect 5341 -1233 5403 -1033
rect 5459 -1233 5521 -1033
rect 5551 -1233 5613 -1033
rect 5669 -1233 5731 -1033
rect 5761 -1233 5823 -1033
rect 5879 -1233 5941 -1033
rect 5971 -1233 6033 -1033
rect 6089 -1233 6151 -1033
rect 6181 -1233 6243 -1033
rect 6299 -1233 6361 -1033
rect 6391 -1233 6453 -1033
rect 6509 -1233 6571 -1033
rect 6601 -1233 6663 -1033
rect 6719 -1233 6781 -1033
rect 6811 -1233 6873 -1033
rect 6929 -1233 6991 -1033
rect 7021 -1233 7083 -1033
rect 7139 -1233 7201 -1033
rect 7231 -1233 7293 -1033
rect 7349 -1233 7411 -1033
rect 7441 -1233 7503 -1033
rect 7559 -1233 7621 -1033
rect 7651 -1233 7713 -1033
rect 7769 -1233 7831 -1033
rect 7861 -1233 7923 -1033
rect 7979 -1233 8041 -1033
rect 8071 -1233 8133 -1033
rect 8189 -1233 8251 -1033
rect 8281 -1233 8343 -1033
rect 8399 -1233 8461 -1033
rect 8491 -1233 8553 -1033
rect 8609 -1233 8671 -1033
rect 8701 -1233 8763 -1033
rect 467 -1271 525 -1265
rect 887 -1271 945 -1265
rect 1307 -1271 1365 -1265
rect 1727 -1271 1785 -1265
rect 2147 -1271 2205 -1265
rect 2567 -1271 2625 -1265
rect 2987 -1271 3045 -1265
rect 3407 -1271 3465 -1265
rect 3827 -1271 3885 -1265
rect 4247 -1271 4305 -1265
rect 4667 -1271 4725 -1265
rect 5087 -1271 5145 -1265
rect 5507 -1271 5565 -1265
rect 5927 -1271 5985 -1265
rect 6347 -1271 6405 -1265
rect 6767 -1271 6825 -1265
rect 7187 -1271 7245 -1265
rect 7607 -1271 7665 -1265
rect 8027 -1271 8085 -1265
rect 8447 -1271 8505 -1265
rect 467 -1305 479 -1271
rect 887 -1305 899 -1271
rect 1307 -1305 1319 -1271
rect 1727 -1305 1739 -1271
rect 2147 -1305 2159 -1271
rect 2567 -1305 2579 -1271
rect 2987 -1305 2999 -1271
rect 3407 -1305 3419 -1271
rect 3827 -1305 3839 -1271
rect 4247 -1305 4259 -1271
rect 4667 -1305 4679 -1271
rect 5087 -1305 5099 -1271
rect 5507 -1305 5519 -1271
rect 5927 -1305 5939 -1271
rect 6347 -1305 6359 -1271
rect 6767 -1305 6779 -1271
rect 7187 -1305 7199 -1271
rect 7607 -1305 7619 -1271
rect 8027 -1305 8039 -1271
rect 8447 -1305 8459 -1271
rect 467 -1311 525 -1305
rect 887 -1311 945 -1305
rect 1307 -1311 1365 -1305
rect 1727 -1311 1785 -1305
rect 2147 -1311 2205 -1305
rect 2567 -1311 2625 -1305
rect 2987 -1311 3045 -1305
rect 3407 -1311 3465 -1305
rect 3827 -1311 3885 -1305
rect 4247 -1311 4305 -1305
rect 4667 -1311 4725 -1305
rect 5087 -1311 5145 -1305
rect 5507 -1311 5565 -1305
rect 5927 -1311 5985 -1305
rect 6347 -1311 6405 -1305
rect 6767 -1311 6825 -1305
rect 7187 -1311 7245 -1305
rect 7607 -1311 7665 -1305
rect 8027 -1311 8085 -1305
rect 8447 -1311 8505 -1305
rect 257 -1401 315 -1395
rect 677 -1401 735 -1395
rect 1097 -1401 1155 -1395
rect 1517 -1401 1575 -1395
rect 1937 -1401 1995 -1395
rect 2357 -1401 2415 -1395
rect 2777 -1401 2835 -1395
rect 3197 -1401 3255 -1395
rect 3617 -1401 3675 -1395
rect 4037 -1401 4095 -1395
rect 4457 -1401 4515 -1395
rect 4877 -1401 4935 -1395
rect 5297 -1401 5355 -1395
rect 5717 -1401 5775 -1395
rect 6137 -1401 6195 -1395
rect 6557 -1401 6615 -1395
rect 6977 -1401 7035 -1395
rect 7397 -1401 7455 -1395
rect 7817 -1401 7875 -1395
rect 8237 -1401 8295 -1395
rect 257 -1435 269 -1401
rect 677 -1435 689 -1401
rect 1097 -1435 1109 -1401
rect 1517 -1435 1529 -1401
rect 1937 -1435 1949 -1401
rect 2357 -1435 2369 -1401
rect 2777 -1435 2789 -1401
rect 3197 -1435 3209 -1401
rect 3617 -1435 3629 -1401
rect 4037 -1435 4049 -1401
rect 4457 -1435 4469 -1401
rect 4877 -1435 4889 -1401
rect 5297 -1435 5309 -1401
rect 5717 -1435 5729 -1401
rect 6137 -1435 6149 -1401
rect 6557 -1435 6569 -1401
rect 6977 -1435 6989 -1401
rect 7397 -1435 7409 -1401
rect 7817 -1435 7829 -1401
rect 8237 -1435 8249 -1401
rect 257 -1441 315 -1435
rect 677 -1441 735 -1435
rect 1097 -1441 1155 -1435
rect 1517 -1441 1575 -1435
rect 1937 -1441 1995 -1435
rect 2357 -1441 2415 -1435
rect 2777 -1441 2835 -1435
rect 3197 -1441 3255 -1435
rect 3617 -1441 3675 -1435
rect 4037 -1441 4095 -1435
rect 4457 -1441 4515 -1435
rect 4877 -1441 4935 -1435
rect 5297 -1441 5355 -1435
rect 5717 -1441 5775 -1435
rect 6137 -1441 6195 -1435
rect 6557 -1441 6615 -1435
rect 6977 -1441 7035 -1435
rect 7397 -1441 7455 -1435
rect 7817 -1441 7875 -1435
rect 8237 -1441 8295 -1435
rect -1 -1673 61 -1473
rect 91 -1673 153 -1473
rect 209 -1673 271 -1473
rect 301 -1673 363 -1473
rect 419 -1673 481 -1473
rect 511 -1673 573 -1473
rect 629 -1673 691 -1473
rect 721 -1673 783 -1473
rect 839 -1673 901 -1473
rect 931 -1673 993 -1473
rect 1049 -1673 1111 -1473
rect 1141 -1673 1203 -1473
rect 1259 -1673 1321 -1473
rect 1351 -1673 1413 -1473
rect 1469 -1673 1531 -1473
rect 1561 -1673 1623 -1473
rect 1679 -1673 1741 -1473
rect 1771 -1673 1833 -1473
rect 1889 -1673 1951 -1473
rect 1981 -1673 2043 -1473
rect 2099 -1673 2161 -1473
rect 2191 -1673 2253 -1473
rect 2309 -1673 2371 -1473
rect 2401 -1673 2463 -1473
rect 2519 -1673 2581 -1473
rect 2611 -1673 2673 -1473
rect 2729 -1673 2791 -1473
rect 2821 -1673 2883 -1473
rect 2939 -1673 3001 -1473
rect 3031 -1673 3093 -1473
rect 3149 -1673 3211 -1473
rect 3241 -1673 3303 -1473
rect 3359 -1673 3421 -1473
rect 3451 -1673 3513 -1473
rect 3569 -1673 3631 -1473
rect 3661 -1673 3723 -1473
rect 3779 -1673 3841 -1473
rect 3871 -1673 3933 -1473
rect 3989 -1673 4051 -1473
rect 4081 -1673 4143 -1473
rect 4199 -1673 4261 -1473
rect 4291 -1673 4353 -1473
rect 4409 -1673 4471 -1473
rect 4501 -1673 4563 -1473
rect 4619 -1673 4681 -1473
rect 4711 -1673 4773 -1473
rect 4829 -1673 4891 -1473
rect 4921 -1673 4983 -1473
rect 5039 -1673 5101 -1473
rect 5131 -1673 5193 -1473
rect 5249 -1673 5311 -1473
rect 5341 -1673 5403 -1473
rect 5459 -1673 5521 -1473
rect 5551 -1673 5613 -1473
rect 5669 -1673 5731 -1473
rect 5761 -1673 5823 -1473
rect 5879 -1673 5941 -1473
rect 5971 -1673 6033 -1473
rect 6089 -1673 6151 -1473
rect 6181 -1673 6243 -1473
rect 6299 -1673 6361 -1473
rect 6391 -1673 6453 -1473
rect 6509 -1673 6571 -1473
rect 6601 -1673 6663 -1473
rect 6719 -1673 6781 -1473
rect 6811 -1673 6873 -1473
rect 6929 -1673 6991 -1473
rect 7021 -1673 7083 -1473
rect 7139 -1673 7201 -1473
rect 7231 -1673 7293 -1473
rect 7349 -1673 7411 -1473
rect 7441 -1673 7503 -1473
rect 7559 -1673 7621 -1473
rect 7651 -1673 7713 -1473
rect 7769 -1673 7831 -1473
rect 7861 -1673 7923 -1473
rect 7979 -1673 8041 -1473
rect 8071 -1673 8133 -1473
rect 8189 -1673 8251 -1473
rect 8281 -1673 8343 -1473
rect 8399 -1673 8461 -1473
rect 8491 -1673 8553 -1473
rect 8609 -1673 8671 -1473
rect 8701 -1673 8763 -1473
rect 467 -1711 525 -1705
rect 887 -1711 945 -1705
rect 1307 -1711 1365 -1705
rect 1727 -1711 1785 -1705
rect 2147 -1711 2205 -1705
rect 2567 -1711 2625 -1705
rect 2987 -1711 3045 -1705
rect 3407 -1711 3465 -1705
rect 3827 -1711 3885 -1705
rect 4247 -1711 4305 -1705
rect 4667 -1711 4725 -1705
rect 5087 -1711 5145 -1705
rect 5507 -1711 5565 -1705
rect 5927 -1711 5985 -1705
rect 6347 -1711 6405 -1705
rect 6767 -1711 6825 -1705
rect 7187 -1711 7245 -1705
rect 7607 -1711 7665 -1705
rect 8027 -1711 8085 -1705
rect 8447 -1711 8505 -1705
rect 467 -1745 479 -1711
rect 887 -1745 899 -1711
rect 1307 -1745 1319 -1711
rect 1727 -1745 1739 -1711
rect 2147 -1745 2159 -1711
rect 2567 -1745 2579 -1711
rect 2987 -1745 2999 -1711
rect 3407 -1745 3419 -1711
rect 3827 -1745 3839 -1711
rect 4247 -1745 4259 -1711
rect 4667 -1745 4679 -1711
rect 5087 -1745 5099 -1711
rect 5507 -1745 5519 -1711
rect 5927 -1745 5939 -1711
rect 6347 -1745 6359 -1711
rect 6767 -1745 6779 -1711
rect 7187 -1745 7199 -1711
rect 7607 -1745 7619 -1711
rect 8027 -1745 8039 -1711
rect 8447 -1745 8459 -1711
rect 467 -1751 525 -1745
rect 887 -1751 945 -1745
rect 1307 -1751 1365 -1745
rect 1727 -1751 1785 -1745
rect 2147 -1751 2205 -1745
rect 2567 -1751 2625 -1745
rect 2987 -1751 3045 -1745
rect 3407 -1751 3465 -1745
rect 3827 -1751 3885 -1745
rect 4247 -1751 4305 -1745
rect 4667 -1751 4725 -1745
rect 5087 -1751 5145 -1745
rect 5507 -1751 5565 -1745
rect 5927 -1751 5985 -1745
rect 6347 -1751 6405 -1745
rect 6767 -1751 6825 -1745
rect 7187 -1751 7245 -1745
rect 7607 -1751 7665 -1745
rect 8027 -1751 8085 -1745
rect 8447 -1751 8505 -1745
rect 257 -1841 315 -1835
rect 677 -1841 735 -1835
rect 1097 -1841 1155 -1835
rect 1517 -1841 1575 -1835
rect 1937 -1841 1995 -1835
rect 2357 -1841 2415 -1835
rect 2777 -1841 2835 -1835
rect 3197 -1841 3255 -1835
rect 3617 -1841 3675 -1835
rect 4037 -1841 4095 -1835
rect 4457 -1841 4515 -1835
rect 4877 -1841 4935 -1835
rect 5297 -1841 5355 -1835
rect 5717 -1841 5775 -1835
rect 6137 -1841 6195 -1835
rect 6557 -1841 6615 -1835
rect 6977 -1841 7035 -1835
rect 7397 -1841 7455 -1835
rect 7817 -1841 7875 -1835
rect 8237 -1841 8295 -1835
rect 257 -1875 269 -1841
rect 677 -1875 689 -1841
rect 1097 -1875 1109 -1841
rect 1517 -1875 1529 -1841
rect 1937 -1875 1949 -1841
rect 2357 -1875 2369 -1841
rect 2777 -1875 2789 -1841
rect 3197 -1875 3209 -1841
rect 3617 -1875 3629 -1841
rect 4037 -1875 4049 -1841
rect 4457 -1875 4469 -1841
rect 4877 -1875 4889 -1841
rect 5297 -1875 5309 -1841
rect 5717 -1875 5729 -1841
rect 6137 -1875 6149 -1841
rect 6557 -1875 6569 -1841
rect 6977 -1875 6989 -1841
rect 7397 -1875 7409 -1841
rect 7817 -1875 7829 -1841
rect 8237 -1875 8249 -1841
rect 257 -1881 315 -1875
rect 677 -1881 735 -1875
rect 1097 -1881 1155 -1875
rect 1517 -1881 1575 -1875
rect 1937 -1881 1995 -1875
rect 2357 -1881 2415 -1875
rect 2777 -1881 2835 -1875
rect 3197 -1881 3255 -1875
rect 3617 -1881 3675 -1875
rect 4037 -1881 4095 -1875
rect 4457 -1881 4515 -1875
rect 4877 -1881 4935 -1875
rect 5297 -1881 5355 -1875
rect 5717 -1881 5775 -1875
rect 6137 -1881 6195 -1875
rect 6557 -1881 6615 -1875
rect 6977 -1881 7035 -1875
rect 7397 -1881 7455 -1875
rect 7817 -1881 7875 -1875
rect 8237 -1881 8295 -1875
rect -1 -2113 61 -1913
rect 91 -2113 153 -1913
rect 209 -2113 271 -1913
rect 301 -2113 363 -1913
rect 419 -2113 481 -1913
rect 511 -2113 573 -1913
rect 629 -2113 691 -1913
rect 721 -2113 783 -1913
rect 839 -2113 901 -1913
rect 931 -2113 993 -1913
rect 1049 -2113 1111 -1913
rect 1141 -2113 1203 -1913
rect 1259 -2113 1321 -1913
rect 1351 -2113 1413 -1913
rect 1469 -2113 1531 -1913
rect 1561 -2113 1623 -1913
rect 1679 -2113 1741 -1913
rect 1771 -2113 1833 -1913
rect 1889 -2113 1951 -1913
rect 1981 -2113 2043 -1913
rect 2099 -2113 2161 -1913
rect 2191 -2113 2253 -1913
rect 2309 -2113 2371 -1913
rect 2401 -2113 2463 -1913
rect 2519 -2113 2581 -1913
rect 2611 -2113 2673 -1913
rect 2729 -2113 2791 -1913
rect 2821 -2113 2883 -1913
rect 2939 -2113 3001 -1913
rect 3031 -2113 3093 -1913
rect 3149 -2113 3211 -1913
rect 3241 -2113 3303 -1913
rect 3359 -2113 3421 -1913
rect 3451 -2113 3513 -1913
rect 3569 -2113 3631 -1913
rect 3661 -2113 3723 -1913
rect 3779 -2113 3841 -1913
rect 3871 -2113 3933 -1913
rect 3989 -2113 4051 -1913
rect 4081 -2113 4143 -1913
rect 4199 -2113 4261 -1913
rect 4291 -2113 4353 -1913
rect 4409 -2113 4471 -1913
rect 4501 -2113 4563 -1913
rect 4619 -2113 4681 -1913
rect 4711 -2113 4773 -1913
rect 4829 -2113 4891 -1913
rect 4921 -2113 4983 -1913
rect 5039 -2113 5101 -1913
rect 5131 -2113 5193 -1913
rect 5249 -2113 5311 -1913
rect 5341 -2113 5403 -1913
rect 5459 -2113 5521 -1913
rect 5551 -2113 5613 -1913
rect 5669 -2113 5731 -1913
rect 5761 -2113 5823 -1913
rect 5879 -2113 5941 -1913
rect 5971 -2113 6033 -1913
rect 6089 -2113 6151 -1913
rect 6181 -2113 6243 -1913
rect 6299 -2113 6361 -1913
rect 6391 -2113 6453 -1913
rect 6509 -2113 6571 -1913
rect 6601 -2113 6663 -1913
rect 6719 -2113 6781 -1913
rect 6811 -2113 6873 -1913
rect 6929 -2113 6991 -1913
rect 7021 -2113 7083 -1913
rect 7139 -2113 7201 -1913
rect 7231 -2113 7293 -1913
rect 7349 -2113 7411 -1913
rect 7441 -2113 7503 -1913
rect 7559 -2113 7621 -1913
rect 7651 -2113 7713 -1913
rect 7769 -2113 7831 -1913
rect 7861 -2113 7923 -1913
rect 7979 -2113 8041 -1913
rect 8071 -2113 8133 -1913
rect 8189 -2113 8251 -1913
rect 8281 -2113 8343 -1913
rect 8399 -2113 8461 -1913
rect 8491 -2113 8553 -1913
rect 8609 -2113 8671 -1913
rect 8701 -2113 8763 -1913
rect 467 -2151 525 -2145
rect 887 -2151 945 -2145
rect 1307 -2151 1365 -2145
rect 1727 -2151 1785 -2145
rect 2147 -2151 2205 -2145
rect 2567 -2151 2625 -2145
rect 2987 -2151 3045 -2145
rect 3407 -2151 3465 -2145
rect 3827 -2151 3885 -2145
rect 4247 -2151 4305 -2145
rect 4667 -2151 4725 -2145
rect 5087 -2151 5145 -2145
rect 5507 -2151 5565 -2145
rect 5927 -2151 5985 -2145
rect 6347 -2151 6405 -2145
rect 6767 -2151 6825 -2145
rect 7187 -2151 7245 -2145
rect 7607 -2151 7665 -2145
rect 8027 -2151 8085 -2145
rect 8447 -2151 8505 -2145
rect 467 -2185 479 -2151
rect 887 -2185 899 -2151
rect 1307 -2185 1319 -2151
rect 1727 -2185 1739 -2151
rect 2147 -2185 2159 -2151
rect 2567 -2185 2579 -2151
rect 2987 -2185 2999 -2151
rect 3407 -2185 3419 -2151
rect 3827 -2185 3839 -2151
rect 4247 -2185 4259 -2151
rect 4667 -2185 4679 -2151
rect 5087 -2185 5099 -2151
rect 5507 -2185 5519 -2151
rect 5927 -2185 5939 -2151
rect 6347 -2185 6359 -2151
rect 6767 -2185 6779 -2151
rect 7187 -2185 7199 -2151
rect 7607 -2185 7619 -2151
rect 8027 -2185 8039 -2151
rect 8447 -2185 8459 -2151
rect 467 -2191 525 -2185
rect 887 -2191 945 -2185
rect 1307 -2191 1365 -2185
rect 1727 -2191 1785 -2185
rect 2147 -2191 2205 -2185
rect 2567 -2191 2625 -2185
rect 2987 -2191 3045 -2185
rect 3407 -2191 3465 -2185
rect 3827 -2191 3885 -2185
rect 4247 -2191 4305 -2185
rect 4667 -2191 4725 -2185
rect 5087 -2191 5145 -2185
rect 5507 -2191 5565 -2185
rect 5927 -2191 5985 -2185
rect 6347 -2191 6405 -2185
rect 6767 -2191 6825 -2185
rect 7187 -2191 7245 -2185
rect 7607 -2191 7665 -2185
rect 8027 -2191 8085 -2185
rect 8447 -2191 8505 -2185
rect 257 -2281 315 -2275
rect 677 -2281 735 -2275
rect 1097 -2281 1155 -2275
rect 1517 -2281 1575 -2275
rect 1937 -2281 1995 -2275
rect 2357 -2281 2415 -2275
rect 2777 -2281 2835 -2275
rect 3197 -2281 3255 -2275
rect 3617 -2281 3675 -2275
rect 4037 -2281 4095 -2275
rect 4457 -2281 4515 -2275
rect 4877 -2281 4935 -2275
rect 5297 -2281 5355 -2275
rect 5717 -2281 5775 -2275
rect 6137 -2281 6195 -2275
rect 6557 -2281 6615 -2275
rect 6977 -2281 7035 -2275
rect 7397 -2281 7455 -2275
rect 7817 -2281 7875 -2275
rect 8237 -2281 8295 -2275
rect 257 -2315 269 -2281
rect 677 -2315 689 -2281
rect 1097 -2315 1109 -2281
rect 1517 -2315 1529 -2281
rect 1937 -2315 1949 -2281
rect 2357 -2315 2369 -2281
rect 2777 -2315 2789 -2281
rect 3197 -2315 3209 -2281
rect 3617 -2315 3629 -2281
rect 4037 -2315 4049 -2281
rect 4457 -2315 4469 -2281
rect 4877 -2315 4889 -2281
rect 5297 -2315 5309 -2281
rect 5717 -2315 5729 -2281
rect 6137 -2315 6149 -2281
rect 6557 -2315 6569 -2281
rect 6977 -2315 6989 -2281
rect 7397 -2315 7409 -2281
rect 7817 -2315 7829 -2281
rect 8237 -2315 8249 -2281
rect 257 -2321 315 -2315
rect 677 -2321 735 -2315
rect 1097 -2321 1155 -2315
rect 1517 -2321 1575 -2315
rect 1937 -2321 1995 -2315
rect 2357 -2321 2415 -2315
rect 2777 -2321 2835 -2315
rect 3197 -2321 3255 -2315
rect 3617 -2321 3675 -2315
rect 4037 -2321 4095 -2315
rect 4457 -2321 4515 -2315
rect 4877 -2321 4935 -2315
rect 5297 -2321 5355 -2315
rect 5717 -2321 5775 -2315
rect 6137 -2321 6195 -2315
rect 6557 -2321 6615 -2315
rect 6977 -2321 7035 -2315
rect 7397 -2321 7455 -2315
rect 7817 -2321 7875 -2315
rect 8237 -2321 8295 -2315
rect -1 -2553 61 -2353
rect 91 -2553 153 -2353
rect 209 -2553 271 -2353
rect 301 -2553 363 -2353
rect 419 -2553 481 -2353
rect 511 -2553 573 -2353
rect 629 -2553 691 -2353
rect 721 -2553 783 -2353
rect 839 -2553 901 -2353
rect 931 -2553 993 -2353
rect 1049 -2553 1111 -2353
rect 1141 -2553 1203 -2353
rect 1259 -2553 1321 -2353
rect 1351 -2553 1413 -2353
rect 1469 -2553 1531 -2353
rect 1561 -2553 1623 -2353
rect 1679 -2553 1741 -2353
rect 1771 -2553 1833 -2353
rect 1889 -2553 1951 -2353
rect 1981 -2553 2043 -2353
rect 2099 -2553 2161 -2353
rect 2191 -2553 2253 -2353
rect 2309 -2553 2371 -2353
rect 2401 -2553 2463 -2353
rect 2519 -2553 2581 -2353
rect 2611 -2553 2673 -2353
rect 2729 -2553 2791 -2353
rect 2821 -2553 2883 -2353
rect 2939 -2553 3001 -2353
rect 3031 -2553 3093 -2353
rect 3149 -2553 3211 -2353
rect 3241 -2553 3303 -2353
rect 3359 -2553 3421 -2353
rect 3451 -2553 3513 -2353
rect 3569 -2553 3631 -2353
rect 3661 -2553 3723 -2353
rect 3779 -2553 3841 -2353
rect 3871 -2553 3933 -2353
rect 3989 -2553 4051 -2353
rect 4081 -2553 4143 -2353
rect 4199 -2553 4261 -2353
rect 4291 -2553 4353 -2353
rect 4409 -2553 4471 -2353
rect 4501 -2553 4563 -2353
rect 4619 -2553 4681 -2353
rect 4711 -2553 4773 -2353
rect 4829 -2553 4891 -2353
rect 4921 -2553 4983 -2353
rect 5039 -2553 5101 -2353
rect 5131 -2553 5193 -2353
rect 5249 -2553 5311 -2353
rect 5341 -2553 5403 -2353
rect 5459 -2553 5521 -2353
rect 5551 -2553 5613 -2353
rect 5669 -2553 5731 -2353
rect 5761 -2553 5823 -2353
rect 5879 -2553 5941 -2353
rect 5971 -2553 6033 -2353
rect 6089 -2553 6151 -2353
rect 6181 -2553 6243 -2353
rect 6299 -2553 6361 -2353
rect 6391 -2553 6453 -2353
rect 6509 -2553 6571 -2353
rect 6601 -2553 6663 -2353
rect 6719 -2553 6781 -2353
rect 6811 -2553 6873 -2353
rect 6929 -2553 6991 -2353
rect 7021 -2553 7083 -2353
rect 7139 -2553 7201 -2353
rect 7231 -2553 7293 -2353
rect 7349 -2553 7411 -2353
rect 7441 -2553 7503 -2353
rect 7559 -2553 7621 -2353
rect 7651 -2553 7713 -2353
rect 7769 -2553 7831 -2353
rect 7861 -2553 7923 -2353
rect 7979 -2553 8041 -2353
rect 8071 -2553 8133 -2353
rect 8189 -2553 8251 -2353
rect 8281 -2553 8343 -2353
rect 8399 -2553 8461 -2353
rect 8491 -2553 8553 -2353
rect 8609 -2553 8671 -2353
rect 8701 -2553 8763 -2353
rect 467 -2591 525 -2585
rect 887 -2591 945 -2585
rect 1307 -2591 1365 -2585
rect 1727 -2591 1785 -2585
rect 2147 -2591 2205 -2585
rect 2567 -2591 2625 -2585
rect 2987 -2591 3045 -2585
rect 3407 -2591 3465 -2585
rect 3827 -2591 3885 -2585
rect 4247 -2591 4305 -2585
rect 4667 -2591 4725 -2585
rect 5087 -2591 5145 -2585
rect 5507 -2591 5565 -2585
rect 5927 -2591 5985 -2585
rect 6347 -2591 6405 -2585
rect 6767 -2591 6825 -2585
rect 7187 -2591 7245 -2585
rect 7607 -2591 7665 -2585
rect 8027 -2591 8085 -2585
rect 8447 -2591 8505 -2585
rect 467 -2625 479 -2591
rect 887 -2625 899 -2591
rect 1307 -2625 1319 -2591
rect 1727 -2625 1739 -2591
rect 2147 -2625 2159 -2591
rect 2567 -2625 2579 -2591
rect 2987 -2625 2999 -2591
rect 3407 -2625 3419 -2591
rect 3827 -2625 3839 -2591
rect 4247 -2625 4259 -2591
rect 4667 -2625 4679 -2591
rect 5087 -2625 5099 -2591
rect 5507 -2625 5519 -2591
rect 5927 -2625 5939 -2591
rect 6347 -2625 6359 -2591
rect 6767 -2625 6779 -2591
rect 7187 -2625 7199 -2591
rect 7607 -2625 7619 -2591
rect 8027 -2625 8039 -2591
rect 8447 -2625 8459 -2591
rect 467 -2631 525 -2625
rect 887 -2631 945 -2625
rect 1307 -2631 1365 -2625
rect 1727 -2631 1785 -2625
rect 2147 -2631 2205 -2625
rect 2567 -2631 2625 -2625
rect 2987 -2631 3045 -2625
rect 3407 -2631 3465 -2625
rect 3827 -2631 3885 -2625
rect 4247 -2631 4305 -2625
rect 4667 -2631 4725 -2625
rect 5087 -2631 5145 -2625
rect 5507 -2631 5565 -2625
rect 5927 -2631 5985 -2625
rect 6347 -2631 6405 -2625
rect 6767 -2631 6825 -2625
rect 7187 -2631 7245 -2625
rect 7607 -2631 7665 -2625
rect 8027 -2631 8085 -2625
rect 8447 -2631 8505 -2625
rect 257 -2721 315 -2715
rect 677 -2721 735 -2715
rect 1097 -2721 1155 -2715
rect 1517 -2721 1575 -2715
rect 1937 -2721 1995 -2715
rect 2357 -2721 2415 -2715
rect 2777 -2721 2835 -2715
rect 3197 -2721 3255 -2715
rect 3617 -2721 3675 -2715
rect 4037 -2721 4095 -2715
rect 4457 -2721 4515 -2715
rect 4877 -2721 4935 -2715
rect 5297 -2721 5355 -2715
rect 5717 -2721 5775 -2715
rect 6137 -2721 6195 -2715
rect 6557 -2721 6615 -2715
rect 6977 -2721 7035 -2715
rect 7397 -2721 7455 -2715
rect 7817 -2721 7875 -2715
rect 8237 -2721 8295 -2715
rect 257 -2755 269 -2721
rect 677 -2755 689 -2721
rect 1097 -2755 1109 -2721
rect 1517 -2755 1529 -2721
rect 1937 -2755 1949 -2721
rect 2357 -2755 2369 -2721
rect 2777 -2755 2789 -2721
rect 3197 -2755 3209 -2721
rect 3617 -2755 3629 -2721
rect 4037 -2755 4049 -2721
rect 4457 -2755 4469 -2721
rect 4877 -2755 4889 -2721
rect 5297 -2755 5309 -2721
rect 5717 -2755 5729 -2721
rect 6137 -2755 6149 -2721
rect 6557 -2755 6569 -2721
rect 6977 -2755 6989 -2721
rect 7397 -2755 7409 -2721
rect 7817 -2755 7829 -2721
rect 8237 -2755 8249 -2721
rect 257 -2761 315 -2755
rect 677 -2761 735 -2755
rect 1097 -2761 1155 -2755
rect 1517 -2761 1575 -2755
rect 1937 -2761 1995 -2755
rect 2357 -2761 2415 -2755
rect 2777 -2761 2835 -2755
rect 3197 -2761 3255 -2755
rect 3617 -2761 3675 -2755
rect 4037 -2761 4095 -2755
rect 4457 -2761 4515 -2755
rect 4877 -2761 4935 -2755
rect 5297 -2761 5355 -2755
rect 5717 -2761 5775 -2755
rect 6137 -2761 6195 -2755
rect 6557 -2761 6615 -2755
rect 6977 -2761 7035 -2755
rect 7397 -2761 7455 -2755
rect 7817 -2761 7875 -2755
rect 8237 -2761 8295 -2755
rect -1 -2993 61 -2793
rect 91 -2993 153 -2793
rect 209 -2993 271 -2793
rect 301 -2993 363 -2793
rect 419 -2993 481 -2793
rect 511 -2993 573 -2793
rect 629 -2993 691 -2793
rect 721 -2993 783 -2793
rect 839 -2993 901 -2793
rect 931 -2993 993 -2793
rect 1049 -2993 1111 -2793
rect 1141 -2993 1203 -2793
rect 1259 -2993 1321 -2793
rect 1351 -2993 1413 -2793
rect 1469 -2993 1531 -2793
rect 1561 -2993 1623 -2793
rect 1679 -2993 1741 -2793
rect 1771 -2993 1833 -2793
rect 1889 -2993 1951 -2793
rect 1981 -2993 2043 -2793
rect 2099 -2993 2161 -2793
rect 2191 -2993 2253 -2793
rect 2309 -2993 2371 -2793
rect 2401 -2993 2463 -2793
rect 2519 -2993 2581 -2793
rect 2611 -2993 2673 -2793
rect 2729 -2993 2791 -2793
rect 2821 -2993 2883 -2793
rect 2939 -2993 3001 -2793
rect 3031 -2993 3093 -2793
rect 3149 -2993 3211 -2793
rect 3241 -2993 3303 -2793
rect 3359 -2993 3421 -2793
rect 3451 -2993 3513 -2793
rect 3569 -2993 3631 -2793
rect 3661 -2993 3723 -2793
rect 3779 -2993 3841 -2793
rect 3871 -2993 3933 -2793
rect 3989 -2993 4051 -2793
rect 4081 -2993 4143 -2793
rect 4199 -2993 4261 -2793
rect 4291 -2993 4353 -2793
rect 4409 -2993 4471 -2793
rect 4501 -2993 4563 -2793
rect 4619 -2993 4681 -2793
rect 4711 -2993 4773 -2793
rect 4829 -2993 4891 -2793
rect 4921 -2993 4983 -2793
rect 5039 -2993 5101 -2793
rect 5131 -2993 5193 -2793
rect 5249 -2993 5311 -2793
rect 5341 -2993 5403 -2793
rect 5459 -2993 5521 -2793
rect 5551 -2993 5613 -2793
rect 5669 -2993 5731 -2793
rect 5761 -2993 5823 -2793
rect 5879 -2993 5941 -2793
rect 5971 -2993 6033 -2793
rect 6089 -2993 6151 -2793
rect 6181 -2993 6243 -2793
rect 6299 -2993 6361 -2793
rect 6391 -2993 6453 -2793
rect 6509 -2993 6571 -2793
rect 6601 -2993 6663 -2793
rect 6719 -2993 6781 -2793
rect 6811 -2993 6873 -2793
rect 6929 -2993 6991 -2793
rect 7021 -2993 7083 -2793
rect 7139 -2993 7201 -2793
rect 7231 -2993 7293 -2793
rect 7349 -2993 7411 -2793
rect 7441 -2993 7503 -2793
rect 7559 -2993 7621 -2793
rect 7651 -2993 7713 -2793
rect 7769 -2993 7831 -2793
rect 7861 -2993 7923 -2793
rect 7979 -2993 8041 -2793
rect 8071 -2993 8133 -2793
rect 8189 -2993 8251 -2793
rect 8281 -2993 8343 -2793
rect 8399 -2993 8461 -2793
rect 8491 -2993 8553 -2793
rect 8609 -2993 8671 -2793
rect 8701 -2993 8763 -2793
rect 467 -3031 525 -3025
rect 887 -3031 945 -3025
rect 1307 -3031 1365 -3025
rect 1727 -3031 1785 -3025
rect 2147 -3031 2205 -3025
rect 2567 -3031 2625 -3025
rect 2987 -3031 3045 -3025
rect 3407 -3031 3465 -3025
rect 3827 -3031 3885 -3025
rect 4247 -3031 4305 -3025
rect 4667 -3031 4725 -3025
rect 5087 -3031 5145 -3025
rect 5507 -3031 5565 -3025
rect 5927 -3031 5985 -3025
rect 6347 -3031 6405 -3025
rect 6767 -3031 6825 -3025
rect 7187 -3031 7245 -3025
rect 7607 -3031 7665 -3025
rect 8027 -3031 8085 -3025
rect 8447 -3031 8505 -3025
rect 467 -3065 479 -3031
rect 887 -3065 899 -3031
rect 1307 -3065 1319 -3031
rect 1727 -3065 1739 -3031
rect 2147 -3065 2159 -3031
rect 2567 -3065 2579 -3031
rect 2987 -3065 2999 -3031
rect 3407 -3065 3419 -3031
rect 3827 -3065 3839 -3031
rect 4247 -3065 4259 -3031
rect 4667 -3065 4679 -3031
rect 5087 -3065 5099 -3031
rect 5507 -3065 5519 -3031
rect 5927 -3065 5939 -3031
rect 6347 -3065 6359 -3031
rect 6767 -3065 6779 -3031
rect 7187 -3065 7199 -3031
rect 7607 -3065 7619 -3031
rect 8027 -3065 8039 -3031
rect 8447 -3065 8459 -3031
rect 467 -3071 525 -3065
rect 887 -3071 945 -3065
rect 1307 -3071 1365 -3065
rect 1727 -3071 1785 -3065
rect 2147 -3071 2205 -3065
rect 2567 -3071 2625 -3065
rect 2987 -3071 3045 -3065
rect 3407 -3071 3465 -3065
rect 3827 -3071 3885 -3065
rect 4247 -3071 4305 -3065
rect 4667 -3071 4725 -3065
rect 5087 -3071 5145 -3065
rect 5507 -3071 5565 -3065
rect 5927 -3071 5985 -3065
rect 6347 -3071 6405 -3065
rect 6767 -3071 6825 -3065
rect 7187 -3071 7245 -3065
rect 7607 -3071 7665 -3065
rect 8027 -3071 8085 -3065
rect 8447 -3071 8505 -3065
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_0
timestamp 1655495960
transform 1 0 4381 0 1 187
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_1
timestamp 1655495960
transform 1 0 4381 0 1 -253
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_2
timestamp 1655495960
transform 1 0 4381 0 1 -693
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_3
timestamp 1655495960
transform 1 0 4381 0 1 -1133
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_4
timestamp 1655495960
transform 1 0 4381 0 1 -1573
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_5
timestamp 1655495960
transform 1 0 4381 0 1 -2013
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_6
timestamp 1655495960
transform 1 0 4381 0 1 -2453
box -4382 -188 4382 188
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_7
timestamp 1655495960
transform 1 0 4381 0 1 -2893
box -4382 -188 4382 188
<< end >>
