magic
tech sky130A
magscale 1 2
timestamp 1652836164
<< nwell >>
rect -53 413 1241 1063
<< pwell >>
rect -53 -51 1241 413
<< nmos >>
rect 147 159 177 265
rect 243 159 273 265
rect 339 159 369 265
rect 435 159 465 265
rect 531 159 561 265
rect 627 159 657 265
rect 723 159 753 265
rect 819 159 849 265
rect 915 159 945 265
rect 1011 159 1041 265
<< pmos >>
rect 147 570 177 844
rect 243 570 273 844
rect 339 570 369 844
rect 435 570 465 844
rect 531 570 561 844
rect 627 570 657 844
rect 723 570 753 844
rect 819 570 849 844
rect 915 570 945 844
rect 1011 570 1041 844
<< ndiff >>
rect 85 253 147 265
rect 85 171 97 253
rect 131 171 147 253
rect 85 159 147 171
rect 177 253 243 265
rect 177 171 193 253
rect 227 171 243 253
rect 177 159 243 171
rect 273 253 339 265
rect 273 171 289 253
rect 323 171 339 253
rect 273 159 339 171
rect 369 253 435 265
rect 369 171 385 253
rect 419 171 435 253
rect 369 159 435 171
rect 465 253 531 265
rect 465 171 481 253
rect 515 171 531 253
rect 465 159 531 171
rect 561 253 627 265
rect 561 171 577 253
rect 611 171 627 253
rect 561 159 627 171
rect 657 253 723 265
rect 657 171 673 253
rect 707 171 723 253
rect 657 159 723 171
rect 753 253 819 265
rect 753 171 769 253
rect 803 171 819 253
rect 753 159 819 171
rect 849 253 915 265
rect 849 171 865 253
rect 899 171 915 253
rect 849 159 915 171
rect 945 253 1011 265
rect 945 171 961 253
rect 995 171 1011 253
rect 945 159 1011 171
rect 1041 253 1103 265
rect 1041 171 1057 253
rect 1091 171 1103 253
rect 1041 159 1103 171
<< pdiff >>
rect 85 832 147 844
rect 85 582 97 832
rect 131 582 147 832
rect 85 570 147 582
rect 177 832 243 844
rect 177 582 193 832
rect 227 582 243 832
rect 177 570 243 582
rect 273 832 339 844
rect 273 582 289 832
rect 323 582 339 832
rect 273 570 339 582
rect 369 832 435 844
rect 369 582 385 832
rect 419 582 435 832
rect 369 570 435 582
rect 465 832 531 844
rect 465 582 481 832
rect 515 582 531 832
rect 465 570 531 582
rect 561 832 627 844
rect 561 582 577 832
rect 611 582 627 832
rect 561 570 627 582
rect 657 832 723 844
rect 657 582 673 832
rect 707 582 723 832
rect 657 570 723 582
rect 753 832 819 844
rect 753 582 769 832
rect 803 582 819 832
rect 753 570 819 582
rect 849 832 915 844
rect 849 582 865 832
rect 899 582 915 832
rect 849 570 915 582
rect 945 832 1011 844
rect 945 582 961 832
rect 995 582 1011 832
rect 945 570 1011 582
rect 1041 832 1103 844
rect 1041 582 1057 832
rect 1091 582 1103 832
rect 1041 570 1103 582
<< ndiffc >>
rect 97 171 131 253
rect 193 171 227 253
rect 289 171 323 253
rect 385 171 419 253
rect 481 171 515 253
rect 577 171 611 253
rect 673 171 707 253
rect 769 171 803 253
rect 865 171 899 253
rect 961 171 995 253
rect 1057 171 1091 253
<< pdiffc >>
rect 97 582 131 832
rect 193 582 227 832
rect 289 582 323 832
rect 385 582 419 832
rect 481 582 515 832
rect 577 582 611 832
rect 673 582 707 832
rect 769 582 803 832
rect 865 582 899 832
rect 961 582 995 832
rect 1057 582 1091 832
<< psubdiff >>
rect -17 343 79 377
rect 1109 343 1205 377
rect -17 281 17 343
rect 1171 281 1205 343
rect -17 19 17 81
rect 1171 19 1205 81
rect -17 -15 79 19
rect 1109 -15 1205 19
<< nsubdiff >>
rect -17 993 79 1027
rect 1109 993 1205 1027
rect -17 931 17 993
rect 1171 931 1205 993
rect -17 483 17 545
rect 1171 483 1205 545
rect -17 449 79 483
rect 1109 449 1205 483
<< psubdiffcont >>
rect 79 343 1109 377
rect -17 81 17 281
rect 1171 81 1205 281
rect 79 -15 1109 19
<< nsubdiffcont >>
rect 79 993 1109 1027
rect -17 545 17 931
rect 1171 545 1205 931
rect 79 449 1109 483
<< poly >>
rect 81 925 1107 941
rect 81 891 97 925
rect 131 891 289 925
rect 323 891 481 925
rect 515 891 673 925
rect 707 891 865 925
rect 899 891 1057 925
rect 1091 891 1107 925
rect 81 875 1107 891
rect 147 844 177 875
rect 243 844 273 875
rect 339 844 369 875
rect 435 844 465 875
rect 531 844 561 875
rect 627 844 657 875
rect 723 844 753 875
rect 819 844 849 875
rect 915 844 945 875
rect 1011 844 1041 875
rect 147 544 177 570
rect 243 544 273 570
rect 339 544 369 570
rect 435 544 465 570
rect 531 544 561 570
rect 627 544 657 570
rect 723 544 753 570
rect 819 544 849 570
rect 915 544 945 570
rect 1011 544 1041 570
rect 147 265 177 291
rect 243 265 273 291
rect 339 265 369 291
rect 435 265 465 291
rect 531 265 561 291
rect 627 265 657 291
rect 723 265 753 291
rect 819 265 849 291
rect 915 265 945 291
rect 1011 265 1041 291
rect 147 137 177 159
rect 243 137 273 159
rect 339 137 369 159
rect 435 137 465 159
rect 531 137 561 159
rect 627 137 657 159
rect 723 137 753 159
rect 819 137 849 159
rect 915 137 945 159
rect 1011 137 1041 159
rect 81 118 1107 137
rect 81 84 97 118
rect 131 84 289 118
rect 323 84 481 118
rect 515 84 673 118
rect 707 84 865 118
rect 899 84 1057 118
rect 1091 84 1107 118
rect 81 71 1107 84
<< polycont >>
rect 97 891 131 925
rect 289 891 323 925
rect 481 891 515 925
rect 673 891 707 925
rect 865 891 899 925
rect 1057 891 1091 925
rect 97 84 131 118
rect 289 84 323 118
rect 481 84 515 118
rect 673 84 707 118
rect 865 84 899 118
rect 1057 84 1091 118
<< locali >>
rect -17 993 79 1027
rect 1109 993 1205 1027
rect -17 931 17 993
rect 1171 931 1205 993
rect 81 891 97 925
rect 131 891 147 925
rect 273 891 289 925
rect 323 891 339 925
rect 465 891 481 925
rect 515 891 531 925
rect 657 891 673 925
rect 707 891 723 925
rect 849 891 865 925
rect 899 891 915 925
rect 1041 891 1057 925
rect 1091 891 1107 925
rect 97 832 131 848
rect 97 566 131 582
rect 193 832 227 848
rect 193 566 227 582
rect 289 832 323 848
rect 289 566 323 582
rect 385 832 419 848
rect 385 566 419 582
rect 481 832 515 848
rect 481 566 515 582
rect 577 832 611 848
rect 577 566 611 582
rect 673 832 707 848
rect 673 566 707 582
rect 769 832 803 848
rect 769 566 803 582
rect 865 832 899 848
rect 865 566 899 582
rect 961 832 995 848
rect 961 566 995 582
rect 1057 832 1091 848
rect 1057 566 1091 582
rect -17 483 17 545
rect 1171 483 1205 545
rect -17 449 79 483
rect 1109 449 1205 483
rect -17 343 79 377
rect 1109 343 1205 377
rect -17 281 17 343
rect 1171 281 1205 343
rect 97 253 131 269
rect 97 155 131 171
rect 193 253 227 269
rect 193 155 227 171
rect 289 253 323 269
rect 289 155 323 171
rect 385 253 419 269
rect 385 155 419 171
rect 481 253 515 269
rect 481 155 515 171
rect 577 253 611 269
rect 577 155 611 171
rect 673 253 707 269
rect 673 155 707 171
rect 769 253 803 269
rect 769 155 803 171
rect 865 253 899 269
rect 865 155 899 171
rect 961 253 995 269
rect 961 155 995 171
rect 1057 253 1091 269
rect 1057 155 1091 171
rect 81 84 97 118
rect 131 84 147 118
rect 273 84 289 118
rect 323 84 339 118
rect 465 84 481 118
rect 515 84 531 118
rect 657 84 673 118
rect 707 84 723 118
rect 849 84 865 118
rect 899 84 915 118
rect 1041 84 1057 118
rect 1091 84 1107 118
rect -17 19 17 81
rect 1171 19 1205 81
rect -17 -15 79 19
rect 1109 -15 1205 19
<< viali >>
rect 97 891 131 925
rect 289 891 323 925
rect 481 891 515 925
rect 673 891 707 925
rect 865 891 899 925
rect 1057 891 1091 925
rect 97 582 131 832
rect 193 582 227 832
rect 289 582 323 832
rect 385 582 419 832
rect 481 582 515 832
rect 577 582 611 832
rect 673 582 707 832
rect 769 582 803 832
rect 865 582 899 832
rect 961 582 995 832
rect 1057 582 1091 832
rect 1171 545 1205 931
rect 97 171 131 253
rect 193 171 227 253
rect 289 171 323 253
rect 385 171 419 253
rect 481 171 515 253
rect 577 171 611 253
rect 673 171 707 253
rect 769 171 803 253
rect 865 171 899 253
rect 961 171 995 253
rect 1057 171 1091 253
rect 97 84 131 118
rect 289 84 323 118
rect 481 84 515 118
rect 673 84 707 118
rect 865 84 899 118
rect 1057 84 1091 118
rect 1171 81 1205 281
<< metal1 >>
rect -87 993 995 1027
rect -216 883 -189 935
rect -137 883 -127 935
rect -87 430 -53 993
rect 78 883 88 935
rect 140 883 150 935
rect 193 844 227 993
rect 271 883 281 935
rect 333 883 343 935
rect 385 844 419 993
rect 462 883 472 935
rect 524 883 534 935
rect 577 844 611 993
rect 654 883 664 935
rect 716 883 726 935
rect 769 844 803 993
rect 846 883 856 935
rect 908 883 918 935
rect 961 844 995 993
rect 1038 883 1048 935
rect 1100 883 1110 935
rect 1165 931 1211 1063
rect 91 832 137 844
rect 91 582 97 832
rect 131 582 137 832
rect 91 570 137 582
rect 187 832 233 844
rect 187 582 193 832
rect 227 582 233 832
rect 187 570 233 582
rect 283 832 329 844
rect 283 582 289 832
rect 323 582 329 832
rect 283 570 329 582
rect 379 832 425 844
rect 379 582 385 832
rect 419 582 425 832
rect 379 570 425 582
rect 475 832 521 844
rect 475 582 481 832
rect 515 582 521 832
rect 475 570 521 582
rect 571 832 617 844
rect 571 582 577 832
rect 611 582 617 832
rect 571 570 617 582
rect 667 832 713 844
rect 667 582 673 832
rect 707 582 713 832
rect 667 570 713 582
rect 763 832 809 844
rect 763 582 769 832
rect 803 582 809 832
rect 763 570 809 582
rect 859 832 905 844
rect 859 582 865 832
rect 899 582 905 832
rect 859 570 905 582
rect 955 832 1001 844
rect 955 582 961 832
rect 995 582 1001 832
rect 955 570 1001 582
rect 1051 832 1097 844
rect 1051 582 1057 832
rect 1091 582 1097 832
rect 1051 570 1097 582
rect -216 396 -53 430
rect -216 76 -189 128
rect -137 76 -127 128
rect -87 19 -53 396
rect 97 430 131 570
rect 289 430 323 570
rect 481 430 515 570
rect 673 430 707 570
rect 865 430 899 570
rect 1057 430 1091 570
rect 1165 545 1171 931
rect 1205 545 1211 931
rect 1165 533 1211 545
rect 97 396 1283 430
rect 97 265 131 396
rect 289 265 323 396
rect 481 265 515 396
rect 673 265 707 396
rect 865 265 899 396
rect 1057 265 1091 396
rect 1165 281 1211 293
rect 91 253 137 265
rect 91 171 97 253
rect 131 171 137 253
rect 91 159 137 171
rect 187 253 233 265
rect 187 171 193 253
rect 227 171 233 253
rect 187 159 233 171
rect 283 253 329 265
rect 283 171 289 253
rect 323 171 329 253
rect 283 159 329 171
rect 379 253 425 265
rect 379 171 385 253
rect 419 171 425 253
rect 379 159 425 171
rect 475 253 521 265
rect 475 171 481 253
rect 515 171 521 253
rect 475 159 521 171
rect 571 253 617 265
rect 571 171 577 253
rect 611 171 617 253
rect 571 159 617 171
rect 667 253 713 265
rect 667 171 673 253
rect 707 171 713 253
rect 667 159 713 171
rect 763 253 809 265
rect 763 171 769 253
rect 803 171 809 253
rect 763 159 809 171
rect 859 253 905 265
rect 859 171 865 253
rect 899 171 905 253
rect 859 159 905 171
rect 955 253 1001 265
rect 955 171 961 253
rect 995 171 1001 253
rect 955 159 1001 171
rect 1051 253 1097 265
rect 1051 171 1057 253
rect 1091 171 1097 253
rect 1051 159 1097 171
rect 81 128 147 131
rect 78 76 88 128
rect 140 76 150 128
rect 81 71 147 76
rect 193 19 227 159
rect 273 128 339 131
rect 269 76 279 128
rect 331 76 341 128
rect 273 71 339 76
rect 385 19 419 159
rect 465 128 531 131
rect 461 76 471 128
rect 523 76 533 128
rect 465 71 531 76
rect 577 19 611 159
rect 657 128 723 131
rect 653 76 663 128
rect 715 76 725 128
rect 657 71 723 76
rect 769 19 803 159
rect 849 127 915 131
rect 846 75 856 127
rect 908 75 918 127
rect 849 71 915 75
rect 961 19 995 159
rect 1041 127 1107 131
rect 1038 75 1048 127
rect 1100 75 1110 127
rect 1165 81 1171 281
rect 1205 81 1211 281
rect 1041 71 1107 75
rect -87 -15 995 19
rect 1165 -51 1211 81
<< via1 >>
rect -189 883 -137 935
rect 88 925 140 935
rect 88 891 97 925
rect 97 891 131 925
rect 131 891 140 925
rect 88 883 140 891
rect 281 925 333 935
rect 281 891 289 925
rect 289 891 323 925
rect 323 891 333 925
rect 281 883 333 891
rect 472 925 524 935
rect 472 891 481 925
rect 481 891 515 925
rect 515 891 524 925
rect 472 883 524 891
rect 664 925 716 935
rect 664 891 673 925
rect 673 891 707 925
rect 707 891 716 925
rect 664 883 716 891
rect 856 925 908 935
rect 856 891 865 925
rect 865 891 899 925
rect 899 891 908 925
rect 856 883 908 891
rect 1048 925 1100 935
rect 1048 891 1057 925
rect 1057 891 1091 925
rect 1091 891 1100 925
rect 1048 883 1100 891
rect -189 76 -137 128
rect 88 118 140 128
rect 88 84 97 118
rect 97 84 131 118
rect 131 84 140 118
rect 88 76 140 84
rect 279 118 331 128
rect 279 84 289 118
rect 289 84 323 118
rect 323 84 331 118
rect 279 76 331 84
rect 471 118 523 128
rect 471 84 481 118
rect 481 84 515 118
rect 515 84 523 118
rect 471 76 523 84
rect 663 118 715 128
rect 663 84 673 118
rect 673 84 707 118
rect 707 84 715 118
rect 663 76 715 84
rect 856 118 908 127
rect 856 84 865 118
rect 865 84 899 118
rect 899 84 908 118
rect 856 75 908 84
rect 1048 118 1100 127
rect 1048 84 1057 118
rect 1057 84 1091 118
rect 1091 84 1100 118
rect 1048 75 1100 84
<< metal2 >>
rect -189 935 -137 945
rect 88 935 140 945
rect 281 935 333 945
rect 472 935 524 945
rect 664 935 716 945
rect 856 935 908 945
rect 1048 935 1100 945
rect -137 883 88 935
rect 140 883 281 935
rect 333 883 472 935
rect 524 883 664 935
rect 716 883 856 935
rect 908 883 1048 935
rect 1100 883 1107 935
rect -189 873 -137 883
rect 88 873 140 883
rect 281 873 333 883
rect 472 873 524 883
rect 664 873 716 883
rect 856 873 908 883
rect 1048 873 1100 883
rect -189 128 -137 138
rect 88 128 140 138
rect 279 128 331 138
rect 471 128 523 138
rect 663 128 715 138
rect 856 128 908 137
rect 1048 128 1100 137
rect -137 76 88 128
rect 140 76 279 128
rect 331 76 471 128
rect 523 76 663 128
rect 715 127 1107 128
rect 715 76 856 127
rect -189 66 -137 76
rect 88 66 140 76
rect 279 66 331 76
rect 471 66 523 76
rect 663 66 715 76
rect 908 76 1048 127
rect 856 65 908 75
rect 1100 76 1107 127
rect 1048 65 1100 75
<< labels >>
flabel metal1 1188 -48 1188 -48 1 FreeSans 400 0 0 0 VSS
port 6 n ground bidirectional
flabel metal1 1188 1058 1188 1058 5 FreeSans 400 0 0 0 VDD
port 5 s power bidirectional
flabel metal1 -211 909 -211 909 3 FreeSans 400 0 0 0 en_b
port 4 e
flabel metal1 -212 413 -212 413 3 FreeSans 400 0 0 0 in
port 1 e
flabel metal1 -212 102 -212 102 3 FreeSans 400 0 0 0 en
port 3 e
flabel metal1 1279 412 1279 412 7 FreeSans 400 0 0 0 out
port 2 w
<< end >>
