magic
tech sky130A
magscale 1 2
timestamp 1653472245
<< nmos >>
rect -936 -140 -816 140
rect -644 -140 -524 140
rect -352 -140 -232 140
rect -60 -140 60 140
rect 232 -140 352 140
rect 524 -140 644 140
rect 816 -140 936 140
<< ndiff >>
rect -994 128 -936 140
rect -994 -128 -982 128
rect -948 -128 -936 128
rect -994 -140 -936 -128
rect -816 128 -758 140
rect -816 -128 -804 128
rect -770 -128 -758 128
rect -816 -140 -758 -128
rect -702 128 -644 140
rect -702 -128 -690 128
rect -656 -128 -644 128
rect -702 -140 -644 -128
rect -524 128 -466 140
rect -524 -128 -512 128
rect -478 -128 -466 128
rect -524 -140 -466 -128
rect -410 128 -352 140
rect -410 -128 -398 128
rect -364 -128 -352 128
rect -410 -140 -352 -128
rect -232 128 -174 140
rect -232 -128 -220 128
rect -186 -128 -174 128
rect -232 -140 -174 -128
rect -118 128 -60 140
rect -118 -128 -106 128
rect -72 -128 -60 128
rect -118 -140 -60 -128
rect 60 128 118 140
rect 60 -128 72 128
rect 106 -128 118 128
rect 60 -140 118 -128
rect 174 128 232 140
rect 174 -128 186 128
rect 220 -128 232 128
rect 174 -140 232 -128
rect 352 128 410 140
rect 352 -128 364 128
rect 398 -128 410 128
rect 352 -140 410 -128
rect 466 128 524 140
rect 466 -128 478 128
rect 512 -128 524 128
rect 466 -140 524 -128
rect 644 128 702 140
rect 644 -128 656 128
rect 690 -128 702 128
rect 644 -140 702 -128
rect 758 128 816 140
rect 758 -128 770 128
rect 804 -128 816 128
rect 758 -140 816 -128
rect 936 128 994 140
rect 936 -128 948 128
rect 982 -128 994 128
rect 936 -140 994 -128
<< ndiffc >>
rect -982 -128 -948 128
rect -804 -128 -770 128
rect -690 -128 -656 128
rect -512 -128 -478 128
rect -398 -128 -364 128
rect -220 -128 -186 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 186 -128 220 128
rect 364 -128 398 128
rect 478 -128 512 128
rect 656 -128 690 128
rect 770 -128 804 128
rect 948 -128 982 128
<< poly >>
rect -914 212 -838 228
rect -914 195 -898 212
rect -936 178 -898 195
rect -854 195 -838 212
rect -622 212 -546 228
rect -622 195 -606 212
rect -854 178 -816 195
rect -936 140 -816 178
rect -644 178 -606 195
rect -562 195 -546 212
rect -330 212 -254 228
rect -330 195 -314 212
rect -562 178 -524 195
rect -644 140 -524 178
rect -352 178 -314 195
rect -270 195 -254 212
rect -38 212 38 228
rect -38 195 -22 212
rect -270 178 -232 195
rect -352 140 -232 178
rect -60 178 -22 195
rect 22 195 38 212
rect 254 212 330 228
rect 254 195 270 212
rect 22 178 60 195
rect -60 140 60 178
rect 232 178 270 195
rect 314 195 330 212
rect 546 212 622 228
rect 546 195 562 212
rect 314 178 352 195
rect 232 140 352 178
rect 524 178 562 195
rect 606 195 622 212
rect 838 212 914 228
rect 838 195 854 212
rect 606 178 644 195
rect 524 140 644 178
rect 816 178 854 195
rect 898 195 914 212
rect 898 178 936 195
rect 816 140 936 178
rect -936 -178 -816 -140
rect -936 -195 -898 -178
rect -914 -212 -898 -195
rect -854 -195 -816 -178
rect -644 -178 -524 -140
rect -644 -195 -606 -178
rect -854 -212 -838 -195
rect -914 -228 -838 -212
rect -622 -212 -606 -195
rect -562 -195 -524 -178
rect -352 -178 -232 -140
rect -352 -195 -314 -178
rect -562 -212 -546 -195
rect -622 -228 -546 -212
rect -330 -212 -314 -195
rect -270 -195 -232 -178
rect -60 -178 60 -140
rect -60 -195 -22 -178
rect -270 -212 -254 -195
rect -330 -228 -254 -212
rect -38 -212 -22 -195
rect 22 -195 60 -178
rect 232 -178 352 -140
rect 232 -195 270 -178
rect 22 -212 38 -195
rect -38 -228 38 -212
rect 254 -212 270 -195
rect 314 -195 352 -178
rect 524 -178 644 -140
rect 524 -195 562 -178
rect 314 -212 330 -195
rect 254 -228 330 -212
rect 546 -212 562 -195
rect 606 -195 644 -178
rect 816 -178 936 -140
rect 816 -195 854 -178
rect 606 -212 622 -195
rect 546 -228 622 -212
rect 838 -212 854 -195
rect 898 -195 936 -178
rect 898 -212 914 -195
rect 838 -228 914 -212
<< polycont >>
rect -898 178 -854 212
rect -606 178 -562 212
rect -314 178 -270 212
rect -22 178 22 212
rect 270 178 314 212
rect 562 178 606 212
rect 854 178 898 212
rect -898 -212 -854 -178
rect -606 -212 -562 -178
rect -314 -212 -270 -178
rect -22 -212 22 -178
rect 270 -212 314 -178
rect 562 -212 606 -178
rect 854 -212 898 -178
<< locali >>
rect -914 178 -898 212
rect -854 178 -838 212
rect -622 178 -606 212
rect -562 178 -546 212
rect -330 178 -314 212
rect -270 178 -254 212
rect -38 178 -22 212
rect 22 178 38 212
rect 254 178 270 212
rect 314 178 330 212
rect 546 178 562 212
rect 606 178 622 212
rect 838 178 854 212
rect 898 178 914 212
rect -982 128 -948 144
rect -982 -144 -948 -128
rect -804 128 -770 144
rect -804 -144 -770 -128
rect -690 128 -656 144
rect -690 -144 -656 -128
rect -512 128 -478 144
rect -512 -144 -478 -128
rect -398 128 -364 144
rect -398 -144 -364 -128
rect -220 128 -186 144
rect -220 -144 -186 -128
rect -106 128 -72 144
rect -106 -144 -72 -128
rect 72 128 106 144
rect 72 -144 106 -128
rect 186 128 220 144
rect 186 -144 220 -128
rect 364 128 398 144
rect 364 -144 398 -128
rect 478 128 512 144
rect 478 -144 512 -128
rect 656 128 690 144
rect 656 -144 690 -128
rect 770 128 804 144
rect 770 -144 804 -128
rect 948 128 982 144
rect 948 -144 982 -128
rect -914 -212 -898 -178
rect -854 -212 -838 -178
rect -622 -212 -606 -178
rect -562 -212 -546 -178
rect -330 -212 -314 -178
rect -270 -212 -254 -178
rect -38 -212 -22 -178
rect 22 -212 38 -178
rect 254 -212 270 -178
rect 314 -212 330 -178
rect 546 -212 562 -178
rect 606 -212 622 -178
rect 838 -212 854 -178
rect 898 -212 914 -178
<< viali >>
rect -898 178 -854 212
rect -606 178 -562 212
rect -314 178 -270 212
rect -22 178 22 212
rect 270 178 314 212
rect 562 178 606 212
rect 854 178 898 212
rect -982 -128 -948 128
rect -804 -128 -770 128
rect -690 -128 -656 128
rect -512 -128 -478 128
rect -398 -128 -364 128
rect -220 -128 -186 128
rect -106 -128 -72 128
rect 72 -128 106 128
rect 186 -128 220 128
rect 364 -128 398 128
rect 478 -128 512 128
rect 656 -128 690 128
rect 770 -128 804 128
rect 948 -128 982 128
rect -898 -212 -854 -178
rect -606 -212 -562 -178
rect -314 -212 -270 -178
rect -22 -212 22 -178
rect 270 -212 314 -178
rect 562 -212 606 -178
rect 854 -212 898 -178
<< metal1 >>
rect -914 212 -838 228
rect -914 178 -898 212
rect -854 178 -838 212
rect -914 172 -838 178
rect -622 212 -546 228
rect -622 178 -606 212
rect -562 178 -546 212
rect -622 172 -546 178
rect -330 212 -254 228
rect -330 178 -314 212
rect -270 178 -254 212
rect -330 172 -254 178
rect -38 212 38 228
rect -38 178 -22 212
rect 22 178 38 212
rect -38 172 38 178
rect 254 212 330 228
rect 254 178 270 212
rect 314 178 330 212
rect 254 172 330 178
rect 546 212 622 228
rect 546 178 562 212
rect 606 178 622 212
rect 546 172 622 178
rect 838 212 914 228
rect 838 178 854 212
rect 898 178 914 212
rect 838 172 914 178
rect -988 128 -942 140
rect -988 -128 -982 128
rect -948 -128 -942 128
rect -988 -140 -942 -128
rect -810 128 -764 140
rect -810 -128 -804 128
rect -770 -128 -764 128
rect -810 -140 -764 -128
rect -696 128 -650 140
rect -696 -128 -690 128
rect -656 -128 -650 128
rect -696 -140 -650 -128
rect -518 128 -472 140
rect -518 -128 -512 128
rect -478 -128 -472 128
rect -518 -140 -472 -128
rect -404 128 -358 140
rect -404 -128 -398 128
rect -364 -128 -358 128
rect -404 -140 -358 -128
rect -226 128 -180 140
rect -226 -128 -220 128
rect -186 -128 -180 128
rect -226 -140 -180 -128
rect -112 128 -66 140
rect -112 -128 -106 128
rect -72 -128 -66 128
rect -112 -140 -66 -128
rect 66 128 112 140
rect 66 -128 72 128
rect 106 -128 112 128
rect 66 -140 112 -128
rect 180 128 226 140
rect 180 -128 186 128
rect 220 -128 226 128
rect 180 -140 226 -128
rect 358 128 404 140
rect 358 -128 364 128
rect 398 -128 404 128
rect 358 -140 404 -128
rect 472 128 518 140
rect 472 -128 478 128
rect 512 -128 518 128
rect 472 -140 518 -128
rect 650 128 696 140
rect 650 -128 656 128
rect 690 -128 696 128
rect 650 -140 696 -128
rect 764 128 810 140
rect 764 -128 770 128
rect 804 -128 810 128
rect 764 -140 810 -128
rect 942 128 988 140
rect 942 -128 948 128
rect 982 -128 988 128
rect 942 -140 988 -128
rect -914 -178 -838 -172
rect -914 -212 -898 -178
rect -854 -212 -838 -178
rect -914 -228 -838 -212
rect -622 -178 -546 -172
rect -622 -212 -606 -178
rect -562 -212 -546 -178
rect -622 -228 -546 -212
rect -330 -178 -254 -172
rect -330 -212 -314 -178
rect -270 -212 -254 -178
rect -330 -228 -254 -212
rect -38 -178 38 -172
rect -38 -212 -22 -178
rect 22 -212 38 -178
rect -38 -228 38 -212
rect 254 -178 330 -172
rect 254 -212 270 -178
rect 314 -212 330 -178
rect 254 -228 330 -212
rect 546 -178 622 -172
rect 546 -212 562 -178
rect 606 -212 622 -178
rect 546 -228 622 -212
rect 838 -178 914 -172
rect 838 -212 854 -178
rect 898 -212 914 -178
rect 838 -228 914 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 7 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
