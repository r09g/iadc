magic
tech sky130A
magscale 1 2
timestamp 1653475687
<< metal1 >>
rect -5059 -1807 -5025 -1423
rect -5945 -1808 -3809 -1807
rect -5945 -1841 -3776 -1808
rect -5945 -2039 -5911 -1841
rect -5877 -1963 -5867 -1910
rect -5814 -1963 -5804 -1910
rect -5699 -1963 -5689 -1910
rect -5636 -1963 -5626 -1910
rect -5520 -1963 -5510 -1910
rect -5457 -1963 -5447 -1910
rect -5343 -1963 -5333 -1910
rect -5280 -1963 -5270 -1910
rect -5165 -1963 -5155 -1910
rect -5102 -1963 -5092 -1910
rect -4986 -1963 -4976 -1910
rect -4923 -1963 -4913 -1910
rect -4809 -1963 -4799 -1910
rect -4746 -1963 -4736 -1910
rect -4631 -1963 -4621 -1910
rect -4568 -1963 -4558 -1910
rect -4453 -1963 -4443 -1910
rect -4390 -1963 -4380 -1910
rect -4275 -1963 -4265 -1910
rect -4212 -1963 -4202 -1910
rect -4096 -1963 -4086 -1910
rect -4033 -1963 -4023 -1910
rect -3919 -1963 -3909 -1910
rect -3856 -1963 -3846 -1910
rect -6302 -2073 -5911 -2039
rect -6302 -2135 -6268 -2073
rect -6126 -2150 -6092 -2073
rect -5945 -2132 -5911 -2073
rect -5857 -2079 -5823 -1963
rect -5679 -2079 -5645 -1963
rect -5501 -2079 -5467 -1963
rect -5322 -2079 -5288 -1963
rect -5145 -2079 -5111 -1963
rect -4967 -2079 -4933 -1963
rect -4789 -2079 -4755 -1963
rect -4611 -2079 -4577 -1963
rect -4433 -2079 -4399 -1963
rect -4255 -2079 -4221 -1963
rect -4077 -2079 -4043 -1963
rect -3898 -2079 -3864 -1963
rect -3810 -2133 -3776 -1841
rect -1119 -1963 -1109 -1910
rect -1056 -1963 -1046 -1910
rect -6508 -2582 -6498 -2529
rect -6445 -2582 -6435 -2529
rect -6635 -3454 -6625 -3401
rect -6572 -3454 -6562 -3401
rect -6625 -5322 -6572 -3454
rect -6498 -3640 -6445 -2582
rect -6054 -2833 -6044 -2780
rect -5991 -2833 -5981 -2780
rect -6302 -2945 -6090 -2911
rect -6302 -3020 -6268 -2945
rect -6124 -3022 -6090 -2945
rect -6035 -2949 -6001 -2833
rect -6124 -3401 -6090 -3259
rect -6144 -3454 -6134 -3401
rect -6081 -3454 -6071 -3401
rect -6508 -3693 -6498 -3640
rect -6445 -3693 -6435 -3640
rect -6498 -4271 -6445 -3693
rect -6302 -3812 -6090 -3778
rect -6302 -3889 -6268 -3812
rect -6124 -3888 -6090 -3812
rect -6035 -3819 -6001 -3311
rect -6508 -4324 -6498 -4271
rect -6445 -4324 -6435 -4271
rect -6498 -5141 -6445 -4324
rect -6124 -4390 -6090 -4128
rect -6144 -4443 -6134 -4390
rect -6081 -4443 -6071 -4390
rect -6302 -4683 -6090 -4649
rect -6302 -4763 -6268 -4683
rect -6124 -4761 -6090 -4683
rect -6035 -4689 -6001 -4181
rect -6508 -5194 -6498 -5141
rect -6445 -5194 -6435 -5141
rect -6635 -5375 -6625 -5322
rect -6572 -5375 -6562 -5322
rect -6498 -6248 -6445 -5194
rect -6124 -5232 -6090 -4998
rect -6144 -5285 -6134 -5232
rect -6081 -5285 -6071 -5232
rect -6301 -5519 -6091 -5518
rect -5946 -5519 -5912 -2388
rect -5856 -2780 -5822 -2447
rect -5768 -2530 -5734 -2389
rect -5787 -2583 -5777 -2530
rect -5724 -2583 -5714 -2530
rect -5876 -2833 -5866 -2780
rect -5813 -2833 -5803 -2780
rect -5856 -2943 -5822 -2833
rect -5679 -2949 -5645 -2447
rect -5857 -3819 -5823 -3311
rect -5768 -3516 -5734 -3258
rect -5787 -3569 -5777 -3516
rect -5724 -3569 -5714 -3516
rect -5679 -3819 -5645 -3311
rect -5857 -4689 -5823 -4181
rect -5768 -4271 -5734 -4128
rect -5788 -4324 -5778 -4271
rect -5725 -4324 -5715 -4271
rect -5679 -4689 -5645 -4181
rect -6301 -5552 -5912 -5519
rect -6301 -5636 -6267 -5552
rect -6125 -5553 -5912 -5552
rect -6125 -5639 -6091 -5553
rect -5946 -5612 -5912 -5553
rect -5857 -5559 -5823 -5051
rect -5768 -5415 -5734 -4999
rect -5787 -5468 -5777 -5415
rect -5724 -5468 -5714 -5415
rect -5679 -5559 -5645 -5051
rect -5590 -5612 -5556 -2388
rect -5501 -2949 -5467 -2441
rect -5412 -2668 -5378 -2388
rect -5431 -2721 -5421 -2668
rect -5368 -2721 -5358 -2668
rect -5323 -2949 -5289 -2441
rect -5501 -3819 -5467 -3311
rect -5412 -3640 -5378 -3258
rect -5432 -3693 -5422 -3640
rect -5369 -3693 -5359 -3640
rect -5323 -3819 -5289 -3311
rect -5501 -4689 -5467 -4181
rect -5412 -4506 -5378 -4128
rect -5432 -4559 -5422 -4506
rect -5369 -4559 -5359 -4506
rect -5323 -4689 -5289 -4181
rect -5501 -5559 -5467 -5051
rect -5412 -5141 -5378 -4998
rect -5432 -5194 -5422 -5141
rect -5369 -5194 -5359 -5141
rect -5323 -5559 -5289 -5051
rect -5234 -5612 -5200 -2388
rect -5145 -2949 -5111 -2441
rect -5056 -2530 -5022 -2388
rect -5076 -2583 -5066 -2530
rect -5013 -2583 -5003 -2530
rect -4967 -2949 -4933 -2441
rect -5145 -3819 -5111 -3311
rect -5056 -3401 -5022 -3259
rect -5076 -3454 -5066 -3401
rect -5013 -3454 -5003 -3401
rect -4967 -3819 -4933 -3311
rect -5145 -4689 -5111 -4181
rect -5056 -4390 -5022 -4127
rect -5076 -4443 -5066 -4390
rect -5013 -4443 -5003 -4390
rect -4967 -4689 -4933 -4181
rect -5145 -5559 -5111 -5051
rect -5056 -5233 -5022 -4998
rect -5076 -5286 -5066 -5233
rect -5013 -5286 -5003 -5233
rect -4967 -5559 -4933 -5051
rect -4878 -5612 -4844 -2388
rect -4789 -2949 -4755 -2441
rect -4700 -2668 -4666 -2388
rect -4720 -2721 -4710 -2668
rect -4657 -2721 -4647 -2668
rect -4611 -2949 -4577 -2441
rect -4789 -3819 -4755 -3311
rect -4700 -3401 -4666 -3258
rect -4720 -3454 -4710 -3401
rect -4657 -3454 -4647 -3401
rect -4611 -3819 -4577 -3311
rect -4789 -4689 -4755 -4181
rect -4700 -4390 -4666 -4128
rect -4719 -4443 -4709 -4390
rect -4656 -4443 -4646 -4390
rect -4611 -4689 -4577 -4181
rect -4789 -5559 -4755 -5051
rect -4700 -5322 -4666 -4998
rect -4720 -5375 -4710 -5322
rect -4657 -5375 -4647 -5322
rect -4611 -5559 -4577 -5051
rect -4522 -5612 -4488 -2388
rect -4433 -2949 -4399 -2441
rect -4344 -2530 -4310 -2388
rect -4364 -2583 -4354 -2530
rect -4301 -2583 -4291 -2530
rect -4255 -2949 -4221 -2441
rect -4433 -3819 -4399 -3311
rect -4344 -3640 -4310 -3258
rect -4363 -3693 -4353 -3640
rect -4300 -3693 -4290 -3640
rect -4254 -3819 -4220 -3311
rect -4433 -4689 -4399 -4181
rect -4344 -4506 -4310 -4128
rect -4363 -4559 -4353 -4506
rect -4300 -4559 -4290 -4506
rect -4255 -4689 -4221 -4181
rect -4433 -5559 -4399 -5051
rect -4344 -5141 -4310 -4998
rect -4363 -5194 -4353 -5141
rect -4300 -5194 -4290 -5141
rect -4255 -5559 -4221 -5051
rect -4166 -5612 -4132 -2388
rect -4077 -2949 -4043 -2441
rect -3988 -2668 -3954 -2388
rect -4008 -2721 -3998 -2668
rect -3945 -2721 -3935 -2668
rect -3899 -2780 -3865 -2441
rect -3810 -2446 -3776 -2388
rect -3633 -2446 -3599 -2364
rect -3454 -2446 -3420 -2370
rect -1099 -2425 -1065 -1963
rect -3810 -2480 -3420 -2446
rect -1119 -2478 -1109 -2425
rect -1056 -2478 -1046 -2425
rect -762 -2478 -752 -2425
rect -699 -2478 -689 -2425
rect -3918 -2833 -3908 -2780
rect -3855 -2833 -3845 -2780
rect -3899 -2949 -3865 -2833
rect -4077 -3819 -4043 -3311
rect -3988 -3516 -3954 -3258
rect -4008 -3569 -3998 -3516
rect -3945 -3569 -3935 -3516
rect -3899 -3819 -3865 -3311
rect -4077 -4689 -4043 -4181
rect -3988 -4271 -3954 -4128
rect -4008 -4324 -3998 -4271
rect -3945 -4324 -3935 -4271
rect -3899 -4689 -3865 -4181
rect -4077 -5559 -4043 -5051
rect -3988 -5415 -3954 -4998
rect -4007 -5468 -3997 -5415
rect -3944 -5468 -3934 -5415
rect -3899 -5559 -3865 -5051
rect -3810 -5612 -3776 -2480
rect -2634 -2611 -2624 -2558
rect -2571 -2611 -2561 -2558
rect -1295 -2611 -1285 -2558
rect -1232 -2611 -1222 -2558
rect -3308 -2721 -3298 -2668
rect -3245 -2721 -3235 -2668
rect -3741 -2833 -3731 -2780
rect -3678 -2833 -3668 -2780
rect -3721 -2949 -3687 -2833
rect -3721 -3819 -3687 -3311
rect -3632 -3316 -3598 -3258
rect -3454 -3316 -3420 -3234
rect -3632 -3350 -3420 -3316
rect -3632 -3401 -3598 -3350
rect -3652 -3454 -3642 -3401
rect -3589 -3454 -3579 -3401
rect -3298 -3516 -3245 -2721
rect -3141 -3454 -3131 -3401
rect -3078 -3454 -3068 -3401
rect -3308 -3569 -3298 -3516
rect -3245 -3569 -3235 -3516
rect -3721 -4689 -3687 -4181
rect -3632 -4186 -3598 -4128
rect -3453 -4186 -3419 -4076
rect -3632 -4220 -3419 -4186
rect -3632 -4390 -3598 -4220
rect -3652 -4443 -3642 -4390
rect -3589 -4443 -3579 -4390
rect -3298 -4506 -3245 -3569
rect -3308 -4559 -3298 -4506
rect -3245 -4559 -3235 -4506
rect -3632 -5056 -3598 -4999
rect -3453 -5056 -3419 -4946
rect -3632 -5090 -3419 -5056
rect -3632 -5319 -3598 -5090
rect -3652 -5372 -3642 -5319
rect -3589 -5372 -3579 -5319
rect -3298 -5416 -3245 -4559
rect -3130 -5233 -3077 -3454
rect -3140 -5286 -3130 -5233
rect -3077 -5286 -3067 -5233
rect -2624 -5324 -2571 -2611
rect -1276 -2885 -1242 -2611
rect -1207 -2718 -1197 -2665
rect -1144 -2718 -1134 -2665
rect -1187 -2825 -1153 -2718
rect -1099 -2884 -1065 -2478
rect -940 -2611 -930 -2558
rect -877 -2611 -867 -2558
rect -1029 -2718 -1019 -2665
rect -966 -2718 -956 -2665
rect -1009 -2831 -975 -2718
rect -920 -2886 -886 -2611
rect -851 -2718 -841 -2665
rect -788 -2718 -778 -2665
rect -831 -2831 -797 -2718
rect -742 -2884 -708 -2478
rect -208 -2605 182 -2571
rect -208 -2883 -174 -2605
rect -139 -2718 -129 -2665
rect -76 -2718 -66 -2665
rect 40 -2718 50 -2665
rect 103 -2718 113 -2665
rect -119 -2831 -85 -2718
rect 59 -2831 93 -2718
rect 148 -2886 182 -2605
rect 217 -2718 227 -2665
rect 280 -2718 290 -2665
rect 237 -2831 271 -2718
rect 594 -2825 628 -1431
rect 1909 -2479 1919 -2426
rect 1972 -2479 1982 -2426
rect 2265 -2479 2275 -2426
rect 2328 -2479 2338 -2426
rect 1038 -2611 1428 -2577
rect 930 -2718 940 -2665
rect 993 -2718 1003 -2665
rect 949 -2831 983 -2718
rect 1038 -2886 1072 -2611
rect 1107 -2718 1117 -2665
rect 1170 -2718 1180 -2665
rect 1285 -2718 1295 -2665
rect 1348 -2718 1358 -2665
rect 1127 -2831 1161 -2718
rect 1305 -2831 1339 -2718
rect -1454 -3282 -1420 -3140
rect -1365 -3282 -1331 -3199
rect -1276 -3282 -1242 -3141
rect -1454 -3316 -1242 -3282
rect -1454 -3317 -1420 -3316
rect -1655 -3510 -1645 -3449
rect -1584 -3510 -1574 -3449
rect -2014 -4465 -2004 -4412
rect -1951 -4465 -1941 -4412
rect -2003 -4517 -1950 -4465
rect -2634 -5377 -2624 -5324
rect -2571 -5377 -2561 -5324
rect -3308 -5469 -3298 -5416
rect -3245 -5469 -3235 -5416
rect -5946 -6016 -5912 -5869
rect -5966 -6069 -5956 -6016
rect -5903 -6069 -5893 -6016
rect -5768 -6131 -5734 -5868
rect -5590 -6016 -5556 -5868
rect -5611 -6069 -5601 -6016
rect -5548 -6069 -5538 -6016
rect -5788 -6184 -5778 -6131
rect -5725 -6184 -5715 -6131
rect -5412 -6248 -5378 -5868
rect -5234 -6016 -5200 -5868
rect -5254 -6069 -5244 -6016
rect -5191 -6069 -5181 -6016
rect -5056 -6131 -5022 -5869
rect -5075 -6184 -5065 -6131
rect -5012 -6184 -5002 -6131
rect -6508 -6301 -6498 -6248
rect -6445 -6301 -6435 -6248
rect -5431 -6301 -5421 -6248
rect -5368 -6301 -5358 -6248
rect -4967 -6376 -4933 -5927
rect -4878 -6016 -4844 -5868
rect -4898 -6069 -4888 -6016
rect -4835 -6069 -4825 -6016
rect -4700 -6248 -4666 -5868
rect -4720 -6301 -4710 -6248
rect -4657 -6301 -4647 -6248
rect -4613 -6376 -4579 -5921
rect -4522 -6016 -4488 -5868
rect -4542 -6069 -4532 -6016
rect -4479 -6069 -4469 -6016
rect -4344 -6131 -4310 -5868
rect -4166 -6016 -4132 -5868
rect -4185 -6069 -4175 -6016
rect -4122 -6069 -4112 -6016
rect -4364 -6184 -4354 -6131
rect -4301 -6184 -4291 -6131
rect -3988 -6247 -3954 -5868
rect -3810 -5928 -3776 -5868
rect -3632 -5928 -3598 -5836
rect -3455 -5928 -3421 -5814
rect -3810 -5962 -3421 -5928
rect -3810 -6016 -3776 -5962
rect -3830 -6069 -3820 -6016
rect -3767 -6069 -3757 -6016
rect -3298 -6131 -3245 -5469
rect -2624 -6007 -2571 -5377
rect -2634 -6060 -2624 -6007
rect -2571 -6060 -2561 -6007
rect -3308 -6184 -3298 -6131
rect -3245 -6184 -3235 -6131
rect -4008 -6300 -3998 -6247
rect -3945 -6300 -3935 -6247
rect -3988 -6301 -3954 -6300
rect -4967 -6378 -4579 -6376
rect -4967 -6410 -4786 -6378
rect -4796 -6431 -4786 -6410
rect -4733 -6410 -4579 -6378
rect -4733 -6431 -4723 -6410
rect -2002 -6714 -1950 -4517
rect -1886 -5285 -1876 -5232
rect -1823 -5285 -1813 -5232
rect -1646 -5278 -1585 -3510
rect -1296 -3624 -1286 -3571
rect -1233 -3624 -1223 -3571
rect -1276 -3784 -1242 -3624
rect -1186 -3724 -1152 -3200
rect -1118 -3509 -1108 -3456
rect -1055 -3509 -1045 -3456
rect -1098 -3784 -1064 -3509
rect -1009 -3724 -975 -3200
rect -939 -3624 -929 -3571
rect -876 -3624 -866 -3571
rect -919 -3784 -885 -3624
rect -831 -3724 -797 -3200
rect -653 -3282 -619 -3199
rect -563 -3282 -529 -3140
rect -474 -3282 -440 -3199
rect -385 -3282 -351 -3140
rect -295 -3282 -261 -3199
rect -653 -3301 -261 -3282
rect -653 -3316 -484 -3301
rect -494 -3354 -484 -3316
rect -431 -3316 -261 -3301
rect -431 -3354 -421 -3316
rect -760 -3509 -750 -3456
rect -697 -3509 -687 -3456
rect -406 -3509 -396 -3456
rect -343 -3509 -333 -3456
rect -742 -3784 -708 -3509
rect -583 -3624 -573 -3571
rect -520 -3624 -510 -3571
rect -564 -3784 -530 -3624
rect -386 -3784 -352 -3509
rect -208 -3571 -174 -3140
rect -227 -3624 -217 -3571
rect -164 -3624 -154 -3571
rect -208 -3784 -174 -3624
rect -119 -3724 -85 -3200
rect -30 -3456 4 -3138
rect 327 -3456 361 -3139
rect 414 -3283 448 -3199
rect 504 -3283 538 -3141
rect 592 -3283 626 -3199
rect 682 -3283 716 -3141
rect 771 -3283 805 -3199
rect 414 -3301 805 -3283
rect 414 -3317 583 -3301
rect 573 -3354 583 -3317
rect 636 -3317 805 -3301
rect 636 -3354 646 -3317
rect -49 -3509 -39 -3456
rect 14 -3509 24 -3456
rect 307 -3509 317 -3456
rect 370 -3509 380 -3456
rect -30 -3784 4 -3509
rect 589 -3598 623 -3354
rect 860 -3456 894 -3139
rect 1216 -3456 1250 -3136
rect 840 -3509 850 -3456
rect 903 -3509 913 -3456
rect 1196 -3509 1206 -3456
rect 1259 -3509 1269 -3456
rect 59 -3632 1160 -3598
rect 59 -3725 93 -3632
rect 149 -3633 271 -3632
rect 149 -3784 183 -3633
rect 237 -3725 271 -3633
rect 948 -3725 982 -3632
rect 1038 -3783 1072 -3632
rect 1126 -3725 1160 -3632
rect 1216 -3802 1250 -3509
rect 1306 -3724 1340 -3200
rect 1394 -3564 1428 -2611
rect 1928 -2885 1962 -2479
rect 2087 -2607 2097 -2554
rect 2150 -2607 2160 -2554
rect 1997 -2718 2007 -2665
rect 2060 -2718 2070 -2665
rect 2017 -2831 2051 -2718
rect 2105 -2881 2139 -2607
rect 2176 -2718 2186 -2665
rect 2239 -2718 2249 -2665
rect 2195 -2831 2229 -2718
rect 2285 -2887 2319 -2479
rect 3183 -2480 3193 -2427
rect 3246 -2480 3256 -2427
rect 2443 -2607 2453 -2554
rect 2506 -2606 2931 -2554
rect 2506 -2607 2516 -2606
rect 2353 -2718 2363 -2665
rect 2416 -2718 2426 -2665
rect 2373 -2831 2407 -2718
rect 2462 -2885 2496 -2607
rect 1482 -3283 1516 -3199
rect 1572 -3283 1606 -3140
rect 1662 -3283 1696 -3199
rect 1750 -3283 1784 -3140
rect 1840 -3283 1874 -3199
rect 1482 -3301 1874 -3283
rect 1482 -3317 1654 -3301
rect 1644 -3354 1654 -3317
rect 1707 -3317 1874 -3301
rect 1707 -3354 1717 -3317
rect 1552 -3509 1562 -3456
rect 1615 -3509 1625 -3456
rect 1909 -3509 1919 -3456
rect 1972 -3509 1982 -3456
rect 1374 -3617 1384 -3564
rect 1437 -3617 1447 -3564
rect 1394 -3809 1428 -3617
rect 1572 -3784 1606 -3509
rect 1731 -3617 1741 -3564
rect 1794 -3617 1804 -3564
rect 1750 -3786 1784 -3617
rect 1929 -3787 1963 -3509
rect 2017 -3724 2051 -3200
rect 2087 -3617 2097 -3564
rect 2150 -3617 2160 -3564
rect 2106 -3785 2140 -3617
rect 2196 -3724 2230 -3200
rect 2265 -3509 2275 -3456
rect 2328 -3509 2338 -3456
rect 2284 -3785 2318 -3509
rect 2373 -3724 2407 -3200
rect 2462 -3284 2496 -3141
rect 2551 -3284 2585 -3199
rect 2641 -3284 2675 -3141
rect 2462 -3318 2675 -3284
rect 2441 -3617 2451 -3564
rect 2504 -3617 2514 -3564
rect 2462 -3786 2496 -3617
rect -1454 -4184 -1420 -4041
rect -1366 -4184 -1332 -4099
rect -1276 -4184 -1242 -4040
rect -1454 -4218 -1242 -4184
rect -1454 -4541 -1242 -4507
rect -1454 -4685 -1420 -4541
rect -1365 -4624 -1331 -4541
rect -1276 -4706 -1242 -4541
rect -1187 -4625 -1153 -4101
rect -1009 -4624 -975 -4100
rect -831 -4192 -797 -4100
rect -653 -4192 -619 -4101
rect -474 -4192 -440 -4101
rect -297 -4192 -263 -4100
rect -851 -4245 -841 -4192
rect -788 -4245 -778 -4192
rect -672 -4245 -662 -4192
rect -609 -4245 -599 -4192
rect -493 -4245 -483 -4192
rect -430 -4245 -420 -4192
rect -316 -4245 -306 -4192
rect -253 -4245 -243 -4192
rect -831 -4624 -797 -4245
rect -653 -4625 -619 -4245
rect -474 -4625 -440 -4245
rect -297 -4624 -263 -4245
rect -119 -4624 -85 -4100
rect -1277 -5097 -1243 -4939
rect -1297 -5150 -1287 -5097
rect -1234 -5150 -1224 -5097
rect -1876 -5337 -1823 -5285
rect -1875 -6364 -1823 -5337
rect -1656 -5339 -1646 -5278
rect -1585 -5339 -1575 -5278
rect -1454 -5442 -1242 -5408
rect -1454 -5585 -1420 -5442
rect -1363 -5524 -1329 -5442
rect -1276 -5592 -1242 -5442
rect -1187 -5525 -1153 -4995
rect -1097 -5213 -1063 -4938
rect -1115 -5266 -1105 -5213
rect -1052 -5266 -1042 -5213
rect -1009 -5524 -975 -4994
rect -919 -5097 -885 -4937
rect -939 -5150 -929 -5097
rect -876 -5150 -866 -5097
rect -830 -5524 -796 -4994
rect -741 -5213 -707 -4937
rect -563 -5097 -529 -4940
rect -582 -5150 -572 -5097
rect -519 -5150 -509 -5097
rect -386 -5213 -352 -4937
rect -208 -5097 -174 -4910
rect -228 -5150 -218 -5097
rect -165 -5150 -155 -5097
rect -761 -5266 -751 -5213
rect -698 -5266 -688 -5213
rect -406 -5266 -396 -5213
rect -343 -5266 -333 -5213
rect -654 -5434 -262 -5400
rect -654 -5523 -620 -5434
rect -563 -5604 -529 -5434
rect -474 -5524 -440 -5434
rect -385 -5612 -351 -5434
rect -296 -5524 -262 -5434
rect -1274 -6364 -1240 -5839
rect -1886 -6417 -1876 -6364
rect -1823 -6417 -1813 -6364
rect -1292 -6417 -1282 -6364
rect -1229 -6417 -1219 -6364
rect -1099 -6479 -1065 -5845
rect -919 -6365 -885 -5833
rect -938 -6417 -928 -6365
rect -876 -6417 -866 -6365
rect -742 -6479 -708 -5839
rect -1120 -6532 -1110 -6479
rect -1057 -6532 -1047 -6479
rect -762 -6532 -752 -6479
rect -699 -6532 -689 -6479
rect -476 -6493 -442 -5901
rect -208 -6077 -174 -5150
rect -119 -5380 -85 -4994
rect -30 -5213 4 -4938
rect 59 -5091 93 -4992
rect 148 -5091 182 -3952
rect 326 -4304 360 -4040
rect 416 -4192 450 -4094
rect 397 -4245 407 -4192
rect 460 -4245 470 -4192
rect 307 -4357 317 -4304
rect 370 -4357 380 -4304
rect 326 -4706 360 -4357
rect 416 -4624 450 -4245
rect 504 -4412 538 -4040
rect 593 -4192 627 -4101
rect 573 -4245 583 -4192
rect 636 -4245 646 -4192
rect 485 -4465 495 -4412
rect 548 -4465 558 -4412
rect 504 -4703 538 -4465
rect 593 -4625 627 -4245
rect 682 -4304 716 -4040
rect 771 -4192 805 -4100
rect 751 -4245 761 -4192
rect 814 -4245 824 -4192
rect 663 -4357 673 -4304
rect 726 -4357 736 -4304
rect 682 -4687 716 -4357
rect 771 -4624 805 -4245
rect 860 -4412 894 -4040
rect 840 -4465 850 -4412
rect 903 -4465 913 -4412
rect 860 -4716 894 -4465
rect 236 -5091 270 -4999
rect 948 -5091 982 -5000
rect 1039 -5091 1073 -3989
rect 1305 -4624 1339 -4094
rect 1484 -4192 1518 -4094
rect 1661 -4192 1695 -4094
rect 1839 -4192 1873 -4094
rect 2017 -4192 2051 -4094
rect 1464 -4245 1474 -4192
rect 1527 -4245 1537 -4192
rect 1642 -4245 1652 -4192
rect 1705 -4245 1715 -4192
rect 1820 -4245 1830 -4192
rect 1883 -4245 1893 -4192
rect 1998 -4245 2008 -4192
rect 2061 -4245 2071 -4192
rect 1484 -4624 1518 -4245
rect 1661 -4624 1695 -4245
rect 1839 -4624 1873 -4245
rect 2017 -4624 2051 -4245
rect 2195 -4625 2229 -4095
rect 2373 -4624 2407 -4094
rect 2463 -4182 2497 -4038
rect 2552 -4182 2586 -4104
rect 2640 -4180 2674 -4020
rect 2640 -4182 2792 -4180
rect 2463 -4214 2792 -4182
rect 2463 -4216 2674 -4214
rect 2528 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect 2550 -4506 2584 -4327
rect 2758 -4446 2792 -4214
rect 2462 -4540 2674 -4506
rect 2736 -4507 2746 -4446
rect 2807 -4507 2817 -4446
rect 2758 -4508 2792 -4507
rect 2462 -4683 2496 -4540
rect 2550 -4623 2584 -4540
rect 2640 -4713 2674 -4540
rect 1128 -5091 1162 -5002
rect 59 -5125 1162 -5091
rect -51 -5266 -41 -5213
rect 12 -5266 22 -5213
rect 306 -5266 316 -5213
rect 369 -5266 379 -5213
rect -138 -5433 -128 -5380
rect -75 -5433 -65 -5380
rect -119 -5524 -85 -5433
rect -30 -5603 4 -5266
rect 40 -5433 50 -5380
rect 103 -5433 113 -5380
rect 218 -5433 228 -5380
rect 281 -5433 291 -5380
rect 59 -5524 93 -5433
rect 238 -5524 272 -5433
rect 326 -5586 360 -5266
rect 593 -5315 627 -5125
rect 1216 -5213 1250 -4940
rect 840 -5266 850 -5213
rect 903 -5266 913 -5213
rect 1197 -5266 1207 -5213
rect 1260 -5266 1270 -5213
rect 415 -5349 804 -5315
rect 415 -5524 449 -5349
rect 505 -5620 539 -5349
rect 592 -5523 626 -5349
rect 681 -5606 715 -5349
rect 770 -5524 804 -5349
rect 860 -5585 894 -5266
rect 930 -5434 940 -5381
rect 993 -5434 1003 -5381
rect 1109 -5433 1119 -5380
rect 1172 -5433 1182 -5380
rect 949 -5524 983 -5434
rect 1128 -5524 1162 -5433
rect 1216 -5623 1250 -5266
rect 1306 -5380 1340 -4994
rect 1394 -5093 1428 -4913
rect 1375 -5146 1385 -5093
rect 1438 -5146 1448 -5093
rect 1286 -5433 1296 -5380
rect 1349 -5433 1359 -5380
rect 1306 -5524 1340 -5433
rect 149 -6077 183 -5822
rect -208 -6111 183 -6077
rect 237 -6250 271 -5901
rect 217 -6303 227 -6250
rect 280 -6303 290 -6250
rect 594 -6493 628 -5899
rect 951 -6250 985 -5899
rect 1038 -6081 1072 -5808
rect 1394 -6081 1428 -5146
rect 1572 -5213 1606 -4938
rect 1750 -5093 1784 -4938
rect 1730 -5146 1740 -5093
rect 1793 -5146 1803 -5093
rect 1927 -5213 1961 -4940
rect 1553 -5266 1563 -5213
rect 1616 -5266 1626 -5213
rect 1907 -5266 1917 -5213
rect 1970 -5266 1980 -5213
rect 1482 -5433 1874 -5399
rect 1482 -5523 1516 -5433
rect 1573 -5607 1607 -5433
rect 1661 -5523 1695 -5433
rect 1749 -5604 1783 -5433
rect 1840 -5523 1874 -5433
rect 2018 -5523 2052 -4993
rect 2106 -5093 2140 -4939
rect 2086 -5146 2096 -5093
rect 2149 -5146 2159 -5093
rect 2195 -5525 2229 -4995
rect 2284 -5213 2318 -4939
rect 2264 -5266 2274 -5213
rect 2327 -5266 2337 -5213
rect 2373 -5525 2407 -4995
rect 2462 -5093 2496 -4937
rect 2443 -5146 2453 -5093
rect 2506 -5146 2516 -5093
rect 2463 -5442 2674 -5408
rect 2463 -5585 2497 -5442
rect 2550 -5525 2584 -5442
rect 2640 -5587 2674 -5442
rect 1038 -6115 1428 -6081
rect 932 -6303 942 -6250
rect 995 -6303 1005 -6250
rect 1662 -6493 1696 -5901
rect 1928 -6124 1962 -5839
rect 2106 -6007 2140 -5842
rect 2086 -6060 2096 -6007
rect 2149 -6060 2159 -6007
rect 2284 -6124 2318 -5841
rect 2462 -6007 2496 -5839
rect 2442 -6060 2452 -6007
rect 2505 -6060 2515 -6007
rect 1908 -6177 1918 -6124
rect 1971 -6177 1981 -6124
rect 2265 -6177 2275 -6124
rect 2328 -6177 2338 -6124
rect 2879 -6365 2931 -2606
rect 3194 -4805 3246 -2480
rect 3184 -4857 3194 -4805
rect 3246 -4857 3256 -4805
rect 4761 -4857 4771 -4805
rect 4823 -4857 4833 -4805
rect 2869 -6417 2879 -6365
rect 2931 -6417 2941 -6365
rect -476 -6527 1696 -6493
rect -742 -6598 -708 -6532
rect 4771 -6597 4823 -4857
rect 5027 -5059 5037 -5006
rect 5090 -5059 5100 -5006
rect 4895 -5265 4905 -5212
rect 4958 -5265 4968 -5212
rect -763 -6651 -753 -6598
rect -700 -6651 -690 -6598
rect 4762 -6650 4772 -6597
rect 4825 -6650 4835 -6597
rect -3884 -6806 -3874 -6753
rect -3821 -6806 -3811 -6753
rect -2013 -6767 -2003 -6714
rect -1950 -6767 -1940 -6714
rect -3864 -7447 -3830 -6806
rect -3741 -6956 -3731 -6903
rect -3678 -6956 -3668 -6903
rect -5629 -7481 -3830 -7447
rect -5628 -7625 -5594 -7481
rect -5544 -7574 -5500 -7481
rect -5450 -7625 -5416 -7481
rect -5366 -7580 -5322 -7481
rect -5188 -7580 -5144 -7481
rect -5094 -7626 -5060 -7481
rect -5010 -7580 -4966 -7481
rect -4832 -7580 -4788 -7481
rect -4738 -7626 -4704 -7481
rect -4654 -7580 -4610 -7481
rect -4476 -7580 -4432 -7481
rect -4382 -7626 -4348 -7481
rect -4298 -7580 -4254 -7481
rect -3722 -7540 -3688 -6956
rect -3551 -7440 -3541 -7388
rect -3489 -7440 -3479 -7388
rect -4026 -7574 -3688 -7540
rect -4026 -7630 -3992 -7574
rect -5628 -10924 -5594 -7880
rect -5544 -8090 -5500 -7964
rect -5544 -8640 -5500 -8514
rect -5544 -9190 -5500 -9064
rect -5544 -9740 -5500 -9614
rect -5544 -10290 -5500 -10164
rect -5544 -10840 -5500 -10714
rect -5450 -10924 -5416 -7880
rect -5366 -8090 -5322 -7964
rect -5366 -8640 -5322 -8514
rect -5366 -9190 -5322 -9064
rect -5366 -9740 -5322 -9614
rect -5366 -10290 -5322 -10164
rect -5366 -10840 -5322 -10714
rect -5272 -10924 -5238 -7880
rect -5188 -8090 -5144 -7964
rect -5188 -8640 -5144 -8514
rect -5188 -9190 -5144 -9064
rect -5188 -9740 -5144 -9614
rect -5188 -10290 -5144 -10164
rect -5188 -10840 -5144 -10714
rect -5094 -10924 -5060 -7881
rect -5010 -8091 -4966 -7965
rect -5010 -8640 -4966 -8514
rect -5010 -9190 -4966 -9064
rect -5010 -9740 -4966 -9614
rect -5010 -10290 -4966 -10164
rect -5010 -10840 -4966 -10714
rect -4916 -10924 -4882 -7880
rect -4832 -8090 -4788 -7964
rect -4832 -8640 -4788 -8514
rect -4832 -9190 -4788 -9064
rect -4832 -9740 -4788 -9614
rect -4832 -10290 -4788 -10164
rect -4832 -10840 -4788 -10714
rect -4738 -10924 -4704 -7880
rect -4654 -8090 -4610 -7964
rect -4654 -8640 -4610 -8514
rect -4654 -9190 -4610 -9064
rect -4654 -9740 -4610 -9614
rect -4654 -10290 -4610 -10164
rect -4654 -10840 -4610 -10714
rect -4560 -10924 -4526 -7880
rect -4476 -8090 -4432 -7964
rect -4476 -8640 -4432 -8514
rect -4476 -9190 -4432 -9064
rect -4476 -9740 -4432 -9614
rect -4476 -10290 -4432 -10164
rect -4476 -10840 -4432 -10714
rect -4382 -10924 -4348 -7880
rect -4298 -8090 -4254 -7964
rect -4298 -8640 -4254 -8514
rect -4298 -9190 -4254 -9064
rect -4298 -9740 -4254 -9614
rect -4298 -10290 -4254 -10164
rect -4298 -10840 -4254 -10714
rect -4204 -10924 -4170 -7880
rect -4120 -8090 -4076 -7964
rect -4120 -8640 -4076 -8514
rect -4120 -9190 -4076 -9064
rect -4120 -9740 -4076 -9614
rect -4120 -10290 -4076 -10164
rect -4120 -10840 -4076 -10714
rect -4026 -10924 -3992 -7880
rect -5272 -11320 -5238 -11181
rect -4916 -11320 -4882 -11180
rect -4560 -11320 -4526 -11180
rect -4204 -11320 -4170 -11180
rect -4120 -11320 -4076 -11264
rect -4026 -11320 -3992 -11180
rect -5272 -11354 -3611 -11320
rect -5512 -11524 -5502 -11471
rect -5449 -11524 -5439 -11471
rect -6976 -11765 -6077 -11712
rect -6024 -11765 -6014 -11712
rect -5636 -11765 -5626 -11712
rect -5573 -11765 -5563 -11712
rect -6233 -12315 -6223 -12262
rect -6170 -12315 -6160 -12262
rect -6976 -13105 -6426 -13052
rect -6373 -13105 -6363 -13052
rect -6223 -13255 -6170 -12315
rect -6077 -12945 -6024 -11765
rect -5922 -11828 -5877 -11812
rect -5922 -11900 -5876 -11828
rect -5817 -11868 -5778 -11812
rect -5617 -11862 -5583 -11765
rect -5824 -11900 -5778 -11868
rect -5492 -11900 -5458 -11524
rect -5010 -11525 -5000 -11472
rect -4947 -11525 -4937 -11472
rect -4512 -11524 -4502 -11471
rect -4449 -11524 -4439 -11471
rect -5386 -11641 -5376 -11588
rect -5323 -11641 -5313 -11588
rect -5137 -11641 -5127 -11588
rect -5074 -11641 -5064 -11588
rect -5367 -11868 -5333 -11641
rect -5117 -11868 -5083 -11641
rect -4992 -11900 -4958 -11525
rect -4887 -11765 -4877 -11712
rect -4824 -11765 -4814 -11712
rect -4637 -11765 -4627 -11712
rect -4574 -11765 -4564 -11712
rect -4867 -11868 -4833 -11765
rect -4617 -11868 -4583 -11765
rect -4492 -11900 -4458 -11524
rect -4387 -11641 -4377 -11588
rect -4324 -11641 -4314 -11588
rect -4367 -11868 -4333 -11641
rect -3938 -11642 -3928 -11589
rect -3875 -11642 -3865 -11589
rect -4172 -11900 -4126 -11812
rect -5824 -11940 -5626 -11900
rect -5574 -11940 -5376 -11900
rect -5324 -11940 -5126 -11900
rect -5074 -11940 -4876 -11900
rect -4823 -11940 -4625 -11900
rect -4574 -11940 -4376 -11900
rect -4324 -11940 -4126 -11900
rect -4074 -11912 -4028 -11812
rect -5818 -12140 -5632 -12100
rect -5574 -12140 -5376 -12100
rect -5324 -12140 -5126 -12100
rect -5074 -12140 -4876 -12100
rect -4825 -12140 -4627 -12100
rect -4574 -12140 -4376 -12100
rect -4324 -12140 -4126 -12100
rect -5744 -12262 -5704 -12140
rect -5761 -12315 -5751 -12262
rect -5698 -12315 -5688 -12262
rect -5495 -12580 -5455 -12140
rect -5245 -12389 -5205 -12140
rect -5261 -12442 -5251 -12389
rect -5198 -12442 -5188 -12389
rect -4995 -12580 -4955 -12140
rect -4746 -12262 -4706 -12140
rect -4762 -12315 -4752 -12262
rect -4699 -12315 -4689 -12262
rect -4495 -12580 -4455 -12140
rect -4244 -12389 -4204 -12140
rect -4261 -12442 -4251 -12389
rect -4198 -12442 -4188 -12389
rect -5824 -12620 -5626 -12580
rect -5574 -12620 -5376 -12580
rect -5324 -12620 -5126 -12580
rect -5074 -12620 -4876 -12580
rect -4824 -12620 -4626 -12580
rect -4574 -12620 -4376 -12580
rect -4324 -12620 -4126 -12580
rect -5922 -12908 -5876 -12808
rect -5824 -12820 -5626 -12780
rect -5574 -12820 -5376 -12780
rect -5324 -12820 -5126 -12780
rect -5074 -12820 -4876 -12780
rect -4824 -12820 -4626 -12780
rect -4574 -12820 -4376 -12780
rect -4324 -12820 -4126 -12780
rect -5824 -12908 -5778 -12820
rect -6087 -12998 -6077 -12945
rect -6024 -12998 -6014 -12945
rect -5720 -13157 -5686 -12820
rect -5617 -13052 -5583 -12852
rect -5367 -12945 -5333 -12852
rect -5386 -12998 -5376 -12945
rect -5323 -12998 -5313 -12945
rect -5636 -13105 -5626 -13052
rect -5573 -13105 -5563 -13052
rect -5740 -13210 -5730 -13157
rect -5677 -13210 -5667 -13157
rect -5240 -13255 -5206 -12820
rect -5117 -12945 -5083 -12852
rect -5136 -12998 -5126 -12945
rect -5073 -12998 -5063 -12945
rect -4867 -13052 -4833 -12852
rect -4887 -13105 -4877 -13052
rect -4824 -13105 -4814 -13052
rect -4742 -13157 -4708 -12820
rect -4617 -13052 -4583 -12852
rect -4367 -12945 -4333 -12852
rect -4386 -12998 -4376 -12945
rect -4323 -12998 -4313 -12945
rect -4637 -13105 -4627 -13052
rect -4574 -13105 -4564 -13052
rect -4762 -13210 -4752 -13157
rect -4699 -13210 -4689 -13157
rect -4240 -13255 -4206 -12820
rect -4172 -12908 -4126 -12820
rect -4074 -12908 -4028 -12808
rect -3928 -13052 -3875 -11642
rect -3798 -12442 -3788 -12389
rect -3735 -12442 -3725 -12389
rect -3938 -13105 -3928 -13052
rect -3875 -13105 -3865 -13052
rect -3928 -13106 -3875 -13105
rect -3788 -13157 -3735 -12442
rect -3798 -13210 -3788 -13157
rect -3735 -13210 -3725 -13157
rect -6233 -13308 -6223 -13255
rect -6170 -13308 -6160 -13255
rect -5260 -13308 -5250 -13255
rect -5197 -13308 -5187 -13255
rect -4260 -13308 -4250 -13255
rect -4197 -13308 -4187 -13255
rect -6965 -13460 -4303 -13426
rect -6028 -13594 -5994 -13460
rect -5939 -13550 -5905 -13460
rect -5850 -13594 -5816 -13460
rect -5761 -13550 -5727 -13460
rect -5583 -13550 -5549 -13460
rect -5405 -13550 -5371 -13460
rect -5227 -13550 -5193 -13460
rect -5049 -13550 -5015 -13460
rect -4871 -13550 -4837 -13460
rect -4693 -13550 -4659 -13460
rect -4515 -13550 -4481 -13460
rect -4337 -13550 -4303 -13460
rect -4248 -13460 -4036 -13426
rect -4248 -13594 -4214 -13460
rect -4159 -13544 -4125 -13460
rect -4070 -13594 -4036 -13460
rect -5850 -13995 -5816 -13851
rect -6169 -14048 -6159 -13995
rect -6106 -14048 -6096 -13995
rect -5870 -14048 -5860 -13995
rect -5807 -14048 -5797 -13995
rect -6159 -14682 -6106 -14048
rect -6028 -14159 -5816 -14125
rect -6027 -14293 -5993 -14159
rect -5939 -14250 -5905 -14159
rect -5850 -14294 -5816 -14159
rect -5761 -14210 -5727 -13900
rect -5672 -14294 -5638 -13850
rect -5583 -14235 -5549 -13919
rect -5494 -14101 -5460 -13850
rect -5514 -14154 -5504 -14101
rect -5451 -14154 -5441 -14101
rect -5405 -14233 -5371 -13917
rect -6169 -14735 -6159 -14682
rect -6106 -14735 -6096 -14682
rect -6159 -15393 -6106 -14735
rect -5850 -14788 -5816 -14550
rect -5870 -14841 -5860 -14788
rect -5807 -14841 -5797 -14788
rect -5761 -14917 -5727 -14601
rect -5672 -15003 -5638 -14550
rect -5583 -14924 -5549 -14608
rect -5494 -14681 -5460 -14550
rect -5514 -14734 -5504 -14681
rect -5451 -14734 -5441 -14681
rect -5405 -14931 -5371 -14615
rect -6028 -15385 -5994 -15249
rect -5939 -15385 -5905 -15294
rect -5850 -15385 -5816 -15250
rect -6169 -15446 -6159 -15393
rect -6106 -15446 -6096 -15393
rect -6028 -15419 -5816 -15385
rect -6159 -16207 -6106 -15446
rect -5850 -15494 -5816 -15419
rect -5870 -15547 -5860 -15494
rect -5807 -15547 -5797 -15494
rect -5761 -15626 -5727 -15310
rect -5672 -15694 -5638 -15250
rect -5583 -15628 -5549 -15312
rect -5494 -15393 -5460 -15250
rect -5514 -15446 -5504 -15393
rect -5451 -15446 -5441 -15393
rect -5405 -15627 -5371 -15311
rect -5316 -15694 -5282 -13850
rect -5227 -14232 -5193 -13916
rect -5138 -13995 -5104 -13851
rect -5157 -14048 -5147 -13995
rect -5094 -14048 -5084 -13995
rect -5049 -14232 -5015 -13916
rect -5227 -14929 -5193 -14613
rect -5138 -14789 -5104 -14550
rect -5158 -14842 -5148 -14789
rect -5095 -14842 -5085 -14789
rect -5049 -14930 -5015 -14614
rect -5227 -15627 -5193 -15311
rect -5138 -15494 -5104 -15251
rect -5158 -15547 -5148 -15494
rect -5095 -15547 -5085 -15494
rect -5049 -15627 -5015 -15311
rect -4960 -15694 -4926 -13850
rect -4871 -14231 -4837 -13915
rect -4782 -14101 -4748 -13850
rect -4801 -14154 -4791 -14101
rect -4738 -14154 -4728 -14101
rect -4693 -14230 -4659 -13914
rect -4871 -14930 -4837 -14614
rect -4782 -14681 -4748 -14550
rect -4802 -14734 -4792 -14681
rect -4739 -14734 -4729 -14681
rect -4693 -14929 -4659 -14613
rect -4871 -15627 -4837 -15311
rect -4782 -15393 -4748 -15250
rect -4802 -15446 -4792 -15393
rect -4739 -15446 -4729 -15393
rect -4693 -15627 -4659 -15311
rect -4604 -15694 -4570 -13850
rect -4515 -14230 -4481 -13914
rect -4426 -13995 -4392 -13850
rect -4446 -14048 -4436 -13995
rect -4383 -14048 -4373 -13995
rect -4337 -14228 -4303 -13912
rect -4248 -14125 -4214 -13850
rect -4159 -13950 -4125 -13900
rect -3664 -14101 -3611 -11354
rect -3541 -12337 -3489 -7440
rect -3392 -7586 -3382 -7533
rect -3329 -7586 -3319 -7533
rect -1392 -7575 -1382 -7522
rect -1329 -7575 -1319 -7522
rect -3542 -12389 -3489 -12337
rect -3552 -12442 -3542 -12389
rect -3489 -12442 -3479 -12389
rect -3382 -13255 -3329 -7586
rect -1372 -7680 -1338 -7575
rect -1213 -7576 -1203 -7523
rect -1150 -7576 -1140 -7523
rect -1035 -7575 -1025 -7522
rect -972 -7575 -962 -7522
rect -858 -7575 -848 -7522
rect -795 -7575 -785 -7522
rect -680 -7575 -670 -7522
rect -617 -7575 -607 -7522
rect -500 -7575 -490 -7522
rect -437 -7575 -427 -7522
rect 745 -7575 755 -7522
rect 808 -7575 818 -7522
rect 922 -7575 932 -7522
rect 985 -7575 995 -7522
rect 1102 -7575 1112 -7522
rect 1165 -7575 1175 -7522
rect -1194 -7681 -1160 -7576
rect -1016 -7681 -982 -7575
rect -838 -7681 -804 -7575
rect -660 -7681 -626 -7575
rect -481 -7681 -447 -7575
rect 765 -7682 799 -7575
rect 942 -7681 976 -7575
rect 1121 -7681 1155 -7575
rect 1279 -7576 1289 -7523
rect 1342 -7576 1352 -7523
rect 1457 -7575 1467 -7522
rect 1520 -7575 1530 -7522
rect 1634 -7575 1644 -7522
rect 1697 -7575 1707 -7522
rect 2880 -7575 2890 -7522
rect 2943 -7575 2953 -7522
rect 3059 -7575 3069 -7522
rect 3122 -7575 3132 -7522
rect 3237 -7575 3247 -7522
rect 3300 -7575 3310 -7522
rect 3414 -7575 3424 -7522
rect 3477 -7575 3487 -7522
rect 1298 -7682 1332 -7576
rect 1476 -7681 1510 -7575
rect 1654 -7681 1688 -7575
rect 2900 -7681 2934 -7575
rect 3078 -7682 3112 -7575
rect 3256 -7681 3290 -7575
rect 3434 -7681 3468 -7575
rect 3593 -7576 3603 -7523
rect 3656 -7576 3666 -7523
rect 3768 -7575 3778 -7522
rect 3831 -7575 3841 -7522
rect 3612 -7681 3646 -7576
rect 3790 -7681 3824 -7575
rect 4198 -7576 4208 -7523
rect 4261 -7576 4271 -7523
rect -2171 -8040 -2137 -7958
rect -1995 -8040 -1961 -7989
rect -2171 -8074 -1961 -8040
rect -1995 -8367 -1961 -8074
rect -1906 -8134 -1872 -8038
rect -1926 -8187 -1916 -8134
rect -1863 -8187 -1853 -8134
rect -1817 -8253 -1783 -7989
rect -1729 -8134 -1695 -8038
rect -1749 -8187 -1739 -8134
rect -1686 -8187 -1676 -8134
rect -1836 -8306 -1826 -8253
rect -1773 -8306 -1763 -8253
rect -2457 -8420 -2447 -8367
rect -2394 -8420 -2384 -8367
rect -2015 -8420 -2005 -8367
rect -1952 -8420 -1942 -8367
rect -2447 -11472 -2394 -8420
rect -2174 -9039 -2140 -8960
rect -1995 -9039 -1961 -8420
rect -2174 -9073 -1961 -9039
rect -2325 -9578 -2315 -9525
rect -2262 -9578 -2252 -9525
rect -2457 -11525 -2447 -11472
rect -2394 -11525 -2384 -11472
rect -3392 -13308 -3382 -13255
rect -3329 -13308 -3319 -13255
rect -4248 -14159 -4036 -14125
rect -3946 -14154 -3936 -14101
rect -3883 -14154 -3611 -14101
rect -4515 -14927 -4481 -14611
rect -4426 -14789 -4392 -14551
rect -4445 -14841 -4435 -14789
rect -4383 -14841 -4373 -14789
rect -4337 -14927 -4303 -14611
rect -4515 -15627 -4481 -15311
rect -4426 -15494 -4392 -15250
rect -4446 -15547 -4436 -15494
rect -4383 -15547 -4373 -15494
rect -4337 -15627 -4303 -15311
rect -4248 -15385 -4214 -14159
rect -4159 -14250 -4125 -14159
rect -4070 -14294 -4036 -14159
rect -3936 -14206 -3883 -14154
rect -3935 -14789 -3883 -14206
rect -3945 -14841 -3935 -14789
rect -3883 -14841 -3873 -14789
rect -4159 -15385 -4125 -15294
rect -4070 -15385 -4036 -15250
rect -4248 -15419 -4036 -15385
rect -4248 -15694 -4214 -15419
rect -3935 -15495 -3883 -14841
rect -2447 -15421 -2394 -11525
rect -2315 -14143 -2262 -9578
rect -1995 -9649 -1961 -9073
rect -1906 -9146 -1872 -9041
rect -1926 -9199 -1916 -9146
rect -1863 -9199 -1853 -9146
rect -1926 -9578 -1916 -9525
rect -1863 -9578 -1853 -9525
rect -2175 -9683 -1961 -9649
rect -1906 -9682 -1872 -9578
rect -2175 -9774 -2141 -9683
rect -1995 -9863 -1961 -9683
rect -1817 -9795 -1783 -8306
rect -1639 -8367 -1605 -7978
rect -1549 -8134 -1515 -8039
rect -1568 -8187 -1558 -8134
rect -1505 -8187 -1495 -8134
rect -1461 -8253 -1427 -7980
rect -1392 -8187 -1382 -8134
rect -1329 -8187 -1319 -8134
rect -1480 -8306 -1470 -8253
rect -1417 -8306 -1407 -8253
rect -1658 -8420 -1648 -8367
rect -1595 -8420 -1585 -8367
rect -1728 -9146 -1694 -9039
rect -1748 -9199 -1738 -9146
rect -1685 -9199 -1675 -9146
rect -1748 -9579 -1738 -9526
rect -1685 -9579 -1675 -9526
rect -1728 -9681 -1694 -9579
rect -1639 -9853 -1605 -8420
rect -1549 -9146 -1515 -9038
rect -1568 -9199 -1558 -9146
rect -1505 -9199 -1495 -9146
rect -1570 -9578 -1560 -9525
rect -1507 -9578 -1497 -9525
rect -1550 -9681 -1516 -9578
rect -1461 -9800 -1427 -8306
rect -1372 -8681 -1338 -8187
rect -1283 -8367 -1249 -7981
rect -1213 -8187 -1203 -8134
rect -1150 -8187 -1140 -8134
rect -1303 -8420 -1293 -8367
rect -1240 -8420 -1230 -8367
rect -1372 -9524 -1338 -9039
rect -1392 -9577 -1382 -9524
rect -1329 -9577 -1319 -9524
rect -1283 -9856 -1249 -8420
rect -1193 -8681 -1159 -8187
rect -1105 -8253 -1071 -7970
rect -1036 -8187 -1026 -8134
rect -973 -8187 -963 -8134
rect -1125 -8306 -1115 -8253
rect -1062 -8306 -1052 -8253
rect -1105 -9808 -1071 -8306
rect -1016 -8681 -982 -8187
rect -927 -8367 -893 -7982
rect -858 -8187 -848 -8134
rect -795 -8187 -785 -8134
rect -946 -8420 -936 -8367
rect -883 -8420 -873 -8367
rect -927 -9857 -893 -8420
rect -838 -8680 -804 -8187
rect -749 -8253 -715 -7968
rect -680 -8187 -670 -8134
rect -617 -8187 -607 -8134
rect -768 -8306 -758 -8253
rect -705 -8306 -695 -8253
rect -749 -9780 -715 -8306
rect -660 -8682 -626 -8187
rect -571 -8366 -537 -7973
rect -501 -8187 -491 -8134
rect -438 -8187 -428 -8134
rect -590 -8419 -580 -8366
rect -527 -8419 -517 -8366
rect -571 -9848 -537 -8419
rect -482 -8681 -448 -8187
rect -393 -8253 -359 -7958
rect -304 -8134 -270 -8039
rect -324 -8187 -314 -8134
rect -261 -8187 -251 -8134
rect -412 -8306 -402 -8253
rect -349 -8306 -339 -8253
rect -393 -9780 -359 -8306
rect -215 -8367 -181 -7971
rect -126 -8134 -92 -8039
rect -146 -8187 -136 -8134
rect -83 -8187 -73 -8134
rect -37 -8253 -3 -7953
rect 52 -8134 86 -8038
rect 32 -8187 42 -8134
rect 95 -8187 105 -8134
rect -57 -8306 -47 -8253
rect 6 -8306 16 -8253
rect -235 -8420 -225 -8367
rect -172 -8420 -162 -8367
rect -303 -9146 -269 -9040
rect -322 -9199 -312 -9146
rect -259 -9199 -249 -9146
rect -324 -9578 -314 -9525
rect -261 -9578 -251 -9525
rect -304 -9682 -270 -9578
rect -215 -9846 -181 -8420
rect -126 -9145 -92 -9038
rect -146 -9198 -136 -9145
rect -83 -9198 -73 -9145
rect -146 -9579 -136 -9526
rect -83 -9579 -73 -9526
rect -126 -9681 -92 -9579
rect -37 -9784 -3 -8306
rect 141 -8368 175 -7980
rect 230 -8134 264 -8040
rect 211 -8187 221 -8134
rect 274 -8187 284 -8134
rect 319 -8253 353 -7962
rect 408 -8134 442 -8040
rect 388 -8187 398 -8134
rect 451 -8187 461 -8134
rect 300 -8306 310 -8253
rect 363 -8306 373 -8253
rect 122 -8421 132 -8368
rect 185 -8421 195 -8368
rect 52 -9146 86 -9040
rect 32 -9199 42 -9146
rect 95 -9199 105 -9146
rect 33 -9578 43 -9525
rect 96 -9578 106 -9525
rect 52 -9682 86 -9578
rect 141 -9855 175 -8421
rect 231 -9145 265 -9039
rect 212 -9198 222 -9145
rect 275 -9198 285 -9145
rect 210 -9578 220 -9525
rect 273 -9578 283 -9525
rect 230 -9681 264 -9578
rect 319 -9794 353 -8306
rect 497 -8366 531 -7970
rect 586 -8134 620 -8039
rect 567 -8187 577 -8134
rect 630 -8187 640 -8134
rect 675 -8253 709 -7965
rect 744 -8187 754 -8134
rect 807 -8187 817 -8134
rect 656 -8306 666 -8253
rect 719 -8306 729 -8253
rect 479 -8419 489 -8366
rect 542 -8419 552 -8366
rect 408 -9146 442 -9038
rect 389 -9199 399 -9146
rect 452 -9199 462 -9146
rect 388 -9578 398 -9525
rect 451 -9578 461 -9525
rect 408 -9682 442 -9578
rect 497 -9845 531 -8419
rect 587 -9146 621 -9040
rect 567 -9199 577 -9146
rect 630 -9199 640 -9146
rect 566 -9578 576 -9525
rect 629 -9578 639 -9525
rect 586 -9682 620 -9578
rect 675 -9789 709 -8306
rect 764 -8682 798 -8187
rect 853 -8366 887 -7969
rect 922 -8187 932 -8134
rect 985 -8187 995 -8134
rect 833 -8419 843 -8366
rect 896 -8419 906 -8366
rect 853 -8791 887 -8419
rect 942 -8681 976 -8187
rect 1031 -8253 1065 -7966
rect 1101 -8187 1111 -8134
rect 1164 -8187 1174 -8134
rect 1012 -8306 1022 -8253
rect 1075 -8306 1085 -8253
rect 1031 -9813 1065 -8306
rect 1120 -8681 1154 -8187
rect 1209 -8367 1243 -7964
rect 1279 -8187 1289 -8134
rect 1342 -8187 1352 -8134
rect 1191 -8420 1201 -8367
rect 1254 -8420 1264 -8367
rect 1209 -9839 1243 -8420
rect 1298 -8681 1332 -8187
rect 1387 -8253 1421 -7965
rect 1456 -8187 1466 -8134
rect 1519 -8187 1529 -8134
rect 1367 -8306 1377 -8253
rect 1430 -8306 1440 -8253
rect 1387 -9813 1421 -8306
rect 1476 -8681 1510 -8187
rect 1565 -8367 1599 -7972
rect 1634 -8187 1644 -8134
rect 1697 -8187 1707 -8134
rect 1546 -8420 1556 -8367
rect 1609 -8420 1619 -8367
rect 1565 -9847 1599 -8420
rect 1654 -8681 1688 -8187
rect 1743 -8253 1777 -7963
rect 1832 -8134 1866 -8039
rect 1812 -8187 1822 -8134
rect 1875 -8187 1885 -8134
rect 1723 -8306 1733 -8253
rect 1786 -8306 1796 -8253
rect 1743 -9781 1777 -8306
rect 1921 -8367 1955 -7972
rect 2010 -8134 2044 -8039
rect 1990 -8187 2000 -8134
rect 2053 -8187 2063 -8134
rect 2099 -8253 2133 -7968
rect 2188 -8134 2222 -8039
rect 2168 -8187 2178 -8134
rect 2231 -8187 2241 -8134
rect 2080 -8306 2090 -8253
rect 2143 -8306 2153 -8253
rect 1901 -8420 1911 -8367
rect 1964 -8420 1974 -8367
rect 1832 -9682 1866 -9026
rect 1921 -9847 1955 -8420
rect 2010 -9682 2044 -9026
rect 2099 -9809 2133 -8306
rect 2277 -8367 2311 -7972
rect 2367 -8134 2401 -8039
rect 2347 -8187 2357 -8134
rect 2410 -8187 2420 -8134
rect 2455 -8253 2489 -7970
rect 2544 -8134 2578 -8039
rect 2524 -8187 2534 -8134
rect 2587 -8187 2597 -8134
rect 2436 -8306 2446 -8253
rect 2499 -8306 2509 -8253
rect 2257 -8420 2267 -8367
rect 2320 -8420 2330 -8367
rect 2188 -9147 2222 -9026
rect 2168 -9200 2178 -9147
rect 2231 -9200 2241 -9147
rect 2188 -9682 2222 -9200
rect 2277 -9847 2311 -8420
rect 2366 -9146 2400 -9040
rect 2347 -9199 2357 -9146
rect 2410 -9199 2420 -9146
rect 2346 -9578 2356 -9525
rect 2409 -9578 2419 -9525
rect 2366 -9682 2400 -9578
rect 2455 -9786 2489 -8306
rect 2633 -8367 2667 -7975
rect 2722 -8134 2756 -8040
rect 2702 -8187 2712 -8134
rect 2765 -8187 2775 -8134
rect 2811 -8253 2845 -7974
rect 2880 -8187 2890 -8134
rect 2943 -8187 2953 -8134
rect 2792 -8306 2802 -8253
rect 2855 -8306 2865 -8253
rect 2614 -8420 2624 -8367
rect 2677 -8420 2687 -8367
rect 2544 -9146 2578 -9041
rect 2524 -9199 2534 -9146
rect 2587 -9199 2597 -9146
rect 2524 -9578 2534 -9525
rect 2587 -9578 2597 -9525
rect 2544 -9681 2578 -9578
rect 2633 -9850 2667 -8420
rect 2722 -9146 2756 -9041
rect 2703 -9199 2713 -9146
rect 2766 -9199 2776 -9146
rect 2702 -9579 2712 -9526
rect 2765 -9579 2775 -9526
rect 2722 -9681 2756 -9579
rect 2811 -9805 2845 -8306
rect 2900 -8682 2934 -8187
rect 2989 -8367 3023 -7976
rect 3058 -8187 3068 -8134
rect 3121 -8187 3131 -8134
rect 2970 -8420 2980 -8367
rect 3033 -8420 3043 -8367
rect 2881 -9578 2891 -9525
rect 2944 -9578 2954 -9525
rect 2900 -9680 2934 -9578
rect 2989 -9851 3023 -8420
rect 3078 -8682 3112 -8187
rect 3167 -8253 3201 -7962
rect 3236 -8187 3246 -8134
rect 3299 -8187 3309 -8134
rect 3148 -8306 3158 -8253
rect 3211 -8306 3221 -8253
rect 3059 -9578 3069 -9525
rect 3122 -9578 3132 -9525
rect 3078 -9680 3112 -9578
rect 3167 -9776 3201 -8306
rect 3256 -8681 3290 -8187
rect 3345 -8367 3379 -7974
rect 3414 -8187 3424 -8134
rect 3477 -8187 3487 -8134
rect 3326 -8420 3336 -8367
rect 3389 -8420 3399 -8367
rect 3256 -9525 3290 -9043
rect 3236 -9578 3246 -9525
rect 3299 -9578 3309 -9525
rect 3256 -9681 3290 -9578
rect 3345 -9849 3379 -8420
rect 3434 -8682 3468 -8187
rect 3523 -8253 3557 -7965
rect 3592 -8187 3602 -8134
rect 3655 -8187 3665 -8134
rect 3503 -8306 3513 -8253
rect 3566 -8306 3576 -8253
rect 3523 -9790 3557 -8306
rect 3612 -8682 3646 -8187
rect 3701 -8367 3735 -7976
rect 3879 -8040 3913 -7965
rect 4056 -8040 4090 -7960
rect 3879 -8074 4090 -8040
rect 3771 -8187 3781 -8134
rect 3834 -8187 3844 -8134
rect 3682 -8420 3692 -8367
rect 3745 -8420 3755 -8367
rect 3701 -9851 3735 -8420
rect 3790 -8681 3824 -8187
rect 3879 -8253 3913 -8074
rect 3859 -8306 3869 -8253
rect 3922 -8306 3932 -8253
rect 3879 -9039 3913 -8306
rect 4056 -9039 4090 -8961
rect 3879 -9073 4090 -9039
rect 3879 -9647 3913 -9073
rect 4208 -9146 4261 -7576
rect 4771 -8862 4823 -6650
rect 4771 -8914 4824 -8862
rect 4761 -8967 4771 -8914
rect 4824 -8967 4834 -8914
rect 4198 -9199 4208 -9146
rect 4261 -9199 4271 -9146
rect 3879 -9681 4092 -9647
rect 3879 -9805 3913 -9681
rect 4058 -9774 4092 -9681
rect -1837 -10561 -1827 -10508
rect -1774 -10561 -1764 -10508
rect -1480 -10561 -1470 -10508
rect -1417 -10561 -1407 -10508
rect -2172 -11039 -2138 -10945
rect -1995 -11039 -1961 -10789
rect -2172 -11073 -1961 -11039
rect -1995 -11237 -1961 -11073
rect -2014 -11290 -2004 -11237
rect -1951 -11290 -1941 -11237
rect -1995 -11647 -1961 -11290
rect -1905 -11519 -1871 -11045
rect -1925 -11572 -1915 -11519
rect -1862 -11572 -1852 -11519
rect -2176 -11681 -1961 -11647
rect -2176 -11771 -2142 -11681
rect -1995 -12142 -1961 -11681
rect -1905 -11683 -1871 -11572
rect -2015 -12195 -2005 -12142
rect -1952 -12195 -1942 -12142
rect -1995 -12646 -1961 -12195
rect -2174 -12680 -1961 -12646
rect -1906 -12677 -1872 -12039
rect -2174 -12765 -2140 -12680
rect -1995 -12800 -1961 -12680
rect -1818 -12820 -1784 -10561
rect -1728 -11519 -1694 -11047
rect -1639 -11128 -1605 -10974
rect -1659 -11181 -1649 -11128
rect -1596 -11181 -1586 -11128
rect -1549 -11519 -1515 -11047
rect -1748 -11572 -1738 -11519
rect -1685 -11572 -1675 -11519
rect -1569 -11572 -1559 -11519
rect -1506 -11572 -1496 -11519
rect -1728 -11681 -1694 -11572
rect -1549 -11681 -1515 -11572
rect -1728 -12680 -1694 -12042
rect -1639 -12142 -1605 -11986
rect -1659 -12195 -1649 -12142
rect -1596 -12195 -1586 -12142
rect -1549 -12679 -1515 -12041
rect -1461 -12828 -1427 -10561
rect -1372 -10681 -1338 -10038
rect -1193 -10681 -1159 -10032
rect -1124 -10561 -1114 -10508
rect -1061 -10561 -1051 -10508
rect -1372 -11519 -1338 -11048
rect -1283 -11126 -1249 -10973
rect -1284 -11128 -1249 -11126
rect -1303 -11181 -1293 -11128
rect -1240 -11181 -1230 -11128
rect -1391 -11572 -1381 -11519
rect -1328 -11572 -1318 -11519
rect -1372 -11680 -1338 -11572
rect -1372 -12680 -1338 -12042
rect -1284 -12254 -1250 -11181
rect -1194 -11519 -1160 -11048
rect -1213 -11572 -1203 -11519
rect -1150 -11572 -1140 -11519
rect -1194 -11681 -1160 -11572
rect -1304 -12307 -1294 -12254
rect -1241 -12307 -1231 -12254
rect -1194 -12679 -1160 -12041
rect -1105 -12802 -1071 -10561
rect -1016 -10681 -982 -10032
rect -838 -10682 -804 -10033
rect -768 -10561 -758 -10508
rect -705 -10561 -695 -10508
rect -1016 -11519 -982 -11048
rect -927 -11128 -893 -10967
rect -947 -11181 -937 -11128
rect -884 -11181 -874 -11128
rect -838 -11519 -804 -11048
rect -1035 -11572 -1025 -11519
rect -972 -11572 -962 -11519
rect -858 -11572 -848 -11519
rect -795 -11572 -785 -11519
rect -1016 -11680 -982 -11572
rect -838 -11681 -804 -11572
rect -1016 -12680 -982 -12042
rect -927 -12383 -893 -11989
rect -947 -12436 -937 -12383
rect -884 -12436 -874 -12383
rect -927 -12774 -893 -12436
rect -838 -12679 -804 -12041
rect -749 -12822 -715 -10561
rect -659 -10681 -625 -10032
rect -482 -10681 -448 -10032
rect 853 -10038 887 -9968
rect 941 -10038 975 -10031
rect 1031 -10038 1065 -9960
rect 759 -10072 1159 -10038
rect 941 -10508 975 -10072
rect -412 -10561 -402 -10508
rect -349 -10561 -339 -10508
rect -56 -10561 -46 -10508
rect 7 -10561 17 -10508
rect 299 -10561 309 -10508
rect 362 -10561 372 -10508
rect 655 -10561 665 -10508
rect 718 -10561 728 -10508
rect 921 -10561 931 -10508
rect 984 -10561 994 -10508
rect 1189 -10561 1199 -10508
rect 1252 -10561 1262 -10508
rect -660 -11519 -626 -11048
rect -571 -11237 -537 -10988
rect -590 -11290 -580 -11237
rect -527 -11290 -517 -11237
rect -482 -11519 -448 -11048
rect -680 -11572 -670 -11519
rect -617 -11572 -607 -11519
rect -502 -11572 -492 -11519
rect -439 -11572 -429 -11519
rect -660 -11681 -626 -11572
rect -482 -11681 -448 -11572
rect -660 -12681 -626 -12043
rect -571 -12253 -537 -11987
rect -592 -12306 -582 -12253
rect -529 -12306 -519 -12253
rect -482 -12681 -448 -12043
rect -393 -12807 -359 -10561
rect -304 -11519 -270 -11048
rect -215 -11357 -181 -10985
rect -234 -11410 -224 -11357
rect -171 -11410 -161 -11357
rect -324 -11572 -314 -11519
rect -261 -11572 -251 -11519
rect -304 -11680 -270 -11572
rect -304 -12682 -270 -12044
rect -215 -12383 -181 -11410
rect -126 -11519 -92 -11048
rect -146 -11572 -136 -11519
rect -83 -11572 -73 -11519
rect -126 -11679 -92 -11572
rect -234 -12436 -224 -12383
rect -171 -12436 -161 -12383
rect -126 -12681 -92 -12043
rect -36 -12799 -2 -10561
rect 52 -11519 86 -11048
rect 141 -11357 175 -10987
rect 121 -11410 131 -11357
rect 184 -11410 194 -11357
rect 141 -11411 175 -11410
rect 230 -11519 264 -11048
rect 32 -11572 42 -11519
rect 95 -11572 105 -11519
rect 210 -11572 220 -11519
rect 273 -11572 283 -11519
rect 52 -11681 86 -11572
rect 230 -11680 264 -11572
rect 52 -12680 86 -12042
rect 141 -12253 175 -11984
rect 120 -12306 130 -12253
rect 183 -12306 193 -12253
rect -1995 -13145 -1961 -12983
rect -2014 -13198 -2004 -13145
rect -1951 -13198 -1941 -13145
rect -1905 -13682 -1871 -13044
rect -1728 -13681 -1694 -13043
rect -1638 -13272 -1604 -12985
rect -1658 -13325 -1648 -13272
rect -1595 -13325 -1585 -13272
rect -1550 -13682 -1516 -13044
rect -1282 -13272 -1248 -12983
rect -927 -13272 -893 -12987
rect -571 -13145 -537 -12985
rect -591 -13198 -581 -13145
rect -528 -13198 -518 -13145
rect -1301 -13325 -1291 -13272
rect -1238 -13325 -1228 -13272
rect -947 -13325 -937 -13272
rect -884 -13325 -874 -13272
rect -927 -13326 -893 -13325
rect -304 -13681 -270 -13037
rect -216 -13394 -182 -12986
rect -235 -13447 -225 -13394
rect -172 -13447 -162 -13394
rect -125 -13682 -91 -13038
rect 52 -13681 86 -13037
rect 141 -13394 175 -12306
rect 230 -12680 264 -12042
rect 319 -12807 353 -10561
rect 408 -11519 442 -11048
rect 497 -11357 531 -10980
rect 477 -11410 487 -11357
rect 540 -11410 550 -11357
rect 389 -11572 399 -11519
rect 452 -11572 462 -11519
rect 408 -11681 442 -11572
rect 408 -12682 442 -12044
rect 496 -12384 530 -11410
rect 586 -11519 620 -11048
rect 567 -11572 577 -11519
rect 630 -11572 640 -11519
rect 586 -11681 620 -11572
rect 476 -12437 486 -12384
rect 539 -12437 549 -12384
rect 587 -12682 621 -12044
rect 675 -12831 709 -10561
rect 941 -10680 975 -10561
rect 853 -11038 887 -10962
rect 942 -11038 976 -11032
rect 1031 -11038 1065 -10957
rect 757 -11072 1159 -11038
rect 764 -11681 798 -11632
rect 942 -11681 976 -11072
rect 1120 -11680 1154 -11632
rect 852 -12038 886 -11953
rect 942 -12038 976 -12032
rect 1031 -12038 1065 -11977
rect 759 -12072 1160 -12038
rect 942 -12648 976 -12072
rect 761 -12682 1160 -12648
rect 852 -12754 886 -12682
rect 1032 -12765 1066 -12682
rect 1209 -12812 1243 -10561
rect 1299 -10681 1333 -10032
rect 1477 -10681 1511 -10032
rect 1546 -10561 1556 -10508
rect 1609 -10561 1619 -10508
rect 1298 -11519 1332 -11048
rect 1387 -11128 1421 -10989
rect 1367 -11181 1377 -11128
rect 1430 -11181 1440 -11128
rect 1477 -11519 1511 -11048
rect 1278 -11572 1288 -11519
rect 1341 -11572 1351 -11519
rect 1458 -11572 1468 -11519
rect 1521 -11572 1531 -11519
rect 1298 -11680 1332 -11572
rect 1477 -11681 1511 -11572
rect 1299 -12681 1333 -12043
rect 1388 -12383 1422 -11989
rect 1368 -12436 1378 -12383
rect 1431 -12436 1441 -12383
rect 1388 -12787 1422 -12436
rect 1476 -12681 1510 -12043
rect 1566 -12817 1600 -10561
rect 1653 -10680 1687 -10031
rect 1832 -10682 1866 -10033
rect 1903 -10561 1913 -10508
rect 1966 -10561 1976 -10508
rect 1654 -11520 1688 -11048
rect 1743 -11128 1777 -10986
rect 1723 -11181 1733 -11128
rect 1786 -11181 1796 -11128
rect 1634 -11573 1644 -11520
rect 1697 -11573 1707 -11520
rect 1654 -11680 1688 -11573
rect 1655 -12682 1689 -12044
rect 1744 -12254 1778 -11181
rect 1832 -11519 1866 -11048
rect 1813 -11572 1823 -11519
rect 1876 -11572 1886 -11519
rect 1832 -11681 1866 -11572
rect 1725 -12307 1735 -12254
rect 1788 -12307 1798 -12254
rect 1833 -12681 1867 -12043
rect 1922 -12787 1956 -10561
rect 2010 -10681 2044 -10032
rect 2188 -10681 2222 -10032
rect 2258 -10561 2268 -10508
rect 2321 -10561 2331 -10508
rect 2613 -10561 2623 -10508
rect 2676 -10561 2686 -10508
rect 2970 -10561 2980 -10508
rect 3033 -10561 3043 -10508
rect 3325 -10561 3335 -10508
rect 3388 -10561 3398 -10508
rect 2010 -11519 2044 -11048
rect 2099 -11128 2133 -10980
rect 2079 -11181 2089 -11128
rect 2142 -11181 2152 -11128
rect 2188 -11519 2222 -11048
rect 1990 -11572 2000 -11519
rect 2053 -11572 2063 -11519
rect 2168 -11572 2178 -11519
rect 2231 -11572 2241 -11519
rect 2010 -11679 2044 -11572
rect 2188 -11679 2222 -11572
rect 2009 -12679 2043 -12041
rect 2098 -12382 2132 -11975
rect 2078 -12435 2088 -12382
rect 2141 -12435 2151 -12382
rect 2098 -12793 2132 -12435
rect 2188 -12679 2222 -12041
rect 2277 -12799 2311 -10561
rect 2366 -11519 2400 -11048
rect 2456 -11237 2490 -10986
rect 2436 -11290 2446 -11237
rect 2499 -11290 2509 -11237
rect 2544 -11519 2578 -11048
rect 2347 -11572 2357 -11519
rect 2410 -11572 2420 -11519
rect 2524 -11572 2534 -11519
rect 2587 -11572 2597 -11519
rect 2366 -11683 2400 -11572
rect 2544 -11681 2578 -11572
rect 2366 -12682 2400 -12044
rect 2455 -12253 2489 -11985
rect 2435 -12306 2445 -12253
rect 2498 -12306 2508 -12253
rect 2544 -12682 2578 -12044
rect 2633 -12804 2667 -10561
rect 2722 -11519 2756 -11048
rect 2810 -11357 2844 -10987
rect 2790 -11410 2800 -11357
rect 2853 -11410 2863 -11357
rect 2703 -11572 2713 -11519
rect 2766 -11572 2776 -11519
rect 2722 -11680 2756 -11572
rect 2722 -12679 2756 -12041
rect 2811 -12382 2845 -11410
rect 2900 -11519 2934 -11048
rect 2880 -11572 2890 -11519
rect 2943 -11572 2953 -11519
rect 2900 -11680 2934 -11572
rect 2791 -12435 2801 -12382
rect 2854 -12435 2864 -12382
rect 2900 -12682 2934 -12044
rect 2989 -12812 3023 -10561
rect 3078 -11519 3112 -11048
rect 3166 -11357 3200 -10984
rect 3147 -11410 3157 -11357
rect 3210 -11410 3220 -11357
rect 3256 -11519 3290 -11048
rect 3058 -11572 3068 -11519
rect 3121 -11572 3131 -11519
rect 3237 -11572 3247 -11519
rect 3300 -11572 3310 -11519
rect 3078 -11681 3112 -11572
rect 3256 -11680 3290 -11572
rect 3078 -12681 3112 -12043
rect 3167 -12250 3201 -11987
rect 3166 -12252 3201 -12250
rect 3148 -12305 3158 -12252
rect 3211 -12305 3221 -12252
rect 123 -13447 133 -13394
rect 186 -13447 196 -13394
rect 230 -13681 264 -13037
rect 408 -13681 442 -13037
rect 496 -13395 530 -12985
rect 477 -13448 487 -13395
rect 540 -13448 550 -13395
rect 587 -13681 621 -13037
rect 942 -13648 976 -13030
rect 1388 -13272 1422 -12980
rect 1743 -13272 1777 -12982
rect 2100 -13272 2134 -12982
rect 1369 -13325 1379 -13272
rect 1432 -13325 1442 -13272
rect 1722 -13325 1732 -13272
rect 1785 -13325 1795 -13272
rect 2081 -13325 2091 -13272
rect 2144 -13325 2154 -13272
rect 762 -13682 1159 -13648
rect 2366 -13681 2400 -13032
rect 2455 -13145 2489 -12988
rect 2436 -13198 2446 -13145
rect 2499 -13198 2509 -13145
rect 2544 -13681 2578 -13032
rect 2723 -13682 2757 -13033
rect 2812 -13394 2846 -12979
rect 2792 -13447 2802 -13394
rect 2855 -13447 2865 -13394
rect 2901 -13681 2935 -13032
rect 3078 -13682 3112 -13033
rect 3166 -13395 3200 -12305
rect 3256 -12682 3290 -12044
rect 3345 -12823 3379 -10561
rect 3434 -10682 3468 -10033
rect 3613 -10682 3647 -10033
rect 3682 -10561 3692 -10508
rect 3745 -10561 3755 -10508
rect 3434 -11519 3468 -11048
rect 3522 -11357 3556 -10969
rect 3503 -11410 3513 -11357
rect 3566 -11410 3576 -11357
rect 3612 -11519 3646 -11048
rect 3415 -11572 3425 -11519
rect 3478 -11572 3488 -11519
rect 3593 -11572 3603 -11519
rect 3656 -11572 3666 -11519
rect 3434 -11681 3468 -11572
rect 3612 -11680 3646 -11572
rect 3434 -12680 3468 -12042
rect 3524 -12142 3558 -11986
rect 3504 -12195 3514 -12142
rect 3567 -12195 3577 -12142
rect 3613 -12680 3647 -12042
rect 3701 -12813 3735 -10561
rect 3791 -10681 3825 -10032
rect 3881 -11037 3915 -10832
rect 4056 -11037 4090 -10965
rect 3790 -11519 3824 -11048
rect 3881 -11071 4090 -11037
rect 3881 -11238 3915 -11071
rect 3861 -11291 3871 -11238
rect 3924 -11291 3934 -11238
rect 3771 -11572 3781 -11519
rect 3834 -11572 3844 -11519
rect 3790 -11679 3824 -11572
rect 3881 -12036 3915 -11291
rect 4058 -12036 4092 -11963
rect 3790 -12680 3824 -12042
rect 3881 -12070 4092 -12036
rect 3881 -12142 3915 -12070
rect 3861 -12195 3871 -12142
rect 3924 -12195 3934 -12142
rect 3881 -12647 3915 -12195
rect 3881 -12681 4090 -12647
rect 3881 -12792 3915 -12681
rect 4056 -12765 4090 -12681
rect 3147 -13448 3157 -13395
rect 3210 -13448 3220 -13395
rect 3257 -13680 3291 -13031
rect 3523 -13394 3557 -12936
rect 3879 -13145 3913 -12987
rect 3860 -13198 3870 -13145
rect 3923 -13198 3933 -13145
rect 3502 -13447 3512 -13394
rect 3565 -13447 3575 -13394
rect 3523 -13448 3557 -13447
rect 853 -13760 887 -13682
rect 1032 -13764 1066 -13682
rect -2173 -14041 -2139 -13961
rect -1995 -14041 -1961 -13828
rect -2173 -14075 -1961 -14041
rect -2325 -14196 -2315 -14143
rect -2262 -14196 -2252 -14143
rect -1995 -14645 -1961 -14075
rect -2176 -14679 -1961 -14645
rect -2176 -14763 -2142 -14679
rect -2457 -15474 -2447 -15421
rect -2394 -15474 -2384 -15421
rect -1995 -15422 -1961 -14679
rect -2015 -15475 -2005 -15422
rect -1952 -15475 -1942 -15422
rect -3945 -15547 -3935 -15495
rect -3883 -15547 -3873 -15495
rect -6028 -16086 -5994 -15950
rect -5939 -16086 -5905 -15994
rect -5850 -16086 -5816 -15950
rect -5672 -16086 -5638 -15950
rect -6028 -16120 -5816 -16086
rect -5850 -16207 -5816 -16120
rect -5692 -16139 -5682 -16086
rect -5629 -16139 -5619 -16086
rect -6169 -16260 -6159 -16207
rect -6106 -16260 -6096 -16207
rect -5869 -16260 -5859 -16207
rect -5806 -16260 -5796 -16207
rect -5494 -16318 -5460 -15951
rect -5316 -16086 -5282 -15950
rect -5336 -16139 -5326 -16086
rect -5273 -16139 -5263 -16086
rect -5138 -16207 -5104 -15951
rect -4960 -16086 -4926 -15951
rect -4980 -16139 -4970 -16086
rect -4917 -16139 -4907 -16086
rect -5158 -16260 -5148 -16207
rect -5095 -16260 -5085 -16207
rect -5514 -16371 -5504 -16318
rect -5451 -16371 -5441 -16318
rect -4970 -16749 -4917 -16139
rect -4782 -16318 -4748 -15951
rect -4604 -16086 -4570 -15951
rect -4624 -16139 -4614 -16086
rect -4561 -16139 -4551 -16086
rect -4426 -16207 -4392 -15950
rect -4248 -16086 -4214 -15950
rect -4159 -16086 -4125 -15994
rect -4070 -16086 -4036 -15950
rect -4268 -16139 -4258 -16086
rect -4205 -16139 -4036 -16086
rect -4447 -16260 -4437 -16207
rect -4384 -16260 -4374 -16207
rect -3935 -16318 -3883 -15547
rect -1995 -15650 -1961 -15475
rect -1906 -15533 -1872 -15041
rect -1925 -15586 -1915 -15533
rect -1862 -15586 -1852 -15533
rect -2173 -15684 -1961 -15650
rect -2173 -15756 -2139 -15684
rect -1995 -15732 -1961 -15684
rect -1906 -16142 -1872 -16038
rect -1927 -16195 -1917 -16142
rect -1864 -16195 -1854 -16142
rect -1817 -16265 -1783 -13909
rect -1728 -15533 -1694 -15038
rect -1639 -15422 -1605 -13831
rect -1659 -15475 -1649 -15422
rect -1596 -15475 -1586 -15422
rect -1748 -15586 -1738 -15533
rect -1685 -15586 -1675 -15533
rect -1639 -15735 -1605 -15475
rect -1550 -15533 -1516 -15038
rect -1570 -15586 -1560 -15533
rect -1507 -15586 -1497 -15533
rect -1728 -16142 -1694 -16040
rect -1550 -16141 -1516 -16039
rect -1748 -16195 -1738 -16142
rect -1685 -16195 -1675 -16142
rect -1571 -16194 -1561 -16141
rect -1508 -16194 -1498 -16141
rect -1837 -16318 -1827 -16265
rect -1774 -16318 -1764 -16265
rect -1461 -16266 -1427 -13909
rect -1371 -14143 -1337 -14038
rect -1391 -14196 -1381 -14143
rect -1328 -14196 -1318 -14143
rect -1371 -14676 -1337 -14196
rect -1372 -15533 -1338 -15040
rect -1283 -15422 -1249 -13834
rect -1194 -14143 -1160 -14038
rect -1214 -14196 -1204 -14143
rect -1151 -14196 -1141 -14143
rect -1303 -15475 -1293 -15422
rect -1240 -15475 -1230 -15422
rect -1392 -15586 -1382 -15533
rect -1329 -15586 -1319 -15533
rect -1283 -15738 -1249 -15475
rect -1194 -15533 -1160 -15038
rect -1214 -15586 -1204 -15533
rect -1151 -15586 -1141 -15533
rect -1372 -16143 -1338 -16040
rect -1194 -16142 -1160 -16040
rect -1391 -16196 -1381 -16143
rect -1328 -16196 -1318 -16143
rect -1214 -16195 -1204 -16142
rect -1151 -16195 -1141 -16142
rect -1104 -16265 -1070 -13912
rect -1016 -14143 -982 -14039
rect -1036 -14196 -1026 -14143
rect -973 -14196 -963 -14143
rect -1015 -15533 -981 -15039
rect -927 -15422 -893 -13831
rect -838 -14143 -804 -14038
rect -858 -14196 -848 -14143
rect -795 -14196 -785 -14143
rect -857 -14579 -847 -14526
rect -794 -14579 -784 -14526
rect -838 -14681 -804 -14579
rect -947 -15475 -937 -15422
rect -884 -15475 -874 -15422
rect -1035 -15586 -1025 -15533
rect -972 -15586 -962 -15533
rect -927 -15735 -893 -15475
rect -857 -15586 -847 -15533
rect -794 -15586 -784 -15533
rect -838 -15680 -804 -15586
rect -1016 -16142 -982 -16039
rect -1036 -16195 -1026 -16142
rect -973 -16195 -963 -16142
rect -749 -16264 -715 -13910
rect -659 -14143 -625 -14040
rect -679 -14196 -669 -14143
rect -616 -14196 -606 -14143
rect -679 -14579 -669 -14526
rect -616 -14579 -606 -14526
rect -660 -14681 -626 -14579
rect -571 -15422 -537 -13831
rect -482 -14143 -448 -14039
rect -501 -14196 -491 -14143
rect -438 -14196 -428 -14143
rect -501 -14579 -491 -14526
rect -438 -14579 -428 -14526
rect -481 -14681 -447 -14579
rect -591 -15475 -581 -15422
rect -528 -15475 -518 -15422
rect -680 -15586 -670 -15533
rect -617 -15586 -607 -15533
rect -660 -15682 -626 -15586
rect -571 -15735 -537 -15475
rect -501 -15586 -491 -15533
rect -438 -15586 -428 -15533
rect -482 -15681 -448 -15586
rect -4802 -16371 -4792 -16318
rect -4739 -16371 -4729 -16318
rect -3945 -16370 -3935 -16318
rect -3883 -16370 -3873 -16318
rect -1481 -16319 -1471 -16266
rect -1418 -16319 -1408 -16266
rect -1124 -16318 -1114 -16265
rect -1061 -16318 -1051 -16265
rect -769 -16317 -759 -16264
rect -706 -16317 -696 -16264
rect -393 -16265 -359 -13906
rect -304 -14527 -270 -14037
rect -324 -14580 -314 -14527
rect -261 -14580 -251 -14527
rect -304 -14681 -270 -14580
rect -215 -15422 -181 -13830
rect -126 -14526 -92 -14040
rect -147 -14579 -137 -14526
rect -84 -14579 -74 -14526
rect -126 -14681 -92 -14579
rect -235 -15475 -225 -15422
rect -172 -15475 -162 -15422
rect -323 -15586 -313 -15533
rect -260 -15586 -250 -15533
rect -304 -15680 -270 -15586
rect -215 -15734 -181 -15475
rect -146 -15586 -136 -15533
rect -83 -15586 -73 -15533
rect -126 -15680 -92 -15586
rect -37 -16265 -3 -13912
rect 52 -14526 86 -14045
rect 33 -14579 43 -14526
rect 96 -14579 106 -14526
rect 52 -14681 86 -14579
rect 141 -15421 175 -13831
rect 122 -15474 132 -15421
rect 185 -15474 195 -15421
rect 33 -15586 43 -15533
rect 96 -15586 106 -15533
rect 52 -15680 86 -15586
rect 141 -15735 175 -15474
rect 230 -15533 264 -15039
rect 211 -15586 221 -15533
rect 274 -15586 284 -15533
rect 230 -16142 264 -16038
rect 210 -16195 220 -16142
rect 273 -16195 283 -16142
rect -413 -16318 -403 -16265
rect -350 -16318 -340 -16265
rect -57 -16318 -47 -16265
rect 6 -16318 16 -16265
rect 319 -16266 353 -13907
rect 408 -15533 442 -15039
rect 497 -15422 531 -13831
rect 477 -15475 487 -15422
rect 540 -15475 550 -15422
rect 388 -15586 398 -15533
rect 451 -15586 461 -15533
rect 497 -15735 531 -15475
rect 585 -15533 619 -15039
rect 565 -15586 575 -15533
rect 628 -15586 638 -15533
rect 408 -16142 442 -16039
rect 586 -16142 620 -16039
rect 387 -16195 397 -16142
rect 450 -16195 460 -16142
rect 566 -16195 576 -16142
rect 629 -16195 639 -16142
rect 675 -16265 709 -13907
rect 764 -15533 798 -15038
rect 853 -15422 887 -14940
rect 833 -15475 843 -15422
rect 896 -15475 906 -15422
rect 745 -15586 755 -15533
rect 808 -15586 818 -15533
rect 853 -15736 887 -15475
rect 941 -15533 975 -15039
rect 921 -15586 931 -15533
rect 984 -15586 994 -15533
rect 765 -16142 799 -16038
rect 943 -16142 977 -16039
rect 745 -16195 755 -16142
rect 808 -16195 818 -16142
rect 923 -16195 933 -16142
rect 986 -16195 996 -16142
rect 1031 -16265 1065 -13908
rect 1120 -15533 1154 -15040
rect 1209 -15422 1243 -13831
rect 1298 -14143 1332 -14039
rect 1278 -14196 1288 -14143
rect 1341 -14196 1351 -14143
rect 1279 -14580 1289 -14527
rect 1342 -14580 1352 -14527
rect 1298 -14681 1332 -14580
rect 1191 -15475 1201 -15422
rect 1254 -15475 1264 -15422
rect 1100 -15586 1110 -15533
rect 1163 -15586 1173 -15533
rect 1209 -15735 1243 -15475
rect 1279 -15586 1289 -15533
rect 1342 -15586 1352 -15533
rect 1298 -15681 1332 -15586
rect 1120 -16142 1154 -16039
rect 1101 -16195 1111 -16142
rect 1164 -16195 1174 -16142
rect 1387 -16265 1421 -13907
rect 1477 -14143 1511 -14039
rect 1456 -14196 1466 -14143
rect 1519 -14196 1529 -14143
rect 1457 -14579 1467 -14526
rect 1520 -14579 1530 -14526
rect 1476 -14681 1510 -14579
rect 1565 -15422 1599 -13831
rect 1654 -14143 1688 -14038
rect 1634 -14196 1644 -14143
rect 1697 -14196 1707 -14143
rect 1634 -14579 1644 -14526
rect 1697 -14579 1707 -14526
rect 1654 -14682 1688 -14579
rect 1545 -15475 1555 -15422
rect 1608 -15475 1618 -15422
rect 1456 -15586 1466 -15533
rect 1519 -15586 1529 -15533
rect 1476 -15682 1510 -15586
rect 1565 -15735 1599 -15475
rect 1633 -15586 1643 -15533
rect 1696 -15586 1706 -15533
rect 1653 -15681 1687 -15586
rect 1744 -16265 1778 -13912
rect 1832 -14142 1866 -14038
rect 1813 -14195 1823 -14142
rect 1876 -14195 1886 -14142
rect 1812 -14579 1822 -14526
rect 1875 -14579 1885 -14526
rect 1833 -14681 1867 -14579
rect 1921 -15422 1955 -13831
rect 2010 -14143 2044 -14038
rect 1990 -14196 2000 -14143
rect 2053 -14196 2063 -14143
rect 1989 -14579 1999 -14526
rect 2052 -14579 2062 -14526
rect 2010 -14682 2044 -14579
rect 1900 -15475 1910 -15422
rect 1963 -15475 1973 -15422
rect 1812 -15586 1822 -15533
rect 1875 -15586 1885 -15533
rect 1832 -15680 1866 -15586
rect 1921 -15735 1955 -15475
rect 1990 -15586 2000 -15533
rect 2053 -15586 2063 -15533
rect 2010 -15681 2044 -15586
rect 2100 -16264 2134 -13913
rect 2188 -14143 2222 -14039
rect 2168 -14196 2178 -14143
rect 2231 -14196 2241 -14143
rect 2170 -14579 2180 -14526
rect 2233 -14579 2243 -14526
rect 2189 -14681 2223 -14579
rect 2277 -15422 2311 -13831
rect 2257 -15475 2267 -15422
rect 2320 -15475 2330 -15422
rect 2169 -15586 2179 -15533
rect 2232 -15586 2242 -15533
rect 2189 -15681 2223 -15586
rect 2277 -15735 2311 -15475
rect 2366 -15533 2400 -15040
rect 2346 -15586 2356 -15533
rect 2409 -15586 2419 -15533
rect 2366 -16142 2400 -16039
rect 2346 -16195 2356 -16142
rect 2409 -16195 2419 -16142
rect 299 -16319 309 -16266
rect 362 -16319 372 -16266
rect 655 -16318 665 -16265
rect 718 -16318 728 -16265
rect 835 -16318 845 -16265
rect 898 -16318 908 -16265
rect 1011 -16318 1021 -16265
rect 1074 -16318 1084 -16265
rect 1367 -16318 1377 -16265
rect 1430 -16318 1440 -16265
rect 1725 -16318 1735 -16265
rect 1788 -16318 1798 -16265
rect 2080 -16317 2090 -16264
rect 2143 -16317 2153 -16264
rect 2455 -16265 2489 -13911
rect 2544 -15533 2578 -15040
rect 2633 -15422 2667 -13832
rect 2614 -15475 2624 -15422
rect 2677 -15475 2687 -15422
rect 2524 -15586 2534 -15533
rect 2587 -15586 2597 -15533
rect 2633 -15736 2667 -15475
rect 2722 -15533 2756 -15040
rect 2702 -15586 2712 -15533
rect 2765 -15586 2775 -15533
rect 2544 -16142 2578 -16039
rect 2722 -16141 2756 -16041
rect 2524 -16195 2534 -16142
rect 2587 -16195 2597 -16142
rect 2703 -16194 2713 -16141
rect 2766 -16194 2776 -16141
rect 2811 -16265 2845 -13910
rect 2900 -15533 2934 -15039
rect 2989 -15422 3023 -13831
rect 2969 -15475 2979 -15422
rect 3032 -15475 3042 -15422
rect 2881 -15586 2891 -15533
rect 2944 -15586 2954 -15533
rect 2989 -15735 3023 -15475
rect 3078 -15533 3112 -15038
rect 3058 -15586 3068 -15533
rect 3121 -15586 3131 -15533
rect 2901 -16142 2935 -16041
rect 3079 -16142 3113 -16039
rect 2881 -16195 2891 -16142
rect 2944 -16195 2954 -16142
rect 3060 -16195 3070 -16142
rect 3123 -16195 3133 -16142
rect 3167 -16264 3201 -13915
rect 3236 -14197 3246 -14144
rect 3299 -14197 3309 -14144
rect 3256 -14680 3290 -14197
rect 3256 -15533 3290 -15039
rect 3345 -15422 3379 -13831
rect 3434 -14143 3468 -14039
rect 3414 -14196 3424 -14143
rect 3477 -14196 3487 -14143
rect 3415 -14579 3425 -14526
rect 3478 -14579 3488 -14526
rect 3434 -14681 3468 -14579
rect 3325 -15475 3335 -15422
rect 3388 -15475 3398 -15422
rect 3237 -15586 3247 -15533
rect 3300 -15586 3310 -15533
rect 3345 -15735 3379 -15475
rect 3414 -15586 3424 -15533
rect 3477 -15586 3487 -15533
rect 3434 -15681 3468 -15586
rect 3257 -16142 3291 -16040
rect 3239 -16195 3249 -16142
rect 3302 -16195 3312 -16142
rect 2435 -16318 2445 -16265
rect 2498 -16318 2508 -16265
rect 2791 -16318 2801 -16265
rect 2854 -16318 2864 -16265
rect 3147 -16317 3157 -16264
rect 3210 -16317 3220 -16264
rect 3524 -16266 3558 -13910
rect 3612 -14143 3646 -14039
rect 3592 -14196 3602 -14143
rect 3655 -14196 3665 -14143
rect 3593 -14579 3603 -14526
rect 3656 -14579 3666 -14526
rect 3612 -14682 3646 -14579
rect 3701 -15422 3735 -13832
rect 3879 -14039 3913 -13907
rect 4057 -14039 4091 -13957
rect 3791 -14143 3825 -14039
rect 3879 -14073 4091 -14039
rect 3771 -14196 3781 -14143
rect 3834 -14196 3844 -14143
rect 3770 -14579 3780 -14526
rect 3833 -14579 3843 -14526
rect 3790 -14682 3824 -14579
rect 3879 -14647 3913 -14073
rect 4905 -14145 4958 -5265
rect 5037 -12896 5090 -5059
rect 5174 -6767 5184 -6714
rect 5237 -6767 5247 -6714
rect 5184 -6819 5237 -6767
rect 5185 -8235 5237 -6819
rect 5175 -8287 5185 -8235
rect 5237 -8287 5247 -8235
rect 11647 -8316 11681 -8315
rect 6690 -8360 6815 -8326
rect 6690 -8507 6724 -8360
rect 6781 -8444 6815 -8360
rect 11044 -8369 11054 -8316
rect 11107 -8369 11117 -8316
rect 11335 -8369 11345 -8316
rect 11398 -8369 11408 -8316
rect 11628 -8369 11638 -8316
rect 11691 -8369 11701 -8316
rect 11922 -8369 11932 -8316
rect 11985 -8369 11995 -8316
rect 12212 -8369 12222 -8316
rect 12275 -8369 12285 -8316
rect 9004 -8442 9395 -8408
rect 6513 -8801 6547 -8725
rect 6689 -8801 6723 -8554
rect 6513 -8835 6723 -8801
rect 6779 -8914 6813 -8798
rect 6759 -8967 6769 -8914
rect 6822 -8967 6832 -8914
rect 6669 -9198 6679 -9145
rect 6732 -9198 6742 -9145
rect 6513 -9699 6547 -9617
rect 6690 -9699 6724 -9198
rect 6779 -9340 6813 -8967
rect 6513 -9733 6724 -9699
rect 6690 -9913 6724 -9733
rect 6670 -9966 6680 -9913
rect 6733 -9966 6743 -9913
rect 6868 -10067 6902 -8642
rect 6957 -8915 6991 -8797
rect 6937 -8968 6947 -8915
rect 7000 -8968 7010 -8915
rect 6957 -9221 6991 -8968
rect 7046 -9221 7080 -8646
rect 7135 -8915 7169 -8798
rect 7116 -8968 7126 -8915
rect 7179 -8968 7189 -8915
rect 6957 -9255 7080 -9221
rect 6957 -9343 6991 -9255
rect 6848 -10120 6858 -10067
rect 6911 -10120 6921 -10067
rect 6510 -10603 6544 -10510
rect 6688 -10603 6722 -10520
rect 6868 -10603 6902 -10120
rect 6958 -10243 6992 -9697
rect 6510 -10637 6902 -10603
rect 6511 -11500 6545 -11423
rect 6688 -11500 6722 -11419
rect 6868 -11500 6902 -10637
rect 6958 -11144 6992 -10595
rect 7046 -10966 7080 -9255
rect 7135 -9344 7169 -8968
rect 7136 -10243 7170 -9697
rect 7224 -10066 7258 -8649
rect 7313 -8913 7347 -8797
rect 7293 -8966 7303 -8913
rect 7356 -8966 7366 -8913
rect 7313 -9343 7347 -8966
rect 7204 -10119 7214 -10066
rect 7267 -10119 7277 -10066
rect 7027 -11019 7037 -10966
rect 7090 -11019 7100 -10966
rect 7046 -11271 7080 -11019
rect 7135 -11143 7169 -10594
rect 6511 -11534 6902 -11500
rect 6868 -11640 6902 -11534
rect 7224 -11640 7258 -10119
rect 7313 -10244 7347 -9698
rect 7313 -11142 7347 -10593
rect 7402 -10966 7436 -8648
rect 7491 -8913 7525 -8798
rect 7472 -8966 7482 -8913
rect 7535 -8966 7545 -8913
rect 7491 -9344 7525 -8966
rect 7492 -10243 7526 -9697
rect 7580 -10066 7614 -8651
rect 7669 -8915 7703 -8798
rect 7649 -8968 7659 -8915
rect 7712 -8968 7722 -8915
rect 7669 -9344 7703 -8968
rect 7561 -10119 7571 -10066
rect 7624 -10119 7634 -10066
rect 7383 -11019 7393 -10966
rect 7446 -11019 7456 -10966
rect 7402 -11273 7436 -11019
rect 7491 -11142 7525 -10593
rect 7580 -11640 7614 -10119
rect 7669 -10244 7703 -9698
rect 7669 -11142 7703 -10593
rect 7758 -10967 7792 -8654
rect 7847 -8914 7881 -8798
rect 7827 -8967 7837 -8914
rect 7890 -8967 7900 -8914
rect 7847 -9344 7881 -8967
rect 7847 -10243 7881 -9697
rect 7936 -10066 7970 -8651
rect 8025 -8915 8059 -8798
rect 8005 -8968 8015 -8915
rect 8068 -8968 8078 -8915
rect 8025 -9344 8059 -8968
rect 7917 -10119 7927 -10066
rect 7980 -10119 7990 -10066
rect 7738 -11020 7748 -10967
rect 7801 -11020 7811 -10967
rect 7758 -11279 7792 -11020
rect 7848 -11142 7882 -10593
rect 7936 -11640 7970 -10119
rect 8025 -10243 8059 -9697
rect 8024 -11143 8058 -10594
rect 8113 -10966 8147 -8656
rect 8203 -8914 8237 -8798
rect 8184 -8967 8194 -8914
rect 8247 -8967 8257 -8914
rect 8203 -9344 8237 -8967
rect 8203 -10242 8237 -9696
rect 8292 -10067 8326 -8660
rect 8381 -8914 8415 -8798
rect 8361 -8967 8371 -8914
rect 8424 -8967 8434 -8914
rect 8381 -9344 8415 -8967
rect 8273 -10120 8283 -10067
rect 8336 -10120 8346 -10067
rect 8093 -11019 8103 -10966
rect 8156 -11019 8166 -10966
rect 8113 -11281 8147 -11019
rect 8203 -11144 8237 -10595
rect 8292 -11640 8326 -10120
rect 8382 -10244 8416 -9698
rect 8381 -11143 8415 -10594
rect 8470 -10966 8504 -8656
rect 8559 -8914 8593 -8798
rect 8539 -8967 8549 -8914
rect 8602 -8967 8612 -8914
rect 8559 -9344 8593 -8967
rect 8559 -10242 8593 -9696
rect 8648 -10066 8682 -8664
rect 8737 -8915 8771 -8798
rect 8717 -8968 8727 -8915
rect 8780 -8968 8790 -8915
rect 8737 -9344 8771 -8968
rect 8628 -10119 8638 -10066
rect 8691 -10119 8701 -10066
rect 8451 -11019 8461 -10966
rect 8514 -11019 8524 -10966
rect 8470 -11281 8504 -11019
rect 8559 -11143 8593 -10594
rect 8648 -11640 8682 -10119
rect 8737 -10244 8771 -9698
rect 8737 -11143 8771 -10594
rect 8826 -10966 8860 -8663
rect 9004 -8668 9038 -8442
rect 9183 -8526 9217 -8442
rect 9361 -8523 9395 -8442
rect 8915 -8914 8949 -8798
rect 8896 -8967 8906 -8914
rect 8959 -8967 8969 -8914
rect 8915 -9344 8949 -8967
rect 9004 -9309 9038 -8713
rect 11063 -8745 11097 -8369
rect 11354 -8586 11388 -8369
rect 11647 -8581 11681 -8369
rect 11941 -8611 11975 -8369
rect 12231 -8440 12265 -8369
rect 12231 -8474 12738 -8440
rect 12231 -8613 12265 -8474
rect 12522 -8547 12556 -8474
rect 12704 -8553 12738 -8474
rect 10968 -8752 11097 -8745
rect 10772 -8830 10806 -8756
rect 10950 -8779 11097 -8752
rect 10950 -8830 10984 -8779
rect 10772 -8864 10984 -8830
rect 10861 -9238 10895 -8864
rect 11063 -8987 11097 -8779
rect 11154 -8974 11188 -8859
rect 11134 -8987 11144 -8974
rect 11063 -9021 11144 -8987
rect 11134 -9027 11144 -9021
rect 11197 -9027 11207 -8974
rect 11154 -9242 11188 -9027
rect 9004 -9343 9394 -9309
rect 11242 -9316 11276 -8780
rect 11445 -8975 11479 -8852
rect 11426 -9028 11436 -8975
rect 11489 -9028 11499 -8975
rect 11445 -9235 11479 -9028
rect 11534 -9306 11568 -8770
rect 11738 -8975 11772 -8856
rect 11718 -9028 11728 -8975
rect 11781 -9028 11791 -8975
rect 11738 -9239 11772 -9028
rect 11825 -9311 11859 -8775
rect 12030 -8976 12064 -8851
rect 12010 -9029 12020 -8976
rect 12073 -9029 12083 -8976
rect 12030 -9234 12064 -9029
rect 12118 -9304 12152 -8768
rect 12321 -8975 12355 -8852
rect 12302 -9028 12312 -8975
rect 12365 -9028 12375 -8975
rect 12321 -9235 12355 -9028
rect 12410 -9318 12444 -8782
rect 12613 -9210 12647 -8828
rect 12525 -9244 12736 -9210
rect 12525 -9337 12559 -9244
rect 12702 -9331 12736 -9244
rect 8915 -10243 8949 -9697
rect 9004 -10067 9038 -9343
rect 9182 -9424 9216 -9343
rect 9360 -9433 9394 -9343
rect 10773 -9601 10807 -9526
rect 10951 -9601 10985 -9512
rect 10773 -9635 10985 -9601
rect 9161 -9967 9171 -9914
rect 9224 -9967 9234 -9914
rect 8985 -10120 8995 -10067
rect 9048 -10120 9058 -10067
rect 8807 -11019 8817 -10966
rect 8870 -11019 8880 -10966
rect 8826 -11288 8860 -11019
rect 8915 -11143 8949 -10594
rect 9004 -11279 9038 -10120
rect 9181 -10214 9215 -9967
rect 10862 -9980 10896 -9635
rect 10772 -10014 10986 -9980
rect 10772 -10085 10806 -10014
rect 10952 -10107 10986 -10014
rect 11063 -10090 11097 -9554
rect 11153 -10000 11187 -9617
rect 11356 -10081 11390 -9541
rect 11446 -10000 11480 -9617
rect 11648 -10086 11682 -9546
rect 11737 -10000 11771 -9617
rect 11940 -10082 11974 -9542
rect 12028 -9999 12062 -9616
rect 12232 -10088 12266 -9548
rect 12320 -9998 12354 -9615
rect 12613 -10013 12647 -9599
rect 9181 -10248 9393 -10214
rect 9181 -10295 9215 -10248
rect 9359 -10326 9393 -10248
rect 9093 -11141 9127 -10605
rect 10772 -10749 10806 -10748
rect 10860 -10749 10894 -10385
rect 10772 -10783 10986 -10749
rect 11152 -10775 11186 -10392
rect 10772 -10853 10806 -10783
rect 10952 -10868 10986 -10783
rect 11244 -10860 11278 -10320
rect 11446 -10771 11480 -10388
rect 11534 -10858 11568 -10318
rect 11737 -10773 11771 -10390
rect 11826 -10860 11860 -10320
rect 12029 -10772 12063 -10389
rect 12118 -10863 12152 -10323
rect 12322 -10771 12356 -10388
rect 12410 -10863 12444 -10323
rect 12525 -10372 12559 -10249
rect 12613 -10372 12647 -10370
rect 12700 -10372 12734 -10281
rect 12525 -10406 12734 -10372
rect 12613 -10784 12647 -10406
rect 9182 -11144 9394 -11110
rect 8912 -11585 8946 -11500
rect 9095 -11585 9129 -11500
rect 9182 -11585 9216 -11144
rect 9360 -11233 9394 -11144
rect 11063 -11274 11097 -10983
rect 11043 -11327 11053 -11274
rect 11106 -11327 11116 -11274
rect 11356 -11275 11390 -11017
rect 11648 -11274 11682 -11002
rect 11940 -11274 11974 -11005
rect 12233 -11274 12267 -11003
rect 12525 -11141 12559 -10996
rect 12701 -11141 12735 -11060
rect 12525 -11175 12735 -11141
rect 11337 -11328 11347 -11275
rect 11400 -11328 11410 -11275
rect 11628 -11327 11638 -11274
rect 11691 -11327 11701 -11274
rect 11921 -11327 11931 -11274
rect 11984 -11327 11994 -11274
rect 12213 -11327 12223 -11274
rect 12276 -11327 12286 -11274
rect 8912 -11619 9216 -11585
rect 6868 -11674 8682 -11640
rect 5027 -12949 5037 -12896
rect 5090 -12949 5100 -12896
rect 5524 -12949 5534 -12896
rect 5587 -12949 5597 -12896
rect 5021 -13086 5031 -13033
rect 5084 -13086 5094 -13033
rect 4895 -14198 4905 -14145
rect 4958 -14198 4968 -14145
rect 4229 -14579 4239 -14526
rect 4292 -14579 4302 -14526
rect 3879 -14681 4091 -14647
rect 3682 -15475 3692 -15422
rect 3745 -15475 3755 -15422
rect 3593 -15586 3603 -15533
rect 3656 -15586 3666 -15533
rect 3612 -15680 3646 -15586
rect 3701 -15736 3735 -15475
rect 3770 -15586 3780 -15533
rect 3833 -15586 3843 -15533
rect 3790 -15680 3824 -15586
rect 3879 -15647 3913 -14681
rect 4057 -14769 4091 -14681
rect 4238 -15139 4291 -14579
rect 4228 -15192 4238 -15139
rect 4291 -15192 4301 -15139
rect 5031 -15140 5084 -13086
rect 5390 -13198 5400 -13145
rect 5453 -13198 5463 -13145
rect 5132 -13447 5142 -13394
rect 5195 -13447 5205 -13394
rect 5142 -14258 5195 -13447
rect 5133 -14311 5143 -14258
rect 5196 -14311 5206 -14258
rect 3879 -15681 4090 -15647
rect 3879 -16265 3913 -15681
rect 4056 -15770 4090 -15681
rect 4238 -16142 4291 -15192
rect 5021 -15193 5031 -15140
rect 5084 -15193 5094 -15140
rect 4228 -16195 4238 -16142
rect 4291 -16195 4301 -16142
rect 846 -16774 899 -16318
rect 3504 -16319 3514 -16266
rect 3567 -16319 3577 -16266
rect 3858 -16318 3868 -16265
rect 3921 -16318 3931 -16265
rect 5031 -16382 5084 -15193
rect 5400 -15253 5453 -13198
rect 5534 -13272 5587 -12949
rect 5524 -13325 5534 -13272
rect 5587 -13325 5597 -13272
rect 6912 -13522 6946 -11674
rect 8940 -13086 8950 -13033
rect 9003 -13086 9013 -13033
rect 9295 -13086 9305 -13033
rect 9358 -13086 9368 -13033
rect 8762 -13209 8772 -13156
rect 8825 -13209 8835 -13156
rect 7516 -13325 7526 -13272
rect 7579 -13325 7589 -13272
rect 7338 -13449 7348 -13396
rect 7401 -13449 7411 -13396
rect 5823 -13575 5833 -13522
rect 5886 -13575 5896 -13522
rect 6003 -13575 6013 -13522
rect 6066 -13575 6076 -13522
rect 5577 -13682 5790 -13648
rect 5843 -13678 5877 -13575
rect 6022 -13680 6056 -13575
rect 6180 -13576 6190 -13523
rect 6243 -13576 6253 -13523
rect 6359 -13575 6369 -13522
rect 6422 -13575 6432 -13522
rect 6200 -13680 6234 -13576
rect 6378 -13680 6412 -13575
rect 6537 -13576 6547 -13523
rect 6600 -13576 6610 -13523
rect 6715 -13575 6725 -13522
rect 6778 -13575 6788 -13522
rect 6892 -13575 6902 -13522
rect 6955 -13575 6965 -13522
rect 6556 -13680 6590 -13576
rect 6734 -13681 6768 -13575
rect 6912 -13679 6946 -13575
rect 7103 -13682 7297 -13648
rect 5577 -13764 5611 -13682
rect 5756 -14145 5790 -13682
rect 7179 -13761 7213 -13682
rect 5736 -14198 5746 -14145
rect 5799 -14198 5809 -14145
rect 5575 -14681 5789 -14647
rect 5843 -14675 5877 -14042
rect 5933 -14258 5967 -13988
rect 5914 -14311 5924 -14258
rect 5977 -14311 5987 -14258
rect 6022 -14680 6056 -14047
rect 6111 -14145 6145 -13992
rect 6091 -14198 6101 -14145
rect 6154 -14198 6164 -14145
rect 6200 -14679 6234 -14046
rect 6289 -14258 6323 -13987
rect 6269 -14311 6279 -14258
rect 6332 -14311 6342 -14258
rect 6378 -14681 6412 -14048
rect 6468 -14145 6502 -13988
rect 6449 -14198 6459 -14145
rect 6512 -14198 6522 -14145
rect 6557 -14681 6591 -14048
rect 6645 -14258 6679 -13987
rect 6823 -14145 6857 -13987
rect 6803 -14198 6813 -14145
rect 6866 -14198 6876 -14145
rect 7000 -14258 7034 -13997
rect 6626 -14311 6636 -14258
rect 6689 -14311 6699 -14258
rect 6981 -14311 6991 -14258
rect 7044 -14311 7054 -14258
rect 7179 -14349 7213 -13987
rect 6822 -14383 7213 -14349
rect 5575 -14772 5609 -14681
rect 5755 -15139 5789 -14681
rect 5735 -15192 5745 -15139
rect 5798 -15192 5808 -15139
rect 5390 -15306 5400 -15253
rect 5453 -15306 5463 -15253
rect 5400 -16267 5453 -15306
rect 5737 -15403 5747 -15350
rect 5800 -15403 5810 -15350
rect 5576 -16038 5610 -15953
rect 5756 -16038 5790 -15403
rect 5844 -15681 5878 -15048
rect 5933 -15252 5967 -14976
rect 5913 -15305 5923 -15252
rect 5976 -15305 5986 -15252
rect 5911 -15601 5921 -15548
rect 5974 -15601 5984 -15548
rect 5931 -15733 5965 -15601
rect 6022 -15682 6056 -15049
rect 6111 -15139 6145 -14980
rect 6091 -15192 6101 -15139
rect 6154 -15192 6164 -15139
rect 6091 -15402 6101 -15349
rect 6154 -15402 6164 -15349
rect 6112 -15736 6146 -15402
rect 6201 -15682 6235 -15049
rect 6289 -15252 6323 -14964
rect 6269 -15305 6279 -15252
rect 6332 -15305 6342 -15252
rect 6269 -15601 6279 -15548
rect 6332 -15601 6342 -15548
rect 6288 -15737 6322 -15601
rect 6379 -15681 6413 -15048
rect 6468 -15139 6502 -14975
rect 6448 -15192 6458 -15139
rect 6511 -15192 6521 -15139
rect 6446 -15403 6456 -15350
rect 6509 -15403 6519 -15350
rect 6467 -15737 6501 -15403
rect 6556 -15681 6590 -15048
rect 6645 -15252 6679 -14957
rect 6822 -14968 6856 -14383
rect 7357 -14424 7391 -13449
rect 7427 -13575 7437 -13522
rect 7490 -13575 7500 -13522
rect 7446 -13681 7480 -13575
rect 6983 -14477 6993 -14424
rect 7046 -14477 7056 -14424
rect 7337 -14477 7347 -14424
rect 7400 -14477 7410 -14424
rect 6822 -15038 6857 -14968
rect 6748 -15072 6942 -15038
rect 6625 -15305 6635 -15252
rect 6688 -15305 6698 -15252
rect 6703 -15404 6713 -15351
rect 6766 -15404 6776 -15351
rect 6624 -15601 6634 -15548
rect 6687 -15601 6697 -15548
rect 6734 -15556 6768 -15404
rect 6822 -15451 6856 -15072
rect 6803 -15504 6813 -15451
rect 6866 -15504 6876 -15451
rect 7002 -15551 7036 -14477
rect 7070 -14576 7080 -14523
rect 7133 -14576 7143 -14523
rect 7090 -14680 7124 -14576
rect 7250 -14577 7260 -14524
rect 7313 -14577 7323 -14524
rect 7269 -14680 7303 -14577
rect 7357 -14782 7391 -14477
rect 7447 -14523 7481 -14048
rect 7429 -14576 7439 -14523
rect 7492 -14576 7502 -14523
rect 7447 -14681 7481 -14576
rect 7535 -14763 7569 -13325
rect 7872 -13326 7882 -13273
rect 7935 -13326 7945 -13273
rect 8228 -13324 8238 -13271
rect 8291 -13324 8301 -13271
rect 7694 -13448 7704 -13395
rect 7757 -13448 7767 -13395
rect 7605 -13575 7615 -13522
rect 7668 -13575 7678 -13522
rect 7624 -13680 7658 -13575
rect 7713 -13730 7747 -13448
rect 7783 -13576 7793 -13523
rect 7846 -13576 7856 -13523
rect 7802 -13681 7836 -13576
rect 7892 -13724 7926 -13326
rect 8051 -13449 8061 -13396
rect 8114 -13449 8124 -13396
rect 7960 -13575 7970 -13522
rect 8023 -13575 8033 -13522
rect 7980 -13681 8014 -13575
rect 8069 -13734 8103 -13449
rect 8138 -13575 8148 -13522
rect 8201 -13575 8211 -13522
rect 8158 -13681 8192 -13575
rect 8248 -13737 8282 -13324
rect 8405 -13449 8415 -13396
rect 8468 -13449 8478 -13396
rect 8316 -13575 8326 -13522
rect 8379 -13575 8389 -13522
rect 8336 -13680 8370 -13575
rect 8425 -13742 8459 -13449
rect 8529 -13682 8723 -13648
rect 8603 -13765 8637 -13682
rect 8781 -13729 8815 -13209
rect 8851 -13575 8861 -13522
rect 8914 -13575 8924 -13522
rect 8871 -13681 8905 -13575
rect 8960 -13731 8994 -13086
rect 9117 -13209 9127 -13156
rect 9180 -13209 9190 -13156
rect 9028 -13575 9038 -13522
rect 9091 -13575 9101 -13522
rect 9048 -13681 9082 -13575
rect 9137 -13734 9171 -13209
rect 9207 -13575 9217 -13522
rect 9270 -13575 9280 -13522
rect 9227 -13681 9261 -13575
rect 9315 -13730 9349 -13086
rect 9473 -13209 9483 -13156
rect 9536 -13209 9546 -13156
rect 9384 -13575 9394 -13522
rect 9447 -13575 9457 -13522
rect 9404 -13681 9438 -13575
rect 9493 -13732 9527 -13209
rect 11432 -13325 11442 -13272
rect 11495 -13325 11505 -13272
rect 11788 -13325 11798 -13272
rect 11851 -13325 11861 -13272
rect 11254 -13449 11264 -13396
rect 11317 -13449 11327 -13396
rect 9919 -13576 9929 -13523
rect 9982 -13576 9992 -13523
rect 10098 -13575 10108 -13522
rect 10161 -13575 10171 -13522
rect 9594 -13682 9788 -13648
rect 9938 -13681 9972 -13576
rect 10117 -13682 10151 -13575
rect 10274 -13576 10284 -13523
rect 10337 -13576 10347 -13523
rect 10452 -13576 10462 -13523
rect 10515 -13576 10525 -13523
rect 10630 -13575 10640 -13522
rect 10693 -13575 10703 -13522
rect 10294 -13682 10328 -13576
rect 10472 -13681 10506 -13576
rect 10650 -13681 10684 -13575
rect 10809 -13576 10819 -13523
rect 10872 -13576 10882 -13523
rect 10828 -13681 10862 -13576
rect 11018 -13682 11212 -13648
rect 9671 -13759 9705 -13682
rect 11095 -13758 11129 -13682
rect 7625 -14681 7659 -14048
rect 7694 -14478 7704 -14425
rect 7757 -14478 7767 -14425
rect 7714 -14735 7748 -14478
rect 7802 -14681 7836 -14048
rect 8226 -14198 8236 -14145
rect 8289 -14198 8299 -14145
rect 8050 -14474 8060 -14421
rect 8113 -14474 8123 -14421
rect 7179 -15350 7213 -14984
rect 7159 -15403 7169 -15350
rect 7222 -15403 7232 -15350
rect 7159 -15505 7169 -15452
rect 7222 -15505 7232 -15452
rect 6734 -15590 6858 -15556
rect 6644 -15745 6678 -15601
rect 6824 -15763 6858 -15590
rect 6984 -15604 6994 -15551
rect 7047 -15604 7057 -15551
rect 7002 -15873 7036 -15604
rect 7178 -16038 7212 -15505
rect 7447 -15680 7481 -15047
rect 7536 -15349 7570 -14982
rect 7516 -15402 7526 -15349
rect 7579 -15402 7589 -15349
rect 7516 -15606 7526 -15553
rect 7579 -15606 7589 -15553
rect 7535 -15747 7569 -15606
rect 7624 -15681 7658 -15048
rect 7803 -15681 7837 -15048
rect 7891 -15349 7925 -14969
rect 8069 -15038 8103 -14474
rect 8000 -15072 8194 -15038
rect 7872 -15402 7882 -15349
rect 7935 -15402 7945 -15349
rect 8069 -15451 8103 -15072
rect 8050 -15504 8060 -15451
rect 8113 -15504 8123 -15451
rect 8247 -15552 8281 -14198
rect 8336 -14523 8370 -14048
rect 8407 -14310 8417 -14257
rect 8470 -14310 8480 -14257
rect 8317 -14576 8327 -14523
rect 8380 -14576 8390 -14523
rect 8336 -14681 8370 -14576
rect 7871 -15605 7881 -15552
rect 7934 -15605 7944 -15552
rect 8227 -15605 8237 -15552
rect 8290 -15605 8300 -15552
rect 7891 -15767 7925 -15605
rect 8247 -15821 8281 -15605
rect 8336 -15680 8370 -15047
rect 5576 -16072 5790 -16038
rect 6557 -16144 6591 -16041
rect 6735 -16144 6769 -16040
rect 6538 -16197 6548 -16144
rect 6601 -16197 6611 -16144
rect 6716 -16197 6726 -16144
rect 6779 -16197 6789 -16144
rect 6912 -16145 6946 -16042
rect 7101 -16072 7295 -16038
rect 6893 -16198 6903 -16145
rect 6956 -16198 6966 -16145
rect 5389 -16320 5399 -16267
rect 5452 -16320 5462 -16267
rect 5021 -16435 5031 -16382
rect 5084 -16435 5094 -16382
rect 7357 -16490 7391 -15942
rect 7713 -16490 7747 -15945
rect 7980 -16145 8014 -16053
rect 7960 -16198 7970 -16145
rect 8023 -16198 8033 -16145
rect 8069 -16490 8103 -15982
rect 8158 -16144 8192 -16045
rect 8139 -16197 8149 -16144
rect 8202 -16197 8212 -16144
rect 8426 -16490 8460 -14310
rect 8514 -14406 8548 -14038
rect 8585 -14198 8595 -14145
rect 8648 -14198 8658 -14145
rect 8494 -14459 8504 -14406
rect 8557 -14459 8567 -14406
rect 8514 -14471 8548 -14459
rect 8495 -14577 8505 -14524
rect 8558 -14577 8568 -14524
rect 8514 -14680 8548 -14577
rect 8604 -14736 8638 -14198
rect 8762 -14311 8772 -14258
rect 8825 -14311 8835 -14258
rect 8692 -14524 8726 -14523
rect 8673 -14577 8683 -14524
rect 8736 -14577 8746 -14524
rect 8692 -14680 8726 -14577
rect 8781 -14748 8815 -14311
rect 8870 -14681 8904 -14048
rect 8940 -14199 8950 -14146
rect 9003 -14199 9013 -14146
rect 8960 -14739 8994 -14199
rect 9048 -14681 9082 -14048
rect 9117 -14312 9127 -14259
rect 9180 -14312 9190 -14259
rect 9137 -14740 9171 -14312
rect 9226 -14681 9260 -14048
rect 9294 -14198 9304 -14145
rect 9357 -14198 9367 -14145
rect 9314 -14744 9348 -14198
rect 9404 -14681 9438 -14048
rect 9651 -14198 9661 -14145
rect 9714 -14198 9724 -14145
rect 9473 -14311 9483 -14258
rect 9536 -14311 9546 -14258
rect 9493 -14735 9527 -14311
rect 9562 -14576 9572 -14523
rect 9625 -14576 9635 -14523
rect 9582 -14677 9616 -14576
rect 9671 -14739 9705 -14198
rect 9763 -14406 9797 -14053
rect 9848 -14259 9882 -13983
rect 9827 -14312 9837 -14259
rect 9890 -14312 9900 -14259
rect 9743 -14459 9753 -14406
rect 9806 -14459 9816 -14406
rect 9763 -14471 9797 -14459
rect 9740 -14576 9750 -14523
rect 9803 -14576 9813 -14523
rect 9760 -14678 9794 -14576
rect 9848 -14800 9882 -14312
rect 9939 -14523 9973 -14049
rect 10026 -14145 10060 -13984
rect 10006 -14198 10016 -14145
rect 10069 -14198 10079 -14145
rect 9919 -14576 9929 -14523
rect 9982 -14576 9992 -14523
rect 9939 -14682 9973 -14576
rect 10026 -14816 10060 -14198
rect 10205 -14258 10239 -13985
rect 10383 -14146 10417 -13985
rect 10363 -14199 10373 -14146
rect 10426 -14199 10436 -14146
rect 10186 -14311 10196 -14258
rect 10249 -14311 10259 -14258
rect 10185 -14475 10195 -14422
rect 10248 -14475 10258 -14422
rect 10205 -15038 10239 -14475
rect 10472 -14681 10506 -14048
rect 10560 -14258 10594 -13983
rect 10540 -14311 10550 -14258
rect 10603 -14311 10613 -14258
rect 10542 -14468 10552 -14415
rect 10605 -14468 10615 -14415
rect 10561 -14736 10595 -14468
rect 10650 -14681 10684 -14048
rect 10738 -14145 10772 -13983
rect 10719 -14198 10729 -14145
rect 10782 -14198 10792 -14145
rect 10828 -14523 10862 -14048
rect 10917 -14258 10951 -13987
rect 11096 -14258 11130 -13934
rect 10898 -14311 10908 -14258
rect 10961 -14311 10971 -14258
rect 11077 -14311 11087 -14258
rect 11140 -14311 11150 -14258
rect 10898 -14466 10908 -14413
rect 10961 -14466 10971 -14413
rect 11273 -14415 11307 -13449
rect 11343 -13575 11353 -13522
rect 11406 -13575 11416 -13522
rect 11362 -13681 11396 -13575
rect 11452 -13733 11486 -13325
rect 11610 -13450 11620 -13397
rect 11673 -13450 11683 -13397
rect 11520 -13575 11530 -13522
rect 11583 -13575 11593 -13522
rect 11540 -13680 11574 -13575
rect 11630 -13735 11664 -13450
rect 11699 -13575 11709 -13522
rect 11762 -13575 11772 -13522
rect 11719 -13681 11753 -13575
rect 11807 -13733 11841 -13325
rect 12142 -13326 12152 -13273
rect 12205 -13326 12215 -13273
rect 12499 -13325 12509 -13272
rect 12562 -13325 12572 -13272
rect 11967 -13449 11977 -13396
rect 12030 -13449 12040 -13396
rect 11876 -13576 11886 -13523
rect 11939 -13576 11949 -13523
rect 11895 -13680 11929 -13576
rect 11986 -13731 12020 -13449
rect 12054 -13575 12064 -13522
rect 12117 -13575 12127 -13522
rect 12073 -13682 12107 -13575
rect 12162 -13737 12196 -13326
rect 12324 -13449 12334 -13396
rect 12387 -13449 12397 -13396
rect 12232 -13576 12242 -13523
rect 12295 -13576 12305 -13523
rect 12252 -13681 12286 -13576
rect 12342 -13733 12376 -13449
rect 12410 -13575 12420 -13522
rect 12473 -13575 12483 -13522
rect 12430 -13681 12464 -13575
rect 12519 -13648 12553 -13325
rect 12519 -13682 12731 -13648
rect 12519 -13734 12553 -13682
rect 12697 -13754 12731 -13682
rect 11430 -14309 11440 -14256
rect 11493 -14309 11503 -14256
rect 10809 -14576 10819 -14523
rect 10872 -14576 10882 -14523
rect 10828 -14681 10862 -14576
rect 8583 -15505 8593 -15452
rect 8646 -15505 8656 -15452
rect 8603 -16038 8637 -15505
rect 8870 -15680 8904 -15047
rect 9049 -15681 9083 -15048
rect 9226 -15680 9260 -15047
rect 9404 -15680 9438 -15047
rect 9653 -15505 9663 -15452
rect 9716 -15505 9726 -15452
rect 8519 -16072 8713 -16038
rect 8781 -16266 8815 -15986
rect 8761 -16319 8771 -16266
rect 8824 -16319 8834 -16266
rect 8960 -16382 8994 -15989
rect 9138 -16266 9172 -15983
rect 9118 -16319 9128 -16266
rect 9181 -16319 9191 -16266
rect 9315 -16382 9349 -15993
rect 9493 -16266 9527 -15980
rect 9672 -16038 9706 -15505
rect 9939 -15681 9973 -15048
rect 10122 -15072 10316 -15038
rect 10205 -15452 10239 -15072
rect 10383 -15351 10417 -14949
rect 10363 -15404 10373 -15351
rect 10426 -15404 10436 -15351
rect 10184 -15505 10194 -15452
rect 10247 -15505 10257 -15452
rect 10472 -15680 10506 -15047
rect 10650 -15680 10684 -15047
rect 10739 -15350 10773 -14959
rect 10720 -15403 10730 -15350
rect 10783 -15403 10793 -15350
rect 10739 -15838 10773 -15403
rect 10828 -15680 10862 -15047
rect 10916 -15815 10950 -14466
rect 11254 -14468 11264 -14415
rect 11317 -14468 11327 -14415
rect 10986 -14576 10996 -14523
rect 11049 -14576 11059 -14523
rect 11165 -14576 11175 -14523
rect 11228 -14576 11238 -14523
rect 11006 -14661 11040 -14576
rect 11184 -14663 11218 -14576
rect 11273 -14789 11307 -14468
rect 11095 -15350 11129 -14948
rect 11451 -15038 11485 -14309
rect 11717 -14678 11751 -14039
rect 11897 -14679 11931 -14040
rect 12075 -14679 12109 -14040
rect 12253 -14681 12287 -14042
rect 12430 -14681 12464 -14042
rect 12520 -14683 12730 -14649
rect 11390 -15072 11584 -15038
rect 11076 -15403 11086 -15350
rect 11139 -15403 11149 -15350
rect 11451 -15441 11485 -15072
rect 11629 -15252 11663 -14992
rect 11609 -15305 11619 -15252
rect 11672 -15305 11682 -15252
rect 11629 -15306 11663 -15305
rect 11074 -15505 11084 -15452
rect 11137 -15505 11147 -15452
rect 11430 -15494 11440 -15441
rect 11493 -15494 11503 -15441
rect 11451 -15502 11485 -15494
rect 9595 -16072 9789 -16038
rect 9474 -16319 9484 -16266
rect 9537 -16319 9547 -16266
rect 8940 -16435 8950 -16382
rect 9003 -16435 9013 -16382
rect 9295 -16435 9305 -16382
rect 9358 -16435 9368 -16382
rect 7337 -16543 7347 -16490
rect 7400 -16543 7410 -16490
rect 7694 -16543 7704 -16490
rect 7757 -16543 7767 -16490
rect 8050 -16543 8060 -16490
rect 8113 -16543 8123 -16490
rect 8406 -16543 8416 -16490
rect 8469 -16543 8479 -16490
rect 9672 -16883 9706 -16072
rect 9848 -16266 9882 -15949
rect 9938 -16144 9972 -16058
rect 9919 -16197 9929 -16144
rect 9982 -16197 9992 -16144
rect 9828 -16319 9838 -16266
rect 9891 -16319 9901 -16266
rect 10028 -16381 10062 -15983
rect 10117 -16145 10151 -16056
rect 10097 -16198 10107 -16145
rect 10160 -16198 10170 -16145
rect 10205 -16265 10239 -15934
rect 10296 -16145 10330 -16058
rect 10277 -16198 10287 -16145
rect 10340 -16198 10350 -16145
rect 10185 -16318 10195 -16265
rect 10248 -16318 10258 -16265
rect 10383 -16381 10417 -15977
rect 10561 -16265 10595 -15952
rect 10540 -16318 10550 -16265
rect 10603 -16318 10613 -16265
rect 10739 -16379 10773 -15959
rect 10917 -16265 10951 -15977
rect 11094 -16037 11128 -15505
rect 11431 -15605 11441 -15552
rect 11494 -15605 11504 -15552
rect 11451 -15738 11485 -15605
rect 11718 -15681 11752 -15048
rect 11808 -15140 11842 -14994
rect 11788 -15193 11798 -15140
rect 11851 -15193 11861 -15140
rect 11787 -15605 11797 -15552
rect 11850 -15605 11860 -15552
rect 11806 -15736 11840 -15605
rect 11897 -15681 11931 -15048
rect 11985 -15252 12019 -14987
rect 11965 -15305 11975 -15252
rect 12028 -15305 12038 -15252
rect 12074 -15680 12108 -15047
rect 12165 -15139 12199 -14972
rect 12145 -15192 12155 -15139
rect 12208 -15192 12218 -15139
rect 12144 -15605 12154 -15552
rect 12207 -15605 12217 -15552
rect 12163 -15736 12197 -15605
rect 12252 -15681 12286 -15048
rect 12342 -15252 12376 -14986
rect 12322 -15305 12332 -15252
rect 12385 -15305 12395 -15252
rect 12431 -15681 12465 -15048
rect 12520 -15139 12554 -14683
rect 12696 -14754 12730 -14683
rect 12501 -15192 12511 -15139
rect 12564 -15192 12574 -15139
rect 12501 -15605 12511 -15552
rect 12564 -15605 12574 -15552
rect 11019 -16071 11213 -16037
rect 10897 -16318 10907 -16265
rect 10960 -16318 10970 -16265
rect 10007 -16434 10017 -16381
rect 10070 -16434 10080 -16381
rect 10364 -16434 10374 -16381
rect 10427 -16434 10437 -16381
rect 10721 -16432 10731 -16379
rect 10784 -16432 10794 -16379
rect 11273 -16490 11307 -15940
rect 11362 -16145 11396 -16055
rect 11342 -16198 11352 -16145
rect 11405 -16198 11415 -16145
rect 11540 -16146 11574 -16053
rect 11520 -16199 11530 -16146
rect 11583 -16199 11593 -16146
rect 11630 -16490 11664 -15962
rect 11718 -16145 11752 -16057
rect 11699 -16198 11709 -16145
rect 11762 -16198 11772 -16145
rect 11985 -16489 12019 -15953
rect 12340 -16489 12374 -15980
rect 12520 -16040 12554 -15605
rect 12698 -16040 12732 -15956
rect 12520 -16074 12732 -16040
rect 11253 -16543 11263 -16490
rect 11316 -16543 11326 -16490
rect 11610 -16543 11620 -16490
rect 11673 -16543 11683 -16490
rect 11965 -16542 11975 -16489
rect 12028 -16542 12038 -16489
rect 12321 -16542 12331 -16489
rect 12384 -16542 12394 -16489
<< via1 >>
rect -5867 -1963 -5814 -1910
rect -5689 -1963 -5636 -1910
rect -5510 -1963 -5457 -1910
rect -5333 -1963 -5280 -1910
rect -5155 -1963 -5102 -1910
rect -4976 -1963 -4923 -1910
rect -4799 -1963 -4746 -1910
rect -4621 -1963 -4568 -1910
rect -4443 -1963 -4390 -1910
rect -4265 -1963 -4212 -1910
rect -4086 -1963 -4033 -1910
rect -3909 -1963 -3856 -1910
rect -1109 -1963 -1056 -1910
rect -6498 -2582 -6445 -2529
rect -6625 -3454 -6572 -3401
rect -6044 -2833 -5991 -2780
rect -6134 -3454 -6081 -3401
rect -6498 -3693 -6445 -3640
rect -6498 -4324 -6445 -4271
rect -6134 -4443 -6081 -4390
rect -6498 -5194 -6445 -5141
rect -6625 -5375 -6572 -5322
rect -6134 -5285 -6081 -5232
rect -5777 -2583 -5724 -2530
rect -5866 -2833 -5813 -2780
rect -5777 -3569 -5724 -3516
rect -5778 -4324 -5725 -4271
rect -5777 -5468 -5724 -5415
rect -5421 -2721 -5368 -2668
rect -5422 -3693 -5369 -3640
rect -5422 -4559 -5369 -4506
rect -5422 -5194 -5369 -5141
rect -5066 -2583 -5013 -2530
rect -5066 -3454 -5013 -3401
rect -5066 -4443 -5013 -4390
rect -5066 -5286 -5013 -5233
rect -4710 -2721 -4657 -2668
rect -4710 -3454 -4657 -3401
rect -4709 -4443 -4656 -4390
rect -4710 -5375 -4657 -5322
rect -4354 -2583 -4301 -2530
rect -4353 -3693 -4300 -3640
rect -4353 -4559 -4300 -4506
rect -4353 -5194 -4300 -5141
rect -3998 -2721 -3945 -2668
rect -1109 -2478 -1056 -2425
rect -752 -2478 -699 -2425
rect -3908 -2833 -3855 -2780
rect -3998 -3569 -3945 -3516
rect -3998 -4324 -3945 -4271
rect -3997 -5468 -3944 -5415
rect -2624 -2611 -2571 -2558
rect -1285 -2611 -1232 -2558
rect -3298 -2721 -3245 -2668
rect -3731 -2833 -3678 -2780
rect -3642 -3454 -3589 -3401
rect -3131 -3454 -3078 -3401
rect -3298 -3569 -3245 -3516
rect -3642 -4443 -3589 -4390
rect -3298 -4559 -3245 -4506
rect -3642 -5372 -3589 -5319
rect -3130 -5286 -3077 -5233
rect -1197 -2718 -1144 -2665
rect -930 -2611 -877 -2558
rect -1019 -2718 -966 -2665
rect -841 -2718 -788 -2665
rect -129 -2718 -76 -2665
rect 50 -2718 103 -2665
rect 227 -2718 280 -2665
rect 1919 -2479 1972 -2426
rect 2275 -2479 2328 -2426
rect 940 -2718 993 -2665
rect 1117 -2718 1170 -2665
rect 1295 -2718 1348 -2665
rect -1645 -3510 -1584 -3449
rect -2004 -4465 -1951 -4412
rect -2624 -5377 -2571 -5324
rect -3298 -5469 -3245 -5416
rect -5956 -6069 -5903 -6016
rect -5601 -6069 -5548 -6016
rect -5778 -6184 -5725 -6131
rect -5244 -6069 -5191 -6016
rect -5065 -6184 -5012 -6131
rect -6498 -6301 -6445 -6248
rect -5421 -6301 -5368 -6248
rect -4888 -6069 -4835 -6016
rect -4710 -6301 -4657 -6248
rect -4532 -6069 -4479 -6016
rect -4175 -6069 -4122 -6016
rect -4354 -6184 -4301 -6131
rect -3820 -6069 -3767 -6016
rect -2624 -6060 -2571 -6007
rect -3298 -6184 -3245 -6131
rect -3998 -6300 -3945 -6247
rect -4786 -6431 -4733 -6378
rect -1876 -5285 -1823 -5232
rect -1286 -3624 -1233 -3571
rect -1108 -3509 -1055 -3456
rect -929 -3624 -876 -3571
rect -484 -3354 -431 -3301
rect -750 -3509 -697 -3456
rect -396 -3509 -343 -3456
rect -573 -3624 -520 -3571
rect -217 -3624 -164 -3571
rect 583 -3354 636 -3301
rect -39 -3509 14 -3456
rect 317 -3509 370 -3456
rect 850 -3509 903 -3456
rect 1206 -3509 1259 -3456
rect 2097 -2607 2150 -2554
rect 2007 -2718 2060 -2665
rect 2186 -2718 2239 -2665
rect 3193 -2480 3246 -2427
rect 2453 -2607 2506 -2554
rect 2363 -2718 2416 -2665
rect 1654 -3354 1707 -3301
rect 1562 -3509 1615 -3456
rect 1919 -3509 1972 -3456
rect 1384 -3617 1437 -3564
rect 1741 -3617 1794 -3564
rect 2097 -3617 2150 -3564
rect 2275 -3509 2328 -3456
rect 2451 -3617 2504 -3564
rect -841 -4245 -788 -4192
rect -662 -4245 -609 -4192
rect -483 -4245 -430 -4192
rect -306 -4245 -253 -4192
rect -1287 -5150 -1234 -5097
rect -1646 -5339 -1585 -5278
rect -1105 -5266 -1052 -5213
rect -929 -5150 -876 -5097
rect -572 -5150 -519 -5097
rect -218 -5150 -165 -5097
rect -751 -5266 -698 -5213
rect -396 -5266 -343 -5213
rect -1876 -6417 -1823 -6364
rect -1282 -6417 -1229 -6364
rect -928 -6417 -876 -6365
rect -1110 -6532 -1057 -6479
rect -752 -6532 -699 -6479
rect 407 -4245 460 -4192
rect 317 -4357 370 -4304
rect 583 -4245 636 -4192
rect 495 -4465 548 -4412
rect 761 -4245 814 -4192
rect 673 -4357 726 -4304
rect 850 -4465 903 -4412
rect 1474 -4245 1527 -4192
rect 1652 -4245 1705 -4192
rect 1830 -4245 1883 -4192
rect 2008 -4245 2061 -4192
rect 2538 -4327 2599 -4266
rect 2746 -4507 2807 -4446
rect -41 -5266 12 -5213
rect 316 -5266 369 -5213
rect -128 -5433 -75 -5380
rect 50 -5433 103 -5380
rect 228 -5433 281 -5380
rect 850 -5266 903 -5213
rect 1207 -5266 1260 -5213
rect 940 -5434 993 -5381
rect 1119 -5433 1172 -5380
rect 1385 -5146 1438 -5093
rect 1296 -5433 1349 -5380
rect 227 -6303 280 -6250
rect 1740 -5146 1793 -5093
rect 1563 -5266 1616 -5213
rect 1917 -5266 1970 -5213
rect 2096 -5146 2149 -5093
rect 2274 -5266 2327 -5213
rect 2453 -5146 2506 -5093
rect 942 -6303 995 -6250
rect 2096 -6060 2149 -6007
rect 2452 -6060 2505 -6007
rect 1918 -6177 1971 -6124
rect 2275 -6177 2328 -6124
rect 3194 -4857 3246 -4805
rect 4771 -4857 4823 -4805
rect 2879 -6417 2931 -6365
rect 5037 -5059 5090 -5006
rect 4905 -5265 4958 -5212
rect -753 -6651 -700 -6598
rect 4772 -6650 4825 -6597
rect -3874 -6806 -3821 -6753
rect -2003 -6767 -1950 -6714
rect -3731 -6956 -3678 -6903
rect -3541 -7440 -3489 -7388
rect -5502 -11524 -5449 -11471
rect -6077 -11765 -6024 -11712
rect -5626 -11765 -5573 -11712
rect -6223 -12315 -6170 -12262
rect -6426 -13105 -6373 -13052
rect -5000 -11525 -4947 -11472
rect -4502 -11524 -4449 -11471
rect -5376 -11641 -5323 -11588
rect -5127 -11641 -5074 -11588
rect -4877 -11765 -4824 -11712
rect -4627 -11765 -4574 -11712
rect -4377 -11641 -4324 -11588
rect -3928 -11642 -3875 -11589
rect -5751 -12315 -5698 -12262
rect -5251 -12442 -5198 -12389
rect -4752 -12315 -4699 -12262
rect -4251 -12442 -4198 -12389
rect -6077 -12998 -6024 -12945
rect -5376 -12998 -5323 -12945
rect -5626 -13105 -5573 -13052
rect -5730 -13210 -5677 -13157
rect -5126 -12998 -5073 -12945
rect -4877 -13105 -4824 -13052
rect -4376 -12998 -4323 -12945
rect -4627 -13105 -4574 -13052
rect -4752 -13210 -4699 -13157
rect -3788 -12442 -3735 -12389
rect -3928 -13105 -3875 -13052
rect -3788 -13210 -3735 -13157
rect -6223 -13308 -6170 -13255
rect -5250 -13308 -5197 -13255
rect -4250 -13308 -4197 -13255
rect -6159 -14048 -6106 -13995
rect -5860 -14048 -5807 -13995
rect -5504 -14154 -5451 -14101
rect -6159 -14735 -6106 -14682
rect -5860 -14841 -5807 -14788
rect -5504 -14734 -5451 -14681
rect -6159 -15446 -6106 -15393
rect -5860 -15547 -5807 -15494
rect -5504 -15446 -5451 -15393
rect -5147 -14048 -5094 -13995
rect -5148 -14842 -5095 -14789
rect -5148 -15547 -5095 -15494
rect -4791 -14154 -4738 -14101
rect -4792 -14734 -4739 -14681
rect -4792 -15446 -4739 -15393
rect -4436 -14048 -4383 -13995
rect -3382 -7586 -3329 -7533
rect -1382 -7575 -1329 -7522
rect -3542 -12442 -3489 -12389
rect -1203 -7576 -1150 -7523
rect -1025 -7575 -972 -7522
rect -848 -7575 -795 -7522
rect -670 -7575 -617 -7522
rect -490 -7575 -437 -7522
rect 755 -7575 808 -7522
rect 932 -7575 985 -7522
rect 1112 -7575 1165 -7522
rect 1289 -7576 1342 -7523
rect 1467 -7575 1520 -7522
rect 1644 -7575 1697 -7522
rect 2890 -7575 2943 -7522
rect 3069 -7575 3122 -7522
rect 3247 -7575 3300 -7522
rect 3424 -7575 3477 -7522
rect 3603 -7576 3656 -7523
rect 3778 -7575 3831 -7522
rect 4208 -7576 4261 -7523
rect -1916 -8187 -1863 -8134
rect -1739 -8187 -1686 -8134
rect -1826 -8306 -1773 -8253
rect -2447 -8420 -2394 -8367
rect -2005 -8420 -1952 -8367
rect -2315 -9578 -2262 -9525
rect -2447 -11525 -2394 -11472
rect -3382 -13308 -3329 -13255
rect -3936 -14154 -3883 -14101
rect -4435 -14841 -4383 -14789
rect -4436 -15547 -4383 -15494
rect -3935 -14841 -3883 -14789
rect -1916 -9199 -1863 -9146
rect -1916 -9578 -1863 -9525
rect -1558 -8187 -1505 -8134
rect -1382 -8187 -1329 -8134
rect -1470 -8306 -1417 -8253
rect -1648 -8420 -1595 -8367
rect -1738 -9199 -1685 -9146
rect -1738 -9579 -1685 -9526
rect -1558 -9199 -1505 -9146
rect -1560 -9578 -1507 -9525
rect -1203 -8187 -1150 -8134
rect -1293 -8420 -1240 -8367
rect -1382 -9577 -1329 -9524
rect -1026 -8187 -973 -8134
rect -1115 -8306 -1062 -8253
rect -848 -8187 -795 -8134
rect -936 -8420 -883 -8367
rect -670 -8187 -617 -8134
rect -758 -8306 -705 -8253
rect -491 -8187 -438 -8134
rect -580 -8419 -527 -8366
rect -314 -8187 -261 -8134
rect -402 -8306 -349 -8253
rect -136 -8187 -83 -8134
rect 42 -8187 95 -8134
rect -47 -8306 6 -8253
rect -225 -8420 -172 -8367
rect -312 -9199 -259 -9146
rect -314 -9578 -261 -9525
rect -136 -9198 -83 -9145
rect -136 -9579 -83 -9526
rect 221 -8187 274 -8134
rect 398 -8187 451 -8134
rect 310 -8306 363 -8253
rect 132 -8421 185 -8368
rect 42 -9199 95 -9146
rect 43 -9578 96 -9525
rect 222 -9198 275 -9145
rect 220 -9578 273 -9525
rect 577 -8187 630 -8134
rect 754 -8187 807 -8134
rect 666 -8306 719 -8253
rect 489 -8419 542 -8366
rect 399 -9199 452 -9146
rect 398 -9578 451 -9525
rect 577 -9199 630 -9146
rect 576 -9578 629 -9525
rect 932 -8187 985 -8134
rect 843 -8419 896 -8366
rect 1111 -8187 1164 -8134
rect 1022 -8306 1075 -8253
rect 1289 -8187 1342 -8134
rect 1201 -8420 1254 -8367
rect 1466 -8187 1519 -8134
rect 1377 -8306 1430 -8253
rect 1644 -8187 1697 -8134
rect 1556 -8420 1609 -8367
rect 1822 -8187 1875 -8134
rect 1733 -8306 1786 -8253
rect 2000 -8187 2053 -8134
rect 2178 -8187 2231 -8134
rect 2090 -8306 2143 -8253
rect 1911 -8420 1964 -8367
rect 2357 -8187 2410 -8134
rect 2534 -8187 2587 -8134
rect 2446 -8306 2499 -8253
rect 2267 -8420 2320 -8367
rect 2178 -9200 2231 -9147
rect 2357 -9199 2410 -9146
rect 2356 -9578 2409 -9525
rect 2712 -8187 2765 -8134
rect 2890 -8187 2943 -8134
rect 2802 -8306 2855 -8253
rect 2624 -8420 2677 -8367
rect 2534 -9199 2587 -9146
rect 2534 -9578 2587 -9525
rect 2713 -9199 2766 -9146
rect 2712 -9579 2765 -9526
rect 3068 -8187 3121 -8134
rect 2980 -8420 3033 -8367
rect 2891 -9578 2944 -9525
rect 3246 -8187 3299 -8134
rect 3158 -8306 3211 -8253
rect 3069 -9578 3122 -9525
rect 3424 -8187 3477 -8134
rect 3336 -8420 3389 -8367
rect 3246 -9578 3299 -9525
rect 3602 -8187 3655 -8134
rect 3513 -8306 3566 -8253
rect 3781 -8187 3834 -8134
rect 3692 -8420 3745 -8367
rect 3869 -8306 3922 -8253
rect 4771 -8967 4824 -8914
rect 4208 -9199 4261 -9146
rect -1827 -10561 -1774 -10508
rect -1470 -10561 -1417 -10508
rect -2004 -11290 -1951 -11237
rect -1915 -11572 -1862 -11519
rect -2005 -12195 -1952 -12142
rect -1649 -11181 -1596 -11128
rect -1738 -11572 -1685 -11519
rect -1559 -11572 -1506 -11519
rect -1649 -12195 -1596 -12142
rect -1114 -10561 -1061 -10508
rect -1293 -11181 -1240 -11128
rect -1381 -11572 -1328 -11519
rect -1203 -11572 -1150 -11519
rect -1294 -12307 -1241 -12254
rect -758 -10561 -705 -10508
rect -937 -11181 -884 -11128
rect -1025 -11572 -972 -11519
rect -848 -11572 -795 -11519
rect -937 -12436 -884 -12383
rect -402 -10561 -349 -10508
rect -46 -10561 7 -10508
rect 309 -10561 362 -10508
rect 665 -10561 718 -10508
rect 931 -10561 984 -10508
rect 1199 -10561 1252 -10508
rect -580 -11290 -527 -11237
rect -670 -11572 -617 -11519
rect -492 -11572 -439 -11519
rect -582 -12306 -529 -12253
rect -224 -11410 -171 -11357
rect -314 -11572 -261 -11519
rect -136 -11572 -83 -11519
rect -224 -12436 -171 -12383
rect 131 -11410 184 -11357
rect 42 -11572 95 -11519
rect 220 -11572 273 -11519
rect 130 -12306 183 -12253
rect -2004 -13198 -1951 -13145
rect -1648 -13325 -1595 -13272
rect -581 -13198 -528 -13145
rect -1291 -13325 -1238 -13272
rect -937 -13325 -884 -13272
rect -225 -13447 -172 -13394
rect 487 -11410 540 -11357
rect 399 -11572 452 -11519
rect 577 -11572 630 -11519
rect 486 -12437 539 -12384
rect 1556 -10561 1609 -10508
rect 1377 -11181 1430 -11128
rect 1288 -11572 1341 -11519
rect 1468 -11572 1521 -11519
rect 1378 -12436 1431 -12383
rect 1913 -10561 1966 -10508
rect 1733 -11181 1786 -11128
rect 1644 -11573 1697 -11520
rect 1823 -11572 1876 -11519
rect 1735 -12307 1788 -12254
rect 2268 -10561 2321 -10508
rect 2623 -10561 2676 -10508
rect 2980 -10561 3033 -10508
rect 3335 -10561 3388 -10508
rect 2089 -11181 2142 -11128
rect 2000 -11572 2053 -11519
rect 2178 -11572 2231 -11519
rect 2088 -12435 2141 -12382
rect 2446 -11290 2499 -11237
rect 2357 -11572 2410 -11519
rect 2534 -11572 2587 -11519
rect 2445 -12306 2498 -12253
rect 2800 -11410 2853 -11357
rect 2713 -11572 2766 -11519
rect 2890 -11572 2943 -11519
rect 2801 -12435 2854 -12382
rect 3157 -11410 3210 -11357
rect 3068 -11572 3121 -11519
rect 3247 -11572 3300 -11519
rect 3158 -12305 3211 -12252
rect 133 -13447 186 -13394
rect 487 -13448 540 -13395
rect 1379 -13325 1432 -13272
rect 1732 -13325 1785 -13272
rect 2091 -13325 2144 -13272
rect 2446 -13198 2499 -13145
rect 2802 -13447 2855 -13394
rect 3692 -10561 3745 -10508
rect 3513 -11410 3566 -11357
rect 3425 -11572 3478 -11519
rect 3603 -11572 3656 -11519
rect 3514 -12195 3567 -12142
rect 3871 -11291 3924 -11238
rect 3781 -11572 3834 -11519
rect 3871 -12195 3924 -12142
rect 3157 -13448 3210 -13395
rect 3870 -13198 3923 -13145
rect 3512 -13447 3565 -13394
rect -2315 -14196 -2262 -14143
rect -2447 -15474 -2394 -15421
rect -2005 -15475 -1952 -15422
rect -3935 -15547 -3883 -15495
rect -5682 -16139 -5629 -16086
rect -6159 -16260 -6106 -16207
rect -5859 -16260 -5806 -16207
rect -5326 -16139 -5273 -16086
rect -4970 -16139 -4917 -16086
rect -5148 -16260 -5095 -16207
rect -5504 -16371 -5451 -16318
rect -4614 -16139 -4561 -16086
rect -4258 -16139 -4205 -16086
rect -4437 -16260 -4384 -16207
rect -1915 -15586 -1862 -15533
rect -1917 -16195 -1864 -16142
rect -1649 -15475 -1596 -15422
rect -1738 -15586 -1685 -15533
rect -1560 -15586 -1507 -15533
rect -1738 -16195 -1685 -16142
rect -1561 -16194 -1508 -16141
rect -1827 -16318 -1774 -16265
rect -1381 -14196 -1328 -14143
rect -1204 -14196 -1151 -14143
rect -1293 -15475 -1240 -15422
rect -1382 -15586 -1329 -15533
rect -1204 -15586 -1151 -15533
rect -1381 -16196 -1328 -16143
rect -1204 -16195 -1151 -16142
rect -1026 -14196 -973 -14143
rect -848 -14196 -795 -14143
rect -847 -14579 -794 -14526
rect -937 -15475 -884 -15422
rect -1025 -15586 -972 -15533
rect -847 -15586 -794 -15533
rect -1026 -16195 -973 -16142
rect -669 -14196 -616 -14143
rect -669 -14579 -616 -14526
rect -491 -14196 -438 -14143
rect -491 -14579 -438 -14526
rect -581 -15475 -528 -15422
rect -670 -15586 -617 -15533
rect -491 -15586 -438 -15533
rect -4792 -16371 -4739 -16318
rect -3935 -16370 -3883 -16318
rect -1471 -16319 -1418 -16266
rect -1114 -16318 -1061 -16265
rect -759 -16317 -706 -16264
rect -314 -14580 -261 -14527
rect -137 -14579 -84 -14526
rect -225 -15475 -172 -15422
rect -313 -15586 -260 -15533
rect -136 -15586 -83 -15533
rect 43 -14579 96 -14526
rect 132 -15474 185 -15421
rect 43 -15586 96 -15533
rect 221 -15586 274 -15533
rect 220 -16195 273 -16142
rect -403 -16318 -350 -16265
rect -47 -16318 6 -16265
rect 487 -15475 540 -15422
rect 398 -15586 451 -15533
rect 575 -15586 628 -15533
rect 397 -16195 450 -16142
rect 576 -16195 629 -16142
rect 843 -15475 896 -15422
rect 755 -15586 808 -15533
rect 931 -15586 984 -15533
rect 755 -16195 808 -16142
rect 933 -16195 986 -16142
rect 1288 -14196 1341 -14143
rect 1289 -14580 1342 -14527
rect 1201 -15475 1254 -15422
rect 1110 -15586 1163 -15533
rect 1289 -15586 1342 -15533
rect 1111 -16195 1164 -16142
rect 1466 -14196 1519 -14143
rect 1467 -14579 1520 -14526
rect 1644 -14196 1697 -14143
rect 1644 -14579 1697 -14526
rect 1555 -15475 1608 -15422
rect 1466 -15586 1519 -15533
rect 1643 -15586 1696 -15533
rect 1823 -14195 1876 -14142
rect 1822 -14579 1875 -14526
rect 2000 -14196 2053 -14143
rect 1999 -14579 2052 -14526
rect 1910 -15475 1963 -15422
rect 1822 -15586 1875 -15533
rect 2000 -15586 2053 -15533
rect 2178 -14196 2231 -14143
rect 2180 -14579 2233 -14526
rect 2267 -15475 2320 -15422
rect 2179 -15586 2232 -15533
rect 2356 -15586 2409 -15533
rect 2356 -16195 2409 -16142
rect 309 -16319 362 -16266
rect 665 -16318 718 -16265
rect 845 -16318 898 -16265
rect 1021 -16318 1074 -16265
rect 1377 -16318 1430 -16265
rect 1735 -16318 1788 -16265
rect 2090 -16317 2143 -16264
rect 2624 -15475 2677 -15422
rect 2534 -15586 2587 -15533
rect 2712 -15586 2765 -15533
rect 2534 -16195 2587 -16142
rect 2713 -16194 2766 -16141
rect 2979 -15475 3032 -15422
rect 2891 -15586 2944 -15533
rect 3068 -15586 3121 -15533
rect 2891 -16195 2944 -16142
rect 3070 -16195 3123 -16142
rect 3246 -14197 3299 -14144
rect 3424 -14196 3477 -14143
rect 3425 -14579 3478 -14526
rect 3335 -15475 3388 -15422
rect 3247 -15586 3300 -15533
rect 3424 -15586 3477 -15533
rect 3249 -16195 3302 -16142
rect 2445 -16318 2498 -16265
rect 2801 -16318 2854 -16265
rect 3157 -16317 3210 -16264
rect 3602 -14196 3655 -14143
rect 3603 -14579 3656 -14526
rect 3781 -14196 3834 -14143
rect 3780 -14579 3833 -14526
rect 5184 -6767 5237 -6714
rect 5185 -8287 5237 -8235
rect 11054 -8369 11107 -8316
rect 11345 -8369 11398 -8316
rect 11638 -8369 11691 -8316
rect 11932 -8369 11985 -8316
rect 12222 -8369 12275 -8316
rect 6769 -8967 6822 -8914
rect 6679 -9198 6732 -9145
rect 6680 -9966 6733 -9913
rect 6947 -8968 7000 -8915
rect 7126 -8968 7179 -8915
rect 6858 -10120 6911 -10067
rect 7303 -8966 7356 -8913
rect 7214 -10119 7267 -10066
rect 7037 -11019 7090 -10966
rect 7482 -8966 7535 -8913
rect 7659 -8968 7712 -8915
rect 7571 -10119 7624 -10066
rect 7393 -11019 7446 -10966
rect 7837 -8967 7890 -8914
rect 8015 -8968 8068 -8915
rect 7927 -10119 7980 -10066
rect 7748 -11020 7801 -10967
rect 8194 -8967 8247 -8914
rect 8371 -8967 8424 -8914
rect 8283 -10120 8336 -10067
rect 8103 -11019 8156 -10966
rect 8549 -8967 8602 -8914
rect 8727 -8968 8780 -8915
rect 8638 -10119 8691 -10066
rect 8461 -11019 8514 -10966
rect 8906 -8967 8959 -8914
rect 11144 -9027 11197 -8974
rect 11436 -9028 11489 -8975
rect 11728 -9028 11781 -8975
rect 12020 -9029 12073 -8976
rect 12312 -9028 12365 -8975
rect 9171 -9967 9224 -9914
rect 8995 -10120 9048 -10067
rect 8817 -11019 8870 -10966
rect 11053 -11327 11106 -11274
rect 11347 -11328 11400 -11275
rect 11638 -11327 11691 -11274
rect 11931 -11327 11984 -11274
rect 12223 -11327 12276 -11274
rect 5037 -12949 5090 -12896
rect 5534 -12949 5587 -12896
rect 5031 -13086 5084 -13033
rect 4905 -14198 4958 -14145
rect 4239 -14579 4292 -14526
rect 3692 -15475 3745 -15422
rect 3603 -15586 3656 -15533
rect 3780 -15586 3833 -15533
rect 4238 -15192 4291 -15139
rect 5400 -13198 5453 -13145
rect 5142 -13447 5195 -13394
rect 5143 -14311 5196 -14258
rect 5031 -15193 5084 -15140
rect 4238 -16195 4291 -16142
rect 3514 -16319 3567 -16266
rect 3868 -16318 3921 -16265
rect 5534 -13325 5587 -13272
rect 8950 -13086 9003 -13033
rect 9305 -13086 9358 -13033
rect 8772 -13209 8825 -13156
rect 7526 -13325 7579 -13272
rect 7348 -13449 7401 -13396
rect 5833 -13575 5886 -13522
rect 6013 -13575 6066 -13522
rect 6190 -13576 6243 -13523
rect 6369 -13575 6422 -13522
rect 6547 -13576 6600 -13523
rect 6725 -13575 6778 -13522
rect 6902 -13575 6955 -13522
rect 5746 -14198 5799 -14145
rect 5924 -14311 5977 -14258
rect 6101 -14198 6154 -14145
rect 6279 -14311 6332 -14258
rect 6459 -14198 6512 -14145
rect 6813 -14198 6866 -14145
rect 6636 -14311 6689 -14258
rect 6991 -14311 7044 -14258
rect 5745 -15192 5798 -15139
rect 5400 -15306 5453 -15253
rect 5747 -15403 5800 -15350
rect 5923 -15305 5976 -15252
rect 5921 -15601 5974 -15548
rect 6101 -15192 6154 -15139
rect 6101 -15402 6154 -15349
rect 6279 -15305 6332 -15252
rect 6279 -15601 6332 -15548
rect 6458 -15192 6511 -15139
rect 6456 -15403 6509 -15350
rect 7437 -13575 7490 -13522
rect 6993 -14477 7046 -14424
rect 7347 -14477 7400 -14424
rect 6635 -15305 6688 -15252
rect 6713 -15404 6766 -15351
rect 6634 -15601 6687 -15548
rect 6813 -15504 6866 -15451
rect 7080 -14576 7133 -14523
rect 7260 -14577 7313 -14524
rect 7439 -14576 7492 -14523
rect 7882 -13326 7935 -13273
rect 8238 -13324 8291 -13271
rect 7704 -13448 7757 -13395
rect 7615 -13575 7668 -13522
rect 7793 -13576 7846 -13523
rect 8061 -13449 8114 -13396
rect 7970 -13575 8023 -13522
rect 8148 -13575 8201 -13522
rect 8415 -13449 8468 -13396
rect 8326 -13575 8379 -13522
rect 8861 -13575 8914 -13522
rect 9127 -13209 9180 -13156
rect 9038 -13575 9091 -13522
rect 9217 -13575 9270 -13522
rect 9483 -13209 9536 -13156
rect 9394 -13575 9447 -13522
rect 11442 -13325 11495 -13272
rect 11798 -13325 11851 -13272
rect 11264 -13449 11317 -13396
rect 9929 -13576 9982 -13523
rect 10108 -13575 10161 -13522
rect 10284 -13576 10337 -13523
rect 10462 -13576 10515 -13523
rect 10640 -13575 10693 -13522
rect 10819 -13576 10872 -13523
rect 7704 -14478 7757 -14425
rect 8236 -14198 8289 -14145
rect 8060 -14474 8113 -14421
rect 7169 -15403 7222 -15350
rect 7169 -15505 7222 -15452
rect 6994 -15604 7047 -15551
rect 7526 -15402 7579 -15349
rect 7526 -15606 7579 -15553
rect 7882 -15402 7935 -15349
rect 8060 -15504 8113 -15451
rect 8417 -14310 8470 -14257
rect 8327 -14576 8380 -14523
rect 7881 -15605 7934 -15552
rect 8237 -15605 8290 -15552
rect 6548 -16197 6601 -16144
rect 6726 -16197 6779 -16144
rect 6903 -16198 6956 -16145
rect 5399 -16320 5452 -16267
rect 5031 -16435 5084 -16382
rect 7970 -16198 8023 -16145
rect 8149 -16197 8202 -16144
rect 8595 -14198 8648 -14145
rect 8504 -14459 8557 -14406
rect 8505 -14577 8558 -14524
rect 8772 -14311 8825 -14258
rect 8683 -14577 8736 -14524
rect 8950 -14199 9003 -14146
rect 9127 -14312 9180 -14259
rect 9304 -14198 9357 -14145
rect 9661 -14198 9714 -14145
rect 9483 -14311 9536 -14258
rect 9572 -14576 9625 -14523
rect 9837 -14312 9890 -14259
rect 9753 -14459 9806 -14406
rect 9750 -14576 9803 -14523
rect 10016 -14198 10069 -14145
rect 9929 -14576 9982 -14523
rect 10373 -14199 10426 -14146
rect 10196 -14311 10249 -14258
rect 10195 -14475 10248 -14422
rect 10550 -14311 10603 -14258
rect 10552 -14468 10605 -14415
rect 10729 -14198 10782 -14145
rect 10908 -14311 10961 -14258
rect 11087 -14311 11140 -14258
rect 10908 -14466 10961 -14413
rect 11353 -13575 11406 -13522
rect 11620 -13450 11673 -13397
rect 11530 -13575 11583 -13522
rect 11709 -13575 11762 -13522
rect 12152 -13326 12205 -13273
rect 12509 -13325 12562 -13272
rect 11977 -13449 12030 -13396
rect 11886 -13576 11939 -13523
rect 12064 -13575 12117 -13522
rect 12334 -13449 12387 -13396
rect 12242 -13576 12295 -13523
rect 12420 -13575 12473 -13522
rect 11440 -14309 11493 -14256
rect 10819 -14576 10872 -14523
rect 8593 -15505 8646 -15452
rect 9663 -15505 9716 -15452
rect 8771 -16319 8824 -16266
rect 9128 -16319 9181 -16266
rect 10373 -15404 10426 -15351
rect 10194 -15505 10247 -15452
rect 10730 -15403 10783 -15350
rect 11264 -14468 11317 -14415
rect 10996 -14576 11049 -14523
rect 11175 -14576 11228 -14523
rect 11086 -15403 11139 -15350
rect 11619 -15305 11672 -15252
rect 11084 -15505 11137 -15452
rect 11440 -15494 11493 -15441
rect 9484 -16319 9537 -16266
rect 8950 -16435 9003 -16382
rect 9305 -16435 9358 -16382
rect 7347 -16543 7400 -16490
rect 7704 -16543 7757 -16490
rect 8060 -16543 8113 -16490
rect 8416 -16543 8469 -16490
rect 9929 -16197 9982 -16144
rect 9838 -16319 9891 -16266
rect 10107 -16198 10160 -16145
rect 10287 -16198 10340 -16145
rect 10195 -16318 10248 -16265
rect 10550 -16318 10603 -16265
rect 11441 -15605 11494 -15552
rect 11798 -15193 11851 -15140
rect 11797 -15605 11850 -15552
rect 11975 -15305 12028 -15252
rect 12155 -15192 12208 -15139
rect 12154 -15605 12207 -15552
rect 12332 -15305 12385 -15252
rect 12511 -15192 12564 -15139
rect 12511 -15605 12564 -15552
rect 10907 -16318 10960 -16265
rect 10017 -16434 10070 -16381
rect 10374 -16434 10427 -16381
rect 10731 -16432 10784 -16379
rect 11352 -16198 11405 -16145
rect 11530 -16199 11583 -16146
rect 11709 -16198 11762 -16145
rect 11263 -16543 11316 -16490
rect 11620 -16543 11673 -16490
rect 11975 -16542 12028 -16489
rect 12331 -16542 12384 -16489
<< metal2 >>
rect -5867 -1910 -5814 -1900
rect -5689 -1910 -5636 -1900
rect -5510 -1910 -5457 -1900
rect -5333 -1910 -5280 -1900
rect -5155 -1910 -5102 -1900
rect -4976 -1910 -4923 -1900
rect -4799 -1910 -4746 -1900
rect -4621 -1910 -4568 -1900
rect -4443 -1910 -4390 -1900
rect -4265 -1910 -4212 -1900
rect -4086 -1910 -4033 -1900
rect -3909 -1910 -3856 -1900
rect -1109 -1910 -1056 -1900
rect -5814 -1963 -5689 -1910
rect -5636 -1963 -5510 -1910
rect -5457 -1963 -5333 -1910
rect -5280 -1963 -5155 -1910
rect -5102 -1963 -4976 -1910
rect -4923 -1963 -4799 -1910
rect -4746 -1963 -4621 -1910
rect -4568 -1963 -4443 -1910
rect -4390 -1963 -4265 -1910
rect -4212 -1963 -4086 -1910
rect -4033 -1963 -3909 -1910
rect -3856 -1963 -1109 -1910
rect -5867 -1973 -5814 -1963
rect -5689 -1973 -5636 -1963
rect -5510 -1973 -5457 -1963
rect -5333 -1973 -5280 -1963
rect -5155 -1973 -5102 -1963
rect -4976 -1973 -4923 -1963
rect -4799 -1973 -4746 -1963
rect -4621 -1973 -4568 -1963
rect -4443 -1973 -4390 -1963
rect -4265 -1973 -4212 -1963
rect -4086 -1973 -4033 -1963
rect -3909 -1973 -3856 -1963
rect -1109 -1973 -1056 -1963
rect -1109 -2425 -1056 -2415
rect -752 -2425 -699 -2415
rect -1056 -2478 -752 -2425
rect -1109 -2488 -1056 -2478
rect -752 -2488 -699 -2478
rect 1919 -2426 1972 -2416
rect 2275 -2426 2328 -2416
rect 3193 -2426 3246 -2417
rect 1972 -2479 2275 -2426
rect 2328 -2427 3246 -2426
rect 2328 -2479 3193 -2427
rect 1919 -2489 1972 -2479
rect 2275 -2489 2328 -2479
rect 3193 -2490 3246 -2480
rect -6498 -2529 -6445 -2519
rect -5777 -2529 -5724 -2520
rect -6445 -2530 -5724 -2529
rect -5066 -2530 -5013 -2520
rect -4354 -2530 -4301 -2520
rect -6445 -2582 -5777 -2530
rect -6498 -2592 -6445 -2582
rect -5724 -2583 -5066 -2530
rect -5013 -2583 -4354 -2530
rect -5777 -2593 -5724 -2583
rect -5066 -2593 -5013 -2583
rect -4354 -2593 -4301 -2583
rect -2624 -2558 -2571 -2548
rect -1285 -2558 -1232 -2548
rect -930 -2558 -877 -2548
rect -2571 -2611 -1285 -2558
rect -1232 -2611 -930 -2558
rect -2624 -2621 -2571 -2611
rect -1285 -2621 -1232 -2611
rect -930 -2621 -877 -2611
rect 2097 -2554 2150 -2544
rect 2453 -2554 2506 -2544
rect 2150 -2607 2453 -2554
rect 2097 -2617 2150 -2607
rect 2453 -2617 2506 -2607
rect -5421 -2668 -5368 -2658
rect -4710 -2668 -4657 -2658
rect -3998 -2668 -3945 -2658
rect -3298 -2668 -3245 -2658
rect -5368 -2721 -4710 -2668
rect -4657 -2721 -3998 -2668
rect -3945 -2721 -3298 -2668
rect -5421 -2731 -5368 -2721
rect -4710 -2731 -4657 -2721
rect -3998 -2731 -3945 -2721
rect -3298 -2731 -3245 -2721
rect -1197 -2665 -1144 -2655
rect -1019 -2665 -966 -2655
rect -841 -2665 -788 -2655
rect -129 -2665 -76 -2655
rect 50 -2665 103 -2655
rect 227 -2665 280 -2655
rect 940 -2665 993 -2655
rect 1117 -2665 1170 -2655
rect 1295 -2665 1348 -2655
rect 2007 -2665 2060 -2655
rect 2186 -2665 2239 -2655
rect 2363 -2665 2416 -2655
rect -1144 -2718 -1019 -2665
rect -966 -2718 -841 -2665
rect -788 -2718 -129 -2665
rect -76 -2718 50 -2665
rect 103 -2718 227 -2665
rect 280 -2718 940 -2665
rect 993 -2718 1117 -2665
rect 1170 -2718 1295 -2665
rect 1348 -2718 2007 -2665
rect 2060 -2718 2186 -2665
rect 2239 -2718 2363 -2665
rect -1197 -2728 -1144 -2718
rect -1019 -2728 -966 -2718
rect -841 -2728 -788 -2718
rect -129 -2728 -76 -2718
rect 50 -2728 103 -2718
rect 227 -2728 280 -2718
rect 940 -2728 993 -2718
rect 1117 -2728 1170 -2718
rect 1295 -2728 1348 -2718
rect 2007 -2728 2060 -2718
rect 2186 -2728 2239 -2718
rect 2363 -2728 2416 -2718
rect -6044 -2780 -5991 -2770
rect -5866 -2780 -5813 -2770
rect -5991 -2833 -5866 -2780
rect -6044 -2843 -5991 -2833
rect -5866 -2843 -5813 -2833
rect -3908 -2780 -3855 -2770
rect -3731 -2780 -3678 -2770
rect -3855 -2833 -3731 -2780
rect -3908 -2843 -3855 -2833
rect -3731 -2843 -3678 -2833
rect -484 -3301 -431 -3291
rect 583 -3301 636 -3291
rect 1654 -3301 1707 -3291
rect -431 -3354 583 -3301
rect 636 -3354 1654 -3301
rect -484 -3364 -431 -3354
rect 583 -3364 636 -3354
rect 1654 -3364 1707 -3354
rect -6625 -3401 -6572 -3391
rect -6134 -3401 -6081 -3391
rect -5066 -3401 -5013 -3391
rect -6572 -3454 -6134 -3401
rect -6081 -3454 -5066 -3401
rect -6625 -3464 -6572 -3454
rect -6134 -3464 -6081 -3454
rect -5066 -3464 -5013 -3454
rect -4710 -3401 -4657 -3391
rect -3642 -3401 -3589 -3391
rect -3131 -3401 -3078 -3391
rect -4657 -3454 -3642 -3401
rect -3589 -3454 -3131 -3401
rect -4710 -3464 -4657 -3454
rect -3642 -3464 -3589 -3454
rect -3131 -3464 -3078 -3454
rect -1645 -3449 -1584 -3439
rect -5777 -3516 -5724 -3506
rect -3998 -3516 -3945 -3506
rect -3298 -3516 -3245 -3506
rect -5724 -3569 -3998 -3516
rect -3945 -3569 -3298 -3516
rect -1108 -3456 -1055 -3446
rect -750 -3456 -697 -3446
rect -396 -3456 -343 -3446
rect -39 -3456 14 -3446
rect 317 -3456 370 -3446
rect -1584 -3509 -1108 -3456
rect -1055 -3509 -750 -3456
rect -697 -3509 -396 -3456
rect -343 -3509 -39 -3456
rect 14 -3509 317 -3456
rect -1645 -3520 -1584 -3510
rect -1108 -3519 -1055 -3509
rect -750 -3519 -697 -3509
rect -396 -3519 -343 -3509
rect -39 -3519 14 -3509
rect 317 -3519 370 -3509
rect 850 -3456 903 -3446
rect 1206 -3456 1259 -3446
rect 1562 -3456 1615 -3446
rect 1919 -3456 1972 -3446
rect 2275 -3456 2328 -3446
rect 3019 -3452 3080 -3442
rect 903 -3509 1206 -3456
rect 1259 -3509 1562 -3456
rect 1615 -3509 1919 -3456
rect 1972 -3509 2275 -3456
rect 2328 -3509 3019 -3456
rect 850 -3519 903 -3509
rect 1206 -3519 1259 -3509
rect 1562 -3519 1615 -3509
rect 1919 -3519 1972 -3509
rect 2275 -3519 2328 -3509
rect 3080 -3509 3891 -3456
rect 3019 -3523 3080 -3513
rect -5777 -3579 -5724 -3569
rect -3998 -3579 -3945 -3569
rect -3298 -3579 -3245 -3569
rect -1286 -3571 -1233 -3561
rect -929 -3571 -876 -3561
rect -573 -3571 -520 -3561
rect -217 -3571 -164 -3561
rect -1702 -3624 -1286 -3571
rect -1233 -3624 -929 -3571
rect -876 -3624 -573 -3571
rect -520 -3624 -217 -3571
rect -6498 -3640 -6445 -3630
rect -5422 -3640 -5369 -3630
rect -4353 -3640 -4300 -3630
rect -1702 -3640 -1649 -3624
rect -1286 -3634 -1233 -3624
rect -929 -3634 -876 -3624
rect -573 -3634 -520 -3624
rect -217 -3634 -164 -3624
rect 1384 -3564 1437 -3554
rect 1741 -3564 1794 -3554
rect 2097 -3564 2150 -3554
rect 2451 -3564 2504 -3554
rect 1437 -3617 1741 -3564
rect 1794 -3617 2097 -3564
rect 2150 -3617 2451 -3564
rect 1384 -3627 1437 -3617
rect 1741 -3627 1794 -3617
rect 2097 -3627 2150 -3617
rect 2451 -3627 2504 -3617
rect -6445 -3693 -5422 -3640
rect -5369 -3693 -4353 -3640
rect -4300 -3693 -1649 -3640
rect -6498 -3703 -6445 -3693
rect -5422 -3703 -5369 -3693
rect -4353 -3703 -4300 -3693
rect -2546 -3928 -2485 -3693
rect -2546 -3999 -2485 -3989
rect -841 -4192 -788 -4182
rect -662 -4192 -609 -4182
rect -483 -4192 -430 -4182
rect -306 -4192 -253 -4182
rect 407 -4192 460 -4182
rect 583 -4192 636 -4182
rect 761 -4192 814 -4182
rect 1474 -4192 1527 -4182
rect 1652 -4192 1705 -4182
rect 1830 -4192 1883 -4182
rect 2008 -4192 2061 -4182
rect -788 -4245 -662 -4192
rect -609 -4245 -483 -4192
rect -430 -4245 -306 -4192
rect -253 -4245 407 -4192
rect 460 -4245 583 -4192
rect 636 -4245 761 -4192
rect 814 -4245 1474 -4192
rect 1527 -4245 1652 -4192
rect 1705 -4245 1830 -4192
rect 1883 -4245 2008 -4192
rect -841 -4255 -788 -4245
rect -662 -4255 -609 -4245
rect -483 -4255 -430 -4245
rect -306 -4255 -253 -4245
rect 407 -4255 460 -4245
rect 583 -4255 636 -4245
rect 761 -4255 814 -4245
rect 1474 -4255 1527 -4245
rect 1652 -4255 1705 -4245
rect 1830 -4255 1883 -4245
rect 2008 -4255 2061 -4245
rect -6498 -4271 -6445 -4261
rect -5778 -4271 -5725 -4261
rect -3998 -4271 -3945 -4261
rect -6445 -4324 -5778 -4271
rect -5725 -4324 -3998 -4271
rect 2538 -4266 2599 -4256
rect 317 -4304 370 -4294
rect 673 -4304 726 -4294
rect -6498 -4334 -6445 -4324
rect -5778 -4334 -5725 -4324
rect -3998 -4334 -3945 -4324
rect -2357 -4357 317 -4304
rect 370 -4357 673 -4304
rect 2538 -4337 2599 -4327
rect -6134 -4390 -6081 -4380
rect -5066 -4390 -5013 -4380
rect -4709 -4390 -4656 -4380
rect -3642 -4390 -3589 -4380
rect -2357 -4390 -2304 -4357
rect 317 -4367 370 -4357
rect 673 -4367 726 -4357
rect -6081 -4443 -5066 -4390
rect -5013 -4443 -4709 -4390
rect -4656 -4443 -3642 -4390
rect -3589 -4443 -2304 -4390
rect -2004 -4412 -1951 -4402
rect 495 -4412 548 -4402
rect 850 -4412 903 -4402
rect -6134 -4453 -6081 -4443
rect -5066 -4453 -5013 -4443
rect -4709 -4453 -4656 -4443
rect -3642 -4453 -3589 -4443
rect -1951 -4465 495 -4412
rect 548 -4465 850 -4412
rect -2004 -4475 -1951 -4465
rect 495 -4475 548 -4465
rect 850 -4475 903 -4465
rect 2746 -4446 2807 -4436
rect -5422 -4506 -5369 -4496
rect -4353 -4506 -4300 -4496
rect -3298 -4506 -3245 -4496
rect -2385 -4505 -2324 -4495
rect -5369 -4559 -4353 -4506
rect -4300 -4559 -3298 -4506
rect -3245 -4559 -2385 -4506
rect -5422 -4569 -5369 -4559
rect -4353 -4569 -4300 -4559
rect -3298 -4569 -3245 -4559
rect 2746 -4517 2807 -4507
rect -2385 -4576 -2324 -4566
rect 3194 -4805 3246 -4795
rect 4771 -4805 4823 -4795
rect 3246 -4857 4771 -4805
rect 3194 -4867 3246 -4857
rect 4771 -4867 4823 -4857
rect 3021 -5002 3082 -4992
rect 5037 -5006 5090 -4996
rect 4985 -5007 5037 -5006
rect 3082 -5059 5037 -5007
rect 3021 -5073 3082 -5063
rect 5037 -5069 5090 -5059
rect -2385 -5093 -2324 -5083
rect -6498 -5141 -6445 -5131
rect -5422 -5141 -5369 -5131
rect -6445 -5187 -5422 -5147
rect -6498 -5204 -6445 -5194
rect -4353 -5141 -4300 -5131
rect -5369 -5188 -4353 -5148
rect -5422 -5204 -5369 -5194
rect -1287 -5097 -1234 -5087
rect -929 -5097 -876 -5087
rect -572 -5097 -519 -5087
rect -218 -5097 -165 -5087
rect -2324 -5150 -1287 -5097
rect -1234 -5150 -929 -5097
rect -876 -5150 -572 -5097
rect -519 -5150 -218 -5097
rect 1385 -5093 1438 -5083
rect 1740 -5093 1793 -5083
rect 2096 -5093 2149 -5083
rect 2453 -5093 2506 -5083
rect -2385 -5164 -2324 -5154
rect -1287 -5160 -1234 -5150
rect -929 -5160 -876 -5150
rect -572 -5160 -519 -5150
rect -218 -5160 -165 -5150
rect 311 -5148 372 -5138
rect -4353 -5204 -4300 -5194
rect -1105 -5213 -1052 -5203
rect -751 -5213 -698 -5203
rect -396 -5213 -343 -5203
rect -41 -5213 12 -5203
rect 1438 -5146 1740 -5093
rect 1793 -5146 2096 -5093
rect 2149 -5146 2453 -5093
rect 1385 -5156 1438 -5146
rect 1740 -5156 1793 -5146
rect 2096 -5156 2149 -5146
rect 2453 -5156 2506 -5146
rect 311 -5213 372 -5209
rect -6134 -5232 -6081 -5222
rect -5066 -5233 -5013 -5223
rect -6081 -5279 -5066 -5239
rect -6134 -5295 -6081 -5285
rect -3130 -5233 -3077 -5223
rect -5013 -5279 -3130 -5239
rect -5066 -5296 -5013 -5286
rect -1876 -5232 -1823 -5222
rect -3077 -5279 -1876 -5239
rect -3130 -5296 -3077 -5286
rect -1052 -5266 -751 -5213
rect -698 -5266 -396 -5213
rect -343 -5266 -41 -5213
rect 12 -5266 316 -5213
rect 369 -5219 372 -5213
rect 846 -5213 903 -5203
rect 1207 -5213 1260 -5203
rect 1563 -5213 1616 -5203
rect 1917 -5213 1970 -5203
rect 2274 -5213 2327 -5203
rect 4905 -5212 4958 -5202
rect -1876 -5295 -1823 -5285
rect -1646 -5278 -1585 -5268
rect -1105 -5276 -1052 -5266
rect -751 -5276 -698 -5266
rect -396 -5276 -343 -5266
rect -41 -5276 12 -5266
rect 316 -5276 369 -5266
rect 846 -5266 850 -5213
rect 903 -5266 1207 -5213
rect 1260 -5266 1563 -5213
rect 1616 -5266 1917 -5213
rect 1970 -5266 2274 -5213
rect 2327 -5265 4905 -5213
rect 2327 -5266 4958 -5265
rect -6625 -5322 -6572 -5312
rect -4710 -5322 -4657 -5312
rect -6572 -5369 -4710 -5329
rect -6625 -5385 -6572 -5375
rect -3642 -5319 -3589 -5309
rect -4657 -5369 -3642 -5329
rect -4710 -5385 -4657 -5375
rect -2624 -5324 -2571 -5314
rect -3589 -5369 -2624 -5329
rect -3642 -5382 -3589 -5372
rect -1646 -5349 -1585 -5339
rect 846 -5278 907 -5266
rect 1207 -5276 1260 -5266
rect 1563 -5276 1616 -5266
rect 1917 -5276 1970 -5266
rect 2274 -5276 2327 -5266
rect 4905 -5275 4958 -5266
rect 846 -5349 907 -5339
rect -2624 -5387 -2571 -5377
rect -128 -5380 -75 -5370
rect 50 -5380 103 -5370
rect 228 -5380 281 -5370
rect 940 -5380 993 -5371
rect 1119 -5380 1172 -5370
rect 1296 -5380 1349 -5370
rect -5777 -5415 -5724 -5405
rect -3997 -5415 -3944 -5405
rect -5724 -5462 -3997 -5422
rect -5777 -5478 -5724 -5468
rect -3298 -5416 -3245 -5406
rect -3944 -5462 -3298 -5422
rect -3997 -5478 -3944 -5468
rect -75 -5433 50 -5380
rect 103 -5433 228 -5380
rect 281 -5381 1119 -5380
rect 281 -5433 940 -5381
rect -128 -5443 -75 -5433
rect 50 -5443 103 -5433
rect 228 -5443 281 -5433
rect 993 -5433 1119 -5381
rect 1172 -5433 1296 -5380
rect 940 -5444 993 -5434
rect 1119 -5443 1172 -5433
rect 1296 -5443 1349 -5433
rect -3298 -5479 -3245 -5469
rect -5956 -6016 -5903 -6006
rect -5601 -6016 -5548 -6006
rect -5244 -6016 -5191 -6006
rect -4888 -6016 -4835 -6006
rect -4532 -6016 -4479 -6006
rect -4175 -6016 -4122 -6006
rect -3820 -6016 -3767 -6006
rect -5903 -6069 -5601 -6016
rect -5548 -6069 -5244 -6016
rect -5191 -6069 -4888 -6016
rect -4835 -6069 -4532 -6016
rect -4479 -6069 -4175 -6016
rect -4122 -6069 -3820 -6016
rect -5956 -6079 -5903 -6069
rect -5601 -6079 -5548 -6069
rect -5244 -6079 -5191 -6069
rect -4888 -6079 -4835 -6069
rect -4532 -6079 -4479 -6069
rect -4175 -6079 -4122 -6069
rect -3820 -6079 -3767 -6069
rect -2624 -6007 -2571 -5997
rect 2096 -6007 2149 -5997
rect 2452 -6007 2505 -5997
rect -2571 -6060 2096 -6007
rect 2149 -6060 2452 -6007
rect -2624 -6070 -2571 -6060
rect 2096 -6070 2149 -6060
rect 2452 -6070 2505 -6060
rect -5778 -6131 -5725 -6121
rect -5065 -6131 -5012 -6121
rect -4354 -6131 -4301 -6121
rect -3298 -6131 -3245 -6121
rect 1918 -6124 1971 -6114
rect 2275 -6124 2328 -6114
rect -2821 -6125 1918 -6124
rect -5725 -6184 -5065 -6131
rect -5012 -6184 -4354 -6131
rect -4301 -6184 -3298 -6131
rect -5778 -6194 -5725 -6184
rect -5065 -6194 -5012 -6184
rect -4354 -6194 -4301 -6184
rect -3298 -6194 -3245 -6184
rect -2856 -6177 1918 -6125
rect 1971 -6177 2275 -6124
rect -6498 -6248 -6445 -6238
rect -5421 -6248 -5368 -6238
rect -4710 -6248 -4657 -6238
rect -3998 -6247 -3945 -6237
rect -6445 -6301 -5421 -6248
rect -5368 -6301 -4710 -6248
rect -4657 -6300 -3998 -6248
rect -4657 -6301 -3945 -6300
rect -6498 -6311 -6445 -6301
rect -5421 -6311 -5368 -6301
rect -4710 -6311 -4657 -6301
rect -3998 -6310 -3945 -6301
rect -4786 -6378 -4733 -6368
rect -2856 -6401 -2803 -6177
rect 1918 -6187 1971 -6177
rect 2275 -6187 2328 -6177
rect -3874 -6408 -2803 -6401
rect -4733 -6431 -2803 -6408
rect -4786 -6454 -2803 -6431
rect -2702 -6250 -2649 -6249
rect 227 -6250 280 -6240
rect 942 -6250 995 -6240
rect -2702 -6303 227 -6250
rect 280 -6303 942 -6250
rect -4786 -6461 -3820 -6454
rect -3874 -6753 -3821 -6461
rect -2702 -6542 -2649 -6303
rect 227 -6313 280 -6303
rect 942 -6313 995 -6303
rect -1876 -6364 -1823 -6354
rect -1282 -6364 -1229 -6354
rect -1823 -6417 -1282 -6364
rect -1229 -6365 -1177 -6364
rect -928 -6365 -876 -6355
rect 2879 -6365 2931 -6355
rect -1229 -6417 -928 -6365
rect -876 -6417 2879 -6365
rect -1876 -6427 -1823 -6417
rect -1282 -6427 -1229 -6417
rect -928 -6427 -876 -6417
rect 2879 -6427 2931 -6417
rect -1110 -6479 -1057 -6469
rect -752 -6479 -699 -6469
rect -1057 -6532 -752 -6479
rect -1110 -6542 -1057 -6532
rect -752 -6542 -699 -6532
rect -3874 -6816 -3821 -6806
rect -3731 -6595 -2649 -6542
rect -3731 -6903 -3678 -6595
rect -753 -6598 -700 -6588
rect 4772 -6597 4825 -6587
rect -700 -6650 4772 -6598
rect -700 -6651 4825 -6650
rect -753 -6661 -700 -6651
rect 4772 -6660 4825 -6651
rect -2003 -6714 -1950 -6704
rect 5184 -6714 5237 -6704
rect -1950 -6767 5184 -6714
rect -2003 -6777 -1950 -6767
rect 5184 -6777 5237 -6767
rect -3545 -6806 -3484 -6796
rect -3545 -6877 -3484 -6867
rect -3731 -6966 -3678 -6956
rect -3541 -7388 -3489 -6877
rect -3386 -6979 -3325 -6969
rect -3386 -7050 -3325 -7040
rect -3541 -7450 -3489 -7440
rect -3382 -7533 -3329 -7050
rect -1382 -7522 -1329 -7512
rect -1203 -7522 -1150 -7513
rect -1025 -7522 -972 -7512
rect -848 -7522 -795 -7512
rect -670 -7522 -617 -7512
rect -490 -7522 -437 -7512
rect 755 -7522 808 -7512
rect 932 -7522 985 -7512
rect 1112 -7522 1165 -7512
rect 1289 -7522 1342 -7513
rect 1467 -7522 1520 -7512
rect 1644 -7522 1697 -7512
rect 2890 -7522 2943 -7512
rect 3069 -7522 3122 -7512
rect 3247 -7522 3300 -7512
rect 3424 -7522 3477 -7512
rect 3603 -7522 3656 -7513
rect 3778 -7522 3831 -7512
rect -1329 -7523 -1025 -7522
rect -1329 -7575 -1203 -7523
rect -1382 -7585 -1329 -7575
rect -1150 -7575 -1025 -7523
rect -972 -7575 -848 -7522
rect -795 -7575 -670 -7522
rect -617 -7575 -490 -7522
rect -437 -7575 755 -7522
rect 808 -7575 932 -7522
rect 985 -7575 1112 -7522
rect 1165 -7523 1467 -7522
rect 1165 -7575 1289 -7523
rect -1203 -7586 -1150 -7576
rect -1025 -7585 -972 -7575
rect -848 -7585 -795 -7575
rect -670 -7585 -617 -7575
rect -490 -7585 -437 -7575
rect 755 -7585 808 -7575
rect 932 -7585 985 -7575
rect 1112 -7585 1165 -7575
rect 1342 -7575 1467 -7523
rect 1520 -7575 1644 -7522
rect 1697 -7575 2890 -7522
rect 2943 -7575 3069 -7522
rect 3122 -7575 3247 -7522
rect 3300 -7575 3424 -7522
rect 3477 -7523 3778 -7522
rect 3477 -7575 3603 -7523
rect 1289 -7586 1342 -7576
rect 1467 -7585 1520 -7575
rect 1644 -7585 1697 -7575
rect 2890 -7585 2943 -7575
rect 3069 -7585 3122 -7575
rect 3247 -7585 3300 -7575
rect 3424 -7585 3477 -7575
rect 3656 -7575 3778 -7523
rect 4208 -7523 4261 -7513
rect 3831 -7575 4208 -7523
rect 3603 -7586 3656 -7576
rect 3778 -7576 4208 -7575
rect 3778 -7585 3831 -7576
rect 4208 -7586 4261 -7576
rect -3382 -7596 -3329 -7586
rect -1916 -8134 -1863 -8124
rect -1739 -8134 -1686 -8124
rect -1558 -8134 -1505 -8124
rect -1382 -8134 -1329 -8124
rect -1203 -8134 -1150 -8124
rect -1026 -8134 -973 -8124
rect -848 -8134 -795 -8124
rect -670 -8134 -617 -8124
rect -491 -8134 -438 -8124
rect -314 -8134 -261 -8124
rect -136 -8134 -83 -8124
rect 42 -8134 95 -8124
rect 221 -8134 274 -8124
rect 398 -8134 451 -8124
rect 577 -8134 630 -8124
rect 754 -8134 807 -8124
rect 932 -8134 985 -8124
rect 1111 -8134 1164 -8124
rect 1289 -8134 1342 -8124
rect 1466 -8134 1519 -8124
rect 1644 -8134 1697 -8124
rect 1822 -8134 1875 -8124
rect 2000 -8134 2053 -8124
rect 2178 -8134 2231 -8124
rect 2357 -8134 2410 -8124
rect 2534 -8134 2587 -8124
rect 2712 -8134 2765 -8124
rect 2890 -8134 2943 -8124
rect 3068 -8134 3121 -8124
rect 3246 -8134 3299 -8124
rect 3424 -8134 3477 -8124
rect 3602 -8134 3655 -8124
rect 3781 -8134 3834 -8124
rect -1863 -8187 -1739 -8134
rect -1686 -8187 -1558 -8134
rect -1505 -8187 -1382 -8134
rect -1329 -8187 -1203 -8134
rect -1150 -8187 -1026 -8134
rect -973 -8187 -848 -8134
rect -795 -8187 -670 -8134
rect -617 -8187 -491 -8134
rect -438 -8187 -314 -8134
rect -261 -8187 -136 -8134
rect -83 -8187 42 -8134
rect 95 -8187 221 -8134
rect 274 -8187 398 -8134
rect 451 -8187 577 -8134
rect 630 -8187 754 -8134
rect 807 -8187 932 -8134
rect 985 -8187 1111 -8134
rect 1164 -8187 1289 -8134
rect 1342 -8187 1466 -8134
rect 1519 -8187 1644 -8134
rect 1697 -8187 1822 -8134
rect 1875 -8187 2000 -8134
rect 2053 -8187 2178 -8134
rect 2231 -8187 2357 -8134
rect 2410 -8187 2534 -8134
rect 2587 -8187 2712 -8134
rect 2765 -8187 2890 -8134
rect 2943 -8187 3068 -8134
rect 3121 -8187 3246 -8134
rect 3299 -8187 3424 -8134
rect 3477 -8187 3602 -8134
rect 3655 -8187 3781 -8134
rect -1916 -8197 -1863 -8187
rect -1739 -8197 -1686 -8187
rect -1558 -8197 -1505 -8187
rect -1382 -8197 -1329 -8187
rect -1203 -8197 -1150 -8187
rect -1026 -8197 -973 -8187
rect -848 -8197 -795 -8187
rect -670 -8197 -617 -8187
rect -491 -8197 -438 -8187
rect -314 -8197 -261 -8187
rect -136 -8197 -83 -8187
rect 42 -8197 95 -8187
rect 221 -8197 274 -8187
rect 398 -8197 451 -8187
rect 577 -8197 630 -8187
rect 754 -8197 807 -8187
rect 932 -8197 985 -8187
rect 1111 -8197 1164 -8187
rect 1289 -8197 1342 -8187
rect 1466 -8197 1519 -8187
rect 1644 -8197 1697 -8187
rect 1822 -8197 1875 -8187
rect 2000 -8197 2053 -8187
rect 2178 -8197 2231 -8187
rect 2357 -8197 2410 -8187
rect 2534 -8197 2587 -8187
rect 2712 -8197 2765 -8187
rect 2890 -8197 2943 -8187
rect 3068 -8197 3121 -8187
rect 3246 -8197 3299 -8187
rect 3424 -8197 3477 -8187
rect 3602 -8197 3655 -8187
rect 3781 -8197 3834 -8187
rect 5185 -8233 5237 -8225
rect 5185 -8235 10564 -8233
rect -1826 -8253 -1773 -8243
rect -1470 -8253 -1417 -8243
rect -1115 -8253 -1062 -8243
rect -758 -8253 -705 -8243
rect -402 -8253 -349 -8243
rect -47 -8253 6 -8243
rect 310 -8253 363 -8243
rect 666 -8253 719 -8243
rect 1022 -8253 1075 -8243
rect 1377 -8253 1430 -8243
rect 1733 -8253 1786 -8243
rect 2090 -8253 2143 -8243
rect 2446 -8253 2499 -8243
rect 2802 -8253 2855 -8243
rect 3158 -8253 3211 -8243
rect 3513 -8253 3566 -8243
rect 3869 -8253 3922 -8243
rect -1773 -8306 -1470 -8253
rect -1417 -8306 -1115 -8253
rect -1062 -8306 -758 -8253
rect -705 -8306 -402 -8253
rect -349 -8306 -47 -8253
rect 6 -8306 310 -8253
rect 363 -8306 666 -8253
rect 719 -8306 1022 -8253
rect 1075 -8306 1377 -8253
rect 1430 -8306 1733 -8253
rect 1786 -8306 2090 -8253
rect 2143 -8306 2446 -8253
rect 2499 -8306 2802 -8253
rect 2855 -8306 3158 -8253
rect 3211 -8306 3513 -8253
rect 3566 -8306 3869 -8253
rect 5237 -8285 10564 -8235
rect 5185 -8297 5237 -8287
rect -1826 -8316 -1773 -8306
rect -1470 -8316 -1417 -8306
rect -1115 -8316 -1062 -8306
rect -758 -8316 -705 -8306
rect -402 -8316 -349 -8306
rect -47 -8316 6 -8306
rect 310 -8316 363 -8306
rect 666 -8316 719 -8306
rect 1022 -8316 1075 -8306
rect 1377 -8316 1430 -8306
rect 1733 -8316 1786 -8306
rect 2090 -8316 2143 -8306
rect 2446 -8316 2499 -8306
rect 2802 -8316 2855 -8306
rect 3158 -8316 3211 -8306
rect 3513 -8316 3566 -8306
rect 3869 -8316 3922 -8306
rect 10512 -8316 10564 -8285
rect 11054 -8316 11107 -8306
rect 11345 -8316 11398 -8306
rect 11638 -8316 11691 -8306
rect 11932 -8316 11985 -8306
rect 12222 -8316 12275 -8306
rect -2447 -8367 -2394 -8357
rect -2005 -8367 -1952 -8357
rect -1648 -8367 -1595 -8357
rect -1293 -8367 -1240 -8357
rect -936 -8367 -883 -8357
rect -580 -8366 -527 -8356
rect -2394 -8420 -2005 -8367
rect -1952 -8420 -1648 -8367
rect -1595 -8420 -1293 -8367
rect -1240 -8420 -936 -8367
rect -883 -8419 -580 -8367
rect -225 -8367 -172 -8357
rect 132 -8367 185 -8358
rect 489 -8366 542 -8356
rect -527 -8419 -225 -8367
rect -883 -8420 -225 -8419
rect -172 -8368 489 -8367
rect -172 -8420 132 -8368
rect -2447 -8430 -2394 -8420
rect -2005 -8430 -1952 -8420
rect -1648 -8430 -1595 -8420
rect -1293 -8430 -1240 -8420
rect -936 -8430 -883 -8420
rect -580 -8429 -527 -8420
rect -225 -8430 -172 -8420
rect 185 -8419 489 -8368
rect 843 -8366 896 -8356
rect 542 -8419 843 -8367
rect 1201 -8367 1254 -8357
rect 1556 -8367 1609 -8357
rect 1911 -8367 1964 -8357
rect 2267 -8367 2320 -8357
rect 2624 -8367 2677 -8357
rect 2980 -8367 3033 -8357
rect 3336 -8367 3389 -8357
rect 3692 -8367 3745 -8357
rect 896 -8419 1201 -8367
rect 185 -8420 1201 -8419
rect 1254 -8420 1556 -8367
rect 1609 -8420 1911 -8367
rect 1964 -8420 2267 -8367
rect 2320 -8420 2624 -8367
rect 2677 -8420 2980 -8367
rect 3033 -8420 3336 -8367
rect 3389 -8420 3692 -8367
rect 10512 -8368 11054 -8316
rect 10584 -8369 11054 -8368
rect 11107 -8369 11345 -8316
rect 11398 -8369 11638 -8316
rect 11691 -8369 11932 -8316
rect 11985 -8369 12222 -8316
rect 11054 -8379 11107 -8369
rect 11345 -8379 11398 -8369
rect 11638 -8379 11691 -8369
rect 11932 -8379 11985 -8369
rect 12222 -8379 12275 -8369
rect 132 -8431 185 -8421
rect 489 -8429 542 -8420
rect 843 -8429 896 -8420
rect 1201 -8430 1254 -8420
rect 1556 -8430 1609 -8420
rect 1911 -8430 1964 -8420
rect 2267 -8430 2320 -8420
rect 2624 -8430 2677 -8420
rect 2980 -8430 3033 -8420
rect 3336 -8430 3389 -8420
rect 3692 -8430 3745 -8420
rect 4771 -8914 4824 -8904
rect 6769 -8914 6822 -8904
rect 6947 -8914 7000 -8905
rect 7126 -8914 7179 -8905
rect 7303 -8913 7356 -8903
rect 4824 -8967 6769 -8914
rect 6822 -8915 7303 -8914
rect 6822 -8967 6947 -8915
rect 4771 -8977 4824 -8967
rect 6769 -8977 6822 -8967
rect 7000 -8967 7126 -8915
rect 6947 -8978 7000 -8968
rect 7179 -8966 7303 -8915
rect 7482 -8913 7535 -8903
rect 7356 -8966 7482 -8914
rect 7659 -8914 7712 -8905
rect 7837 -8914 7890 -8904
rect 8015 -8914 8068 -8905
rect 8194 -8914 8247 -8904
rect 8371 -8914 8424 -8904
rect 8549 -8914 8602 -8904
rect 8727 -8914 8780 -8905
rect 8906 -8914 8959 -8904
rect 7535 -8915 7837 -8914
rect 7535 -8966 7659 -8915
rect 7179 -8967 7659 -8966
rect 7126 -8978 7179 -8968
rect 7303 -8976 7356 -8967
rect 7482 -8976 7535 -8967
rect 7712 -8967 7837 -8915
rect 7890 -8915 8194 -8914
rect 7890 -8967 8015 -8915
rect 7659 -8978 7712 -8968
rect 7837 -8977 7890 -8967
rect 8068 -8967 8194 -8915
rect 8247 -8967 8371 -8914
rect 8424 -8967 8549 -8914
rect 8602 -8915 8906 -8914
rect 8602 -8967 8727 -8915
rect 8015 -8978 8068 -8968
rect 8194 -8977 8247 -8967
rect 8371 -8977 8424 -8967
rect 8549 -8977 8602 -8967
rect 8780 -8967 8906 -8915
rect 8727 -8978 8780 -8968
rect 8906 -8977 8959 -8967
rect 11144 -8974 11197 -8964
rect 11436 -8975 11489 -8965
rect 11728 -8975 11781 -8965
rect 12020 -8975 12073 -8966
rect 12312 -8975 12365 -8965
rect 11197 -9027 11436 -8975
rect 11144 -9028 11436 -9027
rect 11489 -9028 11728 -8975
rect 11781 -8976 12312 -8975
rect 11781 -9028 12020 -8976
rect 11144 -9037 11197 -9028
rect 11436 -9038 11489 -9028
rect 11728 -9038 11781 -9028
rect 12073 -9028 12312 -8976
rect 12020 -9039 12073 -9029
rect 12312 -9038 12365 -9028
rect -1916 -9146 -1863 -9136
rect -1738 -9146 -1685 -9136
rect -1558 -9146 -1505 -9136
rect -312 -9146 -259 -9136
rect -136 -9145 -83 -9135
rect -1863 -9199 -1738 -9146
rect -1685 -9199 -1558 -9146
rect -1505 -9199 -312 -9146
rect -259 -9198 -136 -9146
rect 42 -9146 95 -9136
rect 222 -9145 275 -9135
rect -83 -9198 42 -9146
rect -259 -9199 42 -9198
rect 95 -9198 222 -9146
rect 399 -9146 452 -9136
rect 577 -9146 630 -9136
rect 2178 -9146 2231 -9137
rect 2357 -9146 2410 -9136
rect 2534 -9146 2587 -9136
rect 2713 -9146 2766 -9136
rect 4208 -9146 4261 -9136
rect 6679 -9145 6732 -9135
rect 275 -9198 399 -9146
rect 95 -9199 399 -9198
rect 452 -9199 577 -9146
rect 630 -9147 2357 -9146
rect 630 -9199 2178 -9147
rect -1916 -9209 -1863 -9199
rect -1738 -9209 -1685 -9199
rect -1558 -9209 -1505 -9199
rect -312 -9209 -259 -9199
rect -136 -9208 -83 -9199
rect 42 -9209 95 -9199
rect 222 -9208 275 -9199
rect 399 -9209 452 -9199
rect 577 -9209 630 -9199
rect 2231 -9199 2357 -9147
rect 2410 -9199 2534 -9146
rect 2587 -9199 2713 -9146
rect 2766 -9199 4208 -9146
rect 4261 -9198 6679 -9146
rect 4261 -9199 6732 -9198
rect 2178 -9210 2231 -9200
rect 2357 -9209 2410 -9199
rect 2534 -9209 2587 -9199
rect 2713 -9209 2766 -9199
rect 4208 -9209 4261 -9199
rect 6679 -9208 6732 -9199
rect -2315 -9525 -2262 -9515
rect -1916 -9525 -1863 -9515
rect -1738 -9525 -1685 -9516
rect -1560 -9525 -1507 -9515
rect -1382 -9524 -1329 -9514
rect -2262 -9578 -1916 -9525
rect -1863 -9526 -1560 -9525
rect -1863 -9578 -1738 -9526
rect -2315 -9588 -2262 -9578
rect -1916 -9588 -1863 -9578
rect -1685 -9578 -1560 -9526
rect -1507 -9577 -1382 -9525
rect -314 -9525 -261 -9515
rect -136 -9525 -83 -9516
rect 43 -9525 96 -9515
rect 220 -9525 273 -9515
rect 398 -9525 451 -9515
rect 576 -9525 629 -9515
rect 2356 -9525 2409 -9515
rect 2534 -9525 2587 -9515
rect 2712 -9525 2765 -9516
rect 2891 -9525 2944 -9515
rect 3069 -9525 3122 -9515
rect 3246 -9525 3299 -9515
rect -1329 -9577 -314 -9525
rect -1507 -9578 -314 -9577
rect -261 -9526 43 -9525
rect -261 -9578 -136 -9526
rect -1738 -9589 -1685 -9579
rect -1560 -9588 -1507 -9578
rect -1382 -9587 -1329 -9578
rect -314 -9588 -261 -9578
rect -83 -9578 43 -9526
rect 96 -9578 220 -9525
rect 273 -9578 398 -9525
rect 451 -9578 576 -9525
rect 629 -9578 2356 -9525
rect 2409 -9578 2534 -9525
rect 2587 -9526 2891 -9525
rect 2587 -9578 2712 -9526
rect -136 -9589 -83 -9579
rect 43 -9588 96 -9578
rect 220 -9588 273 -9578
rect 398 -9588 451 -9578
rect 576 -9588 629 -9578
rect 2356 -9588 2409 -9578
rect 2534 -9588 2587 -9578
rect 2765 -9578 2891 -9526
rect 2944 -9578 3069 -9525
rect 3122 -9578 3246 -9525
rect 3299 -9578 5074 -9525
rect 2712 -9589 2765 -9579
rect 2891 -9588 2944 -9578
rect 3069 -9588 3122 -9578
rect 3246 -9588 3299 -9578
rect 6680 -9913 6733 -9903
rect 9171 -9913 9224 -9904
rect 6733 -9914 9224 -9913
rect 6733 -9966 9171 -9914
rect 6680 -9976 6733 -9966
rect 9171 -9977 9224 -9967
rect 6858 -10066 6911 -10057
rect 7214 -10066 7267 -10056
rect 7571 -10066 7624 -10056
rect 7927 -10066 7980 -10056
rect 8283 -10066 8336 -10057
rect 8638 -10066 8691 -10056
rect 8995 -10066 9048 -10057
rect 6858 -10067 7214 -10066
rect 6911 -10119 7214 -10067
rect 7267 -10119 7571 -10066
rect 7624 -10119 7927 -10066
rect 7980 -10067 8638 -10066
rect 7980 -10119 8283 -10067
rect 6858 -10130 6911 -10120
rect 7214 -10129 7267 -10119
rect 7571 -10129 7624 -10119
rect 7927 -10129 7980 -10119
rect 8336 -10119 8638 -10067
rect 8691 -10067 9048 -10066
rect 8691 -10119 8995 -10067
rect 8283 -10130 8336 -10120
rect 8638 -10129 8691 -10119
rect 8995 -10130 9048 -10120
rect -1827 -10508 -1774 -10498
rect -1470 -10508 -1417 -10498
rect -1114 -10508 -1061 -10498
rect -758 -10508 -705 -10498
rect -402 -10508 -349 -10498
rect -46 -10508 7 -10498
rect 309 -10508 362 -10498
rect 665 -10508 718 -10498
rect 931 -10508 984 -10498
rect 1199 -10508 1252 -10498
rect 1556 -10508 1609 -10498
rect 1913 -10508 1966 -10498
rect 2268 -10508 2321 -10498
rect 2623 -10508 2676 -10498
rect 2980 -10508 3033 -10498
rect 3335 -10508 3388 -10498
rect 3692 -10508 3745 -10498
rect -1774 -10561 -1470 -10508
rect -1417 -10561 -1114 -10508
rect -1061 -10561 -758 -10508
rect -705 -10561 -402 -10508
rect -349 -10561 -46 -10508
rect 7 -10561 309 -10508
rect 362 -10561 665 -10508
rect 718 -10561 931 -10508
rect 984 -10561 1199 -10508
rect 1252 -10561 1556 -10508
rect 1609 -10561 1913 -10508
rect 1966 -10561 2268 -10508
rect 2321 -10561 2623 -10508
rect 2676 -10561 2980 -10508
rect 3033 -10561 3335 -10508
rect 3388 -10561 3692 -10508
rect -1827 -10571 -1774 -10561
rect -1470 -10571 -1417 -10561
rect -1114 -10571 -1061 -10561
rect -758 -10571 -705 -10561
rect -402 -10571 -349 -10561
rect -46 -10571 7 -10561
rect 309 -10571 362 -10561
rect 665 -10571 718 -10561
rect 931 -10571 984 -10561
rect 1199 -10571 1252 -10561
rect 1556 -10571 1609 -10561
rect 1913 -10571 1966 -10561
rect 2268 -10571 2321 -10561
rect 2623 -10571 2676 -10561
rect 2980 -10571 3033 -10561
rect 3335 -10571 3388 -10561
rect 3692 -10571 3745 -10561
rect 7037 -10966 7090 -10956
rect 7393 -10966 7446 -10956
rect 7748 -10966 7801 -10957
rect 8103 -10966 8156 -10956
rect 8461 -10966 8514 -10956
rect 8817 -10966 8870 -10956
rect 7090 -11019 7393 -10966
rect 7446 -10967 8103 -10966
rect 7446 -11019 7748 -10967
rect 7037 -11029 7090 -11019
rect 7393 -11029 7446 -11019
rect 7801 -11019 8103 -10967
rect 8156 -11019 8461 -10966
rect 8514 -11019 8817 -10966
rect 7748 -11030 7801 -11020
rect 8103 -11029 8156 -11019
rect 8461 -11029 8514 -11019
rect 8817 -11029 8870 -11019
rect -1649 -11128 -1596 -11118
rect -1293 -11128 -1240 -11118
rect -937 -11128 -884 -11118
rect 1377 -11128 1430 -11118
rect 1733 -11128 1786 -11118
rect 2089 -11128 2142 -11118
rect -1596 -11181 -1293 -11128
rect -1240 -11181 -937 -11128
rect -884 -11181 1377 -11128
rect 1430 -11181 1733 -11128
rect 1786 -11181 2089 -11128
rect -1649 -11191 -1596 -11181
rect -1293 -11191 -1240 -11181
rect -937 -11191 -884 -11181
rect 1377 -11191 1430 -11181
rect 1733 -11191 1786 -11181
rect 2089 -11191 2142 -11181
rect -2004 -11237 -1951 -11227
rect -580 -11237 -527 -11227
rect 2446 -11237 2499 -11227
rect 3871 -11237 3924 -11228
rect -1951 -11290 -580 -11237
rect -527 -11290 2446 -11237
rect 2499 -11238 3924 -11237
rect 2499 -11290 3871 -11238
rect -2004 -11300 -1951 -11290
rect -580 -11300 -527 -11290
rect 2446 -11300 2499 -11290
rect 3871 -11301 3924 -11291
rect 11053 -11274 11106 -11264
rect 11347 -11274 11400 -11265
rect 11638 -11274 11691 -11264
rect 11931 -11274 11984 -11264
rect 12223 -11274 12276 -11264
rect 11106 -11275 11638 -11274
rect 11106 -11327 11347 -11275
rect 11053 -11337 11106 -11327
rect 11400 -11327 11638 -11275
rect 11691 -11327 11931 -11274
rect 11984 -11327 12223 -11274
rect 11347 -11338 11400 -11328
rect 11638 -11337 11691 -11327
rect 11931 -11337 11984 -11327
rect 12223 -11337 12276 -11327
rect -224 -11357 -171 -11347
rect 131 -11357 184 -11347
rect 487 -11357 540 -11347
rect 2800 -11357 2853 -11347
rect 3157 -11357 3210 -11347
rect 3513 -11357 3566 -11347
rect -171 -11410 131 -11357
rect 184 -11410 487 -11357
rect 540 -11410 2800 -11357
rect 2853 -11410 3157 -11357
rect 3210 -11410 3513 -11357
rect -224 -11420 -171 -11410
rect 131 -11420 184 -11410
rect 487 -11420 540 -11410
rect 2800 -11420 2853 -11410
rect 3157 -11420 3210 -11410
rect 3513 -11420 3566 -11410
rect -5502 -11471 -5449 -11461
rect -5000 -11471 -4947 -11462
rect -4502 -11471 -4449 -11461
rect -5449 -11472 -4502 -11471
rect -5449 -11524 -5000 -11472
rect -5502 -11534 -5449 -11524
rect -4947 -11524 -4502 -11472
rect -2447 -11472 -2394 -11462
rect -4449 -11524 -2447 -11472
rect -5000 -11535 -4947 -11525
rect -4502 -11525 -2447 -11524
rect -4502 -11534 -4449 -11525
rect -2447 -11535 -2394 -11525
rect -1915 -11519 -1862 -11509
rect -1738 -11519 -1685 -11509
rect -1559 -11519 -1506 -11509
rect -1381 -11519 -1328 -11509
rect -1203 -11519 -1150 -11509
rect -1025 -11519 -972 -11509
rect -848 -11519 -795 -11509
rect -670 -11519 -617 -11509
rect -492 -11519 -439 -11509
rect -314 -11519 -261 -11509
rect -136 -11519 -83 -11509
rect 42 -11519 95 -11509
rect 220 -11519 273 -11509
rect 399 -11519 452 -11509
rect 577 -11519 630 -11509
rect 1288 -11519 1341 -11509
rect 1468 -11519 1521 -11509
rect 1644 -11519 1697 -11510
rect 1823 -11519 1876 -11509
rect 2000 -11519 2053 -11509
rect 2178 -11519 2231 -11509
rect 2357 -11519 2410 -11509
rect 2534 -11519 2587 -11509
rect 2713 -11519 2766 -11509
rect 2890 -11519 2943 -11509
rect 3068 -11519 3121 -11509
rect 3247 -11519 3300 -11509
rect 3425 -11519 3478 -11509
rect 3603 -11519 3656 -11509
rect 3781 -11519 3834 -11509
rect -1862 -11572 -1738 -11519
rect -1685 -11572 -1559 -11519
rect -1506 -11572 -1381 -11519
rect -1328 -11572 -1203 -11519
rect -1150 -11572 -1025 -11519
rect -972 -11572 -848 -11519
rect -795 -11572 -670 -11519
rect -617 -11572 -492 -11519
rect -439 -11572 -314 -11519
rect -261 -11572 -136 -11519
rect -83 -11572 42 -11519
rect 95 -11572 220 -11519
rect 273 -11572 399 -11519
rect 452 -11572 577 -11519
rect 630 -11572 1288 -11519
rect 1341 -11572 1468 -11519
rect 1521 -11520 1823 -11519
rect 1521 -11572 1644 -11520
rect -5376 -11588 -5323 -11578
rect -5127 -11588 -5074 -11578
rect -4377 -11588 -4324 -11578
rect -3928 -11588 -3875 -11579
rect -1915 -11582 -1862 -11572
rect -1738 -11582 -1685 -11572
rect -1559 -11582 -1506 -11572
rect -1381 -11582 -1328 -11572
rect -1203 -11582 -1150 -11572
rect -1025 -11582 -972 -11572
rect -848 -11582 -795 -11572
rect -670 -11582 -617 -11572
rect -492 -11582 -439 -11572
rect -314 -11582 -261 -11572
rect -136 -11582 -83 -11572
rect 42 -11582 95 -11572
rect 220 -11582 273 -11572
rect 399 -11582 452 -11572
rect 577 -11582 630 -11572
rect 1288 -11582 1341 -11572
rect 1468 -11582 1521 -11572
rect 1697 -11572 1823 -11520
rect 1876 -11572 2000 -11519
rect 2053 -11572 2178 -11519
rect 2231 -11572 2357 -11519
rect 2410 -11572 2534 -11519
rect 2587 -11572 2713 -11519
rect 2766 -11572 2890 -11519
rect 2943 -11572 3068 -11519
rect 3121 -11572 3247 -11519
rect 3300 -11572 3425 -11519
rect 3478 -11572 3603 -11519
rect 3656 -11572 3781 -11519
rect 1644 -11583 1697 -11573
rect 1823 -11582 1876 -11572
rect 2000 -11582 2053 -11572
rect 2178 -11582 2231 -11572
rect 2357 -11582 2410 -11572
rect 2534 -11582 2587 -11572
rect 2713 -11582 2766 -11572
rect 2890 -11582 2943 -11572
rect 3068 -11582 3121 -11572
rect 3247 -11582 3300 -11572
rect 3425 -11582 3478 -11572
rect 3603 -11582 3656 -11572
rect 3781 -11582 3834 -11572
rect -5323 -11641 -5127 -11588
rect -5074 -11641 -4377 -11588
rect -4324 -11589 -3875 -11588
rect -4324 -11641 -3928 -11589
rect -5376 -11651 -5323 -11641
rect -5127 -11651 -5074 -11641
rect -4377 -11651 -4324 -11641
rect -3928 -11652 -3875 -11642
rect -6077 -11712 -6024 -11702
rect -5626 -11712 -5573 -11702
rect -4877 -11712 -4824 -11702
rect -4627 -11712 -4574 -11702
rect -6024 -11765 -5626 -11712
rect -5573 -11765 -4877 -11712
rect -4824 -11765 -4627 -11712
rect -6077 -11775 -6024 -11765
rect -5626 -11775 -5573 -11765
rect -4877 -11775 -4824 -11765
rect -4627 -11775 -4574 -11765
rect -2005 -12142 -1952 -12132
rect -1649 -12142 -1596 -12132
rect 3514 -12142 3567 -12132
rect 3871 -12142 3924 -12132
rect -1952 -12195 -1649 -12142
rect -1596 -12144 -1284 -12142
rect -1250 -12144 3514 -12142
rect -1596 -12195 3514 -12144
rect 3567 -12195 3871 -12142
rect -2005 -12205 -1952 -12195
rect -1649 -12205 -1596 -12195
rect 3514 -12205 3567 -12195
rect 3871 -12205 3924 -12195
rect -6223 -12262 -6170 -12252
rect -5751 -12262 -5698 -12252
rect -4752 -12262 -4699 -12252
rect -6170 -12315 -5751 -12262
rect -5698 -12315 -4752 -12262
rect -6223 -12325 -6170 -12315
rect -5751 -12325 -5698 -12315
rect -4752 -12325 -4699 -12315
rect -1294 -12253 -1241 -12244
rect -582 -12253 -529 -12243
rect 130 -12253 183 -12243
rect 1735 -12253 1788 -12244
rect 2445 -12253 2498 -12243
rect 3158 -12252 3211 -12242
rect -1294 -12254 -582 -12253
rect -1241 -12306 -582 -12254
rect -529 -12306 130 -12253
rect 183 -12254 2445 -12253
rect 183 -12306 1735 -12254
rect -1294 -12317 -1241 -12307
rect -582 -12316 -529 -12306
rect 130 -12316 183 -12306
rect 1788 -12306 2445 -12254
rect 2498 -12305 3158 -12253
rect 2498 -12306 3211 -12305
rect 1735 -12317 1788 -12307
rect 2445 -12316 2498 -12306
rect 3158 -12315 3211 -12306
rect -5251 -12389 -5198 -12379
rect -4251 -12389 -4198 -12379
rect -3788 -12389 -3735 -12379
rect -3542 -12389 -3489 -12379
rect -5198 -12442 -4251 -12389
rect -4198 -12442 -3788 -12389
rect -3735 -12442 -3542 -12389
rect -5251 -12452 -5198 -12442
rect -4251 -12452 -4198 -12442
rect -3788 -12452 -3735 -12442
rect -3542 -12452 -3489 -12442
rect -937 -12383 -884 -12373
rect -224 -12383 -171 -12373
rect 486 -12383 539 -12374
rect 1378 -12383 1431 -12373
rect 2088 -12382 2141 -12372
rect -884 -12436 -224 -12383
rect -171 -12384 1378 -12383
rect -171 -12436 486 -12384
rect -937 -12446 -884 -12436
rect -224 -12446 -171 -12436
rect 539 -12436 1378 -12384
rect 1431 -12435 2088 -12383
rect 2801 -12382 2854 -12372
rect 2141 -12435 2801 -12383
rect 1431 -12436 2854 -12435
rect 486 -12447 539 -12437
rect 1378 -12446 1431 -12436
rect 2088 -12445 2141 -12436
rect 2801 -12445 2854 -12436
rect 5037 -12896 5090 -12886
rect 5534 -12896 5587 -12886
rect -6077 -12945 -6024 -12935
rect -5376 -12945 -5323 -12935
rect -5126 -12945 -5073 -12935
rect -4376 -12945 -4323 -12935
rect -6024 -12998 -5376 -12945
rect -5323 -12998 -5126 -12945
rect -5073 -12998 -4376 -12945
rect 5090 -12949 5534 -12896
rect 5037 -12959 5090 -12949
rect 5534 -12959 5587 -12949
rect -6077 -13008 -6024 -12998
rect -5376 -13008 -5323 -12998
rect -5126 -13008 -5073 -12998
rect -4376 -13008 -4323 -12998
rect 5031 -13033 5084 -13023
rect 8950 -13033 9003 -13023
rect 9305 -13033 9358 -13023
rect -6426 -13052 -6373 -13042
rect -5626 -13052 -5573 -13042
rect -4877 -13052 -4824 -13042
rect -4627 -13052 -4574 -13042
rect -3928 -13052 -3875 -13042
rect -6373 -13105 -5626 -13052
rect -5573 -13105 -4877 -13052
rect -4824 -13105 -4627 -13052
rect -4574 -13105 -3928 -13052
rect 5084 -13086 8950 -13033
rect 9003 -13086 9305 -13033
rect 5031 -13096 5084 -13086
rect 8950 -13096 9003 -13086
rect 9305 -13096 9358 -13086
rect -6426 -13115 -6373 -13105
rect -5626 -13115 -5573 -13105
rect -4877 -13115 -4824 -13105
rect -4627 -13115 -4574 -13105
rect -3928 -13115 -3875 -13105
rect -2004 -13145 -1951 -13135
rect -581 -13145 -528 -13135
rect 2446 -13145 2499 -13135
rect 3870 -13145 3923 -13135
rect 5400 -13145 5453 -13135
rect -5730 -13157 -5677 -13147
rect -4752 -13157 -4699 -13147
rect -3788 -13157 -3735 -13147
rect -5677 -13210 -4752 -13157
rect -4699 -13210 -3788 -13157
rect -1951 -13198 -581 -13145
rect -528 -13198 2446 -13145
rect 2499 -13198 3870 -13145
rect 3923 -13198 5400 -13145
rect 5453 -13156 8828 -13145
rect 9127 -13156 9180 -13146
rect 9483 -13156 9536 -13146
rect 5453 -13198 8772 -13156
rect -2004 -13208 -1951 -13198
rect -581 -13208 -528 -13198
rect 2446 -13208 2499 -13198
rect 3870 -13208 3923 -13198
rect 5400 -13208 5453 -13198
rect -5730 -13220 -5677 -13210
rect -4752 -13220 -4699 -13210
rect -3788 -13220 -3735 -13210
rect 8825 -13209 9127 -13156
rect 9180 -13209 9483 -13156
rect 8772 -13219 8825 -13209
rect 9127 -13219 9180 -13209
rect 9483 -13219 9536 -13209
rect -6223 -13255 -6170 -13245
rect -5250 -13255 -5197 -13245
rect -4250 -13255 -4197 -13245
rect -3382 -13255 -3329 -13245
rect -6170 -13308 -5250 -13255
rect -5197 -13308 -4250 -13255
rect -4197 -13308 -3382 -13255
rect -6223 -13318 -6170 -13308
rect -5250 -13318 -5197 -13308
rect -4250 -13318 -4197 -13308
rect -3382 -13318 -3329 -13308
rect -1648 -13272 -1595 -13262
rect -1291 -13272 -1238 -13262
rect -937 -13272 -884 -13262
rect 1379 -13272 1432 -13262
rect 1732 -13272 1785 -13262
rect 2091 -13272 2144 -13262
rect 5534 -13272 5587 -13262
rect 7526 -13272 7579 -13262
rect 7882 -13272 7935 -13263
rect 8238 -13271 8291 -13261
rect -1595 -13325 -1291 -13272
rect -1238 -13325 -937 -13272
rect -884 -13325 1379 -13272
rect 1432 -13325 1732 -13272
rect 1785 -13325 2091 -13272
rect 2144 -13325 5323 -13272
rect -1648 -13335 -1595 -13325
rect -1291 -13335 -1238 -13325
rect -937 -13335 -884 -13325
rect 1379 -13335 1432 -13325
rect 1732 -13335 1785 -13325
rect 2091 -13335 2144 -13325
rect -225 -13394 -172 -13384
rect 133 -13394 186 -13384
rect 487 -13394 540 -13385
rect 2802 -13394 2855 -13384
rect 3157 -13394 3210 -13385
rect 3512 -13394 3565 -13384
rect 5142 -13394 5195 -13384
rect -172 -13447 133 -13394
rect 186 -13395 2802 -13394
rect 186 -13447 487 -13395
rect -225 -13457 -172 -13447
rect 133 -13457 186 -13447
rect 540 -13447 2802 -13395
rect 2855 -13395 3512 -13394
rect 2855 -13447 3157 -13395
rect 487 -13458 540 -13448
rect 2802 -13457 2855 -13447
rect 3210 -13447 3512 -13395
rect 3565 -13447 5142 -13394
rect 3157 -13458 3210 -13448
rect 3512 -13457 3565 -13447
rect 5142 -13457 5195 -13447
rect 5270 -13396 5323 -13325
rect 5587 -13325 7526 -13272
rect 7579 -13273 8238 -13272
rect 7579 -13325 7882 -13273
rect 5534 -13335 5587 -13325
rect 7526 -13335 7579 -13325
rect 7935 -13324 8238 -13273
rect 11442 -13272 11495 -13262
rect 11798 -13272 11851 -13262
rect 12152 -13272 12205 -13263
rect 12509 -13272 12562 -13262
rect 8291 -13324 11442 -13272
rect 7935 -13325 11442 -13324
rect 11495 -13325 11798 -13272
rect 11851 -13273 12509 -13272
rect 11851 -13325 12152 -13273
rect 7882 -13336 7935 -13326
rect 8238 -13334 8291 -13325
rect 11442 -13335 11495 -13325
rect 11798 -13335 11851 -13325
rect 12205 -13325 12509 -13273
rect 12152 -13336 12205 -13326
rect 12509 -13335 12562 -13325
rect 7348 -13396 7401 -13386
rect 7704 -13395 7757 -13385
rect 5270 -13449 7348 -13396
rect 7401 -13448 7704 -13396
rect 8061 -13396 8114 -13386
rect 8415 -13396 8468 -13386
rect 11264 -13396 11317 -13386
rect 11620 -13396 11673 -13387
rect 11977 -13396 12030 -13386
rect 12334 -13396 12387 -13386
rect 7757 -13448 8061 -13396
rect 7401 -13449 8061 -13448
rect 8114 -13449 8415 -13396
rect 8468 -13449 11264 -13396
rect 11317 -13397 11977 -13396
rect 11317 -13449 11620 -13397
rect 7348 -13459 7401 -13449
rect 7704 -13458 7757 -13449
rect 8061 -13459 8114 -13449
rect 8415 -13459 8468 -13449
rect 11264 -13459 11317 -13449
rect 11673 -13449 11977 -13397
rect 12030 -13449 12334 -13396
rect 11620 -13460 11673 -13450
rect 11977 -13459 12030 -13449
rect 12334 -13459 12387 -13449
rect 5833 -13522 5886 -13512
rect 6013 -13522 6066 -13512
rect 6190 -13522 6243 -13513
rect 6369 -13522 6422 -13512
rect 6547 -13522 6600 -13513
rect 6725 -13522 6778 -13512
rect 6902 -13522 6955 -13512
rect 7437 -13522 7490 -13512
rect 7615 -13522 7668 -13512
rect 7793 -13522 7846 -13513
rect 7970 -13522 8023 -13512
rect 8148 -13522 8201 -13512
rect 8326 -13522 8379 -13512
rect 8861 -13522 8914 -13512
rect 9038 -13522 9091 -13512
rect 9217 -13522 9270 -13512
rect 9394 -13522 9447 -13512
rect 9929 -13522 9982 -13513
rect 10108 -13522 10161 -13512
rect 10284 -13522 10337 -13513
rect 10462 -13522 10515 -13513
rect 10640 -13522 10693 -13512
rect 10819 -13522 10872 -13513
rect 11353 -13522 11406 -13512
rect 11530 -13522 11583 -13512
rect 11709 -13522 11762 -13512
rect 11886 -13522 11939 -13513
rect 12064 -13522 12117 -13512
rect 12242 -13522 12295 -13513
rect 12420 -13522 12473 -13512
rect 5886 -13575 6013 -13522
rect 6066 -13523 6369 -13522
rect 6066 -13575 6190 -13523
rect 5833 -13585 5886 -13575
rect 6013 -13585 6066 -13575
rect 6243 -13575 6369 -13523
rect 6422 -13523 6725 -13522
rect 6422 -13575 6547 -13523
rect 6190 -13586 6243 -13576
rect 6369 -13585 6422 -13575
rect 6600 -13575 6725 -13523
rect 6778 -13575 6902 -13522
rect 6955 -13575 7437 -13522
rect 7490 -13575 7615 -13522
rect 7668 -13523 7970 -13522
rect 7668 -13575 7793 -13523
rect 6547 -13586 6600 -13576
rect 6725 -13585 6778 -13575
rect 6902 -13585 6955 -13575
rect 7437 -13585 7490 -13575
rect 7615 -13585 7668 -13575
rect 7846 -13575 7970 -13523
rect 8023 -13575 8148 -13522
rect 8201 -13575 8326 -13522
rect 8379 -13575 8861 -13522
rect 8914 -13575 9038 -13522
rect 9091 -13575 9217 -13522
rect 9270 -13575 9394 -13522
rect 9447 -13523 10108 -13522
rect 9447 -13575 9929 -13523
rect 7793 -13586 7846 -13576
rect 7970 -13585 8023 -13575
rect 8148 -13585 8201 -13575
rect 8326 -13585 8379 -13575
rect 8861 -13585 8914 -13575
rect 9038 -13585 9091 -13575
rect 9217 -13585 9270 -13575
rect 9394 -13585 9447 -13575
rect 9982 -13575 10108 -13523
rect 10161 -13523 10640 -13522
rect 10161 -13575 10284 -13523
rect 9929 -13586 9982 -13576
rect 10108 -13585 10161 -13575
rect 10337 -13575 10462 -13523
rect 10284 -13586 10337 -13576
rect 10515 -13575 10640 -13523
rect 10693 -13523 11353 -13522
rect 10693 -13575 10819 -13523
rect 10462 -13586 10515 -13576
rect 10640 -13585 10693 -13575
rect 10872 -13575 11353 -13523
rect 11406 -13575 11530 -13522
rect 11583 -13575 11709 -13522
rect 11762 -13523 12064 -13522
rect 11762 -13575 11886 -13523
rect 10819 -13586 10872 -13576
rect 11353 -13585 11406 -13575
rect 11530 -13585 11583 -13575
rect 11709 -13585 11762 -13575
rect 11939 -13575 12064 -13523
rect 12117 -13523 12420 -13522
rect 12117 -13575 12242 -13523
rect 11886 -13586 11939 -13576
rect 12064 -13585 12117 -13575
rect 12295 -13575 12420 -13523
rect 12242 -13586 12295 -13576
rect 12420 -13585 12473 -13575
rect -6159 -13995 -6106 -13985
rect -5860 -13995 -5807 -13985
rect -5147 -13995 -5094 -13985
rect -4436 -13995 -4383 -13985
rect -6106 -14048 -5860 -13995
rect -5807 -14048 -5147 -13995
rect -5094 -14048 -4436 -13995
rect -6159 -14058 -6106 -14048
rect -5860 -14058 -5807 -14048
rect -5147 -14058 -5094 -14048
rect -4436 -14058 -4383 -14048
rect -5504 -14101 -5451 -14091
rect -4791 -14101 -4738 -14091
rect -3936 -14101 -3883 -14091
rect -5451 -14154 -4791 -14101
rect -4738 -14154 -3936 -14101
rect -5504 -14164 -5451 -14154
rect -4791 -14164 -4738 -14154
rect -3936 -14164 -3883 -14154
rect -2315 -14143 -2262 -14133
rect -1381 -14143 -1328 -14133
rect -1204 -14143 -1151 -14133
rect -1026 -14143 -973 -14133
rect -848 -14143 -795 -14133
rect -669 -14143 -616 -14133
rect -491 -14143 -438 -14133
rect 1288 -14143 1341 -14133
rect 1466 -14143 1519 -14133
rect 1644 -14143 1697 -14133
rect 1823 -14142 1876 -14132
rect -2262 -14196 -1381 -14143
rect -1328 -14196 -1204 -14143
rect -1151 -14196 -1026 -14143
rect -973 -14196 -848 -14143
rect -795 -14196 -669 -14143
rect -616 -14196 -491 -14143
rect -438 -14196 1288 -14143
rect 1341 -14196 1466 -14143
rect 1519 -14196 1644 -14143
rect 1697 -14195 1823 -14143
rect 2000 -14143 2053 -14133
rect 2178 -14143 2231 -14133
rect 3246 -14143 3299 -14134
rect 3424 -14143 3477 -14133
rect 3602 -14143 3655 -14133
rect 3781 -14143 3834 -14133
rect 1876 -14195 2000 -14143
rect 1697 -14196 2000 -14195
rect 2053 -14196 2178 -14143
rect 2231 -14144 3424 -14143
rect 2231 -14196 3246 -14144
rect -2315 -14206 -2262 -14196
rect -1381 -14206 -1328 -14196
rect -1204 -14206 -1151 -14196
rect -1026 -14206 -973 -14196
rect -848 -14206 -795 -14196
rect -669 -14206 -616 -14196
rect -491 -14206 -438 -14196
rect 1288 -14206 1341 -14196
rect 1466 -14206 1519 -14196
rect 1644 -14206 1697 -14196
rect 1823 -14205 1876 -14196
rect 2000 -14206 2053 -14196
rect 2178 -14206 2231 -14196
rect 3299 -14196 3424 -14144
rect 3477 -14196 3602 -14143
rect 3655 -14196 3781 -14143
rect 3246 -14207 3299 -14197
rect 3424 -14206 3477 -14196
rect 3602 -14206 3655 -14196
rect 3781 -14206 3834 -14196
rect 4905 -14145 4958 -14135
rect 5746 -14145 5799 -14135
rect 6101 -14145 6154 -14135
rect 6459 -14145 6512 -14135
rect 6813 -14145 6866 -14135
rect 8236 -14145 8289 -14135
rect 8595 -14145 8648 -14135
rect 8950 -14145 9003 -14136
rect 9304 -14145 9357 -14135
rect 9661 -14145 9714 -14135
rect 10016 -14145 10069 -14135
rect 10373 -14145 10426 -14136
rect 10729 -14145 10782 -14135
rect 4958 -14198 5746 -14145
rect 5799 -14198 6101 -14145
rect 6154 -14198 6459 -14145
rect 6512 -14198 6813 -14145
rect 6866 -14198 8236 -14145
rect 8289 -14198 8595 -14145
rect 8648 -14146 9304 -14145
rect 8648 -14198 8950 -14146
rect 4905 -14208 4958 -14198
rect 5746 -14208 5799 -14198
rect 6101 -14208 6154 -14198
rect 6459 -14208 6512 -14198
rect 6813 -14208 6866 -14198
rect 8236 -14208 8289 -14198
rect 8595 -14208 8648 -14198
rect 9003 -14198 9304 -14146
rect 9357 -14198 9661 -14145
rect 9714 -14198 10016 -14145
rect 10069 -14146 10729 -14145
rect 10069 -14198 10373 -14146
rect 8950 -14209 9003 -14199
rect 9304 -14208 9357 -14198
rect 9661 -14208 9714 -14198
rect 10016 -14208 10069 -14198
rect 10426 -14198 10729 -14146
rect 10373 -14209 10426 -14199
rect 10729 -14208 10782 -14198
rect 5143 -14258 5196 -14248
rect 5924 -14258 5977 -14248
rect 6279 -14258 6332 -14248
rect 6636 -14258 6689 -14248
rect 6991 -14258 7044 -14248
rect 8417 -14257 8470 -14247
rect 5196 -14311 5924 -14258
rect 5977 -14311 6279 -14258
rect 6332 -14311 6636 -14258
rect 6689 -14311 6991 -14258
rect 7044 -14310 8417 -14258
rect 8772 -14258 8825 -14248
rect 9127 -14258 9180 -14249
rect 9483 -14258 9536 -14248
rect 9837 -14258 9890 -14249
rect 10196 -14258 10249 -14248
rect 10550 -14258 10603 -14248
rect 10908 -14258 10961 -14248
rect 8470 -14310 8772 -14258
rect 7044 -14311 8772 -14310
rect 8825 -14259 9483 -14258
rect 8825 -14311 9127 -14259
rect 5143 -14321 5196 -14311
rect 5924 -14321 5977 -14311
rect 6279 -14321 6332 -14311
rect 6636 -14321 6689 -14311
rect 6991 -14321 7044 -14311
rect 8417 -14320 8470 -14311
rect 8772 -14321 8825 -14311
rect 9180 -14311 9483 -14259
rect 9536 -14259 10196 -14258
rect 9536 -14311 9837 -14259
rect 9127 -14322 9180 -14312
rect 9483 -14321 9536 -14311
rect 9890 -14311 10196 -14259
rect 10249 -14311 10550 -14258
rect 10603 -14311 10908 -14258
rect 9837 -14322 9890 -14312
rect 10196 -14321 10249 -14311
rect 10550 -14321 10603 -14311
rect 10908 -14321 10961 -14311
rect 11087 -14256 11140 -14248
rect 11440 -14256 11493 -14246
rect 11087 -14258 11440 -14256
rect 11140 -14308 11440 -14258
rect 11140 -14309 11192 -14308
rect 11087 -14321 11140 -14311
rect 11440 -14319 11493 -14309
rect 8504 -14406 8557 -14396
rect 6993 -14424 7046 -14414
rect 7347 -14424 7400 -14414
rect 7704 -14424 7757 -14415
rect 7046 -14477 7347 -14424
rect 7400 -14425 7757 -14424
rect 7400 -14477 7704 -14425
rect 6993 -14487 7046 -14477
rect 7347 -14487 7400 -14477
rect 7704 -14488 7757 -14478
rect 8060 -14421 8113 -14411
rect 8113 -14459 8504 -14421
rect 9753 -14406 9806 -14396
rect 8557 -14459 9753 -14421
rect 10195 -14421 10248 -14412
rect 9806 -14422 10248 -14421
rect 9806 -14459 10195 -14422
rect 8113 -14474 10195 -14459
rect 8060 -14484 8113 -14474
rect 10195 -14485 10248 -14475
rect 10552 -14414 10605 -14405
rect 10908 -14413 10961 -14403
rect 10552 -14415 10908 -14414
rect 10605 -14466 10908 -14415
rect 10961 -14414 11013 -14413
rect 11264 -14414 11317 -14405
rect 10961 -14415 11317 -14414
rect 10961 -14466 11264 -14415
rect 10552 -14478 10605 -14468
rect 10908 -14476 10961 -14466
rect 11264 -14478 11317 -14468
rect -847 -14526 -794 -14516
rect -669 -14526 -616 -14516
rect -491 -14526 -438 -14516
rect -314 -14526 -261 -14517
rect -137 -14526 -84 -14516
rect 43 -14526 96 -14516
rect 1289 -14526 1342 -14517
rect 1467 -14526 1520 -14516
rect 1644 -14526 1697 -14516
rect 1822 -14526 1875 -14516
rect 1999 -14526 2052 -14516
rect 2180 -14526 2233 -14516
rect 3425 -14526 3478 -14516
rect 3603 -14526 3656 -14516
rect 3780 -14526 3833 -14516
rect 4239 -14526 4292 -14516
rect -794 -14579 -669 -14526
rect -616 -14579 -491 -14526
rect -438 -14527 -137 -14526
rect -438 -14579 -314 -14527
rect -847 -14589 -794 -14579
rect -669 -14589 -616 -14579
rect -491 -14589 -438 -14579
rect -261 -14579 -137 -14527
rect -84 -14579 43 -14526
rect 96 -14527 1467 -14526
rect 96 -14579 1289 -14527
rect -314 -14590 -261 -14580
rect -137 -14589 -84 -14579
rect 43 -14589 96 -14579
rect 1342 -14579 1467 -14527
rect 1520 -14579 1644 -14526
rect 1697 -14579 1822 -14526
rect 1875 -14579 1999 -14526
rect 2052 -14579 2180 -14526
rect 2233 -14579 3425 -14526
rect 3478 -14579 3603 -14526
rect 3656 -14579 3780 -14526
rect 3833 -14579 4239 -14526
rect 1289 -14590 1342 -14580
rect 1467 -14589 1520 -14579
rect 1644 -14589 1697 -14579
rect 1822 -14589 1875 -14579
rect 1999 -14589 2052 -14579
rect 2180 -14589 2233 -14579
rect 3425 -14589 3478 -14579
rect 3603 -14589 3656 -14579
rect 3780 -14589 3833 -14579
rect 4239 -14589 4292 -14579
rect 7080 -14523 7133 -14513
rect 7260 -14523 7313 -14514
rect 7439 -14523 7492 -14513
rect 8327 -14523 8380 -14513
rect 8505 -14523 8558 -14514
rect 8683 -14523 8736 -14514
rect 9572 -14523 9625 -14513
rect 9750 -14523 9803 -14513
rect 9929 -14523 9982 -14513
rect 10819 -14523 10872 -14513
rect 10996 -14523 11049 -14513
rect 11175 -14523 11228 -14513
rect 7133 -14524 7439 -14523
rect 7133 -14576 7260 -14524
rect 7080 -14586 7133 -14576
rect 7313 -14576 7439 -14524
rect 7492 -14576 8327 -14523
rect 8380 -14524 9572 -14523
rect 8380 -14576 8505 -14524
rect 7260 -14587 7313 -14577
rect 7439 -14586 7492 -14576
rect 8327 -14586 8380 -14576
rect 8558 -14576 8683 -14524
rect 8505 -14587 8558 -14577
rect 8736 -14576 9572 -14524
rect 9625 -14576 9750 -14523
rect 9803 -14576 9929 -14523
rect 9982 -14576 10819 -14523
rect 10872 -14576 10996 -14523
rect 11049 -14576 11175 -14523
rect 8683 -14587 8736 -14577
rect 9572 -14586 9625 -14576
rect 9750 -14586 9803 -14576
rect 9929 -14586 9982 -14576
rect 10819 -14586 10872 -14576
rect 10996 -14586 11049 -14576
rect 11175 -14586 11228 -14576
rect -6159 -14681 -6106 -14672
rect -5504 -14681 -5451 -14671
rect -4792 -14681 -4739 -14671
rect -6159 -14682 -5504 -14681
rect -6106 -14734 -5504 -14682
rect -5451 -14734 -4792 -14681
rect -6159 -14745 -6106 -14735
rect -5504 -14744 -5451 -14734
rect -4792 -14744 -4739 -14734
rect -5860 -14788 -5807 -14778
rect -5148 -14789 -5095 -14779
rect -4435 -14789 -4383 -14779
rect -3935 -14789 -3883 -14779
rect -5807 -14841 -5148 -14789
rect -5860 -14851 -5807 -14841
rect -5095 -14841 -4435 -14789
rect -4383 -14841 -3935 -14789
rect -5148 -14852 -5095 -14842
rect -4435 -14851 -4383 -14841
rect -3935 -14851 -3883 -14841
rect 4238 -15139 4291 -15129
rect 5031 -15139 5084 -15130
rect 5745 -15139 5798 -15129
rect 6101 -15139 6154 -15129
rect 6458 -15139 6511 -15129
rect 11798 -15139 11851 -15130
rect 12155 -15139 12208 -15129
rect 12511 -15139 12564 -15129
rect 4291 -15140 5745 -15139
rect 4291 -15192 5031 -15140
rect 4238 -15202 4291 -15192
rect 5084 -15192 5745 -15140
rect 5798 -15192 6101 -15139
rect 6154 -15192 6458 -15139
rect 6511 -15140 12155 -15139
rect 6511 -15192 11798 -15140
rect 5031 -15203 5084 -15193
rect 5745 -15202 5798 -15192
rect 6101 -15202 6154 -15192
rect 6458 -15202 6511 -15192
rect 11851 -15192 12155 -15140
rect 12208 -15192 12511 -15139
rect 11798 -15203 11851 -15193
rect 12155 -15202 12208 -15192
rect 12511 -15202 12564 -15192
rect 5400 -15252 5453 -15243
rect 5923 -15252 5976 -15242
rect 6279 -15252 6332 -15242
rect 6635 -15252 6688 -15242
rect 11619 -15252 11672 -15242
rect 11975 -15252 12028 -15242
rect 12332 -15252 12385 -15242
rect 5400 -15253 5923 -15252
rect 5453 -15305 5923 -15253
rect 5976 -15305 6279 -15252
rect 6332 -15305 6635 -15252
rect 6688 -15305 11619 -15252
rect 11672 -15305 11975 -15252
rect 12028 -15305 12332 -15252
rect 5400 -15316 5453 -15306
rect 5923 -15315 5976 -15305
rect 6279 -15315 6332 -15305
rect 6635 -15315 6688 -15305
rect 11619 -15315 11672 -15305
rect 11975 -15315 12028 -15305
rect 12332 -15315 12385 -15305
rect 5747 -15350 5800 -15340
rect 6101 -15349 6154 -15339
rect -6159 -15393 -6106 -15383
rect -5504 -15393 -5451 -15383
rect -4792 -15393 -4739 -15383
rect -6106 -15446 -5504 -15393
rect -5451 -15446 -4792 -15393
rect 5800 -15402 6101 -15350
rect 6456 -15350 6509 -15340
rect 6713 -15350 6766 -15341
rect 7169 -15350 7222 -15340
rect 7526 -15349 7579 -15339
rect 6154 -15402 6456 -15350
rect 5800 -15403 6456 -15402
rect 6509 -15351 7169 -15350
rect 6509 -15403 6713 -15351
rect -6159 -15456 -6106 -15446
rect -5504 -15456 -5451 -15446
rect -4792 -15456 -4739 -15446
rect -2447 -15421 -2394 -15411
rect -2005 -15421 -1952 -15412
rect -2394 -15422 -1952 -15421
rect -1649 -15422 -1596 -15412
rect -1293 -15422 -1240 -15412
rect -937 -15422 -884 -15412
rect -581 -15422 -528 -15412
rect -225 -15422 -172 -15412
rect 132 -15421 185 -15411
rect -2394 -15474 -2005 -15422
rect -2447 -15484 -2394 -15474
rect -1952 -15475 -1649 -15422
rect -1596 -15475 -1293 -15422
rect -1240 -15475 -937 -15422
rect -884 -15475 -581 -15422
rect -528 -15475 -225 -15422
rect -172 -15474 132 -15422
rect 487 -15422 540 -15412
rect 843 -15422 896 -15412
rect 1201 -15422 1254 -15412
rect 1555 -15422 1608 -15412
rect 1910 -15422 1963 -15412
rect 2267 -15422 2320 -15412
rect 2624 -15422 2677 -15412
rect 2979 -15422 3032 -15412
rect 3335 -15422 3388 -15412
rect 3692 -15422 3745 -15412
rect 5747 -15413 5800 -15403
rect 6101 -15412 6154 -15403
rect 6456 -15413 6509 -15403
rect 6766 -15403 7169 -15351
rect 7222 -15402 7526 -15350
rect 7882 -15349 7935 -15339
rect 7579 -15402 7882 -15350
rect 10373 -15350 10426 -15341
rect 10730 -15350 10783 -15340
rect 11086 -15350 11139 -15340
rect 7935 -15351 10730 -15350
rect 7935 -15402 10373 -15351
rect 7222 -15403 10373 -15402
rect 6713 -15414 6766 -15404
rect 7169 -15413 7222 -15403
rect 7526 -15412 7579 -15403
rect 7882 -15412 7935 -15403
rect 10426 -15403 10730 -15351
rect 10783 -15403 11086 -15350
rect 10373 -15414 10426 -15404
rect 10730 -15413 10783 -15403
rect 11086 -15413 11139 -15403
rect 185 -15474 487 -15422
rect -172 -15475 487 -15474
rect 540 -15475 843 -15422
rect 896 -15475 1201 -15422
rect 1254 -15475 1555 -15422
rect 1608 -15475 1910 -15422
rect 1963 -15475 2267 -15422
rect 2320 -15475 2624 -15422
rect 2677 -15475 2979 -15422
rect 3032 -15475 3335 -15422
rect 3388 -15475 3692 -15422
rect 11440 -15441 11493 -15431
rect -5860 -15494 -5807 -15484
rect -5148 -15494 -5095 -15484
rect -4436 -15494 -4383 -15484
rect -2005 -15485 -1952 -15475
rect -1649 -15485 -1596 -15475
rect -1293 -15485 -1240 -15475
rect -937 -15485 -884 -15475
rect -581 -15485 -528 -15475
rect -225 -15485 -172 -15475
rect 132 -15484 185 -15475
rect 487 -15485 540 -15475
rect 843 -15485 896 -15475
rect 1201 -15485 1254 -15475
rect 1555 -15485 1608 -15475
rect 1910 -15485 1963 -15475
rect 2267 -15485 2320 -15475
rect 2624 -15485 2677 -15475
rect 2979 -15485 3032 -15475
rect 3335 -15485 3388 -15475
rect 3692 -15485 3745 -15475
rect 6813 -15451 6866 -15441
rect 7169 -15451 7222 -15442
rect 8060 -15451 8113 -15441
rect 8593 -15451 8646 -15442
rect 9663 -15451 9716 -15442
rect 10194 -15451 10247 -15442
rect 11084 -15451 11137 -15442
rect -3935 -15494 -3883 -15485
rect -5807 -15547 -5148 -15494
rect -5095 -15546 -4436 -15494
rect -5860 -15557 -5807 -15547
rect -5148 -15557 -5095 -15547
rect -4383 -15495 -3883 -15494
rect -4383 -15546 -3935 -15495
rect -4436 -15557 -4383 -15547
rect 6866 -15452 8060 -15451
rect 6866 -15504 7169 -15452
rect 6813 -15514 6866 -15504
rect 7222 -15504 8060 -15452
rect 8113 -15452 11440 -15451
rect 8113 -15504 8593 -15452
rect 7169 -15515 7222 -15505
rect 8060 -15514 8113 -15504
rect 8646 -15504 9663 -15452
rect 8593 -15515 8646 -15505
rect 9716 -15504 10194 -15452
rect 9663 -15515 9716 -15505
rect 10247 -15504 11084 -15452
rect 10194 -15515 10247 -15505
rect 11137 -15494 11440 -15452
rect 11137 -15504 11493 -15494
rect 11084 -15515 11137 -15505
rect -3935 -15557 -3883 -15547
rect -1915 -15533 -1862 -15523
rect -1738 -15533 -1685 -15523
rect -1560 -15533 -1507 -15523
rect -1382 -15533 -1329 -15523
rect -1204 -15533 -1151 -15523
rect -1025 -15533 -972 -15523
rect -847 -15533 -794 -15523
rect -670 -15533 -617 -15523
rect -491 -15533 -438 -15523
rect -313 -15533 -260 -15523
rect -136 -15533 -83 -15523
rect 43 -15533 96 -15523
rect 221 -15533 274 -15523
rect 398 -15533 451 -15523
rect 575 -15533 628 -15523
rect 755 -15533 808 -15523
rect 931 -15533 984 -15523
rect 1110 -15533 1163 -15523
rect 1289 -15533 1342 -15523
rect 1466 -15533 1519 -15523
rect 1643 -15533 1696 -15523
rect 1822 -15533 1875 -15523
rect 2000 -15533 2053 -15523
rect 2179 -15533 2232 -15523
rect 2356 -15533 2409 -15523
rect 2534 -15533 2587 -15523
rect 2712 -15533 2765 -15523
rect 2891 -15533 2944 -15523
rect 3068 -15533 3121 -15523
rect 3247 -15533 3300 -15523
rect 3424 -15533 3477 -15523
rect 3603 -15533 3656 -15523
rect 3780 -15533 3833 -15523
rect -1862 -15586 -1738 -15533
rect -1685 -15586 -1560 -15533
rect -1507 -15586 -1382 -15533
rect -1329 -15586 -1204 -15533
rect -1151 -15586 -1025 -15533
rect -972 -15586 -847 -15533
rect -794 -15586 -670 -15533
rect -617 -15586 -491 -15533
rect -438 -15586 -313 -15533
rect -260 -15586 -136 -15533
rect -83 -15586 43 -15533
rect 96 -15586 221 -15533
rect 274 -15586 398 -15533
rect 451 -15586 575 -15533
rect 628 -15586 755 -15533
rect 808 -15586 931 -15533
rect 984 -15586 1110 -15533
rect 1163 -15586 1289 -15533
rect 1342 -15586 1466 -15533
rect 1519 -15586 1643 -15533
rect 1696 -15586 1822 -15533
rect 1875 -15586 2000 -15533
rect 2053 -15586 2179 -15533
rect 2232 -15586 2356 -15533
rect 2409 -15586 2534 -15533
rect 2587 -15586 2712 -15533
rect 2765 -15586 2891 -15533
rect 2944 -15586 3068 -15533
rect 3121 -15586 3247 -15533
rect 3300 -15586 3424 -15533
rect 3477 -15586 3603 -15533
rect 3656 -15586 3780 -15533
rect -1915 -15596 -1862 -15586
rect -1738 -15596 -1685 -15586
rect -1560 -15596 -1507 -15586
rect -1382 -15596 -1329 -15586
rect -1204 -15596 -1151 -15586
rect -1025 -15596 -972 -15586
rect -847 -15596 -794 -15586
rect -670 -15596 -617 -15586
rect -491 -15596 -438 -15586
rect -313 -15596 -260 -15586
rect -136 -15596 -83 -15586
rect 43 -15596 96 -15586
rect 221 -15596 274 -15586
rect 398 -15596 451 -15586
rect 575 -15596 628 -15586
rect 755 -15596 808 -15586
rect 931 -15596 984 -15586
rect 1110 -15596 1163 -15586
rect 1289 -15596 1342 -15586
rect 1466 -15596 1519 -15586
rect 1643 -15596 1696 -15586
rect 1822 -15596 1875 -15586
rect 2000 -15596 2053 -15586
rect 2179 -15596 2232 -15586
rect 2356 -15596 2409 -15586
rect 2534 -15596 2587 -15586
rect 2712 -15596 2765 -15586
rect 2891 -15596 2944 -15586
rect 3068 -15596 3121 -15586
rect 3247 -15596 3300 -15586
rect 3424 -15596 3477 -15586
rect 3603 -15596 3656 -15586
rect 3780 -15596 3833 -15586
rect 5921 -15547 5974 -15538
rect 6279 -15547 6332 -15538
rect 6634 -15547 6687 -15538
rect 6994 -15547 7047 -15541
rect 5921 -15548 7047 -15547
rect 5974 -15600 6279 -15548
rect 5921 -15611 5974 -15601
rect 6332 -15600 6634 -15548
rect 6279 -15611 6332 -15601
rect 6687 -15551 7047 -15548
rect 6687 -15600 6994 -15551
rect 6634 -15611 6687 -15601
rect 6994 -15614 7047 -15604
rect 7526 -15552 7579 -15543
rect 7881 -15552 7934 -15542
rect 8237 -15552 8290 -15542
rect 11441 -15552 11494 -15542
rect 11797 -15552 11850 -15542
rect 12154 -15552 12207 -15542
rect 12511 -15552 12564 -15542
rect 7526 -15553 7881 -15552
rect 7579 -15605 7881 -15553
rect 7934 -15605 8237 -15552
rect 8290 -15605 11441 -15552
rect 11494 -15605 11797 -15552
rect 11850 -15605 12154 -15552
rect 12207 -15605 12511 -15552
rect 7526 -15616 7579 -15606
rect 7881 -15615 7934 -15605
rect 8237 -15615 8290 -15605
rect 11441 -15615 11494 -15605
rect 11797 -15615 11850 -15605
rect 12154 -15615 12207 -15605
rect 12511 -15615 12564 -15605
rect -5682 -16086 -5629 -16076
rect -5326 -16086 -5273 -16076
rect -4970 -16086 -4917 -16076
rect -4614 -16086 -4561 -16076
rect -4258 -16086 -4205 -16076
rect -5629 -16139 -5326 -16086
rect -5273 -16139 -4970 -16086
rect -4917 -16139 -4614 -16086
rect -4561 -16139 -4258 -16086
rect -5682 -16149 -5629 -16139
rect -5326 -16149 -5273 -16139
rect -4970 -16149 -4917 -16139
rect -4614 -16149 -4561 -16139
rect -4258 -16149 -4205 -16139
rect -1917 -16142 -1864 -16132
rect -1738 -16142 -1685 -16132
rect -1561 -16141 -1508 -16131
rect -1864 -16195 -1738 -16142
rect -1685 -16194 -1561 -16142
rect -1381 -16142 -1328 -16133
rect -1204 -16142 -1151 -16132
rect -1026 -16142 -973 -16132
rect 220 -16142 273 -16132
rect 397 -16142 450 -16132
rect 576 -16142 629 -16132
rect 755 -16142 808 -16132
rect 933 -16142 986 -16132
rect 1111 -16142 1164 -16132
rect 2356 -16142 2409 -16132
rect 2534 -16142 2587 -16132
rect 2713 -16141 2766 -16131
rect -1508 -16143 -1204 -16142
rect -1508 -16194 -1381 -16143
rect -1685 -16195 -1381 -16194
rect -6159 -16207 -6106 -16197
rect -5859 -16207 -5806 -16197
rect -5148 -16207 -5095 -16197
rect -4437 -16207 -4384 -16197
rect -1917 -16205 -1864 -16195
rect -1738 -16205 -1685 -16195
rect -1561 -16204 -1508 -16195
rect -1328 -16195 -1204 -16143
rect -1151 -16195 -1026 -16142
rect -973 -16195 220 -16142
rect 273 -16195 397 -16142
rect 450 -16195 576 -16142
rect 629 -16195 755 -16142
rect 808 -16195 933 -16142
rect 986 -16195 1111 -16142
rect 1164 -16195 2356 -16142
rect 2409 -16195 2534 -16142
rect 2587 -16194 2713 -16142
rect 2891 -16142 2944 -16132
rect 3070 -16142 3123 -16132
rect 3249 -16142 3302 -16132
rect 4238 -16142 4291 -16132
rect 2766 -16194 2891 -16142
rect 2587 -16195 2891 -16194
rect 2944 -16195 3070 -16142
rect 3123 -16195 3249 -16142
rect 3302 -16195 4238 -16142
rect -1381 -16206 -1328 -16196
rect -1204 -16205 -1151 -16195
rect -1026 -16205 -973 -16195
rect 220 -16205 273 -16195
rect 397 -16205 450 -16195
rect 576 -16205 629 -16195
rect 755 -16205 808 -16195
rect 933 -16205 986 -16195
rect 1111 -16205 1164 -16195
rect 2356 -16205 2409 -16195
rect 2534 -16205 2587 -16195
rect 2713 -16204 2766 -16195
rect 2891 -16205 2944 -16195
rect 3070 -16205 3123 -16195
rect 3249 -16205 3302 -16195
rect 4238 -16205 4291 -16195
rect 6548 -16144 6601 -16134
rect 6726 -16144 6779 -16134
rect 6601 -16197 6726 -16145
rect 6903 -16145 6956 -16135
rect 7970 -16145 8023 -16135
rect 8149 -16144 8202 -16134
rect 6779 -16197 6903 -16145
rect 6548 -16198 6903 -16197
rect 6956 -16198 7970 -16145
rect 8023 -16197 8149 -16145
rect 9929 -16144 9982 -16134
rect 8202 -16197 9929 -16145
rect 10107 -16145 10160 -16135
rect 10287 -16145 10340 -16135
rect 11352 -16145 11405 -16135
rect 11530 -16145 11583 -16136
rect 11709 -16145 11762 -16135
rect 9982 -16197 10107 -16145
rect 8023 -16198 10107 -16197
rect 10160 -16198 10287 -16145
rect 10340 -16198 11352 -16145
rect 11405 -16146 11709 -16145
rect 11405 -16198 11530 -16146
rect 6548 -16207 6601 -16198
rect 6726 -16207 6779 -16198
rect -6106 -16260 -5859 -16207
rect -5806 -16260 -5148 -16207
rect -5095 -16260 -4437 -16207
rect 6903 -16208 6956 -16198
rect 7970 -16208 8023 -16198
rect 8149 -16207 8202 -16198
rect 9929 -16207 9982 -16198
rect 10107 -16208 10160 -16198
rect 10287 -16208 10340 -16198
rect 11352 -16208 11405 -16198
rect 11583 -16198 11709 -16146
rect 11530 -16209 11583 -16199
rect 11709 -16208 11762 -16198
rect -6159 -16270 -6106 -16260
rect -5859 -16270 -5806 -16260
rect -5148 -16270 -5095 -16260
rect -4437 -16270 -4384 -16260
rect -1827 -16265 -1774 -16255
rect -1471 -16265 -1418 -16256
rect -1114 -16265 -1061 -16255
rect -759 -16264 -706 -16254
rect -5504 -16318 -5451 -16308
rect -4792 -16318 -4739 -16308
rect -3935 -16318 -3883 -16308
rect -5451 -16370 -4792 -16318
rect -5504 -16381 -5451 -16371
rect -4739 -16370 -3935 -16318
rect -1774 -16266 -1114 -16265
rect -1774 -16318 -1471 -16266
rect -1827 -16328 -1774 -16318
rect -1418 -16318 -1114 -16266
rect -1061 -16317 -759 -16265
rect -403 -16265 -350 -16255
rect -47 -16265 6 -16255
rect 309 -16265 362 -16256
rect 665 -16265 718 -16255
rect 845 -16265 898 -16255
rect 1021 -16265 1074 -16255
rect 1377 -16265 1430 -16255
rect 1735 -16265 1788 -16255
rect 2090 -16264 2143 -16254
rect -706 -16317 -403 -16265
rect -1061 -16318 -403 -16317
rect -350 -16318 -47 -16265
rect 6 -16266 665 -16265
rect 6 -16318 309 -16266
rect -1471 -16329 -1418 -16319
rect -1114 -16328 -1061 -16318
rect -759 -16327 -706 -16318
rect -403 -16328 -350 -16318
rect -47 -16328 6 -16318
rect 362 -16318 665 -16266
rect 718 -16318 845 -16265
rect 898 -16318 1021 -16265
rect 1074 -16318 1377 -16265
rect 1430 -16318 1735 -16265
rect 1788 -16317 2090 -16265
rect 2445 -16265 2498 -16255
rect 2801 -16265 2854 -16255
rect 3157 -16264 3210 -16254
rect 2143 -16317 2445 -16265
rect 1788 -16318 2445 -16317
rect 2498 -16318 2801 -16265
rect 2854 -16317 3157 -16265
rect 3514 -16265 3567 -16256
rect 3868 -16265 3921 -16255
rect 3210 -16266 3868 -16265
rect 3210 -16317 3514 -16266
rect 2854 -16318 3514 -16317
rect 309 -16329 362 -16319
rect 665 -16328 718 -16318
rect 845 -16328 898 -16318
rect 1021 -16328 1074 -16318
rect 1377 -16328 1430 -16318
rect 1735 -16328 1788 -16318
rect 2090 -16327 2143 -16318
rect 2445 -16328 2498 -16318
rect 2801 -16328 2854 -16318
rect 3157 -16327 3210 -16318
rect 3567 -16318 3868 -16266
rect 3514 -16329 3567 -16319
rect 3868 -16328 3921 -16318
rect 5399 -16266 5452 -16257
rect 8771 -16266 8824 -16256
rect 9128 -16266 9181 -16256
rect 9484 -16266 9537 -16256
rect 5399 -16267 8771 -16266
rect 5452 -16319 8771 -16267
rect 8824 -16319 9128 -16266
rect 9181 -16319 9484 -16266
rect 5399 -16330 5452 -16320
rect 8771 -16329 8824 -16319
rect 9128 -16329 9181 -16319
rect 9484 -16329 9537 -16319
rect 9838 -16265 9891 -16256
rect 10195 -16265 10248 -16255
rect 10550 -16265 10603 -16255
rect 10907 -16265 10960 -16255
rect 9838 -16266 10195 -16265
rect 9891 -16318 10195 -16266
rect 10248 -16318 10550 -16265
rect 10603 -16318 10907 -16265
rect 9838 -16329 9891 -16319
rect 10195 -16328 10248 -16318
rect 10550 -16328 10603 -16318
rect 10907 -16328 10960 -16318
rect -4792 -16381 -4739 -16371
rect -3935 -16380 -3883 -16370
rect 5031 -16382 5084 -16372
rect 8950 -16382 9003 -16372
rect 9305 -16382 9358 -16372
rect 5084 -16435 8950 -16382
rect 9003 -16435 9305 -16382
rect 5031 -16445 5084 -16435
rect 8950 -16445 9003 -16435
rect 9305 -16445 9358 -16435
rect 10017 -16380 10070 -16371
rect 10374 -16380 10427 -16371
rect 10731 -16379 10784 -16369
rect 10017 -16381 10731 -16380
rect 10070 -16433 10374 -16381
rect 10017 -16444 10070 -16434
rect 10427 -16432 10731 -16381
rect 10427 -16433 10784 -16432
rect 10374 -16444 10427 -16434
rect 10731 -16442 10784 -16433
rect 7347 -16490 7400 -16480
rect 7704 -16490 7757 -16480
rect 8060 -16490 8113 -16480
rect 8416 -16490 8469 -16480
rect 11263 -16490 11316 -16480
rect 11620 -16490 11673 -16480
rect 11975 -16489 12028 -16479
rect 7400 -16543 7704 -16490
rect 7757 -16543 8060 -16490
rect 8113 -16543 8416 -16490
rect 8469 -16543 11263 -16490
rect 11316 -16543 11620 -16490
rect 11673 -16542 11975 -16490
rect 12331 -16489 12384 -16479
rect 12028 -16542 12331 -16490
rect 11673 -16543 12384 -16542
rect 7347 -16553 7400 -16543
rect 7704 -16553 7757 -16543
rect 8060 -16553 8113 -16543
rect 8416 -16553 8469 -16543
rect 11263 -16553 11316 -16543
rect 11620 -16553 11673 -16543
rect 11975 -16552 12028 -16543
rect 12331 -16552 12384 -16543
<< via2 >>
rect 3019 -3513 3080 -3452
rect -2546 -3989 -2485 -3928
rect 2538 -4327 2599 -4266
rect -2385 -4566 -2324 -4505
rect 2746 -4507 2807 -4446
rect 3021 -5063 3082 -5002
rect -2385 -5154 -2324 -5093
rect 311 -5209 372 -5148
rect -1646 -5339 -1585 -5278
rect 846 -5339 907 -5278
rect -3545 -6867 -3484 -6806
rect -3386 -7040 -3325 -6979
<< metal3 >>
rect 3009 -3452 3090 -3447
rect 3009 -3513 3019 -3452
rect 3080 -3513 3090 -3452
rect 3009 -3518 3090 -3513
rect -2556 -3928 -2475 -3923
rect -2556 -3989 -2546 -3928
rect -2485 -3989 -2475 -3928
rect -2556 -3994 -2475 -3989
rect -2546 -4266 -2485 -3994
rect 2528 -4266 2609 -4261
rect -2546 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect -2546 -6637 -2485 -4327
rect 2528 -4332 2609 -4327
rect 2736 -4446 2817 -4441
rect -2385 -4500 2746 -4446
rect -2395 -4505 2746 -4500
rect -2395 -4566 -2385 -4505
rect -2324 -4507 2746 -4505
rect 2807 -4507 2817 -4446
rect -2324 -4566 -2314 -4507
rect 2736 -4512 2817 -4507
rect -2395 -4571 -2314 -4566
rect -2385 -5088 -2324 -4571
rect 3021 -4997 3082 -3518
rect 3011 -5002 3092 -4997
rect 3011 -5063 3021 -5002
rect 3082 -5063 3092 -5002
rect 3011 -5068 3092 -5063
rect -2395 -5093 -2314 -5088
rect -2395 -5154 -2385 -5093
rect -2324 -5154 -2314 -5093
rect -2395 -5159 -2314 -5154
rect 301 -5147 382 -5143
rect 3021 -5147 3082 -5068
rect 301 -5148 3082 -5147
rect -3545 -6698 -2485 -6637
rect -3545 -6801 -3484 -6698
rect -2385 -6786 -2324 -5159
rect 301 -5209 311 -5148
rect 372 -5208 3082 -5148
rect 372 -5209 382 -5208
rect 301 -5214 382 -5209
rect -1656 -5278 -1575 -5273
rect 836 -5278 917 -5273
rect -1656 -5339 -1646 -5278
rect -1585 -5339 846 -5278
rect 907 -5339 917 -5278
rect -1656 -5344 -1575 -5339
rect 836 -5344 917 -5339
rect -3555 -6806 -3474 -6801
rect -3555 -6867 -3545 -6806
rect -3484 -6867 -3474 -6806
rect -3555 -6872 -3474 -6867
rect -3386 -6847 -2324 -6786
rect -3386 -6974 -3325 -6847
rect -3396 -6979 -3315 -6974
rect -3396 -7040 -3386 -6979
rect -3325 -7040 -3315 -6979
rect -3396 -7045 -3315 -7040
use sky130_fd_pr__nfet_01v8_7P4E2J  sky130_fd_pr__nfet_01v8_7P4E2J_0
timestamp 1653466640
transform 1 0 7953 0 1 -8622
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_7P4E2J  sky130_fd_pr__nfet_01v8_7P4E2J_1
timestamp 1653466640
transform 1 0 7953 0 1 -9522
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_7P4E2J  sky130_fd_pr__nfet_01v8_7P4E2J_2
timestamp 1653466640
transform 1 0 7953 0 1 -10422
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_7P4E2J  sky130_fd_pr__nfet_01v8_7P4E2J_3
timestamp 1653466640
transform 1 0 7953 0 1 -11322
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_0
timestamp 1653033955
transform 1 0 -5032 0 1 -13722
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_1
timestamp 1653033955
transform 1 0 -5032 0 1 -14422
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_2
timestamp 1653033955
transform 1 0 -5032 0 1 -15122
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BASQVB  sky130_fd_pr__nfet_01v8_BASQVB_3
timestamp 1653033955
transform 1 0 -5032 0 1 -15822
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_4
timestamp 1653030110
transform 1 0 959 0 1 -14860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_5
timestamp 1653030110
transform 1 0 959 0 1 -13860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_6
timestamp 1653030110
transform 1 0 959 0 1 -12860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_7
timestamp 1653030110
transform 1 0 959 0 1 -11860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_8
timestamp 1653030110
transform 1 0 959 0 1 -10860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_9
timestamp 1653030110
transform 1 0 959 0 1 -9860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_10
timestamp 1653030110
transform 1 0 959 0 1 -8860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_11
timestamp 1653030110
transform 1 0 959 0 1 -7860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_KEEN2X  sky130_fd_pr__nfet_01v8_KEEN2X_12
timestamp 1653030110
transform 1 0 959 0 1 -15860
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_UFQYRB  sky130_fd_pr__nfet_01v8_UFQYRB_0
timestamp 1653386003
transform 1 0 9154 0 1 -13860
box -3589 -228 3589 228
use sky130_fd_pr__nfet_01v8_UFQYRB  sky130_fd_pr__nfet_01v8_UFQYRB_1
timestamp 1653386003
transform 1 0 9154 0 1 -14860
box -3589 -228 3589 228
use sky130_fd_pr__nfet_01v8_UFQYRB  sky130_fd_pr__nfet_01v8_UFQYRB_2
timestamp 1653386003
transform 1 0 9154 0 1 -15860
box -3589 -228 3589 228
use sky130_fd_pr__nfet_01v8_VJ4JGY  sky130_fd_pr__nfet_01v8_VJ4JGY_0
timestamp 1653472245
transform 1 0 11754 0 1 -8652
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_VJ4JGY  sky130_fd_pr__nfet_01v8_VJ4JGY_1
timestamp 1653472245
transform 1 0 11754 0 1 -9422
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_VJ4JGY  sky130_fd_pr__nfet_01v8_VJ4JGY_2
timestamp 1653472245
transform 1 0 11754 0 1 -10192
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_VJ4JGY  sky130_fd_pr__nfet_01v8_VJ4JGY_3
timestamp 1653472245
transform 1 0 11754 0 1 -10962
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_0
timestamp 1653028559
transform 1 0 -5850 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_1
timestamp 1653028559
transform 1 0 -5850 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_2
timestamp 1653028559
transform 1 0 -5600 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_3
timestamp 1653028559
transform 1 0 -5350 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_4
timestamp 1653028559
transform 1 0 -5100 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_5
timestamp 1653028559
transform 1 0 -4850 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_6
timestamp 1653028559
transform 1 0 -4600 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_7
timestamp 1653028559
transform 1 0 -4350 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_8
timestamp 1653028559
transform 1 0 -4100 0 1 -12700
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_9
timestamp 1653028559
transform 1 0 -5600 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_10
timestamp 1653028559
transform 1 0 -5350 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_11
timestamp 1653028559
transform 1 0 -5100 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_12
timestamp 1653028559
transform 1 0 -4850 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_13
timestamp 1653028559
transform 1 0 -4600 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_14
timestamp 1653028559
transform 1 0 -4350 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_TRAZV8  sky130_fd_pr__nfet_01v8_lvt_TRAZV8_15
timestamp 1653028559
transform 1 0 -4100 0 1 -12020
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_0
timestamp 1653032550
transform 1 0 -4810 0 1 -7752
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_1
timestamp 1653032550
transform 1 0 -4810 0 1 -8302
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_2
timestamp 1653032550
transform 1 0 -4810 0 1 -8852
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_3
timestamp 1653032550
transform 1 0 -4810 0 1 -9402
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_4
timestamp 1653032550
transform 1 0 -4810 0 1 -9952
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_5
timestamp 1653032550
transform 1 0 -4810 0 1 -10502
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_VU7MNH  sky130_fd_pr__nfet_01v8_lvt_VU7MNH_6
timestamp 1653032550
transform 1 0 -4810 0 1 -11052
box -830 -228 830 228
use sky130_fd_pr__pfet_01v8_E4DCBA  sky130_fd_pr__pfet_01v8_E4DCBA_0
timestamp 1653260422
transform 1 0 610 0 1 -3012
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_E4DCBA  sky130_fd_pr__pfet_01v8_E4DCBA_1
timestamp 1653260422
transform 1 0 610 0 1 -3912
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_E4DCBA  sky130_fd_pr__pfet_01v8_E4DCBA_2
timestamp 1653260422
transform 1 0 610 0 1 -4812
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_E4DCBA  sky130_fd_pr__pfet_01v8_E4DCBA_3
timestamp 1653260422
transform 1 0 610 0 1 -5712
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_0
timestamp 1653025074
transform 1 0 -4861 0 1 -2260
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_1
timestamp 1653025074
transform 1 0 -4861 0 1 -3130
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_2
timestamp 1653025074
transform 1 0 -4861 0 1 -4000
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_3
timestamp 1653025074
transform 1 0 -4861 0 1 -4870
box -1489 -240 1489 240
use sky130_fd_pr__pfet_01v8_lvt_6QKDBA  sky130_fd_pr__pfet_01v8_lvt_6QKDBA_4
timestamp 1653025074
transform 1 0 -4861 0 1 -5740
box -1489 -240 1489 240
<< labels >>
flabel metal1 -6957 -13445 -6957 -13445 1 FreeSans 1200 0 0 0 i_bias
flabel metal1 -4277 -7465 -4277 -7465 1 FreeSans 1200 0 0 0 bias_b
flabel metal1 -3636 -11523 -3636 -11523 1 FreeSans 1200 0 0 0 bias_c
flabel metal1 -6950 -11741 -6950 -11741 1 FreeSans 1200 0 0 0 ip
flabel metal1 -6952 -13080 -6952 -13080 1 FreeSans 1200 0 0 0 in
flabel metal2 5049 -9556 5049 -9556 1 FreeSans 1200 0 0 0 cmc
flabel metal1 4262 -15341 4262 -15341 1 FreeSans 1200 0 0 0 bias_a
flabel metal2 3147 -3484 3147 -3484 1 FreeSans 1200 0 0 0 on
flabel metal2 3431 -5243 3431 -5243 1 FreeSans 1200 0 0 0 op
<< end >>
