magic
tech sky130A
timestamp 1654601900
<< error_s >>
rect 129 180 158 183
rect 339 180 368 183
rect 549 180 578 183
rect 759 180 788 183
rect 969 180 998 183
rect 1179 180 1208 183
rect 1389 180 1418 183
rect 1599 180 1628 183
rect 1809 180 1838 183
rect 2019 180 2048 183
rect 2229 180 2258 183
rect 2439 180 2468 183
rect 2649 180 2678 183
rect 2859 180 2888 183
rect 3069 180 3098 183
rect 3279 180 3308 183
rect 3489 180 3518 183
rect 3699 180 3728 183
rect 3909 180 3938 183
rect 4119 180 4148 183
rect 129 163 135 180
rect 339 163 345 180
rect 549 163 555 180
rect 759 163 765 180
rect 969 163 975 180
rect 1179 163 1185 180
rect 1389 163 1395 180
rect 1599 163 1605 180
rect 1809 163 1815 180
rect 2019 163 2025 180
rect 2229 163 2235 180
rect 2439 163 2445 180
rect 2649 163 2655 180
rect 2859 163 2865 180
rect 3069 163 3075 180
rect 3279 163 3285 180
rect 3489 163 3495 180
rect 3699 163 3705 180
rect 3909 163 3915 180
rect 4119 163 4125 180
rect 129 160 158 163
rect 339 160 368 163
rect 549 160 578 163
rect 759 160 788 163
rect 969 160 998 163
rect 1179 160 1208 163
rect 1389 160 1418 163
rect 1599 160 1628 163
rect 1809 160 1838 163
rect 2019 160 2048 163
rect 2229 160 2258 163
rect 2439 160 2468 163
rect 2649 160 2678 163
rect 2859 160 2888 163
rect 3069 160 3098 163
rect 3279 160 3308 163
rect 3489 160 3518 163
rect 3699 160 3728 163
rect 3909 160 3938 163
rect 4119 160 4148 163
rect 234 25 263 28
rect 444 25 473 28
rect 654 25 683 28
rect 864 25 893 28
rect 1074 25 1103 28
rect 1284 25 1313 28
rect 1494 25 1523 28
rect 1704 25 1733 28
rect 1914 25 1943 28
rect 2124 25 2153 28
rect 2334 25 2363 28
rect 2544 25 2573 28
rect 2754 25 2783 28
rect 2964 25 2993 28
rect 3174 25 3203 28
rect 3384 25 3413 28
rect 3594 25 3623 28
rect 3804 25 3833 28
rect 4014 25 4043 28
rect 4224 25 4253 28
rect 234 8 240 25
rect 444 8 450 25
rect 654 8 660 25
rect 864 8 870 25
rect 1074 8 1080 25
rect 1284 8 1290 25
rect 1494 8 1500 25
rect 1704 8 1710 25
rect 1914 8 1920 25
rect 2124 8 2130 25
rect 2334 8 2340 25
rect 2544 8 2550 25
rect 2754 8 2760 25
rect 2964 8 2970 25
rect 3174 8 3180 25
rect 3384 8 3390 25
rect 3594 8 3600 25
rect 3804 8 3810 25
rect 4014 8 4020 25
rect 4224 8 4230 25
rect 234 5 263 8
rect 444 5 473 8
rect 654 5 683 8
rect 864 5 893 8
rect 1074 5 1103 8
rect 1284 5 1313 8
rect 1494 5 1523 8
rect 1704 5 1733 8
rect 1914 5 1943 8
rect 2124 5 2153 8
rect 2334 5 2363 8
rect 2544 5 2573 8
rect 2754 5 2783 8
rect 2964 5 2993 8
rect 3174 5 3203 8
rect 3384 5 3413 8
rect 3594 5 3623 8
rect 3804 5 3833 8
rect 4014 5 4043 8
rect 4224 5 4253 8
rect 129 -40 158 -37
rect 339 -40 368 -37
rect 549 -40 578 -37
rect 759 -40 788 -37
rect 969 -40 998 -37
rect 1179 -40 1208 -37
rect 1389 -40 1418 -37
rect 1599 -40 1628 -37
rect 1809 -40 1838 -37
rect 2019 -40 2048 -37
rect 2229 -40 2258 -37
rect 2439 -40 2468 -37
rect 2649 -40 2678 -37
rect 2859 -40 2888 -37
rect 3069 -40 3098 -37
rect 3279 -40 3308 -37
rect 3489 -40 3518 -37
rect 3699 -40 3728 -37
rect 3909 -40 3938 -37
rect 4119 -40 4148 -37
rect 129 -57 135 -40
rect 339 -57 345 -40
rect 549 -57 555 -40
rect 759 -57 765 -40
rect 969 -57 975 -40
rect 1179 -57 1185 -40
rect 1389 -57 1395 -40
rect 1599 -57 1605 -40
rect 1809 -57 1815 -40
rect 2019 -57 2025 -40
rect 2229 -57 2235 -40
rect 2439 -57 2445 -40
rect 2649 -57 2655 -40
rect 2859 -57 2865 -40
rect 3069 -57 3075 -40
rect 3279 -57 3285 -40
rect 3489 -57 3495 -40
rect 3699 -57 3705 -40
rect 3909 -57 3915 -40
rect 4119 -57 4125 -40
rect 129 -60 158 -57
rect 339 -60 368 -57
rect 549 -60 578 -57
rect 759 -60 788 -57
rect 969 -60 998 -57
rect 1179 -60 1208 -57
rect 1389 -60 1418 -57
rect 1599 -60 1628 -57
rect 1809 -60 1838 -57
rect 2019 -60 2048 -57
rect 2229 -60 2258 -57
rect 2439 -60 2468 -57
rect 2649 -60 2678 -57
rect 2859 -60 2888 -57
rect 3069 -60 3098 -57
rect 3279 -60 3308 -57
rect 3489 -60 3518 -57
rect 3699 -60 3728 -57
rect 3909 -60 3938 -57
rect 4119 -60 4148 -57
rect 234 -195 263 -192
rect 444 -195 473 -192
rect 654 -195 683 -192
rect 864 -195 893 -192
rect 1074 -195 1103 -192
rect 1284 -195 1313 -192
rect 1494 -195 1523 -192
rect 1704 -195 1733 -192
rect 1914 -195 1943 -192
rect 2124 -195 2153 -192
rect 2334 -195 2363 -192
rect 2544 -195 2573 -192
rect 2754 -195 2783 -192
rect 2964 -195 2993 -192
rect 3174 -195 3203 -192
rect 3384 -195 3413 -192
rect 3594 -195 3623 -192
rect 3804 -195 3833 -192
rect 4014 -195 4043 -192
rect 4224 -195 4253 -192
rect 234 -212 240 -195
rect 444 -212 450 -195
rect 654 -212 660 -195
rect 864 -212 870 -195
rect 1074 -212 1080 -195
rect 1284 -212 1290 -195
rect 1494 -212 1500 -195
rect 1704 -212 1710 -195
rect 1914 -212 1920 -195
rect 2124 -212 2130 -195
rect 2334 -212 2340 -195
rect 2544 -212 2550 -195
rect 2754 -212 2760 -195
rect 2964 -212 2970 -195
rect 3174 -212 3180 -195
rect 3384 -212 3390 -195
rect 3594 -212 3600 -195
rect 3804 -212 3810 -195
rect 4014 -212 4020 -195
rect 4224 -212 4230 -195
rect 234 -215 263 -212
rect 444 -215 473 -212
rect 654 -215 683 -212
rect 864 -215 893 -212
rect 1074 -215 1103 -212
rect 1284 -215 1313 -212
rect 1494 -215 1523 -212
rect 1704 -215 1733 -212
rect 1914 -215 1943 -212
rect 2124 -215 2153 -212
rect 2334 -215 2363 -212
rect 2544 -215 2573 -212
rect 2754 -215 2783 -212
rect 2964 -215 2993 -212
rect 3174 -215 3203 -212
rect 3384 -215 3413 -212
rect 3594 -215 3623 -212
rect 3804 -215 3833 -212
rect 4014 -215 4043 -212
rect 4224 -215 4253 -212
rect 129 -260 158 -257
rect 339 -260 368 -257
rect 549 -260 578 -257
rect 759 -260 788 -257
rect 969 -260 998 -257
rect 1179 -260 1208 -257
rect 1389 -260 1418 -257
rect 1599 -260 1628 -257
rect 1809 -260 1838 -257
rect 2019 -260 2048 -257
rect 2229 -260 2258 -257
rect 2439 -260 2468 -257
rect 2649 -260 2678 -257
rect 2859 -260 2888 -257
rect 3069 -260 3098 -257
rect 3279 -260 3308 -257
rect 3489 -260 3518 -257
rect 3699 -260 3728 -257
rect 3909 -260 3938 -257
rect 4119 -260 4148 -257
rect 129 -277 135 -260
rect 339 -277 345 -260
rect 549 -277 555 -260
rect 759 -277 765 -260
rect 969 -277 975 -260
rect 1179 -277 1185 -260
rect 1389 -277 1395 -260
rect 1599 -277 1605 -260
rect 1809 -277 1815 -260
rect 2019 -277 2025 -260
rect 2229 -277 2235 -260
rect 2439 -277 2445 -260
rect 2649 -277 2655 -260
rect 2859 -277 2865 -260
rect 3069 -277 3075 -260
rect 3279 -277 3285 -260
rect 3489 -277 3495 -260
rect 3699 -277 3705 -260
rect 3909 -277 3915 -260
rect 4119 -277 4125 -260
rect 129 -280 158 -277
rect 339 -280 368 -277
rect 549 -280 578 -277
rect 759 -280 788 -277
rect 969 -280 998 -277
rect 1179 -280 1208 -277
rect 1389 -280 1418 -277
rect 1599 -280 1628 -277
rect 1809 -280 1838 -277
rect 2019 -280 2048 -277
rect 2229 -280 2258 -277
rect 2439 -280 2468 -277
rect 2649 -280 2678 -277
rect 2859 -280 2888 -277
rect 3069 -280 3098 -277
rect 3279 -280 3308 -277
rect 3489 -280 3518 -277
rect 3699 -280 3728 -277
rect 3909 -280 3938 -277
rect 4119 -280 4148 -277
rect 234 -415 263 -412
rect 444 -415 473 -412
rect 654 -415 683 -412
rect 864 -415 893 -412
rect 1074 -415 1103 -412
rect 1284 -415 1313 -412
rect 1494 -415 1523 -412
rect 1704 -415 1733 -412
rect 1914 -415 1943 -412
rect 2124 -415 2153 -412
rect 2334 -415 2363 -412
rect 2544 -415 2573 -412
rect 2754 -415 2783 -412
rect 2964 -415 2993 -412
rect 3174 -415 3203 -412
rect 3384 -415 3413 -412
rect 3594 -415 3623 -412
rect 3804 -415 3833 -412
rect 4014 -415 4043 -412
rect 4224 -415 4253 -412
rect 234 -432 240 -415
rect 444 -432 450 -415
rect 654 -432 660 -415
rect 864 -432 870 -415
rect 1074 -432 1080 -415
rect 1284 -432 1290 -415
rect 1494 -432 1500 -415
rect 1704 -432 1710 -415
rect 1914 -432 1920 -415
rect 2124 -432 2130 -415
rect 2334 -432 2340 -415
rect 2544 -432 2550 -415
rect 2754 -432 2760 -415
rect 2964 -432 2970 -415
rect 3174 -432 3180 -415
rect 3384 -432 3390 -415
rect 3594 -432 3600 -415
rect 3804 -432 3810 -415
rect 4014 -432 4020 -415
rect 4224 -432 4230 -415
rect 234 -435 263 -432
rect 444 -435 473 -432
rect 654 -435 683 -432
rect 864 -435 893 -432
rect 1074 -435 1103 -432
rect 1284 -435 1313 -432
rect 1494 -435 1523 -432
rect 1704 -435 1733 -432
rect 1914 -435 1943 -432
rect 2124 -435 2153 -432
rect 2334 -435 2363 -432
rect 2544 -435 2573 -432
rect 2754 -435 2783 -432
rect 2964 -435 2993 -432
rect 3174 -435 3203 -432
rect 3384 -435 3413 -432
rect 3594 -435 3623 -432
rect 3804 -435 3833 -432
rect 4014 -435 4043 -432
rect 4224 -435 4253 -432
rect 129 -480 158 -477
rect 339 -480 368 -477
rect 549 -480 578 -477
rect 759 -480 788 -477
rect 969 -480 998 -477
rect 1179 -480 1208 -477
rect 1389 -480 1418 -477
rect 1599 -480 1628 -477
rect 1809 -480 1838 -477
rect 2019 -480 2048 -477
rect 2229 -480 2258 -477
rect 2439 -480 2468 -477
rect 2649 -480 2678 -477
rect 2859 -480 2888 -477
rect 3069 -480 3098 -477
rect 3279 -480 3308 -477
rect 3489 -480 3518 -477
rect 3699 -480 3728 -477
rect 3909 -480 3938 -477
rect 4119 -480 4148 -477
rect 129 -497 135 -480
rect 339 -497 345 -480
rect 549 -497 555 -480
rect 759 -497 765 -480
rect 969 -497 975 -480
rect 1179 -497 1185 -480
rect 1389 -497 1395 -480
rect 1599 -497 1605 -480
rect 1809 -497 1815 -480
rect 2019 -497 2025 -480
rect 2229 -497 2235 -480
rect 2439 -497 2445 -480
rect 2649 -497 2655 -480
rect 2859 -497 2865 -480
rect 3069 -497 3075 -480
rect 3279 -497 3285 -480
rect 3489 -497 3495 -480
rect 3699 -497 3705 -480
rect 3909 -497 3915 -480
rect 4119 -497 4125 -480
rect 129 -500 158 -497
rect 339 -500 368 -497
rect 549 -500 578 -497
rect 759 -500 788 -497
rect 969 -500 998 -497
rect 1179 -500 1208 -497
rect 1389 -500 1418 -497
rect 1599 -500 1628 -497
rect 1809 -500 1838 -497
rect 2019 -500 2048 -497
rect 2229 -500 2258 -497
rect 2439 -500 2468 -497
rect 2649 -500 2678 -497
rect 2859 -500 2888 -497
rect 3069 -500 3098 -497
rect 3279 -500 3308 -497
rect 3489 -500 3518 -497
rect 3699 -500 3728 -497
rect 3909 -500 3938 -497
rect 4119 -500 4148 -497
rect 234 -635 263 -632
rect 444 -635 473 -632
rect 654 -635 683 -632
rect 864 -635 893 -632
rect 1074 -635 1103 -632
rect 1284 -635 1313 -632
rect 1494 -635 1523 -632
rect 1704 -635 1733 -632
rect 1914 -635 1943 -632
rect 2124 -635 2153 -632
rect 2334 -635 2363 -632
rect 2544 -635 2573 -632
rect 2754 -635 2783 -632
rect 2964 -635 2993 -632
rect 3174 -635 3203 -632
rect 3384 -635 3413 -632
rect 3594 -635 3623 -632
rect 3804 -635 3833 -632
rect 4014 -635 4043 -632
rect 4224 -635 4253 -632
rect 234 -652 240 -635
rect 444 -652 450 -635
rect 654 -652 660 -635
rect 864 -652 870 -635
rect 1074 -652 1080 -635
rect 1284 -652 1290 -635
rect 1494 -652 1500 -635
rect 1704 -652 1710 -635
rect 1914 -652 1920 -635
rect 2124 -652 2130 -635
rect 2334 -652 2340 -635
rect 2544 -652 2550 -635
rect 2754 -652 2760 -635
rect 2964 -652 2970 -635
rect 3174 -652 3180 -635
rect 3384 -652 3390 -635
rect 3594 -652 3600 -635
rect 3804 -652 3810 -635
rect 4014 -652 4020 -635
rect 4224 -652 4230 -635
rect 234 -655 263 -652
rect 444 -655 473 -652
rect 654 -655 683 -652
rect 864 -655 893 -652
rect 1074 -655 1103 -652
rect 1284 -655 1313 -652
rect 1494 -655 1523 -652
rect 1704 -655 1733 -652
rect 1914 -655 1943 -652
rect 2124 -655 2153 -652
rect 2334 -655 2363 -652
rect 2544 -655 2573 -652
rect 2754 -655 2783 -652
rect 2964 -655 2993 -652
rect 3174 -655 3203 -652
rect 3384 -655 3413 -652
rect 3594 -655 3623 -652
rect 3804 -655 3833 -652
rect 4014 -655 4043 -652
rect 4224 -655 4253 -652
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_0
timestamp 1654601900
transform 1 0 2191 0 1 94
box -2191 -94 2191 94
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_1
timestamp 1654601900
transform 1 0 2191 0 1 -126
box -2191 -94 2191 94
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_2
timestamp 1654601900
transform 1 0 2191 0 1 -346
box -2191 -94 2191 94
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_3
timestamp 1654601900
transform 1 0 2191 0 1 -566
box -2191 -94 2191 94
<< end >>
