magic
tech sky130A
timestamp 1653472245
<< nmos >>
rect -468 -70 -408 70
rect -322 -70 -262 70
rect -176 -70 -116 70
rect -30 -70 30 70
rect 116 -70 176 70
rect 262 -70 322 70
rect 408 -70 468 70
<< ndiff >>
rect -497 64 -468 70
rect -497 -64 -491 64
rect -474 -64 -468 64
rect -497 -70 -468 -64
rect -408 64 -379 70
rect -408 -64 -402 64
rect -385 -64 -379 64
rect -408 -70 -379 -64
rect -351 64 -322 70
rect -351 -64 -345 64
rect -328 -64 -322 64
rect -351 -70 -322 -64
rect -262 64 -233 70
rect -262 -64 -256 64
rect -239 -64 -233 64
rect -262 -70 -233 -64
rect -205 64 -176 70
rect -205 -64 -199 64
rect -182 -64 -176 64
rect -205 -70 -176 -64
rect -116 64 -87 70
rect -116 -64 -110 64
rect -93 -64 -87 64
rect -116 -70 -87 -64
rect -59 64 -30 70
rect -59 -64 -53 64
rect -36 -64 -30 64
rect -59 -70 -30 -64
rect 30 64 59 70
rect 30 -64 36 64
rect 53 -64 59 64
rect 30 -70 59 -64
rect 87 64 116 70
rect 87 -64 93 64
rect 110 -64 116 64
rect 87 -70 116 -64
rect 176 64 205 70
rect 176 -64 182 64
rect 199 -64 205 64
rect 176 -70 205 -64
rect 233 64 262 70
rect 233 -64 239 64
rect 256 -64 262 64
rect 233 -70 262 -64
rect 322 64 351 70
rect 322 -64 328 64
rect 345 -64 351 64
rect 322 -70 351 -64
rect 379 64 408 70
rect 379 -64 385 64
rect 402 -64 408 64
rect 379 -70 408 -64
rect 468 64 497 70
rect 468 -64 474 64
rect 491 -64 497 64
rect 468 -70 497 -64
<< ndiffc >>
rect -491 -64 -474 64
rect -402 -64 -385 64
rect -345 -64 -328 64
rect -256 -64 -239 64
rect -199 -64 -182 64
rect -110 -64 -93 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 93 -64 110 64
rect 182 -64 199 64
rect 239 -64 256 64
rect 328 -64 345 64
rect 385 -64 402 64
rect 474 -64 491 64
<< poly >>
rect -457 106 -419 114
rect -457 97 -449 106
rect -468 89 -449 97
rect -427 97 -419 106
rect -311 106 -273 114
rect -311 97 -303 106
rect -427 89 -408 97
rect -468 70 -408 89
rect -322 89 -303 97
rect -281 97 -273 106
rect -165 106 -127 114
rect -165 97 -157 106
rect -281 89 -262 97
rect -322 70 -262 89
rect -176 89 -157 97
rect -135 97 -127 106
rect -19 106 19 114
rect -19 97 -11 106
rect -135 89 -116 97
rect -176 70 -116 89
rect -30 89 -11 97
rect 11 97 19 106
rect 127 106 165 114
rect 127 97 135 106
rect 11 89 30 97
rect -30 70 30 89
rect 116 89 135 97
rect 157 97 165 106
rect 273 106 311 114
rect 273 97 281 106
rect 157 89 176 97
rect 116 70 176 89
rect 262 89 281 97
rect 303 97 311 106
rect 419 106 457 114
rect 419 97 427 106
rect 303 89 322 97
rect 262 70 322 89
rect 408 89 427 97
rect 449 97 457 106
rect 449 89 468 97
rect 408 70 468 89
rect -468 -89 -408 -70
rect -468 -97 -449 -89
rect -457 -106 -449 -97
rect -427 -97 -408 -89
rect -322 -89 -262 -70
rect -322 -97 -303 -89
rect -427 -106 -419 -97
rect -457 -114 -419 -106
rect -311 -106 -303 -97
rect -281 -97 -262 -89
rect -176 -89 -116 -70
rect -176 -97 -157 -89
rect -281 -106 -273 -97
rect -311 -114 -273 -106
rect -165 -106 -157 -97
rect -135 -97 -116 -89
rect -30 -89 30 -70
rect -30 -97 -11 -89
rect -135 -106 -127 -97
rect -165 -114 -127 -106
rect -19 -106 -11 -97
rect 11 -97 30 -89
rect 116 -89 176 -70
rect 116 -97 135 -89
rect 11 -106 19 -97
rect -19 -114 19 -106
rect 127 -106 135 -97
rect 157 -97 176 -89
rect 262 -89 322 -70
rect 262 -97 281 -89
rect 157 -106 165 -97
rect 127 -114 165 -106
rect 273 -106 281 -97
rect 303 -97 322 -89
rect 408 -89 468 -70
rect 408 -97 427 -89
rect 303 -106 311 -97
rect 273 -114 311 -106
rect 419 -106 427 -97
rect 449 -97 468 -89
rect 449 -106 457 -97
rect 419 -114 457 -106
<< polycont >>
rect -449 89 -427 106
rect -303 89 -281 106
rect -157 89 -135 106
rect -11 89 11 106
rect 135 89 157 106
rect 281 89 303 106
rect 427 89 449 106
rect -449 -106 -427 -89
rect -303 -106 -281 -89
rect -157 -106 -135 -89
rect -11 -106 11 -89
rect 135 -106 157 -89
rect 281 -106 303 -89
rect 427 -106 449 -89
<< locali >>
rect -457 89 -449 106
rect -427 89 -419 106
rect -311 89 -303 106
rect -281 89 -273 106
rect -165 89 -157 106
rect -135 89 -127 106
rect -19 89 -11 106
rect 11 89 19 106
rect 127 89 135 106
rect 157 89 165 106
rect 273 89 281 106
rect 303 89 311 106
rect 419 89 427 106
rect 449 89 457 106
rect -491 64 -474 72
rect -491 -72 -474 -64
rect -402 64 -385 72
rect -402 -72 -385 -64
rect -345 64 -328 72
rect -345 -72 -328 -64
rect -256 64 -239 72
rect -256 -72 -239 -64
rect -199 64 -182 72
rect -199 -72 -182 -64
rect -110 64 -93 72
rect -110 -72 -93 -64
rect -53 64 -36 72
rect -53 -72 -36 -64
rect 36 64 53 72
rect 36 -72 53 -64
rect 93 64 110 72
rect 93 -72 110 -64
rect 182 64 199 72
rect 182 -72 199 -64
rect 239 64 256 72
rect 239 -72 256 -64
rect 328 64 345 72
rect 328 -72 345 -64
rect 385 64 402 72
rect 385 -72 402 -64
rect 474 64 491 72
rect 474 -72 491 -64
rect -457 -106 -449 -89
rect -427 -106 -419 -89
rect -311 -106 -303 -89
rect -281 -106 -273 -89
rect -165 -106 -157 -89
rect -135 -106 -127 -89
rect -19 -106 -11 -89
rect 11 -106 19 -89
rect 127 -106 135 -89
rect 157 -106 165 -89
rect 273 -106 281 -89
rect 303 -106 311 -89
rect 419 -106 427 -89
rect 449 -106 457 -89
<< viali >>
rect -449 89 -427 106
rect -303 89 -281 106
rect -157 89 -135 106
rect -11 89 11 106
rect 135 89 157 106
rect 281 89 303 106
rect 427 89 449 106
rect -491 -64 -474 64
rect -402 -64 -385 64
rect -345 -64 -328 64
rect -256 -64 -239 64
rect -199 -64 -182 64
rect -110 -64 -93 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 93 -64 110 64
rect 182 -64 199 64
rect 239 -64 256 64
rect 328 -64 345 64
rect 385 -64 402 64
rect 474 -64 491 64
rect -449 -106 -427 -89
rect -303 -106 -281 -89
rect -157 -106 -135 -89
rect -11 -106 11 -89
rect 135 -106 157 -89
rect 281 -106 303 -89
rect 427 -106 449 -89
<< metal1 >>
rect -457 106 -419 114
rect -457 89 -449 106
rect -427 89 -419 106
rect -457 86 -419 89
rect -311 106 -273 114
rect -311 89 -303 106
rect -281 89 -273 106
rect -311 86 -273 89
rect -165 106 -127 114
rect -165 89 -157 106
rect -135 89 -127 106
rect -165 86 -127 89
rect -19 106 19 114
rect -19 89 -11 106
rect 11 89 19 106
rect -19 86 19 89
rect 127 106 165 114
rect 127 89 135 106
rect 157 89 165 106
rect 127 86 165 89
rect 273 106 311 114
rect 273 89 281 106
rect 303 89 311 106
rect 273 86 311 89
rect 419 106 457 114
rect 419 89 427 106
rect 449 89 457 106
rect 419 86 457 89
rect -494 64 -471 70
rect -494 -64 -491 64
rect -474 -64 -471 64
rect -494 -70 -471 -64
rect -405 64 -382 70
rect -405 -64 -402 64
rect -385 -64 -382 64
rect -405 -70 -382 -64
rect -348 64 -325 70
rect -348 -64 -345 64
rect -328 -64 -325 64
rect -348 -70 -325 -64
rect -259 64 -236 70
rect -259 -64 -256 64
rect -239 -64 -236 64
rect -259 -70 -236 -64
rect -202 64 -179 70
rect -202 -64 -199 64
rect -182 -64 -179 64
rect -202 -70 -179 -64
rect -113 64 -90 70
rect -113 -64 -110 64
rect -93 -64 -90 64
rect -113 -70 -90 -64
rect -56 64 -33 70
rect -56 -64 -53 64
rect -36 -64 -33 64
rect -56 -70 -33 -64
rect 33 64 56 70
rect 33 -64 36 64
rect 53 -64 56 64
rect 33 -70 56 -64
rect 90 64 113 70
rect 90 -64 93 64
rect 110 -64 113 64
rect 90 -70 113 -64
rect 179 64 202 70
rect 179 -64 182 64
rect 199 -64 202 64
rect 179 -70 202 -64
rect 236 64 259 70
rect 236 -64 239 64
rect 256 -64 259 64
rect 236 -70 259 -64
rect 325 64 348 70
rect 325 -64 328 64
rect 345 -64 348 64
rect 325 -70 348 -64
rect 382 64 405 70
rect 382 -64 385 64
rect 402 -64 405 64
rect 382 -70 405 -64
rect 471 64 494 70
rect 471 -64 474 64
rect 491 -64 494 64
rect 471 -70 494 -64
rect -457 -89 -419 -86
rect -457 -106 -449 -89
rect -427 -106 -419 -89
rect -457 -114 -419 -106
rect -311 -89 -273 -86
rect -311 -106 -303 -89
rect -281 -106 -273 -89
rect -311 -114 -273 -106
rect -165 -89 -127 -86
rect -165 -106 -157 -89
rect -135 -106 -127 -89
rect -165 -114 -127 -106
rect -19 -89 19 -86
rect -19 -106 -11 -89
rect 11 -106 19 -89
rect -19 -114 19 -106
rect 127 -89 165 -86
rect 127 -106 135 -89
rect 157 -106 165 -89
rect 127 -114 165 -106
rect 273 -89 311 -86
rect 273 -106 281 -89
rect 303 -106 311 -89
rect 273 -114 311 -106
rect 419 -89 457 -86
rect 419 -106 427 -89
rect 449 -106 457 -89
rect 419 -114 457 -106
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 7 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
