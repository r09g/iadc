magic
tech sky130A
timestamp 1654720150
<< error_p >>
rect -765 286 -736 289
rect -686 286 -657 289
rect -607 286 -578 289
rect -528 286 -499 289
rect -449 286 -420 289
rect -370 286 -341 289
rect -291 286 -262 289
rect -212 286 -183 289
rect -133 286 -104 289
rect -54 286 -25 289
rect 25 286 54 289
rect 104 286 133 289
rect 183 286 212 289
rect 262 286 291 289
rect 341 286 370 289
rect 420 286 449 289
rect 499 286 528 289
rect 578 286 607 289
rect 657 286 686 289
rect 736 286 765 289
rect -765 269 -759 286
rect -686 269 -680 286
rect -607 269 -601 286
rect -528 269 -522 286
rect -449 269 -443 286
rect -370 269 -364 286
rect -291 269 -285 286
rect -212 269 -206 286
rect -133 269 -127 286
rect -54 269 -48 286
rect 25 269 31 286
rect 104 269 110 286
rect 183 269 189 286
rect 262 269 268 286
rect 341 269 347 286
rect 420 269 426 286
rect 499 269 505 286
rect 578 269 584 286
rect 657 269 663 286
rect 736 269 742 286
rect -765 266 -736 269
rect -686 266 -657 269
rect -607 266 -578 269
rect -528 266 -499 269
rect -449 266 -420 269
rect -370 266 -341 269
rect -291 266 -262 269
rect -212 266 -183 269
rect -133 266 -104 269
rect -54 266 -25 269
rect 25 266 54 269
rect 104 266 133 269
rect 183 266 212 269
rect 262 266 291 269
rect 341 266 370 269
rect 420 266 449 269
rect 499 266 528 269
rect 578 266 607 269
rect 657 266 686 269
rect 736 266 765 269
rect -765 -269 -736 -266
rect -686 -269 -657 -266
rect -607 -269 -578 -266
rect -528 -269 -499 -266
rect -449 -269 -420 -266
rect -370 -269 -341 -266
rect -291 -269 -262 -266
rect -212 -269 -183 -266
rect -133 -269 -104 -266
rect -54 -269 -25 -266
rect 25 -269 54 -266
rect 104 -269 133 -266
rect 183 -269 212 -266
rect 262 -269 291 -266
rect 341 -269 370 -266
rect 420 -269 449 -266
rect 499 -269 528 -266
rect 578 -269 607 -266
rect 657 -269 686 -266
rect 736 -269 765 -266
rect -765 -286 -759 -269
rect -686 -286 -680 -269
rect -607 -286 -601 -269
rect -528 -286 -522 -269
rect -449 -286 -443 -269
rect -370 -286 -364 -269
rect -291 -286 -285 -269
rect -212 -286 -206 -269
rect -133 -286 -127 -269
rect -54 -286 -48 -269
rect 25 -286 31 -269
rect 104 -286 110 -269
rect 183 -286 189 -269
rect 262 -286 268 -269
rect 341 -286 347 -269
rect 420 -286 426 -269
rect 499 -286 505 -269
rect 578 -286 584 -269
rect 657 -286 663 -269
rect 736 -286 742 -269
rect -765 -289 -736 -286
rect -686 -289 -657 -286
rect -607 -289 -578 -286
rect -528 -289 -499 -286
rect -449 -289 -420 -286
rect -370 -289 -341 -286
rect -291 -289 -262 -286
rect -212 -289 -183 -286
rect -133 -289 -104 -286
rect -54 -289 -25 -286
rect 25 -289 54 -286
rect 104 -289 133 -286
rect 183 -289 212 -286
rect 262 -289 291 -286
rect 341 -289 370 -286
rect 420 -289 449 -286
rect 499 -289 528 -286
rect 578 -289 607 -286
rect 657 -289 686 -286
rect 736 -289 765 -286
<< pwell >>
rect -889 -379 889 379
<< mvnmos >>
rect -775 -250 -725 250
rect -696 -250 -646 250
rect -617 -250 -567 250
rect -538 -250 -488 250
rect -459 -250 -409 250
rect -380 -250 -330 250
rect -301 -250 -251 250
rect -222 -250 -172 250
rect -143 -250 -93 250
rect -64 -250 -14 250
rect 14 -250 64 250
rect 93 -250 143 250
rect 172 -250 222 250
rect 251 -250 301 250
rect 330 -250 380 250
rect 409 -250 459 250
rect 488 -250 538 250
rect 567 -250 617 250
rect 646 -250 696 250
rect 725 -250 775 250
<< mvndiff >>
rect -804 244 -775 250
rect -804 -244 -798 244
rect -781 -244 -775 244
rect -804 -250 -775 -244
rect -725 244 -696 250
rect -725 -244 -719 244
rect -702 -244 -696 244
rect -725 -250 -696 -244
rect -646 244 -617 250
rect -646 -244 -640 244
rect -623 -244 -617 244
rect -646 -250 -617 -244
rect -567 244 -538 250
rect -567 -244 -561 244
rect -544 -244 -538 244
rect -567 -250 -538 -244
rect -488 244 -459 250
rect -488 -244 -482 244
rect -465 -244 -459 244
rect -488 -250 -459 -244
rect -409 244 -380 250
rect -409 -244 -403 244
rect -386 -244 -380 244
rect -409 -250 -380 -244
rect -330 244 -301 250
rect -330 -244 -324 244
rect -307 -244 -301 244
rect -330 -250 -301 -244
rect -251 244 -222 250
rect -251 -244 -245 244
rect -228 -244 -222 244
rect -251 -250 -222 -244
rect -172 244 -143 250
rect -172 -244 -166 244
rect -149 -244 -143 244
rect -172 -250 -143 -244
rect -93 244 -64 250
rect -93 -244 -87 244
rect -70 -244 -64 244
rect -93 -250 -64 -244
rect -14 244 14 250
rect -14 -244 -8 244
rect 8 -244 14 244
rect -14 -250 14 -244
rect 64 244 93 250
rect 64 -244 70 244
rect 87 -244 93 244
rect 64 -250 93 -244
rect 143 244 172 250
rect 143 -244 149 244
rect 166 -244 172 244
rect 143 -250 172 -244
rect 222 244 251 250
rect 222 -244 228 244
rect 245 -244 251 244
rect 222 -250 251 -244
rect 301 244 330 250
rect 301 -244 307 244
rect 324 -244 330 244
rect 301 -250 330 -244
rect 380 244 409 250
rect 380 -244 386 244
rect 403 -244 409 244
rect 380 -250 409 -244
rect 459 244 488 250
rect 459 -244 465 244
rect 482 -244 488 244
rect 459 -250 488 -244
rect 538 244 567 250
rect 538 -244 544 244
rect 561 -244 567 244
rect 538 -250 567 -244
rect 617 244 646 250
rect 617 -244 623 244
rect 640 -244 646 244
rect 617 -250 646 -244
rect 696 244 725 250
rect 696 -244 702 244
rect 719 -244 725 244
rect 696 -250 725 -244
rect 775 244 804 250
rect 775 -244 781 244
rect 798 -244 804 244
rect 775 -250 804 -244
<< mvndiffc >>
rect -798 -244 -781 244
rect -719 -244 -702 244
rect -640 -244 -623 244
rect -561 -244 -544 244
rect -482 -244 -465 244
rect -403 -244 -386 244
rect -324 -244 -307 244
rect -245 -244 -228 244
rect -166 -244 -149 244
rect -87 -244 -70 244
rect -8 -244 8 244
rect 70 -244 87 244
rect 149 -244 166 244
rect 228 -244 245 244
rect 307 -244 324 244
rect 386 -244 403 244
rect 465 -244 482 244
rect 544 -244 561 244
rect 623 -244 640 244
rect 702 -244 719 244
rect 781 -244 798 244
<< mvpsubdiff >>
rect -871 355 871 361
rect -871 338 -817 355
rect 817 338 871 355
rect -871 332 871 338
rect -871 307 -842 332
rect -871 -307 -865 307
rect -848 -307 -842 307
rect 842 307 871 332
rect -871 -332 -842 -307
rect 842 -307 848 307
rect 865 -307 871 307
rect 842 -332 871 -307
rect -871 -338 871 -332
rect -871 -355 -817 -338
rect 817 -355 871 -338
rect -871 -361 871 -355
<< mvpsubdiffcont >>
rect -817 338 817 355
rect -865 -307 -848 307
rect 848 -307 865 307
rect -817 -355 817 -338
<< poly >>
rect -775 286 -725 294
rect -775 269 -767 286
rect -733 269 -725 286
rect -775 250 -725 269
rect -696 286 -646 294
rect -696 269 -688 286
rect -654 269 -646 286
rect -696 250 -646 269
rect -617 286 -567 294
rect -617 269 -609 286
rect -575 269 -567 286
rect -617 250 -567 269
rect -538 286 -488 294
rect -538 269 -530 286
rect -496 269 -488 286
rect -538 250 -488 269
rect -459 286 -409 294
rect -459 269 -451 286
rect -417 269 -409 286
rect -459 250 -409 269
rect -380 286 -330 294
rect -380 269 -372 286
rect -338 269 -330 286
rect -380 250 -330 269
rect -301 286 -251 294
rect -301 269 -293 286
rect -259 269 -251 286
rect -301 250 -251 269
rect -222 286 -172 294
rect -222 269 -214 286
rect -180 269 -172 286
rect -222 250 -172 269
rect -143 286 -93 294
rect -143 269 -135 286
rect -101 269 -93 286
rect -143 250 -93 269
rect -64 286 -14 294
rect -64 269 -56 286
rect -22 269 -14 286
rect -64 250 -14 269
rect 14 286 64 294
rect 14 269 22 286
rect 56 269 64 286
rect 14 250 64 269
rect 93 286 143 294
rect 93 269 101 286
rect 135 269 143 286
rect 93 250 143 269
rect 172 286 222 294
rect 172 269 180 286
rect 214 269 222 286
rect 172 250 222 269
rect 251 286 301 294
rect 251 269 259 286
rect 293 269 301 286
rect 251 250 301 269
rect 330 286 380 294
rect 330 269 338 286
rect 372 269 380 286
rect 330 250 380 269
rect 409 286 459 294
rect 409 269 417 286
rect 451 269 459 286
rect 409 250 459 269
rect 488 286 538 294
rect 488 269 496 286
rect 530 269 538 286
rect 488 250 538 269
rect 567 286 617 294
rect 567 269 575 286
rect 609 269 617 286
rect 567 250 617 269
rect 646 286 696 294
rect 646 269 654 286
rect 688 269 696 286
rect 646 250 696 269
rect 725 286 775 294
rect 725 269 733 286
rect 767 269 775 286
rect 725 250 775 269
rect -775 -269 -725 -250
rect -775 -286 -767 -269
rect -733 -286 -725 -269
rect -775 -294 -725 -286
rect -696 -269 -646 -250
rect -696 -286 -688 -269
rect -654 -286 -646 -269
rect -696 -294 -646 -286
rect -617 -269 -567 -250
rect -617 -286 -609 -269
rect -575 -286 -567 -269
rect -617 -294 -567 -286
rect -538 -269 -488 -250
rect -538 -286 -530 -269
rect -496 -286 -488 -269
rect -538 -294 -488 -286
rect -459 -269 -409 -250
rect -459 -286 -451 -269
rect -417 -286 -409 -269
rect -459 -294 -409 -286
rect -380 -269 -330 -250
rect -380 -286 -372 -269
rect -338 -286 -330 -269
rect -380 -294 -330 -286
rect -301 -269 -251 -250
rect -301 -286 -293 -269
rect -259 -286 -251 -269
rect -301 -294 -251 -286
rect -222 -269 -172 -250
rect -222 -286 -214 -269
rect -180 -286 -172 -269
rect -222 -294 -172 -286
rect -143 -269 -93 -250
rect -143 -286 -135 -269
rect -101 -286 -93 -269
rect -143 -294 -93 -286
rect -64 -269 -14 -250
rect -64 -286 -56 -269
rect -22 -286 -14 -269
rect -64 -294 -14 -286
rect 14 -269 64 -250
rect 14 -286 22 -269
rect 56 -286 64 -269
rect 14 -294 64 -286
rect 93 -269 143 -250
rect 93 -286 101 -269
rect 135 -286 143 -269
rect 93 -294 143 -286
rect 172 -269 222 -250
rect 172 -286 180 -269
rect 214 -286 222 -269
rect 172 -294 222 -286
rect 251 -269 301 -250
rect 251 -286 259 -269
rect 293 -286 301 -269
rect 251 -294 301 -286
rect 330 -269 380 -250
rect 330 -286 338 -269
rect 372 -286 380 -269
rect 330 -294 380 -286
rect 409 -269 459 -250
rect 409 -286 417 -269
rect 451 -286 459 -269
rect 409 -294 459 -286
rect 488 -269 538 -250
rect 488 -286 496 -269
rect 530 -286 538 -269
rect 488 -294 538 -286
rect 567 -269 617 -250
rect 567 -286 575 -269
rect 609 -286 617 -269
rect 567 -294 617 -286
rect 646 -269 696 -250
rect 646 -286 654 -269
rect 688 -286 696 -269
rect 646 -294 696 -286
rect 725 -269 775 -250
rect 725 -286 733 -269
rect 767 -286 775 -269
rect 725 -294 775 -286
<< polycont >>
rect -767 269 -733 286
rect -688 269 -654 286
rect -609 269 -575 286
rect -530 269 -496 286
rect -451 269 -417 286
rect -372 269 -338 286
rect -293 269 -259 286
rect -214 269 -180 286
rect -135 269 -101 286
rect -56 269 -22 286
rect 22 269 56 286
rect 101 269 135 286
rect 180 269 214 286
rect 259 269 293 286
rect 338 269 372 286
rect 417 269 451 286
rect 496 269 530 286
rect 575 269 609 286
rect 654 269 688 286
rect 733 269 767 286
rect -767 -286 -733 -269
rect -688 -286 -654 -269
rect -609 -286 -575 -269
rect -530 -286 -496 -269
rect -451 -286 -417 -269
rect -372 -286 -338 -269
rect -293 -286 -259 -269
rect -214 -286 -180 -269
rect -135 -286 -101 -269
rect -56 -286 -22 -269
rect 22 -286 56 -269
rect 101 -286 135 -269
rect 180 -286 214 -269
rect 259 -286 293 -269
rect 338 -286 372 -269
rect 417 -286 451 -269
rect 496 -286 530 -269
rect 575 -286 609 -269
rect 654 -286 688 -269
rect 733 -286 767 -269
<< locali >>
rect -865 338 -817 355
rect 817 338 865 355
rect -865 307 -848 338
rect 848 307 865 338
rect -775 269 -767 286
rect -733 269 -725 286
rect -696 269 -688 286
rect -654 269 -646 286
rect -617 269 -609 286
rect -575 269 -567 286
rect -538 269 -530 286
rect -496 269 -488 286
rect -459 269 -451 286
rect -417 269 -409 286
rect -380 269 -372 286
rect -338 269 -330 286
rect -301 269 -293 286
rect -259 269 -251 286
rect -222 269 -214 286
rect -180 269 -172 286
rect -143 269 -135 286
rect -101 269 -93 286
rect -64 269 -56 286
rect -22 269 -14 286
rect 14 269 22 286
rect 56 269 64 286
rect 93 269 101 286
rect 135 269 143 286
rect 172 269 180 286
rect 214 269 222 286
rect 251 269 259 286
rect 293 269 301 286
rect 330 269 338 286
rect 372 269 380 286
rect 409 269 417 286
rect 451 269 459 286
rect 488 269 496 286
rect 530 269 538 286
rect 567 269 575 286
rect 609 269 617 286
rect 646 269 654 286
rect 688 269 696 286
rect 725 269 733 286
rect 767 269 775 286
rect -798 244 -781 252
rect -798 -252 -781 -244
rect -719 244 -702 252
rect -719 -252 -702 -244
rect -640 244 -623 252
rect -640 -252 -623 -244
rect -561 244 -544 252
rect -561 -252 -544 -244
rect -482 244 -465 252
rect -482 -252 -465 -244
rect -403 244 -386 252
rect -403 -252 -386 -244
rect -324 244 -307 252
rect -324 -252 -307 -244
rect -245 244 -228 252
rect -245 -252 -228 -244
rect -166 244 -149 252
rect -166 -252 -149 -244
rect -87 244 -70 252
rect -87 -252 -70 -244
rect -8 244 8 252
rect -8 -252 8 -244
rect 70 244 87 252
rect 70 -252 87 -244
rect 149 244 166 252
rect 149 -252 166 -244
rect 228 244 245 252
rect 228 -252 245 -244
rect 307 244 324 252
rect 307 -252 324 -244
rect 386 244 403 252
rect 386 -252 403 -244
rect 465 244 482 252
rect 465 -252 482 -244
rect 544 244 561 252
rect 544 -252 561 -244
rect 623 244 640 252
rect 623 -252 640 -244
rect 702 244 719 252
rect 702 -252 719 -244
rect 781 244 798 252
rect 781 -252 798 -244
rect -775 -286 -767 -269
rect -733 -286 -725 -269
rect -696 -286 -688 -269
rect -654 -286 -646 -269
rect -617 -286 -609 -269
rect -575 -286 -567 -269
rect -538 -286 -530 -269
rect -496 -286 -488 -269
rect -459 -286 -451 -269
rect -417 -286 -409 -269
rect -380 -286 -372 -269
rect -338 -286 -330 -269
rect -301 -286 -293 -269
rect -259 -286 -251 -269
rect -222 -286 -214 -269
rect -180 -286 -172 -269
rect -143 -286 -135 -269
rect -101 -286 -93 -269
rect -64 -286 -56 -269
rect -22 -286 -14 -269
rect 14 -286 22 -269
rect 56 -286 64 -269
rect 93 -286 101 -269
rect 135 -286 143 -269
rect 172 -286 180 -269
rect 214 -286 222 -269
rect 251 -286 259 -269
rect 293 -286 301 -269
rect 330 -286 338 -269
rect 372 -286 380 -269
rect 409 -286 417 -269
rect 451 -286 459 -269
rect 488 -286 496 -269
rect 530 -286 538 -269
rect 567 -286 575 -269
rect 609 -286 617 -269
rect 646 -286 654 -269
rect 688 -286 696 -269
rect 725 -286 733 -269
rect 767 -286 775 -269
rect -865 -338 -848 -307
rect 848 -338 865 -307
rect -865 -355 -817 -338
rect 817 -355 865 -338
<< viali >>
rect -759 269 -742 286
rect -680 269 -663 286
rect -601 269 -584 286
rect -522 269 -505 286
rect -443 269 -426 286
rect -364 269 -347 286
rect -285 269 -268 286
rect -206 269 -189 286
rect -127 269 -110 286
rect -48 269 -31 286
rect 31 269 48 286
rect 110 269 127 286
rect 189 269 206 286
rect 268 269 285 286
rect 347 269 364 286
rect 426 269 443 286
rect 505 269 522 286
rect 584 269 601 286
rect 663 269 680 286
rect 742 269 759 286
rect -798 -244 -781 244
rect -719 -244 -702 244
rect -640 -244 -623 244
rect -561 -244 -544 244
rect -482 -244 -465 244
rect -403 -244 -386 244
rect -324 -244 -307 244
rect -245 -244 -228 244
rect -166 -244 -149 244
rect -87 -244 -70 244
rect -8 -244 8 244
rect 70 -244 87 244
rect 149 -244 166 244
rect 228 -244 245 244
rect 307 -244 324 244
rect 386 -244 403 244
rect 465 -244 482 244
rect 544 -244 561 244
rect 623 -244 640 244
rect 702 -244 719 244
rect 781 -244 798 244
rect -759 -286 -742 -269
rect -680 -286 -663 -269
rect -601 -286 -584 -269
rect -522 -286 -505 -269
rect -443 -286 -426 -269
rect -364 -286 -347 -269
rect -285 -286 -268 -269
rect -206 -286 -189 -269
rect -127 -286 -110 -269
rect -48 -286 -31 -269
rect 31 -286 48 -269
rect 110 -286 127 -269
rect 189 -286 206 -269
rect 268 -286 285 -269
rect 347 -286 364 -269
rect 426 -286 443 -269
rect 505 -286 522 -269
rect 584 -286 601 -269
rect 663 -286 680 -269
rect 742 -286 759 -269
<< metal1 >>
rect -765 286 -736 289
rect -765 269 -759 286
rect -742 269 -736 286
rect -765 266 -736 269
rect -686 286 -657 289
rect -686 269 -680 286
rect -663 269 -657 286
rect -686 266 -657 269
rect -607 286 -578 289
rect -607 269 -601 286
rect -584 269 -578 286
rect -607 266 -578 269
rect -528 286 -499 289
rect -528 269 -522 286
rect -505 269 -499 286
rect -528 266 -499 269
rect -449 286 -420 289
rect -449 269 -443 286
rect -426 269 -420 286
rect -449 266 -420 269
rect -370 286 -341 289
rect -370 269 -364 286
rect -347 269 -341 286
rect -370 266 -341 269
rect -291 286 -262 289
rect -291 269 -285 286
rect -268 269 -262 286
rect -291 266 -262 269
rect -212 286 -183 289
rect -212 269 -206 286
rect -189 269 -183 286
rect -212 266 -183 269
rect -133 286 -104 289
rect -133 269 -127 286
rect -110 269 -104 286
rect -133 266 -104 269
rect -54 286 -25 289
rect -54 269 -48 286
rect -31 269 -25 286
rect -54 266 -25 269
rect 25 286 54 289
rect 25 269 31 286
rect 48 269 54 286
rect 25 266 54 269
rect 104 286 133 289
rect 104 269 110 286
rect 127 269 133 286
rect 104 266 133 269
rect 183 286 212 289
rect 183 269 189 286
rect 206 269 212 286
rect 183 266 212 269
rect 262 286 291 289
rect 262 269 268 286
rect 285 269 291 286
rect 262 266 291 269
rect 341 286 370 289
rect 341 269 347 286
rect 364 269 370 286
rect 341 266 370 269
rect 420 286 449 289
rect 420 269 426 286
rect 443 269 449 286
rect 420 266 449 269
rect 499 286 528 289
rect 499 269 505 286
rect 522 269 528 286
rect 499 266 528 269
rect 578 286 607 289
rect 578 269 584 286
rect 601 269 607 286
rect 578 266 607 269
rect 657 286 686 289
rect 657 269 663 286
rect 680 269 686 286
rect 657 266 686 269
rect 736 286 765 289
rect 736 269 742 286
rect 759 269 765 286
rect 736 266 765 269
rect -801 244 -778 250
rect -801 -244 -798 244
rect -781 -244 -778 244
rect -801 -250 -778 -244
rect -722 244 -699 250
rect -722 -244 -719 244
rect -702 -244 -699 244
rect -722 -250 -699 -244
rect -643 244 -620 250
rect -643 -244 -640 244
rect -623 -244 -620 244
rect -643 -250 -620 -244
rect -564 244 -541 250
rect -564 -244 -561 244
rect -544 -244 -541 244
rect -564 -250 -541 -244
rect -485 244 -462 250
rect -485 -244 -482 244
rect -465 -244 -462 244
rect -485 -250 -462 -244
rect -406 244 -383 250
rect -406 -244 -403 244
rect -386 -244 -383 244
rect -406 -250 -383 -244
rect -327 244 -304 250
rect -327 -244 -324 244
rect -307 -244 -304 244
rect -327 -250 -304 -244
rect -248 244 -225 250
rect -248 -244 -245 244
rect -228 -244 -225 244
rect -248 -250 -225 -244
rect -169 244 -146 250
rect -169 -244 -166 244
rect -149 -244 -146 244
rect -169 -250 -146 -244
rect -90 244 -67 250
rect -90 -244 -87 244
rect -70 -244 -67 244
rect -90 -250 -67 -244
rect -11 244 11 250
rect -11 -244 -8 244
rect 8 -244 11 244
rect -11 -250 11 -244
rect 67 244 90 250
rect 67 -244 70 244
rect 87 -244 90 244
rect 67 -250 90 -244
rect 146 244 169 250
rect 146 -244 149 244
rect 166 -244 169 244
rect 146 -250 169 -244
rect 225 244 248 250
rect 225 -244 228 244
rect 245 -244 248 244
rect 225 -250 248 -244
rect 304 244 327 250
rect 304 -244 307 244
rect 324 -244 327 244
rect 304 -250 327 -244
rect 383 244 406 250
rect 383 -244 386 244
rect 403 -244 406 244
rect 383 -250 406 -244
rect 462 244 485 250
rect 462 -244 465 244
rect 482 -244 485 244
rect 462 -250 485 -244
rect 541 244 564 250
rect 541 -244 544 244
rect 561 -244 564 244
rect 541 -250 564 -244
rect 620 244 643 250
rect 620 -244 623 244
rect 640 -244 643 244
rect 620 -250 643 -244
rect 699 244 722 250
rect 699 -244 702 244
rect 719 -244 722 244
rect 699 -250 722 -244
rect 778 244 801 250
rect 778 -244 781 244
rect 798 -244 801 244
rect 778 -250 801 -244
rect -765 -269 -736 -266
rect -765 -286 -759 -269
rect -742 -286 -736 -269
rect -765 -289 -736 -286
rect -686 -269 -657 -266
rect -686 -286 -680 -269
rect -663 -286 -657 -269
rect -686 -289 -657 -286
rect -607 -269 -578 -266
rect -607 -286 -601 -269
rect -584 -286 -578 -269
rect -607 -289 -578 -286
rect -528 -269 -499 -266
rect -528 -286 -522 -269
rect -505 -286 -499 -269
rect -528 -289 -499 -286
rect -449 -269 -420 -266
rect -449 -286 -443 -269
rect -426 -286 -420 -269
rect -449 -289 -420 -286
rect -370 -269 -341 -266
rect -370 -286 -364 -269
rect -347 -286 -341 -269
rect -370 -289 -341 -286
rect -291 -269 -262 -266
rect -291 -286 -285 -269
rect -268 -286 -262 -269
rect -291 -289 -262 -286
rect -212 -269 -183 -266
rect -212 -286 -206 -269
rect -189 -286 -183 -269
rect -212 -289 -183 -286
rect -133 -269 -104 -266
rect -133 -286 -127 -269
rect -110 -286 -104 -269
rect -133 -289 -104 -286
rect -54 -269 -25 -266
rect -54 -286 -48 -269
rect -31 -286 -25 -269
rect -54 -289 -25 -286
rect 25 -269 54 -266
rect 25 -286 31 -269
rect 48 -286 54 -269
rect 25 -289 54 -286
rect 104 -269 133 -266
rect 104 -286 110 -269
rect 127 -286 133 -269
rect 104 -289 133 -286
rect 183 -269 212 -266
rect 183 -286 189 -269
rect 206 -286 212 -269
rect 183 -289 212 -286
rect 262 -269 291 -266
rect 262 -286 268 -269
rect 285 -286 291 -269
rect 262 -289 291 -286
rect 341 -269 370 -266
rect 341 -286 347 -269
rect 364 -286 370 -269
rect 341 -289 370 -286
rect 420 -269 449 -266
rect 420 -286 426 -269
rect 443 -286 449 -269
rect 420 -289 449 -286
rect 499 -269 528 -266
rect 499 -286 505 -269
rect 522 -286 528 -269
rect 499 -289 528 -286
rect 578 -269 607 -266
rect 578 -286 584 -269
rect 601 -286 607 -269
rect 578 -289 607 -286
rect 657 -269 686 -266
rect 657 -286 663 -269
rect 680 -286 686 -269
rect 657 -289 686 -286
rect 736 -269 765 -266
rect 736 -286 742 -269
rect 759 -286 765 -269
rect 736 -289 765 -286
<< properties >>
string FIXED_BBOX -857 -346 857 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
