magic
tech sky130A
magscale 1 2
timestamp 1654558272
<< nwell >>
rect -7664 -7309 3823 -1120
<< pwell >>
rect -7664 -17642 13838 -7439
<< psubdiff >>
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect -7605 -17459 -7505 -17268
rect 13619 -7731 13719 -7621
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< nsubdiff >>
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect -7605 -7140 -7512 -6976
rect 3610 -1520 3703 -1353
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
<< psubdiffcont >>
rect -7264 -7621 13443 -7521
rect -7605 -17268 -7505 -7850
rect 13619 -17149 13719 -7731
<< nsubdiffcont >>
rect -7379 -1353 3329 -1260
rect -7605 -6976 -7512 -1507
rect 3610 -6989 3703 -1520
rect -7282 -7233 3426 -7140
<< locali >>
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect -7605 -7140 -7512 -6976
rect 3610 -1520 3703 -1353
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect -7605 -17459 -7505 -17268
rect 13619 -7731 13719 -7621
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< viali >>
rect -7379 -1353 3329 -1260
rect -7323 -17559 13384 -17459
<< metal1 >>
rect 7034 2713 7080 2891
rect 16034 2713 16080 2891
rect 7034 1691 7080 1863
rect 16034 1691 16080 1863
rect 7034 913 7080 1091
rect 16034 913 16080 1091
rect 7034 -109 7080 63
rect 16034 -109 16080 63
rect 7034 -887 7080 -709
rect 16034 -887 16080 -709
rect -7605 -1260 3704 -1200
rect -7605 -1353 -7379 -1260
rect 3329 -1353 3704 -1260
rect -7605 -1467 3704 -1353
rect -5132 -1741 -4948 -1467
rect -5945 -1841 -3776 -1741
rect -5945 -2039 -5911 -1841
rect -5877 -1963 -5867 -1910
rect -5814 -1963 -5804 -1910
rect -5699 -1963 -5689 -1910
rect -5636 -1963 -5626 -1910
rect -5520 -1963 -5510 -1910
rect -5457 -1963 -5447 -1910
rect -5343 -1963 -5333 -1910
rect -5280 -1963 -5270 -1910
rect -5165 -1963 -5155 -1910
rect -5102 -1963 -5092 -1910
rect -4986 -1963 -4976 -1910
rect -4923 -1963 -4913 -1910
rect -4809 -1963 -4799 -1910
rect -4746 -1963 -4736 -1910
rect -4631 -1963 -4621 -1910
rect -4568 -1963 -4558 -1910
rect -4453 -1963 -4443 -1910
rect -4390 -1963 -4380 -1910
rect -4275 -1963 -4265 -1910
rect -4212 -1963 -4202 -1910
rect -4096 -1963 -4086 -1910
rect -4033 -1963 -4023 -1910
rect -3919 -1963 -3909 -1910
rect -3856 -1963 -3846 -1910
rect -6302 -2073 -5911 -2039
rect -6302 -2135 -6268 -2073
rect -6126 -2150 -6092 -2073
rect -5945 -2132 -5911 -2073
rect -5857 -2079 -5823 -1963
rect -5679 -2079 -5645 -1963
rect -5501 -2079 -5467 -1963
rect -5322 -2079 -5288 -1963
rect -5145 -2079 -5111 -1963
rect -4967 -2079 -4933 -1963
rect -4789 -2079 -4755 -1963
rect -4611 -2079 -4577 -1963
rect -4433 -2079 -4399 -1963
rect -4255 -2079 -4221 -1963
rect -4077 -2079 -4043 -1963
rect -3898 -2079 -3864 -1963
rect -3810 -2133 -3776 -1841
rect -1119 -1963 -1109 -1910
rect -1056 -1963 -1046 -1910
rect -6508 -2582 -6498 -2529
rect -6445 -2582 -6435 -2529
rect -6635 -3454 -6625 -3401
rect -6572 -3454 -6562 -3401
rect -6625 -5322 -6572 -3454
rect -6498 -3640 -6445 -2582
rect -6054 -2833 -6044 -2780
rect -5991 -2833 -5981 -2780
rect -6302 -2945 -6090 -2911
rect -6302 -3020 -6268 -2945
rect -6124 -3022 -6090 -2945
rect -6035 -2949 -6001 -2833
rect -6124 -3401 -6090 -3259
rect -6144 -3454 -6134 -3401
rect -6081 -3454 -6071 -3401
rect -6508 -3693 -6498 -3640
rect -6445 -3693 -6435 -3640
rect -6498 -4271 -6445 -3693
rect -6302 -3812 -6090 -3778
rect -6302 -3889 -6268 -3812
rect -6124 -3888 -6090 -3812
rect -6035 -3819 -6001 -3311
rect -6508 -4324 -6498 -4271
rect -6445 -4324 -6435 -4271
rect -6498 -5141 -6445 -4324
rect -6124 -4390 -6090 -4128
rect -6144 -4443 -6134 -4390
rect -6081 -4443 -6071 -4390
rect -6302 -4683 -6090 -4649
rect -6302 -4763 -6268 -4683
rect -6124 -4761 -6090 -4683
rect -6035 -4689 -6001 -4181
rect -6508 -5194 -6498 -5141
rect -6445 -5194 -6435 -5141
rect -6635 -5375 -6625 -5322
rect -6572 -5375 -6562 -5322
rect -6498 -6248 -6445 -5194
rect -6124 -5232 -6090 -4998
rect -6144 -5285 -6134 -5232
rect -6081 -5285 -6071 -5232
rect -6301 -5519 -6091 -5518
rect -5946 -5519 -5912 -2388
rect -5856 -2780 -5822 -2447
rect -5768 -2530 -5734 -2389
rect -5787 -2583 -5777 -2530
rect -5724 -2583 -5714 -2530
rect -5876 -2833 -5866 -2780
rect -5813 -2833 -5803 -2780
rect -5856 -2943 -5822 -2833
rect -5679 -2949 -5645 -2447
rect -5857 -3819 -5823 -3311
rect -5768 -3516 -5734 -3258
rect -5787 -3569 -5777 -3516
rect -5724 -3569 -5714 -3516
rect -5679 -3819 -5645 -3311
rect -5857 -4689 -5823 -4181
rect -5768 -4271 -5734 -4128
rect -5788 -4324 -5778 -4271
rect -5725 -4324 -5715 -4271
rect -5679 -4689 -5645 -4181
rect -6301 -5552 -5912 -5519
rect -6301 -5636 -6267 -5552
rect -6125 -5553 -5912 -5552
rect -6125 -5639 -6091 -5553
rect -5946 -5612 -5912 -5553
rect -5857 -5559 -5823 -5051
rect -5768 -5415 -5734 -4999
rect -5787 -5468 -5777 -5415
rect -5724 -5468 -5714 -5415
rect -5679 -5559 -5645 -5051
rect -5590 -5612 -5556 -2388
rect -5501 -2949 -5467 -2441
rect -5412 -2668 -5378 -2388
rect -5431 -2721 -5421 -2668
rect -5368 -2721 -5358 -2668
rect -5323 -2949 -5289 -2441
rect -5501 -3819 -5467 -3311
rect -5412 -3640 -5378 -3258
rect -5432 -3693 -5422 -3640
rect -5369 -3693 -5359 -3640
rect -5323 -3819 -5289 -3311
rect -5501 -4689 -5467 -4181
rect -5412 -4506 -5378 -4128
rect -5432 -4559 -5422 -4506
rect -5369 -4559 -5359 -4506
rect -5323 -4689 -5289 -4181
rect -5501 -5559 -5467 -5051
rect -5412 -5141 -5378 -4998
rect -5432 -5194 -5422 -5141
rect -5369 -5194 -5359 -5141
rect -5323 -5559 -5289 -5051
rect -5234 -5612 -5200 -2388
rect -5145 -2949 -5111 -2441
rect -5056 -2530 -5022 -2388
rect -5076 -2583 -5066 -2530
rect -5013 -2583 -5003 -2530
rect -4967 -2949 -4933 -2441
rect -5145 -3819 -5111 -3311
rect -5056 -3401 -5022 -3259
rect -5076 -3454 -5066 -3401
rect -5013 -3454 -5003 -3401
rect -4967 -3819 -4933 -3311
rect -5145 -4689 -5111 -4181
rect -5056 -4390 -5022 -4127
rect -5076 -4443 -5066 -4390
rect -5013 -4443 -5003 -4390
rect -4967 -4689 -4933 -4181
rect -5145 -5559 -5111 -5051
rect -5056 -5233 -5022 -4998
rect -5076 -5286 -5066 -5233
rect -5013 -5286 -5003 -5233
rect -4967 -5559 -4933 -5051
rect -4878 -5612 -4844 -2388
rect -4789 -2949 -4755 -2441
rect -4700 -2668 -4666 -2388
rect -4720 -2721 -4710 -2668
rect -4657 -2721 -4647 -2668
rect -4611 -2949 -4577 -2441
rect -4789 -3819 -4755 -3311
rect -4700 -3401 -4666 -3258
rect -4720 -3454 -4710 -3401
rect -4657 -3454 -4647 -3401
rect -4611 -3819 -4577 -3311
rect -4789 -4689 -4755 -4181
rect -4700 -4390 -4666 -4128
rect -4719 -4443 -4709 -4390
rect -4656 -4443 -4646 -4390
rect -4611 -4689 -4577 -4181
rect -4789 -5559 -4755 -5051
rect -4700 -5322 -4666 -4998
rect -4720 -5375 -4710 -5322
rect -4657 -5375 -4647 -5322
rect -4611 -5559 -4577 -5051
rect -4522 -5612 -4488 -2388
rect -4433 -2949 -4399 -2441
rect -4344 -2530 -4310 -2388
rect -4364 -2583 -4354 -2530
rect -4301 -2583 -4291 -2530
rect -4255 -2949 -4221 -2441
rect -4433 -3819 -4399 -3311
rect -4344 -3640 -4310 -3258
rect -4363 -3693 -4353 -3640
rect -4300 -3693 -4290 -3640
rect -4254 -3819 -4220 -3311
rect -4433 -4689 -4399 -4181
rect -4344 -4506 -4310 -4128
rect -4363 -4559 -4353 -4506
rect -4300 -4559 -4290 -4506
rect -4255 -4689 -4221 -4181
rect -4433 -5559 -4399 -5051
rect -4344 -5141 -4310 -4998
rect -4363 -5194 -4353 -5141
rect -4300 -5194 -4290 -5141
rect -4255 -5559 -4221 -5051
rect -4166 -5612 -4132 -2388
rect -4077 -2949 -4043 -2441
rect -3988 -2668 -3954 -2388
rect -4008 -2721 -3998 -2668
rect -3945 -2721 -3935 -2668
rect -3899 -2780 -3865 -2441
rect -3810 -2446 -3776 -2388
rect -3633 -2446 -3599 -2364
rect -3454 -2446 -3420 -2370
rect -1099 -2425 -1065 -1963
rect -3810 -2480 -3420 -2446
rect -1119 -2478 -1109 -2425
rect -1056 -2478 -1046 -2425
rect -762 -2478 -752 -2425
rect -699 -2478 -689 -2425
rect -3918 -2833 -3908 -2780
rect -3855 -2833 -3845 -2780
rect -3899 -2949 -3865 -2833
rect -4077 -3819 -4043 -3311
rect -3988 -3516 -3954 -3258
rect -4008 -3569 -3998 -3516
rect -3945 -3569 -3935 -3516
rect -3899 -3819 -3865 -3311
rect -4077 -4689 -4043 -4181
rect -3988 -4271 -3954 -4128
rect -4008 -4324 -3998 -4271
rect -3945 -4324 -3935 -4271
rect -3899 -4689 -3865 -4181
rect -4077 -5559 -4043 -5051
rect -3988 -5415 -3954 -4998
rect -4007 -5468 -3997 -5415
rect -3944 -5468 -3934 -5415
rect -3899 -5559 -3865 -5051
rect -3810 -5612 -3776 -2480
rect -2634 -2611 -2624 -2558
rect -2571 -2611 -2561 -2558
rect -1295 -2611 -1285 -2558
rect -1232 -2611 -1222 -2558
rect -3308 -2721 -3298 -2668
rect -3245 -2721 -3235 -2668
rect -3741 -2833 -3731 -2780
rect -3678 -2833 -3668 -2780
rect -3721 -2949 -3687 -2833
rect -3721 -3819 -3687 -3311
rect -3632 -3316 -3598 -3258
rect -3454 -3316 -3420 -3234
rect -3632 -3350 -3420 -3316
rect -3632 -3401 -3598 -3350
rect -3652 -3454 -3642 -3401
rect -3589 -3454 -3579 -3401
rect -3298 -3516 -3245 -2721
rect -3141 -3454 -3131 -3401
rect -3078 -3454 -3068 -3401
rect -3308 -3569 -3298 -3516
rect -3245 -3569 -3235 -3516
rect -3721 -4689 -3687 -4181
rect -3632 -4186 -3598 -4128
rect -3453 -4186 -3419 -4076
rect -3632 -4220 -3419 -4186
rect -3632 -4390 -3598 -4220
rect -3652 -4443 -3642 -4390
rect -3589 -4443 -3579 -4390
rect -3298 -4506 -3245 -3569
rect -3308 -4559 -3298 -4506
rect -3245 -4559 -3235 -4506
rect -3632 -5056 -3598 -4999
rect -3453 -5056 -3419 -4946
rect -3632 -5090 -3419 -5056
rect -3632 -5319 -3598 -5090
rect -3652 -5372 -3642 -5319
rect -3589 -5372 -3579 -5319
rect -3298 -5416 -3245 -4559
rect -3130 -5233 -3077 -3454
rect -3140 -5286 -3130 -5233
rect -3077 -5286 -3067 -5233
rect -2624 -5324 -2571 -2611
rect -1276 -2885 -1242 -2611
rect -1207 -2718 -1197 -2665
rect -1144 -2718 -1134 -2665
rect -1187 -2825 -1153 -2718
rect -1099 -2884 -1065 -2478
rect -940 -2611 -930 -2558
rect -877 -2611 -867 -2558
rect -1029 -2718 -1019 -2665
rect -966 -2718 -956 -2665
rect -1009 -2831 -975 -2718
rect -920 -2886 -886 -2611
rect -851 -2718 -841 -2665
rect -788 -2718 -778 -2665
rect -831 -2831 -797 -2718
rect -742 -2884 -708 -2478
rect -208 -2605 182 -2571
rect -208 -2883 -174 -2605
rect -139 -2718 -129 -2665
rect -76 -2718 -66 -2665
rect 40 -2718 50 -2665
rect 103 -2718 113 -2665
rect -119 -2831 -85 -2718
rect 59 -2831 93 -2718
rect 148 -2886 182 -2605
rect 217 -2718 227 -2665
rect 280 -2718 290 -2665
rect 237 -2831 271 -2718
rect 594 -2825 628 -1467
rect 7034 -1909 7080 -1737
rect 16034 -1909 16080 -1737
rect 5327 -2258 5337 -2205
rect 5390 -2258 5400 -2205
rect 1909 -2479 1919 -2426
rect 1972 -2479 1982 -2426
rect 2265 -2479 2275 -2426
rect 2328 -2479 2338 -2426
rect 1038 -2611 1428 -2577
rect 930 -2718 940 -2665
rect 993 -2718 1003 -2665
rect 949 -2831 983 -2718
rect 1038 -2886 1072 -2611
rect 1107 -2718 1117 -2665
rect 1170 -2718 1180 -2665
rect 1285 -2718 1295 -2665
rect 1348 -2718 1358 -2665
rect 1127 -2831 1161 -2718
rect 1305 -2831 1339 -2718
rect -1454 -3282 -1420 -3140
rect -1365 -3282 -1331 -3199
rect -1276 -3282 -1242 -3141
rect -1454 -3316 -1242 -3282
rect -1454 -3317 -1420 -3316
rect -1655 -3510 -1645 -3449
rect -1584 -3510 -1574 -3449
rect -2014 -4465 -2004 -4412
rect -1951 -4465 -1941 -4412
rect -2003 -4517 -1950 -4465
rect -2634 -5377 -2624 -5324
rect -2571 -5377 -2561 -5324
rect -3308 -5469 -3298 -5416
rect -3245 -5469 -3235 -5416
rect -5946 -6016 -5912 -5869
rect -5966 -6069 -5956 -6016
rect -5903 -6069 -5893 -6016
rect -5768 -6131 -5734 -5868
rect -5590 -6016 -5556 -5868
rect -5611 -6069 -5601 -6016
rect -5548 -6069 -5538 -6016
rect -5788 -6184 -5778 -6131
rect -5725 -6184 -5715 -6131
rect -5412 -6248 -5378 -5868
rect -5234 -6016 -5200 -5868
rect -5254 -6069 -5244 -6016
rect -5191 -6069 -5181 -6016
rect -5056 -6131 -5022 -5869
rect -5075 -6184 -5065 -6131
rect -5012 -6184 -5002 -6131
rect -6508 -6301 -6498 -6248
rect -6445 -6301 -6435 -6248
rect -5431 -6301 -5421 -6248
rect -5368 -6301 -5358 -6248
rect -4967 -6376 -4933 -5927
rect -4878 -6016 -4844 -5868
rect -4898 -6069 -4888 -6016
rect -4835 -6069 -4825 -6016
rect -4700 -6248 -4666 -5868
rect -4720 -6301 -4710 -6248
rect -4657 -6301 -4647 -6248
rect -4613 -6376 -4579 -5921
rect -4522 -6016 -4488 -5868
rect -4542 -6069 -4532 -6016
rect -4479 -6069 -4469 -6016
rect -4344 -6131 -4310 -5868
rect -4166 -6016 -4132 -5868
rect -4185 -6069 -4175 -6016
rect -4122 -6069 -4112 -6016
rect -4364 -6184 -4354 -6131
rect -4301 -6184 -4291 -6131
rect -3988 -6247 -3954 -5868
rect -3810 -5928 -3776 -5868
rect -3632 -5928 -3598 -5836
rect -3455 -5928 -3421 -5814
rect -3810 -5962 -3421 -5928
rect -3810 -6016 -3776 -5962
rect -3830 -6069 -3820 -6016
rect -3767 -6069 -3757 -6016
rect -3298 -6131 -3245 -5469
rect -2624 -6007 -2571 -5377
rect -2634 -6060 -2624 -6007
rect -2571 -6060 -2561 -6007
rect -3308 -6184 -3298 -6131
rect -3245 -6184 -3235 -6131
rect -4008 -6300 -3998 -6247
rect -3945 -6300 -3935 -6247
rect -3988 -6301 -3954 -6300
rect -4967 -6378 -4579 -6376
rect -4967 -6410 -4786 -6378
rect -4796 -6431 -4786 -6410
rect -4733 -6410 -4579 -6378
rect -4733 -6431 -4723 -6410
rect -2002 -6714 -1950 -4517
rect -1886 -5285 -1876 -5232
rect -1823 -5285 -1813 -5232
rect -1646 -5278 -1585 -3510
rect -1296 -3624 -1286 -3571
rect -1233 -3624 -1223 -3571
rect -1276 -3784 -1242 -3624
rect -1186 -3724 -1152 -3200
rect -1118 -3509 -1108 -3456
rect -1055 -3509 -1045 -3456
rect -1098 -3784 -1064 -3509
rect -1009 -3724 -975 -3200
rect -939 -3624 -929 -3571
rect -876 -3624 -866 -3571
rect -919 -3784 -885 -3624
rect -831 -3724 -797 -3200
rect -653 -3282 -619 -3199
rect -563 -3282 -529 -3140
rect -474 -3282 -440 -3199
rect -385 -3282 -351 -3140
rect -295 -3282 -261 -3199
rect -653 -3301 -261 -3282
rect -653 -3316 -484 -3301
rect -494 -3354 -484 -3316
rect -431 -3316 -261 -3301
rect -431 -3354 -421 -3316
rect -760 -3509 -750 -3456
rect -697 -3509 -687 -3456
rect -406 -3509 -396 -3456
rect -343 -3509 -333 -3456
rect -742 -3784 -708 -3509
rect -583 -3624 -573 -3571
rect -520 -3624 -510 -3571
rect -564 -3784 -530 -3624
rect -386 -3784 -352 -3509
rect -208 -3571 -174 -3140
rect -227 -3624 -217 -3571
rect -164 -3624 -154 -3571
rect -208 -3784 -174 -3624
rect -119 -3724 -85 -3200
rect -30 -3456 4 -3138
rect 327 -3456 361 -3139
rect 414 -3283 448 -3199
rect 504 -3283 538 -3141
rect 592 -3283 626 -3199
rect 682 -3283 716 -3141
rect 771 -3283 805 -3199
rect 414 -3301 805 -3283
rect 414 -3317 583 -3301
rect 573 -3354 583 -3317
rect 636 -3317 805 -3301
rect 636 -3354 646 -3317
rect -49 -3509 -39 -3456
rect 14 -3509 24 -3456
rect 307 -3509 317 -3456
rect 370 -3509 380 -3456
rect -30 -3784 4 -3509
rect 589 -3598 623 -3354
rect 860 -3456 894 -3139
rect 1216 -3456 1250 -3136
rect 840 -3509 850 -3456
rect 903 -3509 913 -3456
rect 1196 -3509 1206 -3456
rect 1259 -3509 1269 -3456
rect 59 -3632 1160 -3598
rect 59 -3725 93 -3632
rect 149 -3633 271 -3632
rect 149 -3784 183 -3633
rect 237 -3725 271 -3633
rect 948 -3725 982 -3632
rect 1038 -3783 1072 -3632
rect 1126 -3725 1160 -3632
rect 1216 -3802 1250 -3509
rect 1306 -3724 1340 -3200
rect 1394 -3564 1428 -2611
rect 1928 -2885 1962 -2479
rect 2087 -2607 2097 -2554
rect 2150 -2607 2160 -2554
rect 1997 -2718 2007 -2665
rect 2060 -2718 2070 -2665
rect 2017 -2831 2051 -2718
rect 2105 -2881 2139 -2607
rect 2176 -2718 2186 -2665
rect 2239 -2718 2249 -2665
rect 2195 -2831 2229 -2718
rect 2285 -2887 2319 -2479
rect 3183 -2480 3193 -2427
rect 3246 -2480 3256 -2427
rect 2443 -2607 2453 -2554
rect 2506 -2606 2931 -2554
rect 2506 -2607 2516 -2606
rect 2353 -2718 2363 -2665
rect 2416 -2718 2426 -2665
rect 2373 -2831 2407 -2718
rect 2462 -2885 2496 -2607
rect 1482 -3283 1516 -3199
rect 1572 -3283 1606 -3140
rect 1662 -3283 1696 -3199
rect 1750 -3283 1784 -3140
rect 1840 -3283 1874 -3199
rect 1482 -3301 1874 -3283
rect 1482 -3317 1654 -3301
rect 1644 -3354 1654 -3317
rect 1707 -3317 1874 -3301
rect 1707 -3354 1717 -3317
rect 1552 -3509 1562 -3456
rect 1615 -3509 1625 -3456
rect 1909 -3509 1919 -3456
rect 1972 -3509 1982 -3456
rect 1374 -3617 1384 -3564
rect 1437 -3617 1447 -3564
rect 1394 -3809 1428 -3617
rect 1572 -3784 1606 -3509
rect 1731 -3617 1741 -3564
rect 1794 -3617 1804 -3564
rect 1750 -3786 1784 -3617
rect 1929 -3787 1963 -3509
rect 2017 -3724 2051 -3200
rect 2087 -3617 2097 -3564
rect 2150 -3617 2160 -3564
rect 2106 -3785 2140 -3617
rect 2196 -3724 2230 -3200
rect 2265 -3509 2275 -3456
rect 2328 -3509 2338 -3456
rect 2284 -3785 2318 -3509
rect 2373 -3724 2407 -3200
rect 2462 -3284 2496 -3141
rect 2551 -3284 2585 -3199
rect 2641 -3284 2675 -3141
rect 2462 -3318 2675 -3284
rect 2441 -3617 2451 -3564
rect 2504 -3617 2514 -3564
rect 2462 -3786 2496 -3617
rect -1454 -4184 -1420 -4041
rect -1366 -4184 -1332 -4099
rect -1276 -4184 -1242 -4040
rect -1454 -4218 -1242 -4184
rect -1454 -4541 -1242 -4507
rect -1454 -4685 -1420 -4541
rect -1365 -4624 -1331 -4541
rect -1276 -4706 -1242 -4541
rect -1187 -4625 -1153 -4101
rect -1009 -4624 -975 -4100
rect -831 -4192 -797 -4100
rect -653 -4192 -619 -4101
rect -474 -4192 -440 -4101
rect -297 -4192 -263 -4100
rect -851 -4245 -841 -4192
rect -788 -4245 -778 -4192
rect -672 -4245 -662 -4192
rect -609 -4245 -599 -4192
rect -493 -4245 -483 -4192
rect -430 -4245 -420 -4192
rect -316 -4245 -306 -4192
rect -253 -4245 -243 -4192
rect -831 -4624 -797 -4245
rect -653 -4625 -619 -4245
rect -474 -4625 -440 -4245
rect -297 -4624 -263 -4245
rect -119 -4624 -85 -4100
rect -1277 -5097 -1243 -4939
rect -1297 -5150 -1287 -5097
rect -1234 -5150 -1224 -5097
rect -1876 -5337 -1823 -5285
rect -1875 -6364 -1823 -5337
rect -1656 -5339 -1646 -5278
rect -1585 -5339 -1575 -5278
rect -1454 -5442 -1242 -5408
rect -1454 -5585 -1420 -5442
rect -1363 -5524 -1329 -5442
rect -1276 -5592 -1242 -5442
rect -1187 -5525 -1153 -4995
rect -1097 -5213 -1063 -4938
rect -1115 -5266 -1105 -5213
rect -1052 -5266 -1042 -5213
rect -1009 -5524 -975 -4994
rect -919 -5097 -885 -4937
rect -939 -5150 -929 -5097
rect -876 -5150 -866 -5097
rect -830 -5524 -796 -4994
rect -741 -5213 -707 -4937
rect -563 -5097 -529 -4940
rect -582 -5150 -572 -5097
rect -519 -5150 -509 -5097
rect -386 -5213 -352 -4937
rect -208 -5097 -174 -4910
rect -228 -5150 -218 -5097
rect -165 -5150 -155 -5097
rect -761 -5266 -751 -5213
rect -698 -5266 -688 -5213
rect -406 -5266 -396 -5213
rect -343 -5266 -333 -5213
rect -654 -5434 -262 -5400
rect -654 -5523 -620 -5434
rect -563 -5604 -529 -5434
rect -474 -5524 -440 -5434
rect -385 -5612 -351 -5434
rect -296 -5524 -262 -5434
rect -1274 -6364 -1240 -5839
rect -1886 -6417 -1876 -6364
rect -1823 -6417 -1813 -6364
rect -1292 -6417 -1282 -6364
rect -1229 -6417 -1219 -6364
rect -1099 -6479 -1065 -5845
rect -919 -6365 -885 -5833
rect -938 -6417 -928 -6365
rect -876 -6417 -866 -6365
rect -742 -6479 -708 -5839
rect -1120 -6532 -1110 -6479
rect -1057 -6532 -1047 -6479
rect -762 -6532 -752 -6479
rect -699 -6532 -689 -6479
rect -476 -6493 -442 -5901
rect -208 -6077 -174 -5150
rect -119 -5380 -85 -4994
rect -30 -5213 4 -4938
rect 59 -5091 93 -4992
rect 148 -5091 182 -3952
rect 326 -4304 360 -4040
rect 416 -4192 450 -4094
rect 397 -4245 407 -4192
rect 460 -4245 470 -4192
rect 307 -4357 317 -4304
rect 370 -4357 380 -4304
rect 326 -4706 360 -4357
rect 416 -4624 450 -4245
rect 504 -4412 538 -4040
rect 593 -4192 627 -4101
rect 573 -4245 583 -4192
rect 636 -4245 646 -4192
rect 485 -4465 495 -4412
rect 548 -4465 558 -4412
rect 504 -4703 538 -4465
rect 593 -4625 627 -4245
rect 682 -4304 716 -4040
rect 771 -4192 805 -4100
rect 751 -4245 761 -4192
rect 814 -4245 824 -4192
rect 663 -4357 673 -4304
rect 726 -4357 736 -4304
rect 682 -4687 716 -4357
rect 771 -4624 805 -4245
rect 860 -4412 894 -4040
rect 840 -4465 850 -4412
rect 903 -4465 913 -4412
rect 860 -4716 894 -4465
rect 236 -5091 270 -4999
rect 948 -5091 982 -5000
rect 1039 -5091 1073 -3989
rect 1305 -4624 1339 -4094
rect 1484 -4192 1518 -4094
rect 1661 -4192 1695 -4094
rect 1839 -4192 1873 -4094
rect 2017 -4192 2051 -4094
rect 1464 -4245 1474 -4192
rect 1527 -4245 1537 -4192
rect 1642 -4245 1652 -4192
rect 1705 -4245 1715 -4192
rect 1820 -4245 1830 -4192
rect 1883 -4245 1893 -4192
rect 1998 -4245 2008 -4192
rect 2061 -4245 2071 -4192
rect 1484 -4624 1518 -4245
rect 1661 -4624 1695 -4245
rect 1839 -4624 1873 -4245
rect 2017 -4624 2051 -4245
rect 2195 -4625 2229 -4095
rect 2373 -4624 2407 -4094
rect 2463 -4182 2497 -4038
rect 2552 -4182 2586 -4104
rect 2640 -4180 2674 -4020
rect 2640 -4182 2792 -4180
rect 2463 -4214 2792 -4182
rect 2463 -4216 2674 -4214
rect 2528 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect 2550 -4506 2584 -4327
rect 2758 -4446 2792 -4214
rect 2462 -4540 2674 -4506
rect 2736 -4507 2746 -4446
rect 2807 -4507 2817 -4446
rect 2758 -4508 2792 -4507
rect 2462 -4683 2496 -4540
rect 2550 -4623 2584 -4540
rect 2640 -4713 2674 -4540
rect 1128 -5091 1162 -5002
rect 59 -5125 1162 -5091
rect -51 -5266 -41 -5213
rect 12 -5266 22 -5213
rect 306 -5266 316 -5213
rect 369 -5266 379 -5213
rect -138 -5433 -128 -5380
rect -75 -5433 -65 -5380
rect -119 -5524 -85 -5433
rect -30 -5603 4 -5266
rect 40 -5433 50 -5380
rect 103 -5433 113 -5380
rect 218 -5433 228 -5380
rect 281 -5433 291 -5380
rect 59 -5524 93 -5433
rect 238 -5524 272 -5433
rect 326 -5586 360 -5266
rect 593 -5315 627 -5125
rect 1216 -5213 1250 -4940
rect 840 -5266 850 -5213
rect 903 -5266 913 -5213
rect 1197 -5266 1207 -5213
rect 1260 -5266 1270 -5213
rect 415 -5349 804 -5315
rect 415 -5524 449 -5349
rect 505 -5620 539 -5349
rect 592 -5523 626 -5349
rect 681 -5606 715 -5349
rect 770 -5524 804 -5349
rect 860 -5585 894 -5266
rect 930 -5434 940 -5381
rect 993 -5434 1003 -5381
rect 1109 -5433 1119 -5380
rect 1172 -5433 1182 -5380
rect 949 -5524 983 -5434
rect 1128 -5524 1162 -5433
rect 1216 -5623 1250 -5266
rect 1306 -5380 1340 -4994
rect 1394 -5093 1428 -4913
rect 1375 -5146 1385 -5093
rect 1438 -5146 1448 -5093
rect 1286 -5433 1296 -5380
rect 1349 -5433 1359 -5380
rect 1306 -5524 1340 -5433
rect 149 -6077 183 -5822
rect -208 -6111 183 -6077
rect 237 -6250 271 -5901
rect 217 -6303 227 -6250
rect 280 -6303 290 -6250
rect 594 -6493 628 -5899
rect 951 -6250 985 -5899
rect 1038 -6081 1072 -5808
rect 1394 -6081 1428 -5146
rect 1572 -5213 1606 -4938
rect 1750 -5093 1784 -4938
rect 1730 -5146 1740 -5093
rect 1793 -5146 1803 -5093
rect 1927 -5213 1961 -4940
rect 1553 -5266 1563 -5213
rect 1616 -5266 1626 -5213
rect 1907 -5266 1917 -5213
rect 1970 -5266 1980 -5213
rect 1482 -5433 1874 -5399
rect 1482 -5523 1516 -5433
rect 1573 -5607 1607 -5433
rect 1661 -5523 1695 -5433
rect 1749 -5604 1783 -5433
rect 1840 -5523 1874 -5433
rect 2018 -5523 2052 -4993
rect 2106 -5093 2140 -4939
rect 2086 -5146 2096 -5093
rect 2149 -5146 2159 -5093
rect 2195 -5525 2229 -4995
rect 2284 -5213 2318 -4939
rect 2264 -5266 2274 -5213
rect 2327 -5266 2337 -5213
rect 2373 -5525 2407 -4995
rect 2462 -5093 2496 -4937
rect 2443 -5146 2453 -5093
rect 2506 -5146 2516 -5093
rect 2463 -5442 2674 -5408
rect 2463 -5585 2497 -5442
rect 2550 -5525 2584 -5442
rect 2640 -5587 2674 -5442
rect 1038 -6115 1428 -6081
rect 932 -6303 942 -6250
rect 995 -6303 1005 -6250
rect 1662 -6493 1696 -5901
rect 1928 -6124 1962 -5839
rect 2106 -6007 2140 -5842
rect 2086 -6060 2096 -6007
rect 2149 -6060 2159 -6007
rect 2284 -6124 2318 -5841
rect 2462 -6007 2496 -5839
rect 2442 -6060 2452 -6007
rect 2505 -6060 2515 -6007
rect 1908 -6177 1918 -6124
rect 1971 -6177 1981 -6124
rect 2265 -6177 2275 -6124
rect 2328 -6177 2338 -6124
rect 2879 -6365 2931 -2606
rect 3194 -4805 3246 -2480
rect 3184 -4857 3194 -4805
rect 3246 -4857 3256 -4805
rect 4761 -4857 4771 -4805
rect 4823 -4857 4833 -4805
rect 2869 -6417 2879 -6365
rect 2931 -6417 2941 -6365
rect -476 -6527 1696 -6493
rect -742 -6598 -708 -6532
rect 4771 -6597 4823 -4857
rect 5027 -5059 5037 -5006
rect 5090 -5059 5100 -5006
rect 4895 -5265 4905 -5212
rect 4958 -5265 4968 -5212
rect -763 -6651 -753 -6598
rect -700 -6651 -690 -6598
rect 4762 -6650 4772 -6597
rect 4825 -6650 4835 -6597
rect -2013 -6767 -2003 -6714
rect -1950 -6767 -1940 -6714
rect 4771 -6891 4823 -6650
rect 4905 -6889 4958 -5265
rect 5037 -6887 5090 -5059
rect 5337 -5527 5390 -2258
rect 6670 -2263 6680 -2199
rect 6744 -2263 6754 -2199
rect 7034 -2687 7080 -2509
rect 16034 -2687 16080 -2509
rect 6212 -3515 6222 -3451
rect 6286 -3515 6296 -3451
rect 7034 -3709 7080 -3537
rect 16034 -3709 16080 -3537
rect 7034 -4487 7080 -4309
rect 16034 -4487 16080 -4309
rect 5604 -5271 5614 -5207
rect 5678 -5271 5688 -5207
rect 7034 -5509 7080 -5337
rect 16034 -5509 16080 -5337
rect 5327 -5580 5337 -5527
rect 5390 -5580 5400 -5527
rect 7034 -6287 7080 -6109
rect 16034 -6287 16080 -6109
rect 17826 -6521 17901 -4862
rect 17821 -6585 17831 -6521
rect 17895 -6585 17905 -6521
rect 4760 -6944 4770 -6891
rect 4823 -6944 4833 -6891
rect 4896 -6942 4906 -6889
rect 4959 -6942 4969 -6889
rect 5028 -6940 5038 -6887
rect 5091 -6940 5101 -6887
rect 7034 -7309 7080 -7137
rect 16034 -7309 16080 -7137
rect -3883 -7697 -3873 -7691
rect -5629 -7731 -3873 -7697
rect -5628 -7875 -5594 -7731
rect -5544 -7824 -5500 -7731
rect -5450 -7875 -5416 -7731
rect -5366 -7830 -5322 -7731
rect -5188 -7830 -5144 -7731
rect -5094 -7876 -5060 -7731
rect -5010 -7830 -4966 -7731
rect -4832 -7830 -4788 -7731
rect -4738 -7876 -4704 -7731
rect -4654 -7830 -4610 -7731
rect -4476 -7830 -4432 -7731
rect -4382 -7876 -4348 -7731
rect -4298 -7830 -4254 -7731
rect -3883 -7743 -3873 -7731
rect -3821 -7743 -3811 -7691
rect -3741 -7790 -3731 -7785
rect -4026 -7824 -3731 -7790
rect -4026 -7880 -3992 -7824
rect -3741 -7837 -3731 -7824
rect -3679 -7837 -3669 -7785
rect -3551 -7840 -3541 -7788
rect -3489 -7840 -3479 -7788
rect -5628 -11756 -5594 -8130
rect -5544 -8340 -5500 -8214
rect -5544 -8890 -5500 -8764
rect -5544 -9440 -5500 -9314
rect -5544 -9990 -5500 -9864
rect -5544 -10540 -5500 -10414
rect -5544 -11090 -5500 -10964
rect -5544 -11655 -5500 -11485
rect -5450 -11799 -5416 -8130
rect -5366 -8340 -5322 -8214
rect -5366 -8890 -5322 -8764
rect -5366 -9440 -5322 -9314
rect -5366 -9990 -5322 -9864
rect -5366 -10540 -5322 -10414
rect -5366 -11090 -5322 -10964
rect -5272 -11174 -5238 -8130
rect -5188 -8340 -5144 -8214
rect -5188 -8890 -5144 -8764
rect -5188 -9440 -5144 -9314
rect -5188 -9990 -5144 -9864
rect -5188 -10540 -5144 -10414
rect -5188 -11090 -5144 -10964
rect -5364 -11655 -5320 -11485
rect -5272 -12119 -5238 -11431
rect -5188 -11656 -5144 -11486
rect -5094 -11830 -5060 -8131
rect -5010 -8341 -4966 -8215
rect -5010 -8890 -4966 -8764
rect -5010 -9440 -4966 -9314
rect -5010 -9990 -4966 -9864
rect -5010 -10540 -4966 -10414
rect -5010 -11090 -4966 -10964
rect -4916 -11174 -4882 -8130
rect -4832 -8340 -4788 -8214
rect -4832 -8890 -4788 -8764
rect -4832 -9440 -4788 -9314
rect -4832 -9990 -4788 -9864
rect -4832 -10540 -4788 -10414
rect -4832 -11090 -4788 -10964
rect -5010 -11655 -4966 -11485
rect -4916 -12119 -4882 -11430
rect -4832 -11657 -4788 -11487
rect -4738 -11788 -4704 -8130
rect -4654 -8340 -4610 -8214
rect -4654 -8890 -4610 -8764
rect -4654 -9440 -4610 -9314
rect -4654 -9990 -4610 -9864
rect -4654 -10540 -4610 -10414
rect -4654 -11090 -4610 -10964
rect -4560 -11174 -4526 -8130
rect -4476 -8340 -4432 -8214
rect -4476 -8890 -4432 -8764
rect -4476 -9440 -4432 -9314
rect -4476 -9990 -4432 -9864
rect -4476 -10540 -4432 -10414
rect -4476 -11090 -4432 -10964
rect -4654 -11657 -4610 -11487
rect -4560 -12119 -4526 -11430
rect -4476 -11656 -4432 -11486
rect -4382 -11804 -4348 -8130
rect -4298 -8340 -4254 -8214
rect -4298 -8890 -4254 -8764
rect -4298 -9440 -4254 -9314
rect -4298 -9990 -4254 -9864
rect -4298 -10540 -4254 -10414
rect -4298 -11090 -4254 -10964
rect -4204 -11174 -4170 -8130
rect -4120 -8340 -4076 -8214
rect -4120 -8890 -4076 -8764
rect -4120 -9440 -4076 -9314
rect -4120 -9990 -4076 -9864
rect -4120 -10540 -4076 -10414
rect -4120 -11090 -4076 -10964
rect -4026 -11174 -3992 -8130
rect -4298 -11656 -4254 -11486
rect -4204 -12119 -4170 -11430
rect -4120 -11656 -4076 -11486
rect -4113 -12119 -4079 -12030
rect -4026 -12119 -3992 -11430
rect -5272 -12153 -3611 -12119
rect -5512 -12324 -5502 -12271
rect -5449 -12324 -5439 -12271
rect -6976 -12565 -6077 -12512
rect -6024 -12565 -6014 -12512
rect -5636 -12565 -5626 -12512
rect -5573 -12565 -5563 -12512
rect -6233 -13115 -6223 -13062
rect -6170 -13115 -6160 -13062
rect -6976 -13905 -6426 -13852
rect -6373 -13905 -6363 -13852
rect -6223 -14055 -6170 -13115
rect -6077 -13745 -6024 -12565
rect -5922 -12628 -5877 -12612
rect -5922 -12700 -5876 -12628
rect -5817 -12668 -5778 -12612
rect -5617 -12662 -5583 -12565
rect -5824 -12700 -5778 -12668
rect -5492 -12700 -5458 -12324
rect -5010 -12325 -5000 -12272
rect -4947 -12325 -4937 -12272
rect -4512 -12324 -4502 -12271
rect -4449 -12324 -4439 -12271
rect -5386 -12441 -5376 -12388
rect -5323 -12441 -5313 -12388
rect -5137 -12441 -5127 -12388
rect -5074 -12441 -5064 -12388
rect -5367 -12668 -5333 -12441
rect -5117 -12668 -5083 -12441
rect -4992 -12700 -4958 -12325
rect -4887 -12565 -4877 -12512
rect -4824 -12565 -4814 -12512
rect -4637 -12565 -4627 -12512
rect -4574 -12565 -4564 -12512
rect -4867 -12668 -4833 -12565
rect -4617 -12668 -4583 -12565
rect -4492 -12700 -4458 -12324
rect -4387 -12441 -4377 -12388
rect -4324 -12441 -4314 -12388
rect -4367 -12668 -4333 -12441
rect -3938 -12442 -3928 -12389
rect -3875 -12442 -3865 -12389
rect -4172 -12700 -4126 -12612
rect -5824 -12740 -5626 -12700
rect -5574 -12740 -5376 -12700
rect -5324 -12740 -5126 -12700
rect -5074 -12740 -4876 -12700
rect -4823 -12740 -4625 -12700
rect -4574 -12740 -4376 -12700
rect -4324 -12740 -4126 -12700
rect -4074 -12712 -4028 -12612
rect -5818 -12940 -5632 -12900
rect -5574 -12940 -5376 -12900
rect -5324 -12940 -5126 -12900
rect -5074 -12940 -4876 -12900
rect -4825 -12940 -4627 -12900
rect -4574 -12940 -4376 -12900
rect -4324 -12940 -4126 -12900
rect -5744 -13062 -5704 -12940
rect -5761 -13115 -5751 -13062
rect -5698 -13115 -5688 -13062
rect -5495 -13380 -5455 -12940
rect -5245 -13189 -5205 -12940
rect -5261 -13242 -5251 -13189
rect -5198 -13242 -5188 -13189
rect -4995 -13380 -4955 -12940
rect -4746 -13062 -4706 -12940
rect -4762 -13115 -4752 -13062
rect -4699 -13115 -4689 -13062
rect -4495 -13380 -4455 -12940
rect -4244 -13189 -4204 -12940
rect -4261 -13242 -4251 -13189
rect -4198 -13242 -4188 -13189
rect -5824 -13420 -5626 -13380
rect -5574 -13420 -5376 -13380
rect -5324 -13420 -5126 -13380
rect -5074 -13420 -4876 -13380
rect -4824 -13420 -4626 -13380
rect -4574 -13420 -4376 -13380
rect -4324 -13420 -4126 -13380
rect -5922 -13708 -5876 -13608
rect -5824 -13620 -5626 -13580
rect -5574 -13620 -5376 -13580
rect -5324 -13620 -5126 -13580
rect -5074 -13620 -4876 -13580
rect -4824 -13620 -4626 -13580
rect -4574 -13620 -4376 -13580
rect -4324 -13620 -4126 -13580
rect -5824 -13708 -5778 -13620
rect -6087 -13798 -6077 -13745
rect -6024 -13798 -6014 -13745
rect -5720 -13957 -5686 -13620
rect -5617 -13852 -5583 -13652
rect -5367 -13745 -5333 -13652
rect -5386 -13798 -5376 -13745
rect -5323 -13798 -5313 -13745
rect -5636 -13905 -5626 -13852
rect -5573 -13905 -5563 -13852
rect -5740 -14010 -5730 -13957
rect -5677 -14010 -5667 -13957
rect -5240 -14055 -5206 -13620
rect -5117 -13745 -5083 -13652
rect -5136 -13798 -5126 -13745
rect -5073 -13798 -5063 -13745
rect -4867 -13852 -4833 -13652
rect -4887 -13905 -4877 -13852
rect -4824 -13905 -4814 -13852
rect -4742 -13957 -4708 -13620
rect -4617 -13852 -4583 -13652
rect -4367 -13745 -4333 -13652
rect -4386 -13798 -4376 -13745
rect -4323 -13798 -4313 -13745
rect -4637 -13905 -4627 -13852
rect -4574 -13905 -4564 -13852
rect -4762 -14010 -4752 -13957
rect -4699 -14010 -4689 -13957
rect -4240 -14055 -4206 -13620
rect -4172 -13708 -4126 -13620
rect -4074 -13708 -4028 -13608
rect -3928 -13852 -3875 -12442
rect -3798 -13242 -3788 -13189
rect -3735 -13242 -3725 -13189
rect -3938 -13905 -3928 -13852
rect -3875 -13905 -3865 -13852
rect -3928 -13906 -3875 -13905
rect -3788 -13957 -3735 -13242
rect -3798 -14010 -3788 -13957
rect -3735 -14010 -3725 -13957
rect -6233 -14108 -6223 -14055
rect -6170 -14108 -6160 -14055
rect -5260 -14108 -5250 -14055
rect -5197 -14108 -5187 -14055
rect -4260 -14108 -4250 -14055
rect -4197 -14108 -4187 -14055
rect -6965 -14260 -4303 -14226
rect -6028 -14394 -5994 -14260
rect -5939 -14350 -5905 -14260
rect -5850 -14394 -5816 -14260
rect -5761 -14350 -5727 -14260
rect -5583 -14350 -5549 -14260
rect -5405 -14350 -5371 -14260
rect -5227 -14350 -5193 -14260
rect -5049 -14350 -5015 -14260
rect -4871 -14350 -4837 -14260
rect -4693 -14350 -4659 -14260
rect -4515 -14350 -4481 -14260
rect -4337 -14350 -4303 -14260
rect -4248 -14260 -4036 -14226
rect -4248 -14394 -4214 -14260
rect -4159 -14344 -4125 -14260
rect -4070 -14394 -4036 -14260
rect -5850 -14795 -5816 -14651
rect -6169 -14848 -6159 -14795
rect -6106 -14848 -6096 -14795
rect -5870 -14848 -5860 -14795
rect -5807 -14848 -5797 -14795
rect -6159 -15482 -6106 -14848
rect -6028 -14959 -5816 -14925
rect -6027 -15093 -5993 -14959
rect -5939 -15050 -5905 -14959
rect -5850 -15094 -5816 -14959
rect -5761 -15010 -5727 -14700
rect -5672 -15094 -5638 -14650
rect -5583 -15035 -5549 -14719
rect -5494 -14901 -5460 -14650
rect -5514 -14954 -5504 -14901
rect -5451 -14954 -5441 -14901
rect -5405 -15033 -5371 -14717
rect -6169 -15535 -6159 -15482
rect -6106 -15535 -6096 -15482
rect -6159 -16193 -6106 -15535
rect -5850 -15588 -5816 -15350
rect -5870 -15641 -5860 -15588
rect -5807 -15641 -5797 -15588
rect -5761 -15717 -5727 -15401
rect -5672 -15803 -5638 -15350
rect -5583 -15724 -5549 -15408
rect -5494 -15481 -5460 -15350
rect -5514 -15534 -5504 -15481
rect -5451 -15534 -5441 -15481
rect -5405 -15731 -5371 -15415
rect -6028 -16185 -5994 -16049
rect -5939 -16185 -5905 -16094
rect -5850 -16185 -5816 -16050
rect -6169 -16246 -6159 -16193
rect -6106 -16246 -6096 -16193
rect -6028 -16219 -5816 -16185
rect -6159 -17007 -6106 -16246
rect -5850 -16294 -5816 -16219
rect -5870 -16347 -5860 -16294
rect -5807 -16347 -5797 -16294
rect -5761 -16426 -5727 -16110
rect -5672 -16494 -5638 -16050
rect -5583 -16428 -5549 -16112
rect -5494 -16193 -5460 -16050
rect -5514 -16246 -5504 -16193
rect -5451 -16246 -5441 -16193
rect -5405 -16427 -5371 -16111
rect -5316 -16494 -5282 -14650
rect -5227 -15032 -5193 -14716
rect -5138 -14795 -5104 -14651
rect -5157 -14848 -5147 -14795
rect -5094 -14848 -5084 -14795
rect -5049 -15032 -5015 -14716
rect -5227 -15729 -5193 -15413
rect -5138 -15589 -5104 -15350
rect -5158 -15642 -5148 -15589
rect -5095 -15642 -5085 -15589
rect -5049 -15730 -5015 -15414
rect -5227 -16427 -5193 -16111
rect -5138 -16294 -5104 -16051
rect -5158 -16347 -5148 -16294
rect -5095 -16347 -5085 -16294
rect -5049 -16427 -5015 -16111
rect -4960 -16494 -4926 -14650
rect -4871 -15031 -4837 -14715
rect -4782 -14901 -4748 -14650
rect -4801 -14954 -4791 -14901
rect -4738 -14954 -4728 -14901
rect -4693 -15030 -4659 -14714
rect -4871 -15730 -4837 -15414
rect -4782 -15481 -4748 -15350
rect -4802 -15534 -4792 -15481
rect -4739 -15534 -4729 -15481
rect -4693 -15729 -4659 -15413
rect -4871 -16427 -4837 -16111
rect -4782 -16193 -4748 -16050
rect -4802 -16246 -4792 -16193
rect -4739 -16246 -4729 -16193
rect -4693 -16427 -4659 -16111
rect -4604 -16494 -4570 -14650
rect -4515 -15030 -4481 -14714
rect -4426 -14795 -4392 -14650
rect -4446 -14848 -4436 -14795
rect -4383 -14848 -4373 -14795
rect -4337 -15028 -4303 -14712
rect -4248 -14925 -4214 -14650
rect -4159 -14750 -4125 -14700
rect -3664 -14901 -3611 -12153
rect -3541 -13137 -3489 -7840
rect 4761 -7907 4771 -7854
rect 4824 -7907 4834 -7854
rect 4896 -7905 4906 -7852
rect 4959 -7905 4969 -7852
rect 5027 -7903 5037 -7850
rect 5090 -7903 5100 -7850
rect -3392 -7986 -3382 -7933
rect -3329 -7986 -3319 -7933
rect -1392 -7975 -1382 -7922
rect -1329 -7975 -1319 -7922
rect -3542 -13189 -3489 -13137
rect -3552 -13242 -3542 -13189
rect -3489 -13242 -3479 -13189
rect -3382 -14055 -3329 -7986
rect -1372 -8080 -1338 -7975
rect -1213 -7976 -1203 -7923
rect -1150 -7976 -1140 -7923
rect -1035 -7975 -1025 -7922
rect -972 -7975 -962 -7922
rect -858 -7975 -848 -7922
rect -795 -7975 -785 -7922
rect -680 -7975 -670 -7922
rect -617 -7975 -607 -7922
rect -500 -7975 -490 -7922
rect -437 -7975 -427 -7922
rect 745 -7975 755 -7922
rect 808 -7975 818 -7922
rect 922 -7975 932 -7922
rect 985 -7975 995 -7922
rect 1102 -7975 1112 -7922
rect 1165 -7975 1175 -7922
rect -1194 -8081 -1160 -7976
rect -1016 -8081 -982 -7975
rect -838 -8081 -804 -7975
rect -660 -8081 -626 -7975
rect -481 -8081 -447 -7975
rect 765 -8082 799 -7975
rect 942 -8081 976 -7975
rect 1121 -8081 1155 -7975
rect 1279 -7976 1289 -7923
rect 1342 -7976 1352 -7923
rect 1457 -7975 1467 -7922
rect 1520 -7975 1530 -7922
rect 1634 -7975 1644 -7922
rect 1697 -7975 1707 -7922
rect 2880 -7975 2890 -7922
rect 2943 -7975 2953 -7922
rect 3059 -7975 3069 -7922
rect 3122 -7975 3132 -7922
rect 3237 -7975 3247 -7922
rect 3300 -7975 3310 -7922
rect 3414 -7975 3424 -7922
rect 3477 -7975 3487 -7922
rect 1298 -8082 1332 -7976
rect 1476 -8081 1510 -7975
rect 1654 -8081 1688 -7975
rect 2900 -8081 2934 -7975
rect 3078 -8082 3112 -7975
rect 3256 -8081 3290 -7975
rect 3434 -8081 3468 -7975
rect 3593 -7976 3603 -7923
rect 3656 -7976 3666 -7923
rect 3768 -7975 3778 -7922
rect 3831 -7975 3841 -7922
rect 3612 -8081 3646 -7976
rect 3790 -8081 3824 -7975
rect 4198 -7976 4208 -7923
rect 4261 -7976 4271 -7923
rect -2171 -8440 -2137 -8358
rect -1995 -8440 -1961 -8389
rect -2171 -8474 -1961 -8440
rect -1995 -8767 -1961 -8474
rect -1906 -8534 -1872 -8438
rect -1926 -8587 -1916 -8534
rect -1863 -8587 -1853 -8534
rect -1817 -8653 -1783 -8389
rect -1729 -8534 -1695 -8438
rect -1749 -8587 -1739 -8534
rect -1686 -8587 -1676 -8534
rect -1836 -8706 -1826 -8653
rect -1773 -8706 -1763 -8653
rect -2457 -8820 -2447 -8767
rect -2394 -8820 -2384 -8767
rect -2015 -8820 -2005 -8767
rect -1952 -8820 -1942 -8767
rect -2447 -12272 -2394 -8820
rect -2174 -9439 -2140 -9360
rect -1995 -9439 -1961 -8820
rect -2174 -9473 -1961 -9439
rect -2325 -9978 -2315 -9925
rect -2262 -9978 -2252 -9925
rect -2457 -12325 -2447 -12272
rect -2394 -12325 -2384 -12272
rect -3392 -14108 -3382 -14055
rect -3329 -14108 -3319 -14055
rect -4248 -14959 -4036 -14925
rect -3946 -14954 -3936 -14901
rect -3883 -14954 -3611 -14901
rect -4515 -15727 -4481 -15411
rect -4426 -15589 -4392 -15351
rect -4445 -15641 -4435 -15589
rect -4383 -15641 -4373 -15589
rect -4337 -15727 -4303 -15411
rect -4515 -16427 -4481 -16111
rect -4426 -16294 -4392 -16050
rect -4446 -16347 -4436 -16294
rect -4383 -16347 -4373 -16294
rect -4337 -16427 -4303 -16111
rect -4248 -16185 -4214 -14959
rect -4159 -15050 -4125 -14959
rect -4070 -15094 -4036 -14959
rect -3936 -15006 -3883 -14954
rect -3935 -15589 -3883 -15006
rect -3945 -15641 -3935 -15589
rect -3883 -15641 -3873 -15589
rect -4159 -16185 -4125 -16094
rect -4070 -16185 -4036 -16050
rect -4248 -16219 -4036 -16185
rect -4248 -16494 -4214 -16219
rect -3935 -16295 -3883 -15641
rect -2447 -15821 -2394 -12325
rect -2315 -14543 -2262 -9978
rect -1995 -10049 -1961 -9473
rect -1906 -9546 -1872 -9441
rect -1926 -9599 -1916 -9546
rect -1863 -9599 -1853 -9546
rect -1926 -9978 -1916 -9925
rect -1863 -9978 -1853 -9925
rect -2175 -10083 -1961 -10049
rect -1906 -10082 -1872 -9978
rect -2175 -10174 -2141 -10083
rect -1995 -10263 -1961 -10083
rect -1817 -10195 -1783 -8706
rect -1639 -8767 -1605 -8378
rect -1549 -8534 -1515 -8439
rect -1568 -8587 -1558 -8534
rect -1505 -8587 -1495 -8534
rect -1461 -8653 -1427 -8380
rect -1392 -8587 -1382 -8534
rect -1329 -8587 -1319 -8534
rect -1480 -8706 -1470 -8653
rect -1417 -8706 -1407 -8653
rect -1658 -8820 -1648 -8767
rect -1595 -8820 -1585 -8767
rect -1728 -9546 -1694 -9439
rect -1748 -9599 -1738 -9546
rect -1685 -9599 -1675 -9546
rect -1748 -9979 -1738 -9926
rect -1685 -9979 -1675 -9926
rect -1728 -10081 -1694 -9979
rect -1639 -10253 -1605 -8820
rect -1549 -9546 -1515 -9438
rect -1568 -9599 -1558 -9546
rect -1505 -9599 -1495 -9546
rect -1570 -9978 -1560 -9925
rect -1507 -9978 -1497 -9925
rect -1550 -10081 -1516 -9978
rect -1461 -10200 -1427 -8706
rect -1372 -9081 -1338 -8587
rect -1283 -8767 -1249 -8381
rect -1213 -8587 -1203 -8534
rect -1150 -8587 -1140 -8534
rect -1303 -8820 -1293 -8767
rect -1240 -8820 -1230 -8767
rect -1372 -9924 -1338 -9439
rect -1392 -9977 -1382 -9924
rect -1329 -9977 -1319 -9924
rect -1283 -10256 -1249 -8820
rect -1193 -9081 -1159 -8587
rect -1105 -8653 -1071 -8370
rect -1036 -8587 -1026 -8534
rect -973 -8587 -963 -8534
rect -1125 -8706 -1115 -8653
rect -1062 -8706 -1052 -8653
rect -1105 -10208 -1071 -8706
rect -1016 -9081 -982 -8587
rect -927 -8767 -893 -8382
rect -858 -8587 -848 -8534
rect -795 -8587 -785 -8534
rect -946 -8820 -936 -8767
rect -883 -8820 -873 -8767
rect -927 -10257 -893 -8820
rect -838 -9080 -804 -8587
rect -749 -8653 -715 -8368
rect -680 -8587 -670 -8534
rect -617 -8587 -607 -8534
rect -768 -8706 -758 -8653
rect -705 -8706 -695 -8653
rect -749 -10180 -715 -8706
rect -660 -9082 -626 -8587
rect -571 -8766 -537 -8373
rect -501 -8587 -491 -8534
rect -438 -8587 -428 -8534
rect -590 -8819 -580 -8766
rect -527 -8819 -517 -8766
rect -571 -10248 -537 -8819
rect -482 -9081 -448 -8587
rect -393 -8653 -359 -8358
rect -304 -8534 -270 -8439
rect -324 -8587 -314 -8534
rect -261 -8587 -251 -8534
rect -412 -8706 -402 -8653
rect -349 -8706 -339 -8653
rect -393 -10180 -359 -8706
rect -215 -8767 -181 -8371
rect -126 -8534 -92 -8439
rect -146 -8587 -136 -8534
rect -83 -8587 -73 -8534
rect -37 -8653 -3 -8353
rect 52 -8534 86 -8438
rect 32 -8587 42 -8534
rect 95 -8587 105 -8534
rect -57 -8706 -47 -8653
rect 6 -8706 16 -8653
rect -235 -8820 -225 -8767
rect -172 -8820 -162 -8767
rect -303 -9546 -269 -9440
rect -322 -9599 -312 -9546
rect -259 -9599 -249 -9546
rect -324 -9978 -314 -9925
rect -261 -9978 -251 -9925
rect -304 -10082 -270 -9978
rect -215 -10246 -181 -8820
rect -126 -9545 -92 -9438
rect -146 -9598 -136 -9545
rect -83 -9598 -73 -9545
rect -146 -9979 -136 -9926
rect -83 -9979 -73 -9926
rect -126 -10081 -92 -9979
rect -37 -10184 -3 -8706
rect 141 -8768 175 -8380
rect 230 -8534 264 -8440
rect 211 -8587 221 -8534
rect 274 -8587 284 -8534
rect 319 -8653 353 -8362
rect 408 -8534 442 -8440
rect 388 -8587 398 -8534
rect 451 -8587 461 -8534
rect 300 -8706 310 -8653
rect 363 -8706 373 -8653
rect 122 -8821 132 -8768
rect 185 -8821 195 -8768
rect 52 -9546 86 -9440
rect 32 -9599 42 -9546
rect 95 -9599 105 -9546
rect 33 -9978 43 -9925
rect 96 -9978 106 -9925
rect 52 -10082 86 -9978
rect 141 -10255 175 -8821
rect 231 -9545 265 -9439
rect 212 -9598 222 -9545
rect 275 -9598 285 -9545
rect 210 -9978 220 -9925
rect 273 -9978 283 -9925
rect 230 -10081 264 -9978
rect 319 -10194 353 -8706
rect 497 -8766 531 -8370
rect 586 -8534 620 -8439
rect 567 -8587 577 -8534
rect 630 -8587 640 -8534
rect 675 -8653 709 -8365
rect 744 -8587 754 -8534
rect 807 -8587 817 -8534
rect 656 -8706 666 -8653
rect 719 -8706 729 -8653
rect 479 -8819 489 -8766
rect 542 -8819 552 -8766
rect 408 -9546 442 -9438
rect 389 -9599 399 -9546
rect 452 -9599 462 -9546
rect 388 -9978 398 -9925
rect 451 -9978 461 -9925
rect 408 -10082 442 -9978
rect 497 -10245 531 -8819
rect 587 -9546 621 -9440
rect 567 -9599 577 -9546
rect 630 -9599 640 -9546
rect 566 -9978 576 -9925
rect 629 -9978 639 -9925
rect 586 -10082 620 -9978
rect 675 -10189 709 -8706
rect 764 -9082 798 -8587
rect 853 -8766 887 -8369
rect 922 -8587 932 -8534
rect 985 -8587 995 -8534
rect 833 -8819 843 -8766
rect 896 -8819 906 -8766
rect 853 -9191 887 -8819
rect 942 -9081 976 -8587
rect 1031 -8653 1065 -8366
rect 1101 -8587 1111 -8534
rect 1164 -8587 1174 -8534
rect 1012 -8706 1022 -8653
rect 1075 -8706 1085 -8653
rect 1031 -10213 1065 -8706
rect 1120 -9081 1154 -8587
rect 1209 -8767 1243 -8364
rect 1279 -8587 1289 -8534
rect 1342 -8587 1352 -8534
rect 1191 -8820 1201 -8767
rect 1254 -8820 1264 -8767
rect 1209 -10239 1243 -8820
rect 1298 -9081 1332 -8587
rect 1387 -8653 1421 -8365
rect 1456 -8587 1466 -8534
rect 1519 -8587 1529 -8534
rect 1367 -8706 1377 -8653
rect 1430 -8706 1440 -8653
rect 1387 -10213 1421 -8706
rect 1476 -9081 1510 -8587
rect 1565 -8767 1599 -8372
rect 1634 -8587 1644 -8534
rect 1697 -8587 1707 -8534
rect 1546 -8820 1556 -8767
rect 1609 -8820 1619 -8767
rect 1565 -10247 1599 -8820
rect 1654 -9081 1688 -8587
rect 1743 -8653 1777 -8363
rect 1832 -8534 1866 -8439
rect 1812 -8587 1822 -8534
rect 1875 -8587 1885 -8534
rect 1723 -8706 1733 -8653
rect 1786 -8706 1796 -8653
rect 1743 -10181 1777 -8706
rect 1921 -8767 1955 -8372
rect 2010 -8534 2044 -8439
rect 1990 -8587 2000 -8534
rect 2053 -8587 2063 -8534
rect 2099 -8653 2133 -8368
rect 2188 -8534 2222 -8439
rect 2168 -8587 2178 -8534
rect 2231 -8587 2241 -8534
rect 2080 -8706 2090 -8653
rect 2143 -8706 2153 -8653
rect 1901 -8820 1911 -8767
rect 1964 -8820 1974 -8767
rect 1832 -10082 1866 -9426
rect 1921 -10247 1955 -8820
rect 2010 -10082 2044 -9426
rect 2099 -10209 2133 -8706
rect 2277 -8767 2311 -8372
rect 2367 -8534 2401 -8439
rect 2347 -8587 2357 -8534
rect 2410 -8587 2420 -8534
rect 2455 -8653 2489 -8370
rect 2544 -8534 2578 -8439
rect 2524 -8587 2534 -8534
rect 2587 -8587 2597 -8534
rect 2436 -8706 2446 -8653
rect 2499 -8706 2509 -8653
rect 2257 -8820 2267 -8767
rect 2320 -8820 2330 -8767
rect 2188 -9547 2222 -9426
rect 2168 -9600 2178 -9547
rect 2231 -9600 2241 -9547
rect 2188 -10082 2222 -9600
rect 2277 -10247 2311 -8820
rect 2366 -9546 2400 -9440
rect 2347 -9599 2357 -9546
rect 2410 -9599 2420 -9546
rect 2346 -9978 2356 -9925
rect 2409 -9978 2419 -9925
rect 2366 -10082 2400 -9978
rect 2455 -10186 2489 -8706
rect 2633 -8767 2667 -8375
rect 2722 -8534 2756 -8440
rect 2702 -8587 2712 -8534
rect 2765 -8587 2775 -8534
rect 2811 -8653 2845 -8374
rect 2880 -8587 2890 -8534
rect 2943 -8587 2953 -8534
rect 2792 -8706 2802 -8653
rect 2855 -8706 2865 -8653
rect 2614 -8820 2624 -8767
rect 2677 -8820 2687 -8767
rect 2544 -9546 2578 -9441
rect 2524 -9599 2534 -9546
rect 2587 -9599 2597 -9546
rect 2524 -9978 2534 -9925
rect 2587 -9978 2597 -9925
rect 2544 -10081 2578 -9978
rect 2633 -10250 2667 -8820
rect 2722 -9546 2756 -9441
rect 2703 -9599 2713 -9546
rect 2766 -9599 2776 -9546
rect 2702 -9979 2712 -9926
rect 2765 -9979 2775 -9926
rect 2722 -10081 2756 -9979
rect 2811 -10205 2845 -8706
rect 2900 -9082 2934 -8587
rect 2989 -8767 3023 -8376
rect 3058 -8587 3068 -8534
rect 3121 -8587 3131 -8534
rect 2970 -8820 2980 -8767
rect 3033 -8820 3043 -8767
rect 2881 -9978 2891 -9925
rect 2944 -9978 2954 -9925
rect 2900 -10080 2934 -9978
rect 2989 -10251 3023 -8820
rect 3078 -9082 3112 -8587
rect 3167 -8653 3201 -8362
rect 3236 -8587 3246 -8534
rect 3299 -8587 3309 -8534
rect 3148 -8706 3158 -8653
rect 3211 -8706 3221 -8653
rect 3059 -9978 3069 -9925
rect 3122 -9978 3132 -9925
rect 3078 -10080 3112 -9978
rect 3167 -10176 3201 -8706
rect 3256 -9081 3290 -8587
rect 3345 -8767 3379 -8374
rect 3414 -8587 3424 -8534
rect 3477 -8587 3487 -8534
rect 3326 -8820 3336 -8767
rect 3389 -8820 3399 -8767
rect 3256 -9925 3290 -9443
rect 3236 -9978 3246 -9925
rect 3299 -9978 3309 -9925
rect 3256 -10081 3290 -9978
rect 3345 -10249 3379 -8820
rect 3434 -9082 3468 -8587
rect 3523 -8653 3557 -8365
rect 3592 -8587 3602 -8534
rect 3655 -8587 3665 -8534
rect 3503 -8706 3513 -8653
rect 3566 -8706 3576 -8653
rect 3523 -10190 3557 -8706
rect 3612 -9082 3646 -8587
rect 3701 -8767 3735 -8376
rect 3879 -8440 3913 -8365
rect 4056 -8440 4090 -8360
rect 3879 -8474 4090 -8440
rect 3771 -8587 3781 -8534
rect 3834 -8587 3844 -8534
rect 3682 -8820 3692 -8767
rect 3745 -8820 3755 -8767
rect 3701 -10251 3735 -8820
rect 3790 -9081 3824 -8587
rect 3879 -8653 3913 -8474
rect 3859 -8706 3869 -8653
rect 3922 -8706 3932 -8653
rect 3879 -9439 3913 -8706
rect 4056 -9439 4090 -9361
rect 3879 -9473 4090 -9439
rect 3879 -10047 3913 -9473
rect 4208 -9546 4261 -7976
rect 4771 -9262 4823 -7907
rect 4771 -9314 4824 -9262
rect 4761 -9367 4771 -9314
rect 4824 -9367 4834 -9314
rect 4198 -9599 4208 -9546
rect 4261 -9599 4271 -9546
rect 3879 -10081 4092 -10047
rect 3879 -10205 3913 -10081
rect 4058 -10174 4092 -10081
rect -1837 -10961 -1827 -10908
rect -1774 -10961 -1764 -10908
rect -1480 -10961 -1470 -10908
rect -1417 -10961 -1407 -10908
rect -2172 -11439 -2138 -11345
rect -1995 -11439 -1961 -11189
rect -2172 -11473 -1961 -11439
rect -1995 -11637 -1961 -11473
rect -2014 -11690 -2004 -11637
rect -1951 -11690 -1941 -11637
rect -1995 -12047 -1961 -11690
rect -1905 -11919 -1871 -11445
rect -1925 -11972 -1915 -11919
rect -1862 -11972 -1852 -11919
rect -2176 -12081 -1961 -12047
rect -2176 -12171 -2142 -12081
rect -1995 -12542 -1961 -12081
rect -1905 -12083 -1871 -11972
rect -2015 -12595 -2005 -12542
rect -1952 -12595 -1942 -12542
rect -1995 -13046 -1961 -12595
rect -2174 -13080 -1961 -13046
rect -1906 -13077 -1872 -12439
rect -2174 -13165 -2140 -13080
rect -1995 -13200 -1961 -13080
rect -1818 -13220 -1784 -10961
rect -1728 -11919 -1694 -11447
rect -1639 -11528 -1605 -11374
rect -1659 -11581 -1649 -11528
rect -1596 -11581 -1586 -11528
rect -1549 -11919 -1515 -11447
rect -1748 -11972 -1738 -11919
rect -1685 -11972 -1675 -11919
rect -1569 -11972 -1559 -11919
rect -1506 -11972 -1496 -11919
rect -1728 -12081 -1694 -11972
rect -1549 -12081 -1515 -11972
rect -1728 -13080 -1694 -12442
rect -1639 -12542 -1605 -12386
rect -1659 -12595 -1649 -12542
rect -1596 -12595 -1586 -12542
rect -1549 -13079 -1515 -12441
rect -1461 -13228 -1427 -10961
rect -1372 -11081 -1338 -10438
rect -1193 -11081 -1159 -10432
rect -1124 -10961 -1114 -10908
rect -1061 -10961 -1051 -10908
rect -1372 -11919 -1338 -11448
rect -1283 -11526 -1249 -11373
rect -1284 -11528 -1249 -11526
rect -1303 -11581 -1293 -11528
rect -1240 -11581 -1230 -11528
rect -1391 -11972 -1381 -11919
rect -1328 -11972 -1318 -11919
rect -1372 -12080 -1338 -11972
rect -1372 -13080 -1338 -12442
rect -1284 -12654 -1250 -11581
rect -1194 -11919 -1160 -11448
rect -1213 -11972 -1203 -11919
rect -1150 -11972 -1140 -11919
rect -1194 -12081 -1160 -11972
rect -1304 -12707 -1294 -12654
rect -1241 -12707 -1231 -12654
rect -1194 -13079 -1160 -12441
rect -1105 -13202 -1071 -10961
rect -1016 -11081 -982 -10432
rect -838 -11082 -804 -10433
rect -768 -10961 -758 -10908
rect -705 -10961 -695 -10908
rect -1016 -11919 -982 -11448
rect -927 -11528 -893 -11367
rect -947 -11581 -937 -11528
rect -884 -11581 -874 -11528
rect -838 -11919 -804 -11448
rect -1035 -11972 -1025 -11919
rect -972 -11972 -962 -11919
rect -858 -11972 -848 -11919
rect -795 -11972 -785 -11919
rect -1016 -12080 -982 -11972
rect -838 -12081 -804 -11972
rect -1016 -13080 -982 -12442
rect -927 -12783 -893 -12389
rect -947 -12836 -937 -12783
rect -884 -12836 -874 -12783
rect -927 -13174 -893 -12836
rect -838 -13079 -804 -12441
rect -749 -13222 -715 -10961
rect -659 -11081 -625 -10432
rect -482 -11081 -448 -10432
rect 853 -10438 887 -10368
rect 941 -10438 975 -10431
rect 1031 -10438 1065 -10360
rect 759 -10472 1159 -10438
rect 941 -10908 975 -10472
rect -412 -10961 -402 -10908
rect -349 -10961 -339 -10908
rect -56 -10961 -46 -10908
rect 7 -10961 17 -10908
rect 299 -10961 309 -10908
rect 362 -10961 372 -10908
rect 655 -10961 665 -10908
rect 718 -10961 728 -10908
rect 921 -10961 931 -10908
rect 984 -10961 994 -10908
rect 1189 -10961 1199 -10908
rect 1252 -10961 1262 -10908
rect -660 -11919 -626 -11448
rect -571 -11637 -537 -11388
rect -590 -11690 -580 -11637
rect -527 -11690 -517 -11637
rect -482 -11919 -448 -11448
rect -680 -11972 -670 -11919
rect -617 -11972 -607 -11919
rect -502 -11972 -492 -11919
rect -439 -11972 -429 -11919
rect -660 -12081 -626 -11972
rect -482 -12081 -448 -11972
rect -660 -13081 -626 -12443
rect -571 -12653 -537 -12387
rect -592 -12706 -582 -12653
rect -529 -12706 -519 -12653
rect -482 -13081 -448 -12443
rect -393 -13207 -359 -10961
rect -304 -11919 -270 -11448
rect -215 -11757 -181 -11385
rect -234 -11810 -224 -11757
rect -171 -11810 -161 -11757
rect -324 -11972 -314 -11919
rect -261 -11972 -251 -11919
rect -304 -12080 -270 -11972
rect -304 -13082 -270 -12444
rect -215 -12783 -181 -11810
rect -126 -11919 -92 -11448
rect -146 -11972 -136 -11919
rect -83 -11972 -73 -11919
rect -126 -12079 -92 -11972
rect -234 -12836 -224 -12783
rect -171 -12836 -161 -12783
rect -126 -13081 -92 -12443
rect -36 -13199 -2 -10961
rect 52 -11919 86 -11448
rect 141 -11757 175 -11387
rect 121 -11810 131 -11757
rect 184 -11810 194 -11757
rect 141 -11811 175 -11810
rect 230 -11919 264 -11448
rect 32 -11972 42 -11919
rect 95 -11972 105 -11919
rect 210 -11972 220 -11919
rect 273 -11972 283 -11919
rect 52 -12081 86 -11972
rect 230 -12080 264 -11972
rect 52 -13080 86 -12442
rect 141 -12653 175 -12384
rect 120 -12706 130 -12653
rect 183 -12706 193 -12653
rect -1995 -13545 -1961 -13383
rect -2014 -13598 -2004 -13545
rect -1951 -13598 -1941 -13545
rect -1905 -14082 -1871 -13444
rect -1728 -14081 -1694 -13443
rect -1638 -13672 -1604 -13385
rect -1658 -13725 -1648 -13672
rect -1595 -13725 -1585 -13672
rect -1550 -14082 -1516 -13444
rect -1282 -13672 -1248 -13383
rect -927 -13672 -893 -13387
rect -571 -13545 -537 -13385
rect -591 -13598 -581 -13545
rect -528 -13598 -518 -13545
rect -1301 -13725 -1291 -13672
rect -1238 -13725 -1228 -13672
rect -947 -13725 -937 -13672
rect -884 -13725 -874 -13672
rect -927 -13726 -893 -13725
rect -304 -14081 -270 -13437
rect -216 -13794 -182 -13386
rect -235 -13847 -225 -13794
rect -172 -13847 -162 -13794
rect -125 -14082 -91 -13438
rect 52 -14081 86 -13437
rect 141 -13794 175 -12706
rect 230 -13080 264 -12442
rect 319 -13207 353 -10961
rect 408 -11919 442 -11448
rect 497 -11757 531 -11380
rect 477 -11810 487 -11757
rect 540 -11810 550 -11757
rect 389 -11972 399 -11919
rect 452 -11972 462 -11919
rect 408 -12081 442 -11972
rect 408 -13082 442 -12444
rect 496 -12784 530 -11810
rect 586 -11919 620 -11448
rect 567 -11972 577 -11919
rect 630 -11972 640 -11919
rect 586 -12081 620 -11972
rect 476 -12837 486 -12784
rect 539 -12837 549 -12784
rect 587 -13082 621 -12444
rect 675 -13231 709 -10961
rect 941 -11080 975 -10961
rect 853 -11438 887 -11362
rect 942 -11438 976 -11432
rect 1031 -11438 1065 -11357
rect 757 -11472 1159 -11438
rect 764 -12081 798 -12032
rect 942 -12081 976 -11472
rect 1120 -12080 1154 -12032
rect 852 -12438 886 -12353
rect 942 -12438 976 -12432
rect 1031 -12438 1065 -12377
rect 759 -12472 1160 -12438
rect 942 -13048 976 -12472
rect 761 -13082 1160 -13048
rect 852 -13154 886 -13082
rect 1032 -13165 1066 -13082
rect 1209 -13212 1243 -10961
rect 1299 -11081 1333 -10432
rect 1477 -11081 1511 -10432
rect 1546 -10961 1556 -10908
rect 1609 -10961 1619 -10908
rect 1298 -11919 1332 -11448
rect 1387 -11528 1421 -11389
rect 1367 -11581 1377 -11528
rect 1430 -11581 1440 -11528
rect 1477 -11919 1511 -11448
rect 1278 -11972 1288 -11919
rect 1341 -11972 1351 -11919
rect 1458 -11972 1468 -11919
rect 1521 -11972 1531 -11919
rect 1298 -12080 1332 -11972
rect 1477 -12081 1511 -11972
rect 1299 -13081 1333 -12443
rect 1388 -12783 1422 -12389
rect 1368 -12836 1378 -12783
rect 1431 -12836 1441 -12783
rect 1388 -13187 1422 -12836
rect 1476 -13081 1510 -12443
rect 1566 -13217 1600 -10961
rect 1653 -11080 1687 -10431
rect 1832 -11082 1866 -10433
rect 1903 -10961 1913 -10908
rect 1966 -10961 1976 -10908
rect 1654 -11920 1688 -11448
rect 1743 -11528 1777 -11386
rect 1723 -11581 1733 -11528
rect 1786 -11581 1796 -11528
rect 1634 -11973 1644 -11920
rect 1697 -11973 1707 -11920
rect 1654 -12080 1688 -11973
rect 1655 -13082 1689 -12444
rect 1744 -12654 1778 -11581
rect 1832 -11919 1866 -11448
rect 1813 -11972 1823 -11919
rect 1876 -11972 1886 -11919
rect 1832 -12081 1866 -11972
rect 1725 -12707 1735 -12654
rect 1788 -12707 1798 -12654
rect 1833 -13081 1867 -12443
rect 1922 -13187 1956 -10961
rect 2010 -11081 2044 -10432
rect 2188 -11081 2222 -10432
rect 2258 -10961 2268 -10908
rect 2321 -10961 2331 -10908
rect 2613 -10961 2623 -10908
rect 2676 -10961 2686 -10908
rect 2970 -10961 2980 -10908
rect 3033 -10961 3043 -10908
rect 3325 -10961 3335 -10908
rect 3388 -10961 3398 -10908
rect 2010 -11919 2044 -11448
rect 2099 -11528 2133 -11380
rect 2079 -11581 2089 -11528
rect 2142 -11581 2152 -11528
rect 2188 -11919 2222 -11448
rect 1990 -11972 2000 -11919
rect 2053 -11972 2063 -11919
rect 2168 -11972 2178 -11919
rect 2231 -11972 2241 -11919
rect 2010 -12079 2044 -11972
rect 2188 -12079 2222 -11972
rect 2009 -13079 2043 -12441
rect 2098 -12782 2132 -12375
rect 2078 -12835 2088 -12782
rect 2141 -12835 2151 -12782
rect 2098 -13193 2132 -12835
rect 2188 -13079 2222 -12441
rect 2277 -13199 2311 -10961
rect 2366 -11919 2400 -11448
rect 2456 -11637 2490 -11386
rect 2436 -11690 2446 -11637
rect 2499 -11690 2509 -11637
rect 2544 -11919 2578 -11448
rect 2347 -11972 2357 -11919
rect 2410 -11972 2420 -11919
rect 2524 -11972 2534 -11919
rect 2587 -11972 2597 -11919
rect 2366 -12083 2400 -11972
rect 2544 -12081 2578 -11972
rect 2366 -13082 2400 -12444
rect 2455 -12653 2489 -12385
rect 2435 -12706 2445 -12653
rect 2498 -12706 2508 -12653
rect 2544 -13082 2578 -12444
rect 2633 -13204 2667 -10961
rect 2722 -11919 2756 -11448
rect 2810 -11757 2844 -11387
rect 2790 -11810 2800 -11757
rect 2853 -11810 2863 -11757
rect 2703 -11972 2713 -11919
rect 2766 -11972 2776 -11919
rect 2722 -12080 2756 -11972
rect 2722 -13079 2756 -12441
rect 2811 -12782 2845 -11810
rect 2900 -11919 2934 -11448
rect 2880 -11972 2890 -11919
rect 2943 -11972 2953 -11919
rect 2900 -12080 2934 -11972
rect 2791 -12835 2801 -12782
rect 2854 -12835 2864 -12782
rect 2900 -13082 2934 -12444
rect 2989 -13212 3023 -10961
rect 3078 -11919 3112 -11448
rect 3166 -11757 3200 -11384
rect 3147 -11810 3157 -11757
rect 3210 -11810 3220 -11757
rect 3256 -11919 3290 -11448
rect 3058 -11972 3068 -11919
rect 3121 -11972 3131 -11919
rect 3237 -11972 3247 -11919
rect 3300 -11972 3310 -11919
rect 3078 -12081 3112 -11972
rect 3256 -12080 3290 -11972
rect 3078 -13081 3112 -12443
rect 3167 -12650 3201 -12387
rect 3166 -12652 3201 -12650
rect 3148 -12705 3158 -12652
rect 3211 -12705 3221 -12652
rect 123 -13847 133 -13794
rect 186 -13847 196 -13794
rect 230 -14081 264 -13437
rect 408 -14081 442 -13437
rect 496 -13795 530 -13385
rect 477 -13848 487 -13795
rect 540 -13848 550 -13795
rect 587 -14081 621 -13437
rect 942 -14048 976 -13430
rect 1388 -13672 1422 -13380
rect 1743 -13672 1777 -13382
rect 2100 -13672 2134 -13382
rect 1369 -13725 1379 -13672
rect 1432 -13725 1442 -13672
rect 1722 -13725 1732 -13672
rect 1785 -13725 1795 -13672
rect 2081 -13725 2091 -13672
rect 2144 -13725 2154 -13672
rect 762 -14082 1159 -14048
rect 2366 -14081 2400 -13432
rect 2455 -13545 2489 -13388
rect 2436 -13598 2446 -13545
rect 2499 -13598 2509 -13545
rect 2544 -14081 2578 -13432
rect 2723 -14082 2757 -13433
rect 2812 -13794 2846 -13379
rect 2792 -13847 2802 -13794
rect 2855 -13847 2865 -13794
rect 2901 -14081 2935 -13432
rect 3078 -14082 3112 -13433
rect 3166 -13795 3200 -12705
rect 3256 -13082 3290 -12444
rect 3345 -13223 3379 -10961
rect 3434 -11082 3468 -10433
rect 3613 -11082 3647 -10433
rect 3682 -10961 3692 -10908
rect 3745 -10961 3755 -10908
rect 3434 -11919 3468 -11448
rect 3522 -11757 3556 -11369
rect 3503 -11810 3513 -11757
rect 3566 -11810 3576 -11757
rect 3612 -11919 3646 -11448
rect 3415 -11972 3425 -11919
rect 3478 -11972 3488 -11919
rect 3593 -11972 3603 -11919
rect 3656 -11972 3666 -11919
rect 3434 -12081 3468 -11972
rect 3612 -12080 3646 -11972
rect 3434 -13080 3468 -12442
rect 3524 -12542 3558 -12386
rect 3504 -12595 3514 -12542
rect 3567 -12595 3577 -12542
rect 3613 -13080 3647 -12442
rect 3701 -13213 3735 -10961
rect 3791 -11081 3825 -10432
rect 3881 -11437 3915 -11232
rect 4056 -11437 4090 -11365
rect 3790 -11919 3824 -11448
rect 3881 -11471 4090 -11437
rect 3881 -11638 3915 -11471
rect 3861 -11691 3871 -11638
rect 3924 -11691 3934 -11638
rect 3771 -11972 3781 -11919
rect 3834 -11972 3844 -11919
rect 3790 -12079 3824 -11972
rect 3881 -12436 3915 -11691
rect 4058 -12436 4092 -12363
rect 3790 -13080 3824 -12442
rect 3881 -12470 4092 -12436
rect 3881 -12542 3915 -12470
rect 3861 -12595 3871 -12542
rect 3924 -12595 3934 -12542
rect 3881 -13047 3915 -12595
rect 3881 -13081 4090 -13047
rect 3881 -13192 3915 -13081
rect 4056 -13165 4090 -13081
rect 3147 -13848 3157 -13795
rect 3210 -13848 3220 -13795
rect 3257 -14080 3291 -13431
rect 3523 -13794 3557 -13336
rect 3879 -13545 3913 -13387
rect 3860 -13598 3870 -13545
rect 3923 -13598 3933 -13545
rect 3502 -13847 3512 -13794
rect 3565 -13847 3575 -13794
rect 3523 -13848 3557 -13847
rect 853 -14160 887 -14082
rect 1032 -14164 1066 -14082
rect -2173 -14441 -2139 -14361
rect -1995 -14441 -1961 -14228
rect -2173 -14475 -1961 -14441
rect -2325 -14596 -2315 -14543
rect -2262 -14596 -2252 -14543
rect -1995 -15045 -1961 -14475
rect -2176 -15079 -1961 -15045
rect -2176 -15163 -2142 -15079
rect -2457 -15874 -2447 -15821
rect -2394 -15874 -2384 -15821
rect -1995 -15822 -1961 -15079
rect -2015 -15875 -2005 -15822
rect -1952 -15875 -1942 -15822
rect -1995 -16050 -1961 -15875
rect -1906 -15933 -1872 -15441
rect -1925 -15986 -1915 -15933
rect -1862 -15986 -1852 -15933
rect -2173 -16084 -1961 -16050
rect -2173 -16156 -2139 -16084
rect -1995 -16132 -1961 -16084
rect -3945 -16347 -3935 -16295
rect -3883 -16347 -3873 -16295
rect -6028 -16886 -5994 -16750
rect -5939 -16886 -5905 -16794
rect -5850 -16886 -5816 -16750
rect -5672 -16886 -5638 -16750
rect -6028 -16920 -5816 -16886
rect -5850 -17007 -5816 -16920
rect -5692 -16939 -5682 -16886
rect -5629 -16939 -5619 -16886
rect -6169 -17060 -6159 -17007
rect -6106 -17060 -6096 -17007
rect -5869 -17060 -5859 -17007
rect -5806 -17060 -5796 -17007
rect -5494 -17118 -5460 -16751
rect -5316 -16886 -5282 -16750
rect -5336 -16939 -5326 -16886
rect -5273 -16939 -5263 -16886
rect -5138 -17007 -5104 -16751
rect -4960 -16886 -4926 -16751
rect -4980 -16939 -4970 -16886
rect -4917 -16939 -4907 -16886
rect -5158 -17060 -5148 -17007
rect -5095 -17060 -5085 -17007
rect -5514 -17171 -5504 -17118
rect -5451 -17171 -5441 -17118
rect -7605 -17251 -7329 -17250
rect -4970 -17251 -4917 -16939
rect -4782 -17118 -4748 -16751
rect -4604 -16886 -4570 -16751
rect -4624 -16939 -4614 -16886
rect -4561 -16939 -4551 -16886
rect -4426 -17007 -4392 -16750
rect -4248 -16886 -4214 -16750
rect -4159 -16886 -4125 -16794
rect -4070 -16886 -4036 -16750
rect -4268 -16939 -4258 -16886
rect -4205 -16939 -4036 -16886
rect -4447 -17060 -4437 -17007
rect -4384 -17060 -4374 -17007
rect -3935 -17118 -3883 -16347
rect -1906 -16542 -1872 -16438
rect -1927 -16595 -1917 -16542
rect -1864 -16595 -1854 -16542
rect -1817 -16665 -1783 -14309
rect -1728 -15933 -1694 -15438
rect -1639 -15822 -1605 -14231
rect -1659 -15875 -1649 -15822
rect -1596 -15875 -1586 -15822
rect -1748 -15986 -1738 -15933
rect -1685 -15986 -1675 -15933
rect -1639 -16135 -1605 -15875
rect -1550 -15933 -1516 -15438
rect -1570 -15986 -1560 -15933
rect -1507 -15986 -1497 -15933
rect -1728 -16542 -1694 -16440
rect -1550 -16541 -1516 -16439
rect -1748 -16595 -1738 -16542
rect -1685 -16595 -1675 -16542
rect -1571 -16594 -1561 -16541
rect -1508 -16594 -1498 -16541
rect -1736 -16665 -1528 -16655
rect -1837 -16718 -1827 -16665
rect -1774 -16718 -1764 -16665
rect -1736 -16718 -1720 -16665
rect -1548 -16718 -1528 -16665
rect -1461 -16666 -1427 -14309
rect -1371 -14543 -1337 -14438
rect -1391 -14596 -1381 -14543
rect -1328 -14596 -1318 -14543
rect -1371 -15076 -1337 -14596
rect -1372 -15933 -1338 -15440
rect -1283 -15822 -1249 -14234
rect -1194 -14543 -1160 -14438
rect -1214 -14596 -1204 -14543
rect -1151 -14596 -1141 -14543
rect -1303 -15875 -1293 -15822
rect -1240 -15875 -1230 -15822
rect -1392 -15986 -1382 -15933
rect -1329 -15986 -1319 -15933
rect -1283 -16138 -1249 -15875
rect -1194 -15933 -1160 -15438
rect -1214 -15986 -1204 -15933
rect -1151 -15986 -1141 -15933
rect -1372 -16543 -1338 -16440
rect -1194 -16542 -1160 -16440
rect -1391 -16596 -1381 -16543
rect -1328 -16596 -1318 -16543
rect -1214 -16595 -1204 -16542
rect -1151 -16595 -1141 -16542
rect -1104 -16665 -1070 -14312
rect -1016 -14543 -982 -14439
rect -1036 -14596 -1026 -14543
rect -973 -14596 -963 -14543
rect -1015 -15933 -981 -15439
rect -927 -15822 -893 -14231
rect -838 -14543 -804 -14438
rect -858 -14596 -848 -14543
rect -795 -14596 -785 -14543
rect -857 -14979 -847 -14926
rect -794 -14979 -784 -14926
rect -838 -15081 -804 -14979
rect -947 -15875 -937 -15822
rect -884 -15875 -874 -15822
rect -1035 -15986 -1025 -15933
rect -972 -15986 -962 -15933
rect -927 -16135 -893 -15875
rect -857 -15986 -847 -15933
rect -794 -15986 -784 -15933
rect -838 -16080 -804 -15986
rect -1016 -16542 -982 -16439
rect -1036 -16595 -1026 -16542
rect -973 -16595 -963 -16542
rect -749 -16664 -715 -14310
rect -659 -14543 -625 -14440
rect -679 -14596 -669 -14543
rect -616 -14596 -606 -14543
rect -679 -14979 -669 -14926
rect -616 -14979 -606 -14926
rect -660 -15081 -626 -14979
rect -571 -15822 -537 -14231
rect -482 -14543 -448 -14439
rect -501 -14596 -491 -14543
rect -438 -14596 -428 -14543
rect -501 -14979 -491 -14926
rect -438 -14979 -428 -14926
rect -481 -15081 -447 -14979
rect -591 -15875 -581 -15822
rect -528 -15875 -518 -15822
rect -680 -15986 -670 -15933
rect -617 -15986 -607 -15933
rect -660 -16082 -626 -15986
rect -571 -16135 -537 -15875
rect -501 -15986 -491 -15933
rect -438 -15986 -428 -15933
rect -482 -16081 -448 -15986
rect -4802 -17171 -4792 -17118
rect -4739 -17171 -4729 -17118
rect -3945 -17170 -3935 -17118
rect -3883 -17170 -3873 -17118
rect -1736 -17251 -1528 -16718
rect -1481 -16719 -1471 -16666
rect -1418 -16719 -1408 -16666
rect -1124 -16718 -1114 -16665
rect -1061 -16718 -1051 -16665
rect -769 -16717 -759 -16664
rect -706 -16717 -696 -16664
rect -658 -16665 -450 -16656
rect -393 -16665 -359 -14306
rect -304 -14927 -270 -14437
rect -324 -14980 -314 -14927
rect -261 -14980 -251 -14927
rect -304 -15081 -270 -14980
rect -215 -15822 -181 -14230
rect -126 -14926 -92 -14440
rect -147 -14979 -137 -14926
rect -84 -14979 -74 -14926
rect -126 -15081 -92 -14979
rect -235 -15875 -225 -15822
rect -172 -15875 -162 -15822
rect -323 -15986 -313 -15933
rect -260 -15986 -250 -15933
rect -304 -16080 -270 -15986
rect -215 -16134 -181 -15875
rect -146 -15986 -136 -15933
rect -83 -15986 -73 -15933
rect -126 -16080 -92 -15986
rect -37 -16665 -3 -14312
rect 52 -14926 86 -14445
rect 33 -14979 43 -14926
rect 96 -14979 106 -14926
rect 52 -15081 86 -14979
rect 141 -15821 175 -14231
rect 122 -15874 132 -15821
rect 185 -15874 195 -15821
rect 33 -15986 43 -15933
rect 96 -15986 106 -15933
rect 52 -16080 86 -15986
rect 141 -16135 175 -15874
rect 230 -15933 264 -15439
rect 211 -15986 221 -15933
rect 274 -15986 284 -15933
rect 230 -16542 264 -16438
rect 210 -16595 220 -16542
rect 273 -16595 283 -16542
rect -658 -16718 -646 -16665
rect -471 -16718 -450 -16665
rect -413 -16718 -403 -16665
rect -350 -16718 -340 -16665
rect -57 -16718 -47 -16665
rect 6 -16718 16 -16665
rect 319 -16666 353 -14307
rect 408 -15933 442 -15439
rect 497 -15822 531 -14231
rect 477 -15875 487 -15822
rect 540 -15875 550 -15822
rect 388 -15986 398 -15933
rect 451 -15986 461 -15933
rect 497 -16135 531 -15875
rect 585 -15933 619 -15439
rect 565 -15986 575 -15933
rect 628 -15986 638 -15933
rect 408 -16542 442 -16439
rect 586 -16542 620 -16439
rect 387 -16595 397 -16542
rect 450 -16595 460 -16542
rect 566 -16595 576 -16542
rect 629 -16595 639 -16542
rect 408 -16665 616 -16649
rect 675 -16665 709 -14307
rect 764 -15933 798 -15438
rect 853 -15822 887 -15340
rect 833 -15875 843 -15822
rect 896 -15875 906 -15822
rect 745 -15986 755 -15933
rect 808 -15986 818 -15933
rect 853 -16136 887 -15875
rect 941 -15933 975 -15439
rect 921 -15986 931 -15933
rect 984 -15986 994 -15933
rect 765 -16542 799 -16438
rect 943 -16542 977 -16439
rect 745 -16595 755 -16542
rect 808 -16595 818 -16542
rect 923 -16595 933 -16542
rect 986 -16595 996 -16542
rect 1031 -16665 1065 -14308
rect 1120 -15933 1154 -15440
rect 1209 -15822 1243 -14231
rect 1298 -14543 1332 -14439
rect 1278 -14596 1288 -14543
rect 1341 -14596 1351 -14543
rect 1279 -14980 1289 -14927
rect 1342 -14980 1352 -14927
rect 1298 -15081 1332 -14980
rect 1191 -15875 1201 -15822
rect 1254 -15875 1264 -15822
rect 1100 -15986 1110 -15933
rect 1163 -15986 1173 -15933
rect 1209 -16135 1243 -15875
rect 1279 -15986 1289 -15933
rect 1342 -15986 1352 -15933
rect 1298 -16081 1332 -15986
rect 1120 -16542 1154 -16439
rect 1101 -16595 1111 -16542
rect 1164 -16595 1174 -16542
rect 1387 -16665 1421 -14307
rect 1477 -14543 1511 -14439
rect 1456 -14596 1466 -14543
rect 1519 -14596 1529 -14543
rect 1457 -14979 1467 -14926
rect 1520 -14979 1530 -14926
rect 1476 -15081 1510 -14979
rect 1565 -15822 1599 -14231
rect 1654 -14543 1688 -14438
rect 1634 -14596 1644 -14543
rect 1697 -14596 1707 -14543
rect 1634 -14979 1644 -14926
rect 1697 -14979 1707 -14926
rect 1654 -15082 1688 -14979
rect 1545 -15875 1555 -15822
rect 1608 -15875 1618 -15822
rect 1456 -15986 1466 -15933
rect 1519 -15986 1529 -15933
rect 1476 -16082 1510 -15986
rect 1565 -16135 1599 -15875
rect 1633 -15986 1643 -15933
rect 1696 -15986 1706 -15933
rect 1653 -16081 1687 -15986
rect 1488 -16665 1696 -16658
rect 1744 -16665 1778 -14312
rect 1832 -14542 1866 -14438
rect 1813 -14595 1823 -14542
rect 1876 -14595 1886 -14542
rect 1812 -14979 1822 -14926
rect 1875 -14979 1885 -14926
rect 1833 -15081 1867 -14979
rect 1921 -15822 1955 -14231
rect 2010 -14543 2044 -14438
rect 1990 -14596 2000 -14543
rect 2053 -14596 2063 -14543
rect 1989 -14979 1999 -14926
rect 2052 -14979 2062 -14926
rect 2010 -15082 2044 -14979
rect 1900 -15875 1910 -15822
rect 1963 -15875 1973 -15822
rect 1812 -15986 1822 -15933
rect 1875 -15986 1885 -15933
rect 1832 -16080 1866 -15986
rect 1921 -16135 1955 -15875
rect 1990 -15986 2000 -15933
rect 2053 -15986 2063 -15933
rect 2010 -16081 2044 -15986
rect 2100 -16664 2134 -14313
rect 2188 -14543 2222 -14439
rect 2168 -14596 2178 -14543
rect 2231 -14596 2241 -14543
rect 2170 -14979 2180 -14926
rect 2233 -14979 2243 -14926
rect 2189 -15081 2223 -14979
rect 2277 -15822 2311 -14231
rect 2257 -15875 2267 -15822
rect 2320 -15875 2330 -15822
rect 2169 -15986 2179 -15933
rect 2232 -15986 2242 -15933
rect 2189 -16081 2223 -15986
rect 2277 -16135 2311 -15875
rect 2366 -15933 2400 -15440
rect 2346 -15986 2356 -15933
rect 2409 -15986 2419 -15933
rect 2366 -16542 2400 -16439
rect 2346 -16595 2356 -16542
rect 2409 -16595 2419 -16542
rect -658 -17251 -450 -16718
rect 299 -16719 309 -16666
rect 362 -16719 372 -16666
rect 408 -16718 426 -16665
rect 595 -16718 616 -16665
rect 655 -16718 665 -16665
rect 718 -16718 728 -16665
rect 1011 -16718 1021 -16665
rect 1074 -16718 1084 -16665
rect 1367 -16718 1377 -16665
rect 1430 -16718 1440 -16665
rect 1488 -16718 1501 -16665
rect 1671 -16718 1696 -16665
rect 1725 -16718 1735 -16665
rect 1788 -16718 1798 -16665
rect 2080 -16717 2090 -16664
rect 2143 -16717 2153 -16664
rect 2455 -16665 2489 -14311
rect 2544 -15933 2578 -15440
rect 2633 -15822 2667 -14232
rect 2614 -15875 2624 -15822
rect 2677 -15875 2687 -15822
rect 2524 -15986 2534 -15933
rect 2587 -15986 2597 -15933
rect 2633 -16136 2667 -15875
rect 2722 -15933 2756 -15440
rect 2702 -15986 2712 -15933
rect 2765 -15986 2775 -15933
rect 2544 -16542 2578 -16439
rect 2722 -16541 2756 -16441
rect 2524 -16595 2534 -16542
rect 2587 -16595 2597 -16542
rect 2703 -16594 2713 -16541
rect 2766 -16594 2776 -16541
rect 2547 -16665 2755 -16653
rect 2811 -16665 2845 -14310
rect 2900 -15933 2934 -15439
rect 2989 -15822 3023 -14231
rect 2969 -15875 2979 -15822
rect 3032 -15875 3042 -15822
rect 2881 -15986 2891 -15933
rect 2944 -15986 2954 -15933
rect 2989 -16135 3023 -15875
rect 3078 -15933 3112 -15438
rect 3058 -15986 3068 -15933
rect 3121 -15986 3131 -15933
rect 2901 -16542 2935 -16441
rect 3079 -16542 3113 -16439
rect 2881 -16595 2891 -16542
rect 2944 -16595 2954 -16542
rect 3060 -16595 3070 -16542
rect 3123 -16595 3133 -16542
rect 3167 -16664 3201 -14315
rect 3236 -14597 3246 -14544
rect 3299 -14597 3309 -14544
rect 3256 -15080 3290 -14597
rect 3256 -15933 3290 -15439
rect 3345 -15822 3379 -14231
rect 3434 -14543 3468 -14439
rect 3414 -14596 3424 -14543
rect 3477 -14596 3487 -14543
rect 3415 -14979 3425 -14926
rect 3478 -14979 3488 -14926
rect 3434 -15081 3468 -14979
rect 3325 -15875 3335 -15822
rect 3388 -15875 3398 -15822
rect 3237 -15986 3247 -15933
rect 3300 -15986 3310 -15933
rect 3345 -16135 3379 -15875
rect 3414 -15986 3424 -15933
rect 3477 -15986 3487 -15933
rect 3434 -16081 3468 -15986
rect 3257 -16542 3291 -16440
rect 3239 -16595 3249 -16542
rect 3302 -16595 3312 -16542
rect 2435 -16718 2445 -16665
rect 2498 -16718 2508 -16665
rect 2547 -16718 2568 -16665
rect 2732 -16718 2755 -16665
rect 2791 -16718 2801 -16665
rect 2854 -16718 2864 -16665
rect 3147 -16717 3157 -16664
rect 3210 -16717 3220 -16664
rect 3524 -16666 3558 -14310
rect 3612 -14543 3646 -14439
rect 3592 -14596 3602 -14543
rect 3655 -14596 3665 -14543
rect 3593 -14979 3603 -14926
rect 3656 -14979 3666 -14926
rect 3612 -15082 3646 -14979
rect 3701 -15822 3735 -14232
rect 3879 -14439 3913 -14307
rect 4057 -14439 4091 -14357
rect 3791 -14543 3825 -14439
rect 3879 -14473 4091 -14439
rect 3771 -14596 3781 -14543
rect 3834 -14596 3844 -14543
rect 3770 -14979 3780 -14926
rect 3833 -14979 3843 -14926
rect 3790 -15082 3824 -14979
rect 3879 -15047 3913 -14473
rect 4905 -14545 4958 -7905
rect 5037 -13296 5090 -7903
rect 5174 -7908 5184 -7855
rect 5237 -7908 5247 -7855
rect 5327 -7903 5337 -7850
rect 5390 -7903 5400 -7850
rect 5185 -8635 5237 -7908
rect 5175 -8687 5185 -8635
rect 5237 -8687 5247 -8635
rect 5337 -9925 5390 -7903
rect 11647 -8716 11681 -8715
rect 6690 -8760 6815 -8726
rect 6690 -8907 6724 -8760
rect 6781 -8844 6815 -8760
rect 11044 -8769 11054 -8716
rect 11107 -8769 11117 -8716
rect 11335 -8769 11345 -8716
rect 11398 -8769 11408 -8716
rect 11628 -8769 11638 -8716
rect 11691 -8769 11701 -8716
rect 11922 -8769 11932 -8716
rect 11985 -8769 11995 -8716
rect 12212 -8769 12222 -8716
rect 12275 -8769 12285 -8716
rect 9004 -8842 9395 -8808
rect 6513 -9201 6547 -9125
rect 6689 -9201 6723 -8954
rect 6513 -9235 6723 -9201
rect 6779 -9314 6813 -9198
rect 6759 -9367 6769 -9314
rect 6822 -9367 6832 -9314
rect 6669 -9598 6679 -9545
rect 6732 -9598 6742 -9545
rect 5327 -9978 5337 -9925
rect 5390 -9978 5400 -9925
rect 6513 -10099 6547 -10017
rect 6690 -10099 6724 -9598
rect 6779 -9740 6813 -9367
rect 6513 -10133 6724 -10099
rect 6690 -10313 6724 -10133
rect 6670 -10366 6680 -10313
rect 6733 -10366 6743 -10313
rect 6868 -10467 6902 -9042
rect 6957 -9315 6991 -9197
rect 6937 -9368 6947 -9315
rect 7000 -9368 7010 -9315
rect 6957 -9621 6991 -9368
rect 7046 -9621 7080 -9046
rect 7135 -9315 7169 -9198
rect 7116 -9368 7126 -9315
rect 7179 -9368 7189 -9315
rect 6957 -9655 7080 -9621
rect 6957 -9743 6991 -9655
rect 6848 -10520 6858 -10467
rect 6911 -10520 6921 -10467
rect 6510 -11003 6544 -10910
rect 6688 -11003 6722 -10920
rect 6868 -11003 6902 -10520
rect 6958 -10643 6992 -10097
rect 6510 -11037 6902 -11003
rect 6511 -11900 6545 -11823
rect 6688 -11900 6722 -11819
rect 6868 -11900 6902 -11037
rect 6958 -11544 6992 -10995
rect 7046 -11366 7080 -9655
rect 7135 -9744 7169 -9368
rect 7136 -10643 7170 -10097
rect 7224 -10466 7258 -9049
rect 7313 -9313 7347 -9197
rect 7293 -9366 7303 -9313
rect 7356 -9366 7366 -9313
rect 7313 -9743 7347 -9366
rect 7204 -10519 7214 -10466
rect 7267 -10519 7277 -10466
rect 7027 -11419 7037 -11366
rect 7090 -11419 7100 -11366
rect 7046 -11671 7080 -11419
rect 7135 -11543 7169 -10994
rect 6511 -11934 6902 -11900
rect 6868 -12040 6902 -11934
rect 7224 -12040 7258 -10519
rect 7313 -10644 7347 -10098
rect 7313 -11542 7347 -10993
rect 7402 -11366 7436 -9048
rect 7491 -9313 7525 -9198
rect 7472 -9366 7482 -9313
rect 7535 -9366 7545 -9313
rect 7491 -9744 7525 -9366
rect 7492 -10643 7526 -10097
rect 7580 -10466 7614 -9051
rect 7669 -9315 7703 -9198
rect 7649 -9368 7659 -9315
rect 7712 -9368 7722 -9315
rect 7669 -9744 7703 -9368
rect 7561 -10519 7571 -10466
rect 7624 -10519 7634 -10466
rect 7383 -11419 7393 -11366
rect 7446 -11419 7456 -11366
rect 7402 -11673 7436 -11419
rect 7491 -11542 7525 -10993
rect 7580 -12040 7614 -10519
rect 7669 -10644 7703 -10098
rect 7669 -11542 7703 -10993
rect 7758 -11367 7792 -9054
rect 7847 -9314 7881 -9198
rect 7827 -9367 7837 -9314
rect 7890 -9367 7900 -9314
rect 7847 -9744 7881 -9367
rect 7847 -10643 7881 -10097
rect 7936 -10466 7970 -9051
rect 8025 -9315 8059 -9198
rect 8005 -9368 8015 -9315
rect 8068 -9368 8078 -9315
rect 8025 -9744 8059 -9368
rect 7917 -10519 7927 -10466
rect 7980 -10519 7990 -10466
rect 7738 -11420 7748 -11367
rect 7801 -11420 7811 -11367
rect 7758 -11679 7792 -11420
rect 7848 -11542 7882 -10993
rect 7936 -12040 7970 -10519
rect 8025 -10643 8059 -10097
rect 8024 -11543 8058 -10994
rect 8113 -11366 8147 -9056
rect 8203 -9314 8237 -9198
rect 8184 -9367 8194 -9314
rect 8247 -9367 8257 -9314
rect 8203 -9744 8237 -9367
rect 8203 -10642 8237 -10096
rect 8292 -10467 8326 -9060
rect 8381 -9314 8415 -9198
rect 8361 -9367 8371 -9314
rect 8424 -9367 8434 -9314
rect 8381 -9744 8415 -9367
rect 8273 -10520 8283 -10467
rect 8336 -10520 8346 -10467
rect 8093 -11419 8103 -11366
rect 8156 -11419 8166 -11366
rect 8113 -11681 8147 -11419
rect 8203 -11544 8237 -10995
rect 8292 -12040 8326 -10520
rect 8382 -10644 8416 -10098
rect 8381 -11543 8415 -10994
rect 8470 -11366 8504 -9056
rect 8559 -9314 8593 -9198
rect 8539 -9367 8549 -9314
rect 8602 -9367 8612 -9314
rect 8559 -9744 8593 -9367
rect 8559 -10642 8593 -10096
rect 8648 -10466 8682 -9064
rect 8737 -9315 8771 -9198
rect 8717 -9368 8727 -9315
rect 8780 -9368 8790 -9315
rect 8737 -9744 8771 -9368
rect 8628 -10519 8638 -10466
rect 8691 -10519 8701 -10466
rect 8451 -11419 8461 -11366
rect 8514 -11419 8524 -11366
rect 8470 -11681 8504 -11419
rect 8559 -11543 8593 -10994
rect 8648 -12040 8682 -10519
rect 8737 -10644 8771 -10098
rect 8737 -11543 8771 -10994
rect 8826 -11366 8860 -9063
rect 9004 -9068 9038 -8842
rect 9183 -8926 9217 -8842
rect 9361 -8923 9395 -8842
rect 8915 -9314 8949 -9198
rect 8896 -9367 8906 -9314
rect 8959 -9367 8969 -9314
rect 8915 -9744 8949 -9367
rect 9004 -9709 9038 -9113
rect 11063 -9145 11097 -8769
rect 11354 -8986 11388 -8769
rect 11647 -8981 11681 -8769
rect 11941 -9011 11975 -8769
rect 12231 -8840 12265 -8769
rect 12231 -8874 12738 -8840
rect 12231 -9013 12265 -8874
rect 12522 -8947 12556 -8874
rect 12704 -8953 12738 -8874
rect 10968 -9152 11097 -9145
rect 10772 -9230 10806 -9156
rect 10950 -9179 11097 -9152
rect 10950 -9230 10984 -9179
rect 10772 -9264 10984 -9230
rect 10861 -9638 10895 -9264
rect 11063 -9387 11097 -9179
rect 11154 -9374 11188 -9259
rect 11134 -9387 11144 -9374
rect 11063 -9421 11144 -9387
rect 11134 -9427 11144 -9421
rect 11197 -9427 11207 -9374
rect 11154 -9642 11188 -9427
rect 9004 -9743 9394 -9709
rect 11242 -9716 11276 -9180
rect 11445 -9375 11479 -9252
rect 11426 -9428 11436 -9375
rect 11489 -9428 11499 -9375
rect 11445 -9635 11479 -9428
rect 11534 -9706 11568 -9170
rect 11738 -9375 11772 -9256
rect 11718 -9428 11728 -9375
rect 11781 -9428 11791 -9375
rect 11738 -9639 11772 -9428
rect 11825 -9711 11859 -9175
rect 12030 -9376 12064 -9251
rect 12010 -9429 12020 -9376
rect 12073 -9429 12083 -9376
rect 12030 -9634 12064 -9429
rect 12118 -9704 12152 -9168
rect 12321 -9375 12355 -9252
rect 12302 -9428 12312 -9375
rect 12365 -9428 12375 -9375
rect 12321 -9635 12355 -9428
rect 12410 -9718 12444 -9182
rect 12613 -9610 12647 -9228
rect 12525 -9644 12736 -9610
rect 12525 -9737 12559 -9644
rect 12702 -9731 12736 -9644
rect 8915 -10643 8949 -10097
rect 9004 -10467 9038 -9743
rect 9182 -9824 9216 -9743
rect 9360 -9833 9394 -9743
rect 10773 -10001 10807 -9926
rect 10951 -10001 10985 -9912
rect 10773 -10035 10985 -10001
rect 9161 -10367 9171 -10314
rect 9224 -10367 9234 -10314
rect 8985 -10520 8995 -10467
rect 9048 -10520 9058 -10467
rect 8807 -11419 8817 -11366
rect 8870 -11419 8880 -11366
rect 8826 -11688 8860 -11419
rect 8915 -11543 8949 -10994
rect 9004 -11679 9038 -10520
rect 9181 -10614 9215 -10367
rect 10862 -10380 10896 -10035
rect 10772 -10414 10986 -10380
rect 10772 -10485 10806 -10414
rect 10952 -10507 10986 -10414
rect 11063 -10490 11097 -9954
rect 11153 -10400 11187 -10017
rect 11356 -10481 11390 -9941
rect 11446 -10400 11480 -10017
rect 11648 -10486 11682 -9946
rect 11737 -10400 11771 -10017
rect 11940 -10482 11974 -9942
rect 12028 -10399 12062 -10016
rect 12232 -10488 12266 -9948
rect 12320 -10398 12354 -10015
rect 12613 -10413 12647 -9999
rect 9181 -10648 9393 -10614
rect 9181 -10695 9215 -10648
rect 9359 -10726 9393 -10648
rect 9093 -11541 9127 -11005
rect 10772 -11149 10806 -11148
rect 10860 -11149 10894 -10785
rect 10772 -11183 10986 -11149
rect 11152 -11175 11186 -10792
rect 10772 -11253 10806 -11183
rect 10952 -11268 10986 -11183
rect 11244 -11260 11278 -10720
rect 11446 -11171 11480 -10788
rect 11534 -11258 11568 -10718
rect 11737 -11173 11771 -10790
rect 11826 -11260 11860 -10720
rect 12029 -11172 12063 -10789
rect 12118 -11263 12152 -10723
rect 12322 -11171 12356 -10788
rect 12410 -11263 12444 -10723
rect 12525 -10772 12559 -10649
rect 12613 -10772 12647 -10770
rect 12700 -10772 12734 -10681
rect 12525 -10806 12734 -10772
rect 12613 -11184 12647 -10806
rect 9182 -11544 9394 -11510
rect 8912 -11985 8946 -11900
rect 9095 -11985 9129 -11900
rect 9182 -11985 9216 -11544
rect 9360 -11633 9394 -11544
rect 11063 -11674 11097 -11383
rect 11043 -11727 11053 -11674
rect 11106 -11727 11116 -11674
rect 11356 -11675 11390 -11417
rect 11648 -11674 11682 -11402
rect 11940 -11674 11974 -11405
rect 12233 -11674 12267 -11403
rect 12525 -11541 12559 -11396
rect 12701 -11541 12735 -11460
rect 12525 -11575 12735 -11541
rect 11337 -11728 11347 -11675
rect 11400 -11728 11410 -11675
rect 11628 -11727 11638 -11674
rect 11691 -11727 11701 -11674
rect 11921 -11727 11931 -11674
rect 11984 -11727 11994 -11674
rect 12213 -11727 12223 -11674
rect 12276 -11727 12286 -11674
rect 13012 -11726 13022 -11673
rect 13075 -11726 13085 -11673
rect 8912 -12019 9216 -11985
rect 6868 -12074 8682 -12040
rect 5027 -13349 5037 -13296
rect 5090 -13349 5100 -13296
rect 5524 -13349 5534 -13296
rect 5587 -13349 5597 -13296
rect 5021 -13486 5031 -13433
rect 5084 -13486 5094 -13433
rect 4895 -14598 4905 -14545
rect 4958 -14598 4968 -14545
rect 4229 -14979 4239 -14926
rect 4292 -14979 4302 -14926
rect 3879 -15081 4091 -15047
rect 3682 -15875 3692 -15822
rect 3745 -15875 3755 -15822
rect 3593 -15986 3603 -15933
rect 3656 -15986 3666 -15933
rect 3612 -16080 3646 -15986
rect 3701 -16136 3735 -15875
rect 3770 -15986 3780 -15933
rect 3833 -15986 3843 -15933
rect 3790 -16080 3824 -15986
rect 3879 -16047 3913 -15081
rect 4057 -15169 4091 -15081
rect 4238 -15539 4291 -14979
rect 4228 -15592 4238 -15539
rect 4291 -15592 4301 -15539
rect 5031 -15540 5084 -13486
rect 5390 -13598 5400 -13545
rect 5453 -13598 5463 -13545
rect 5132 -13847 5142 -13794
rect 5195 -13847 5205 -13794
rect 5142 -14658 5195 -13847
rect 5133 -14711 5143 -14658
rect 5196 -14711 5206 -14658
rect 3879 -16081 4090 -16047
rect 3614 -16665 3822 -16658
rect 3879 -16665 3913 -16081
rect 4056 -16170 4090 -16081
rect 4238 -16542 4291 -15592
rect 5021 -15593 5031 -15540
rect 5084 -15593 5094 -15540
rect 4228 -16595 4238 -16542
rect 4291 -16595 4301 -16542
rect 408 -17251 616 -16718
rect 1488 -17251 1696 -16718
rect 2547 -17251 2755 -16718
rect 3504 -16719 3514 -16666
rect 3567 -16719 3577 -16666
rect 3614 -16718 3633 -16665
rect 3804 -16718 3822 -16665
rect 3858 -16718 3868 -16665
rect 3921 -16718 3931 -16665
rect 3614 -17251 3822 -16718
rect 5031 -16782 5084 -15593
rect 5400 -15653 5453 -13598
rect 5534 -13672 5587 -13349
rect 5524 -13725 5534 -13672
rect 5587 -13725 5597 -13672
rect 6912 -13922 6946 -12074
rect 8940 -13486 8950 -13433
rect 9003 -13486 9013 -13433
rect 9295 -13486 9305 -13433
rect 9358 -13486 9368 -13433
rect 8762 -13609 8772 -13556
rect 8825 -13609 8835 -13556
rect 7516 -13725 7526 -13672
rect 7579 -13725 7589 -13672
rect 7338 -13849 7348 -13796
rect 7401 -13849 7411 -13796
rect 5823 -13975 5833 -13922
rect 5886 -13975 5896 -13922
rect 6003 -13975 6013 -13922
rect 6066 -13975 6076 -13922
rect 5577 -14082 5790 -14048
rect 5843 -14078 5877 -13975
rect 6022 -14080 6056 -13975
rect 6180 -13976 6190 -13923
rect 6243 -13976 6253 -13923
rect 6359 -13975 6369 -13922
rect 6422 -13975 6432 -13922
rect 6200 -14080 6234 -13976
rect 6378 -14080 6412 -13975
rect 6537 -13976 6547 -13923
rect 6600 -13976 6610 -13923
rect 6715 -13975 6725 -13922
rect 6778 -13975 6788 -13922
rect 6892 -13975 6902 -13922
rect 6955 -13975 6965 -13922
rect 6556 -14080 6590 -13976
rect 6734 -14081 6768 -13975
rect 6912 -14079 6946 -13975
rect 7103 -14082 7297 -14048
rect 5577 -14164 5611 -14082
rect 5756 -14545 5790 -14082
rect 7179 -14161 7213 -14082
rect 5736 -14598 5746 -14545
rect 5799 -14598 5809 -14545
rect 5575 -15081 5789 -15047
rect 5843 -15075 5877 -14442
rect 5933 -14658 5967 -14388
rect 5914 -14711 5924 -14658
rect 5977 -14711 5987 -14658
rect 6022 -15080 6056 -14447
rect 6111 -14545 6145 -14392
rect 6091 -14598 6101 -14545
rect 6154 -14598 6164 -14545
rect 6200 -15079 6234 -14446
rect 6289 -14658 6323 -14387
rect 6269 -14711 6279 -14658
rect 6332 -14711 6342 -14658
rect 6378 -15081 6412 -14448
rect 6468 -14545 6502 -14388
rect 6449 -14598 6459 -14545
rect 6512 -14598 6522 -14545
rect 6557 -15081 6591 -14448
rect 6645 -14658 6679 -14387
rect 6823 -14545 6857 -14387
rect 6803 -14598 6813 -14545
rect 6866 -14598 6876 -14545
rect 7000 -14658 7034 -14397
rect 6626 -14711 6636 -14658
rect 6689 -14711 6699 -14658
rect 6981 -14711 6991 -14658
rect 7044 -14711 7054 -14658
rect 7179 -14749 7213 -14387
rect 6822 -14783 7213 -14749
rect 5575 -15172 5609 -15081
rect 5755 -15539 5789 -15081
rect 5735 -15592 5745 -15539
rect 5798 -15592 5808 -15539
rect 5390 -15706 5400 -15653
rect 5453 -15706 5463 -15653
rect 5400 -16667 5453 -15706
rect 5737 -15803 5747 -15750
rect 5800 -15803 5810 -15750
rect 5576 -16438 5610 -16353
rect 5756 -16438 5790 -15803
rect 5844 -16081 5878 -15448
rect 5933 -15652 5967 -15376
rect 5913 -15705 5923 -15652
rect 5976 -15705 5986 -15652
rect 5911 -16001 5921 -15948
rect 5974 -16001 5984 -15948
rect 5931 -16133 5965 -16001
rect 6022 -16082 6056 -15449
rect 6111 -15539 6145 -15380
rect 6091 -15592 6101 -15539
rect 6154 -15592 6164 -15539
rect 6091 -15802 6101 -15749
rect 6154 -15802 6164 -15749
rect 6112 -16136 6146 -15802
rect 6201 -16082 6235 -15449
rect 6289 -15652 6323 -15364
rect 6269 -15705 6279 -15652
rect 6332 -15705 6342 -15652
rect 6269 -16001 6279 -15948
rect 6332 -16001 6342 -15948
rect 6288 -16137 6322 -16001
rect 6379 -16081 6413 -15448
rect 6468 -15539 6502 -15375
rect 6448 -15592 6458 -15539
rect 6511 -15592 6521 -15539
rect 6446 -15803 6456 -15750
rect 6509 -15803 6519 -15750
rect 6467 -16137 6501 -15803
rect 6556 -16081 6590 -15448
rect 6645 -15652 6679 -15357
rect 6822 -15368 6856 -14783
rect 7357 -14824 7391 -13849
rect 7427 -13975 7437 -13922
rect 7490 -13975 7500 -13922
rect 7446 -14081 7480 -13975
rect 6983 -14877 6993 -14824
rect 7046 -14877 7056 -14824
rect 7337 -14877 7347 -14824
rect 7400 -14877 7410 -14824
rect 6822 -15438 6857 -15368
rect 6748 -15472 6942 -15438
rect 6625 -15705 6635 -15652
rect 6688 -15705 6698 -15652
rect 6703 -15804 6713 -15751
rect 6766 -15804 6776 -15751
rect 6624 -16001 6634 -15948
rect 6687 -16001 6697 -15948
rect 6734 -15956 6768 -15804
rect 6822 -15851 6856 -15472
rect 6803 -15904 6813 -15851
rect 6866 -15904 6876 -15851
rect 7002 -15951 7036 -14877
rect 7070 -14976 7080 -14923
rect 7133 -14976 7143 -14923
rect 7090 -15080 7124 -14976
rect 7250 -14977 7260 -14924
rect 7313 -14977 7323 -14924
rect 7269 -15080 7303 -14977
rect 7357 -15182 7391 -14877
rect 7447 -14923 7481 -14448
rect 7429 -14976 7439 -14923
rect 7492 -14976 7502 -14923
rect 7447 -15081 7481 -14976
rect 7535 -15163 7569 -13725
rect 7872 -13726 7882 -13673
rect 7935 -13726 7945 -13673
rect 8228 -13724 8238 -13671
rect 8291 -13724 8301 -13671
rect 7694 -13848 7704 -13795
rect 7757 -13848 7767 -13795
rect 7605 -13975 7615 -13922
rect 7668 -13975 7678 -13922
rect 7624 -14080 7658 -13975
rect 7713 -14130 7747 -13848
rect 7783 -13976 7793 -13923
rect 7846 -13976 7856 -13923
rect 7802 -14081 7836 -13976
rect 7892 -14124 7926 -13726
rect 8051 -13849 8061 -13796
rect 8114 -13849 8124 -13796
rect 7960 -13975 7970 -13922
rect 8023 -13975 8033 -13922
rect 7980 -14081 8014 -13975
rect 8069 -14134 8103 -13849
rect 8138 -13975 8148 -13922
rect 8201 -13975 8211 -13922
rect 8158 -14081 8192 -13975
rect 8248 -14137 8282 -13724
rect 8405 -13849 8415 -13796
rect 8468 -13849 8478 -13796
rect 8316 -13975 8326 -13922
rect 8379 -13975 8389 -13922
rect 8336 -14080 8370 -13975
rect 8425 -14142 8459 -13849
rect 8529 -14082 8723 -14048
rect 8603 -14165 8637 -14082
rect 8781 -14129 8815 -13609
rect 8851 -13975 8861 -13922
rect 8914 -13975 8924 -13922
rect 8871 -14081 8905 -13975
rect 8960 -14131 8994 -13486
rect 9117 -13609 9127 -13556
rect 9180 -13609 9190 -13556
rect 9028 -13975 9038 -13922
rect 9091 -13975 9101 -13922
rect 9048 -14081 9082 -13975
rect 9137 -14134 9171 -13609
rect 9207 -13975 9217 -13922
rect 9270 -13975 9280 -13922
rect 9227 -14081 9261 -13975
rect 9315 -14130 9349 -13486
rect 9473 -13609 9483 -13556
rect 9536 -13609 9546 -13556
rect 9384 -13975 9394 -13922
rect 9447 -13975 9457 -13922
rect 9404 -14081 9438 -13975
rect 9493 -14132 9527 -13609
rect 11432 -13725 11442 -13672
rect 11495 -13725 11505 -13672
rect 11788 -13725 11798 -13672
rect 11851 -13725 11861 -13672
rect 11254 -13849 11264 -13796
rect 11317 -13849 11327 -13796
rect 9919 -13976 9929 -13923
rect 9982 -13976 9992 -13923
rect 10098 -13975 10108 -13922
rect 10161 -13975 10171 -13922
rect 9594 -14082 9788 -14048
rect 9938 -14081 9972 -13976
rect 10117 -14082 10151 -13975
rect 10274 -13976 10284 -13923
rect 10337 -13976 10347 -13923
rect 10452 -13976 10462 -13923
rect 10515 -13976 10525 -13923
rect 10630 -13975 10640 -13922
rect 10693 -13975 10703 -13922
rect 10294 -14082 10328 -13976
rect 10472 -14081 10506 -13976
rect 10650 -14081 10684 -13975
rect 10809 -13976 10819 -13923
rect 10872 -13976 10882 -13923
rect 10828 -14081 10862 -13976
rect 11018 -14082 11212 -14048
rect 9671 -14159 9705 -14082
rect 11095 -14158 11129 -14082
rect 7625 -15081 7659 -14448
rect 7694 -14878 7704 -14825
rect 7757 -14878 7767 -14825
rect 7714 -15135 7748 -14878
rect 7802 -15081 7836 -14448
rect 8226 -14598 8236 -14545
rect 8289 -14598 8299 -14545
rect 8050 -14874 8060 -14821
rect 8113 -14874 8123 -14821
rect 7179 -15750 7213 -15384
rect 7159 -15803 7169 -15750
rect 7222 -15803 7232 -15750
rect 7159 -15905 7169 -15852
rect 7222 -15905 7232 -15852
rect 6734 -15990 6858 -15956
rect 6644 -16145 6678 -16001
rect 6824 -16163 6858 -15990
rect 6984 -16004 6994 -15951
rect 7047 -16004 7057 -15951
rect 7002 -16273 7036 -16004
rect 7178 -16438 7212 -15905
rect 7447 -16080 7481 -15447
rect 7536 -15749 7570 -15382
rect 7516 -15802 7526 -15749
rect 7579 -15802 7589 -15749
rect 7516 -16006 7526 -15953
rect 7579 -16006 7589 -15953
rect 7535 -16147 7569 -16006
rect 7624 -16081 7658 -15448
rect 7803 -16081 7837 -15448
rect 7891 -15749 7925 -15369
rect 8069 -15438 8103 -14874
rect 8000 -15472 8194 -15438
rect 7872 -15802 7882 -15749
rect 7935 -15802 7945 -15749
rect 8069 -15851 8103 -15472
rect 8050 -15904 8060 -15851
rect 8113 -15904 8123 -15851
rect 8247 -15952 8281 -14598
rect 8336 -14923 8370 -14448
rect 8407 -14710 8417 -14657
rect 8470 -14710 8480 -14657
rect 8317 -14976 8327 -14923
rect 8380 -14976 8390 -14923
rect 8336 -15081 8370 -14976
rect 7871 -16005 7881 -15952
rect 7934 -16005 7944 -15952
rect 8227 -16005 8237 -15952
rect 8290 -16005 8300 -15952
rect 7891 -16167 7925 -16005
rect 8247 -16221 8281 -16005
rect 8336 -16080 8370 -15447
rect 5576 -16472 5790 -16438
rect 6557 -16544 6591 -16441
rect 6735 -16544 6769 -16440
rect 6538 -16597 6548 -16544
rect 6601 -16597 6611 -16544
rect 6716 -16597 6726 -16544
rect 6779 -16597 6789 -16544
rect 6912 -16545 6946 -16442
rect 7101 -16472 7295 -16438
rect 6893 -16598 6903 -16545
rect 6956 -16598 6966 -16545
rect 5389 -16720 5399 -16667
rect 5452 -16720 5462 -16667
rect 5021 -16835 5031 -16782
rect 5084 -16835 5094 -16782
rect 7357 -16890 7391 -16342
rect 7713 -16890 7747 -16345
rect 7980 -16545 8014 -16453
rect 7960 -16598 7970 -16545
rect 8023 -16598 8033 -16545
rect 8069 -16890 8103 -16382
rect 8158 -16544 8192 -16445
rect 8139 -16597 8149 -16544
rect 8202 -16597 8212 -16544
rect 8426 -16890 8460 -14710
rect 8514 -14806 8548 -14438
rect 8585 -14598 8595 -14545
rect 8648 -14598 8658 -14545
rect 8494 -14859 8504 -14806
rect 8557 -14859 8567 -14806
rect 8514 -14871 8548 -14859
rect 8495 -14977 8505 -14924
rect 8558 -14977 8568 -14924
rect 8514 -15080 8548 -14977
rect 8604 -15136 8638 -14598
rect 8762 -14711 8772 -14658
rect 8825 -14711 8835 -14658
rect 8692 -14924 8726 -14923
rect 8673 -14977 8683 -14924
rect 8736 -14977 8746 -14924
rect 8692 -15080 8726 -14977
rect 8781 -15148 8815 -14711
rect 8870 -15081 8904 -14448
rect 8940 -14599 8950 -14546
rect 9003 -14599 9013 -14546
rect 8960 -15139 8994 -14599
rect 9048 -15081 9082 -14448
rect 9117 -14712 9127 -14659
rect 9180 -14712 9190 -14659
rect 9137 -15140 9171 -14712
rect 9226 -15081 9260 -14448
rect 9294 -14598 9304 -14545
rect 9357 -14598 9367 -14545
rect 9314 -15144 9348 -14598
rect 9404 -15081 9438 -14448
rect 9651 -14598 9661 -14545
rect 9714 -14598 9724 -14545
rect 9473 -14711 9483 -14658
rect 9536 -14711 9546 -14658
rect 9493 -15135 9527 -14711
rect 9562 -14976 9572 -14923
rect 9625 -14976 9635 -14923
rect 9582 -15077 9616 -14976
rect 9671 -15139 9705 -14598
rect 9763 -14806 9797 -14453
rect 9848 -14659 9882 -14383
rect 9827 -14712 9837 -14659
rect 9890 -14712 9900 -14659
rect 9743 -14859 9753 -14806
rect 9806 -14859 9816 -14806
rect 9763 -14871 9797 -14859
rect 9740 -14976 9750 -14923
rect 9803 -14976 9813 -14923
rect 9760 -15078 9794 -14976
rect 9848 -15200 9882 -14712
rect 9939 -14923 9973 -14449
rect 10026 -14545 10060 -14384
rect 10006 -14598 10016 -14545
rect 10069 -14598 10079 -14545
rect 9919 -14976 9929 -14923
rect 9982 -14976 9992 -14923
rect 9939 -15082 9973 -14976
rect 10026 -15216 10060 -14598
rect 10205 -14658 10239 -14385
rect 10383 -14546 10417 -14385
rect 10363 -14599 10373 -14546
rect 10426 -14599 10436 -14546
rect 10186 -14711 10196 -14658
rect 10249 -14711 10259 -14658
rect 10185 -14875 10195 -14822
rect 10248 -14875 10258 -14822
rect 10205 -15438 10239 -14875
rect 10472 -15081 10506 -14448
rect 10560 -14658 10594 -14383
rect 10540 -14711 10550 -14658
rect 10603 -14711 10613 -14658
rect 10542 -14868 10552 -14815
rect 10605 -14868 10615 -14815
rect 10561 -15136 10595 -14868
rect 10650 -15081 10684 -14448
rect 10738 -14545 10772 -14383
rect 10719 -14598 10729 -14545
rect 10782 -14598 10792 -14545
rect 10828 -14923 10862 -14448
rect 10917 -14658 10951 -14387
rect 11096 -14658 11130 -14334
rect 10898 -14711 10908 -14658
rect 10961 -14711 10971 -14658
rect 11077 -14711 11087 -14658
rect 11140 -14711 11150 -14658
rect 10898 -14866 10908 -14813
rect 10961 -14866 10971 -14813
rect 11273 -14815 11307 -13849
rect 11343 -13975 11353 -13922
rect 11406 -13975 11416 -13922
rect 11362 -14081 11396 -13975
rect 11452 -14133 11486 -13725
rect 11610 -13850 11620 -13797
rect 11673 -13850 11683 -13797
rect 11520 -13975 11530 -13922
rect 11583 -13975 11593 -13922
rect 11540 -14080 11574 -13975
rect 11630 -14135 11664 -13850
rect 11699 -13975 11709 -13922
rect 11762 -13975 11772 -13922
rect 11719 -14081 11753 -13975
rect 11807 -14133 11841 -13725
rect 12142 -13726 12152 -13673
rect 12205 -13726 12215 -13673
rect 12499 -13725 12509 -13672
rect 12562 -13725 12572 -13672
rect 11967 -13849 11977 -13796
rect 12030 -13849 12040 -13796
rect 11876 -13976 11886 -13923
rect 11939 -13976 11949 -13923
rect 11895 -14080 11929 -13976
rect 11986 -14131 12020 -13849
rect 12054 -13975 12064 -13922
rect 12117 -13975 12127 -13922
rect 12073 -14082 12107 -13975
rect 12162 -14137 12196 -13726
rect 12324 -13849 12334 -13796
rect 12387 -13849 12397 -13796
rect 12232 -13976 12242 -13923
rect 12295 -13976 12305 -13923
rect 12252 -14081 12286 -13976
rect 12342 -14133 12376 -13849
rect 12410 -13975 12420 -13922
rect 12473 -13975 12483 -13922
rect 12430 -14081 12464 -13975
rect 12519 -14048 12553 -13725
rect 12519 -14082 12731 -14048
rect 12519 -14134 12553 -14082
rect 12697 -14154 12731 -14082
rect 11430 -14709 11440 -14656
rect 11493 -14709 11503 -14656
rect 10809 -14976 10819 -14923
rect 10872 -14976 10882 -14923
rect 10828 -15081 10862 -14976
rect 8583 -15905 8593 -15852
rect 8646 -15905 8656 -15852
rect 8603 -16438 8637 -15905
rect 8870 -16080 8904 -15447
rect 9049 -16081 9083 -15448
rect 9226 -16080 9260 -15447
rect 9404 -16080 9438 -15447
rect 9653 -15905 9663 -15852
rect 9716 -15905 9726 -15852
rect 8519 -16472 8713 -16438
rect 8781 -16666 8815 -16386
rect 8761 -16719 8771 -16666
rect 8824 -16719 8834 -16666
rect 8960 -16782 8994 -16389
rect 9138 -16666 9172 -16383
rect 9118 -16719 9128 -16666
rect 9181 -16719 9191 -16666
rect 9315 -16782 9349 -16393
rect 9493 -16666 9527 -16380
rect 9672 -16438 9706 -15905
rect 9939 -16081 9973 -15448
rect 10122 -15472 10316 -15438
rect 10205 -15852 10239 -15472
rect 10383 -15751 10417 -15349
rect 10363 -15804 10373 -15751
rect 10426 -15804 10436 -15751
rect 10184 -15905 10194 -15852
rect 10247 -15905 10257 -15852
rect 10472 -16080 10506 -15447
rect 10650 -16080 10684 -15447
rect 10739 -15750 10773 -15359
rect 10720 -15803 10730 -15750
rect 10783 -15803 10793 -15750
rect 10739 -16238 10773 -15803
rect 10828 -16080 10862 -15447
rect 10916 -16215 10950 -14866
rect 11254 -14868 11264 -14815
rect 11317 -14868 11327 -14815
rect 10986 -14976 10996 -14923
rect 11049 -14976 11059 -14923
rect 11165 -14976 11175 -14923
rect 11228 -14976 11238 -14923
rect 11006 -15061 11040 -14976
rect 11184 -15063 11218 -14976
rect 11273 -15189 11307 -14868
rect 11095 -15750 11129 -15348
rect 11451 -15438 11485 -14709
rect 11717 -15078 11751 -14439
rect 11897 -15079 11931 -14440
rect 12075 -15079 12109 -14440
rect 12253 -15081 12287 -14442
rect 12430 -15081 12464 -14442
rect 12520 -15083 12730 -15049
rect 11390 -15472 11584 -15438
rect 11076 -15803 11086 -15750
rect 11139 -15803 11149 -15750
rect 11451 -15841 11485 -15472
rect 11629 -15652 11663 -15392
rect 11609 -15705 11619 -15652
rect 11672 -15705 11682 -15652
rect 11629 -15706 11663 -15705
rect 11074 -15905 11084 -15852
rect 11137 -15905 11147 -15852
rect 11430 -15894 11440 -15841
rect 11493 -15894 11503 -15841
rect 11451 -15902 11485 -15894
rect 9595 -16472 9789 -16438
rect 9474 -16719 9484 -16666
rect 9537 -16719 9547 -16666
rect 8940 -16835 8950 -16782
rect 9003 -16835 9013 -16782
rect 9295 -16835 9305 -16782
rect 9358 -16835 9368 -16782
rect 7337 -16943 7347 -16890
rect 7400 -16943 7410 -16890
rect 7694 -16943 7704 -16890
rect 7757 -16943 7767 -16890
rect 8050 -16943 8060 -16890
rect 8113 -16943 8123 -16890
rect 8406 -16943 8416 -16890
rect 8469 -16943 8479 -16890
rect 9672 -17251 9706 -16472
rect 9848 -16666 9882 -16349
rect 9938 -16544 9972 -16458
rect 9919 -16597 9929 -16544
rect 9982 -16597 9992 -16544
rect 9828 -16719 9838 -16666
rect 9891 -16719 9901 -16666
rect 10028 -16781 10062 -16383
rect 10117 -16545 10151 -16456
rect 10097 -16598 10107 -16545
rect 10160 -16598 10170 -16545
rect 10205 -16665 10239 -16334
rect 10296 -16545 10330 -16458
rect 10277 -16598 10287 -16545
rect 10340 -16598 10350 -16545
rect 10185 -16718 10195 -16665
rect 10248 -16718 10258 -16665
rect 10383 -16781 10417 -16377
rect 10561 -16665 10595 -16352
rect 10540 -16718 10550 -16665
rect 10603 -16718 10613 -16665
rect 10739 -16779 10773 -16359
rect 10917 -16665 10951 -16377
rect 11094 -16437 11128 -15905
rect 11431 -16005 11441 -15952
rect 11494 -16005 11504 -15952
rect 11451 -16138 11485 -16005
rect 11718 -16081 11752 -15448
rect 11808 -15540 11842 -15394
rect 11788 -15593 11798 -15540
rect 11851 -15593 11861 -15540
rect 11787 -16005 11797 -15952
rect 11850 -16005 11860 -15952
rect 11806 -16136 11840 -16005
rect 11897 -16081 11931 -15448
rect 11985 -15652 12019 -15387
rect 11965 -15705 11975 -15652
rect 12028 -15705 12038 -15652
rect 12074 -16080 12108 -15447
rect 12165 -15539 12199 -15372
rect 12145 -15592 12155 -15539
rect 12208 -15592 12218 -15539
rect 12144 -16005 12154 -15952
rect 12207 -16005 12217 -15952
rect 12163 -16136 12197 -16005
rect 12252 -16081 12286 -15448
rect 12342 -15652 12376 -15386
rect 12322 -15705 12332 -15652
rect 12385 -15705 12395 -15652
rect 12431 -16081 12465 -15448
rect 12520 -15539 12554 -15083
rect 12696 -15154 12730 -15083
rect 12501 -15592 12511 -15539
rect 12564 -15592 12574 -15539
rect 12501 -16005 12511 -15952
rect 12564 -16005 12574 -15952
rect 11019 -16471 11213 -16437
rect 10897 -16718 10907 -16665
rect 10960 -16718 10970 -16665
rect 10007 -16834 10017 -16781
rect 10070 -16834 10080 -16781
rect 10364 -16834 10374 -16781
rect 10427 -16834 10437 -16781
rect 10721 -16832 10731 -16779
rect 10784 -16832 10794 -16779
rect 11273 -16890 11307 -16340
rect 11362 -16545 11396 -16455
rect 11342 -16598 11352 -16545
rect 11405 -16598 11415 -16545
rect 11540 -16546 11574 -16453
rect 11520 -16599 11530 -16546
rect 11583 -16599 11593 -16546
rect 11630 -16890 11664 -16362
rect 11718 -16545 11752 -16457
rect 11699 -16598 11709 -16545
rect 11762 -16598 11772 -16545
rect 11985 -16889 12019 -16353
rect 12340 -16889 12374 -16380
rect 12520 -16440 12554 -16005
rect 12698 -16440 12732 -16356
rect 12520 -16474 12732 -16440
rect 11253 -16943 11263 -16890
rect 11316 -16943 11326 -16890
rect 11610 -16943 11620 -16890
rect 11673 -16943 11683 -16890
rect 11965 -16942 11975 -16889
rect 12028 -16942 12038 -16889
rect 12321 -16942 12331 -16889
rect 12384 -16942 12394 -16889
rect 13022 -17251 13075 -11726
rect 18337 -13421 18412 -6747
rect 18327 -13496 18337 -13421
rect 18412 -13496 18422 -13421
rect 18337 -13506 18412 -13496
rect -7605 -17459 13720 -17251
rect -7605 -17559 -7323 -17459
rect 13384 -17527 13720 -17459
rect 13384 -17559 13719 -17527
rect -7605 -17587 13719 -17559
<< via1 >>
rect -5867 -1963 -5814 -1910
rect -5689 -1963 -5636 -1910
rect -5510 -1963 -5457 -1910
rect -5333 -1963 -5280 -1910
rect -5155 -1963 -5102 -1910
rect -4976 -1963 -4923 -1910
rect -4799 -1963 -4746 -1910
rect -4621 -1963 -4568 -1910
rect -4443 -1963 -4390 -1910
rect -4265 -1963 -4212 -1910
rect -4086 -1963 -4033 -1910
rect -3909 -1963 -3856 -1910
rect -1109 -1963 -1056 -1910
rect -6498 -2582 -6445 -2529
rect -6625 -3454 -6572 -3401
rect -6044 -2833 -5991 -2780
rect -6134 -3454 -6081 -3401
rect -6498 -3693 -6445 -3640
rect -6498 -4324 -6445 -4271
rect -6134 -4443 -6081 -4390
rect -6498 -5194 -6445 -5141
rect -6625 -5375 -6572 -5322
rect -6134 -5285 -6081 -5232
rect -5777 -2583 -5724 -2530
rect -5866 -2833 -5813 -2780
rect -5777 -3569 -5724 -3516
rect -5778 -4324 -5725 -4271
rect -5777 -5468 -5724 -5415
rect -5421 -2721 -5368 -2668
rect -5422 -3693 -5369 -3640
rect -5422 -4559 -5369 -4506
rect -5422 -5194 -5369 -5141
rect -5066 -2583 -5013 -2530
rect -5066 -3454 -5013 -3401
rect -5066 -4443 -5013 -4390
rect -5066 -5286 -5013 -5233
rect -4710 -2721 -4657 -2668
rect -4710 -3454 -4657 -3401
rect -4709 -4443 -4656 -4390
rect -4710 -5375 -4657 -5322
rect -4354 -2583 -4301 -2530
rect -4353 -3693 -4300 -3640
rect -4353 -4559 -4300 -4506
rect -4353 -5194 -4300 -5141
rect -3998 -2721 -3945 -2668
rect -1109 -2478 -1056 -2425
rect -752 -2478 -699 -2425
rect -3908 -2833 -3855 -2780
rect -3998 -3569 -3945 -3516
rect -3998 -4324 -3945 -4271
rect -3997 -5468 -3944 -5415
rect -2624 -2611 -2571 -2558
rect -1285 -2611 -1232 -2558
rect -3298 -2721 -3245 -2668
rect -3731 -2833 -3678 -2780
rect -3642 -3454 -3589 -3401
rect -3131 -3454 -3078 -3401
rect -3298 -3569 -3245 -3516
rect -3642 -4443 -3589 -4390
rect -3298 -4559 -3245 -4506
rect -3642 -5372 -3589 -5319
rect -3130 -5286 -3077 -5233
rect -1197 -2718 -1144 -2665
rect -930 -2611 -877 -2558
rect -1019 -2718 -966 -2665
rect -841 -2718 -788 -2665
rect -129 -2718 -76 -2665
rect 50 -2718 103 -2665
rect 227 -2718 280 -2665
rect 5337 -2258 5390 -2205
rect 1919 -2479 1972 -2426
rect 2275 -2479 2328 -2426
rect 940 -2718 993 -2665
rect 1117 -2718 1170 -2665
rect 1295 -2718 1348 -2665
rect -1645 -3510 -1584 -3449
rect -2004 -4465 -1951 -4412
rect -2624 -5377 -2571 -5324
rect -3298 -5469 -3245 -5416
rect -5956 -6069 -5903 -6016
rect -5601 -6069 -5548 -6016
rect -5778 -6184 -5725 -6131
rect -5244 -6069 -5191 -6016
rect -5065 -6184 -5012 -6131
rect -6498 -6301 -6445 -6248
rect -5421 -6301 -5368 -6248
rect -4888 -6069 -4835 -6016
rect -4710 -6301 -4657 -6248
rect -4532 -6069 -4479 -6016
rect -4175 -6069 -4122 -6016
rect -4354 -6184 -4301 -6131
rect -3820 -6069 -3767 -6016
rect -2624 -6060 -2571 -6007
rect -3298 -6184 -3245 -6131
rect -3998 -6300 -3945 -6247
rect -4786 -6431 -4733 -6378
rect -1876 -5285 -1823 -5232
rect -1286 -3624 -1233 -3571
rect -1108 -3509 -1055 -3456
rect -929 -3624 -876 -3571
rect -484 -3354 -431 -3301
rect -750 -3509 -697 -3456
rect -396 -3509 -343 -3456
rect -573 -3624 -520 -3571
rect -217 -3624 -164 -3571
rect 583 -3354 636 -3301
rect -39 -3509 14 -3456
rect 317 -3509 370 -3456
rect 850 -3509 903 -3456
rect 1206 -3509 1259 -3456
rect 2097 -2607 2150 -2554
rect 2007 -2718 2060 -2665
rect 2186 -2718 2239 -2665
rect 3193 -2480 3246 -2427
rect 2453 -2607 2506 -2554
rect 2363 -2718 2416 -2665
rect 1654 -3354 1707 -3301
rect 1562 -3509 1615 -3456
rect 1919 -3509 1972 -3456
rect 1384 -3617 1437 -3564
rect 1741 -3617 1794 -3564
rect 2097 -3617 2150 -3564
rect 2275 -3509 2328 -3456
rect 2451 -3617 2504 -3564
rect -841 -4245 -788 -4192
rect -662 -4245 -609 -4192
rect -483 -4245 -430 -4192
rect -306 -4245 -253 -4192
rect -1287 -5150 -1234 -5097
rect -1646 -5339 -1585 -5278
rect -1105 -5266 -1052 -5213
rect -929 -5150 -876 -5097
rect -572 -5150 -519 -5097
rect -218 -5150 -165 -5097
rect -751 -5266 -698 -5213
rect -396 -5266 -343 -5213
rect -1876 -6417 -1823 -6364
rect -1282 -6417 -1229 -6364
rect -928 -6417 -876 -6365
rect -1110 -6532 -1057 -6479
rect -752 -6532 -699 -6479
rect 407 -4245 460 -4192
rect 317 -4357 370 -4304
rect 583 -4245 636 -4192
rect 495 -4465 548 -4412
rect 761 -4245 814 -4192
rect 673 -4357 726 -4304
rect 850 -4465 903 -4412
rect 1474 -4245 1527 -4192
rect 1652 -4245 1705 -4192
rect 1830 -4245 1883 -4192
rect 2008 -4245 2061 -4192
rect 2538 -4327 2599 -4266
rect 2746 -4507 2807 -4446
rect -41 -5266 12 -5213
rect 316 -5266 369 -5213
rect -128 -5433 -75 -5380
rect 50 -5433 103 -5380
rect 228 -5433 281 -5380
rect 850 -5266 903 -5213
rect 1207 -5266 1260 -5213
rect 940 -5434 993 -5381
rect 1119 -5433 1172 -5380
rect 1385 -5146 1438 -5093
rect 1296 -5433 1349 -5380
rect 227 -6303 280 -6250
rect 1740 -5146 1793 -5093
rect 1563 -5266 1616 -5213
rect 1917 -5266 1970 -5213
rect 2096 -5146 2149 -5093
rect 2274 -5266 2327 -5213
rect 2453 -5146 2506 -5093
rect 942 -6303 995 -6250
rect 2096 -6060 2149 -6007
rect 2452 -6060 2505 -6007
rect 1918 -6177 1971 -6124
rect 2275 -6177 2328 -6124
rect 3194 -4857 3246 -4805
rect 4771 -4857 4823 -4805
rect 2879 -6417 2931 -6365
rect 5037 -5059 5090 -5006
rect 4905 -5265 4958 -5212
rect -753 -6651 -700 -6598
rect 4772 -6650 4825 -6597
rect -2003 -6767 -1950 -6714
rect 6680 -2263 6744 -2199
rect 6222 -3515 6286 -3451
rect 5614 -5271 5678 -5207
rect 5337 -5580 5390 -5527
rect 17831 -6585 17895 -6521
rect 4770 -6944 4823 -6891
rect 4906 -6942 4959 -6889
rect 5038 -6940 5091 -6887
rect -3873 -7743 -3821 -7691
rect -3731 -7837 -3679 -7785
rect -3541 -7840 -3489 -7788
rect -5502 -12324 -5449 -12271
rect -6077 -12565 -6024 -12512
rect -5626 -12565 -5573 -12512
rect -6223 -13115 -6170 -13062
rect -6426 -13905 -6373 -13852
rect -5000 -12325 -4947 -12272
rect -4502 -12324 -4449 -12271
rect -5376 -12441 -5323 -12388
rect -5127 -12441 -5074 -12388
rect -4877 -12565 -4824 -12512
rect -4627 -12565 -4574 -12512
rect -4377 -12441 -4324 -12388
rect -3928 -12442 -3875 -12389
rect -5751 -13115 -5698 -13062
rect -5251 -13242 -5198 -13189
rect -4752 -13115 -4699 -13062
rect -4251 -13242 -4198 -13189
rect -6077 -13798 -6024 -13745
rect -5376 -13798 -5323 -13745
rect -5626 -13905 -5573 -13852
rect -5730 -14010 -5677 -13957
rect -5126 -13798 -5073 -13745
rect -4877 -13905 -4824 -13852
rect -4376 -13798 -4323 -13745
rect -4627 -13905 -4574 -13852
rect -4752 -14010 -4699 -13957
rect -3788 -13242 -3735 -13189
rect -3928 -13905 -3875 -13852
rect -3788 -14010 -3735 -13957
rect -6223 -14108 -6170 -14055
rect -5250 -14108 -5197 -14055
rect -4250 -14108 -4197 -14055
rect -6159 -14848 -6106 -14795
rect -5860 -14848 -5807 -14795
rect -5504 -14954 -5451 -14901
rect -6159 -15535 -6106 -15482
rect -5860 -15641 -5807 -15588
rect -5504 -15534 -5451 -15481
rect -6159 -16246 -6106 -16193
rect -5860 -16347 -5807 -16294
rect -5504 -16246 -5451 -16193
rect -5147 -14848 -5094 -14795
rect -5148 -15642 -5095 -15589
rect -5148 -16347 -5095 -16294
rect -4791 -14954 -4738 -14901
rect -4792 -15534 -4739 -15481
rect -4792 -16246 -4739 -16193
rect -4436 -14848 -4383 -14795
rect 4771 -7907 4824 -7854
rect 4906 -7905 4959 -7852
rect 5037 -7903 5090 -7850
rect -3382 -7986 -3329 -7933
rect -1382 -7975 -1329 -7922
rect -3542 -13242 -3489 -13189
rect -1203 -7976 -1150 -7923
rect -1025 -7975 -972 -7922
rect -848 -7975 -795 -7922
rect -670 -7975 -617 -7922
rect -490 -7975 -437 -7922
rect 755 -7975 808 -7922
rect 932 -7975 985 -7922
rect 1112 -7975 1165 -7922
rect 1289 -7976 1342 -7923
rect 1467 -7975 1520 -7922
rect 1644 -7975 1697 -7922
rect 2890 -7975 2943 -7922
rect 3069 -7975 3122 -7922
rect 3247 -7975 3300 -7922
rect 3424 -7975 3477 -7922
rect 3603 -7976 3656 -7923
rect 3778 -7975 3831 -7922
rect 4208 -7976 4261 -7923
rect -1916 -8587 -1863 -8534
rect -1739 -8587 -1686 -8534
rect -1826 -8706 -1773 -8653
rect -2447 -8820 -2394 -8767
rect -2005 -8820 -1952 -8767
rect -2315 -9978 -2262 -9925
rect -2447 -12325 -2394 -12272
rect -3382 -14108 -3329 -14055
rect -3936 -14954 -3883 -14901
rect -4435 -15641 -4383 -15589
rect -4436 -16347 -4383 -16294
rect -3935 -15641 -3883 -15589
rect -1916 -9599 -1863 -9546
rect -1916 -9978 -1863 -9925
rect -1558 -8587 -1505 -8534
rect -1382 -8587 -1329 -8534
rect -1470 -8706 -1417 -8653
rect -1648 -8820 -1595 -8767
rect -1738 -9599 -1685 -9546
rect -1738 -9979 -1685 -9926
rect -1558 -9599 -1505 -9546
rect -1560 -9978 -1507 -9925
rect -1203 -8587 -1150 -8534
rect -1293 -8820 -1240 -8767
rect -1382 -9977 -1329 -9924
rect -1026 -8587 -973 -8534
rect -1115 -8706 -1062 -8653
rect -848 -8587 -795 -8534
rect -936 -8820 -883 -8767
rect -670 -8587 -617 -8534
rect -758 -8706 -705 -8653
rect -491 -8587 -438 -8534
rect -580 -8819 -527 -8766
rect -314 -8587 -261 -8534
rect -402 -8706 -349 -8653
rect -136 -8587 -83 -8534
rect 42 -8587 95 -8534
rect -47 -8706 6 -8653
rect -225 -8820 -172 -8767
rect -312 -9599 -259 -9546
rect -314 -9978 -261 -9925
rect -136 -9598 -83 -9545
rect -136 -9979 -83 -9926
rect 221 -8587 274 -8534
rect 398 -8587 451 -8534
rect 310 -8706 363 -8653
rect 132 -8821 185 -8768
rect 42 -9599 95 -9546
rect 43 -9978 96 -9925
rect 222 -9598 275 -9545
rect 220 -9978 273 -9925
rect 577 -8587 630 -8534
rect 754 -8587 807 -8534
rect 666 -8706 719 -8653
rect 489 -8819 542 -8766
rect 399 -9599 452 -9546
rect 398 -9978 451 -9925
rect 577 -9599 630 -9546
rect 576 -9978 629 -9925
rect 932 -8587 985 -8534
rect 843 -8819 896 -8766
rect 1111 -8587 1164 -8534
rect 1022 -8706 1075 -8653
rect 1289 -8587 1342 -8534
rect 1201 -8820 1254 -8767
rect 1466 -8587 1519 -8534
rect 1377 -8706 1430 -8653
rect 1644 -8587 1697 -8534
rect 1556 -8820 1609 -8767
rect 1822 -8587 1875 -8534
rect 1733 -8706 1786 -8653
rect 2000 -8587 2053 -8534
rect 2178 -8587 2231 -8534
rect 2090 -8706 2143 -8653
rect 1911 -8820 1964 -8767
rect 2357 -8587 2410 -8534
rect 2534 -8587 2587 -8534
rect 2446 -8706 2499 -8653
rect 2267 -8820 2320 -8767
rect 2178 -9600 2231 -9547
rect 2357 -9599 2410 -9546
rect 2356 -9978 2409 -9925
rect 2712 -8587 2765 -8534
rect 2890 -8587 2943 -8534
rect 2802 -8706 2855 -8653
rect 2624 -8820 2677 -8767
rect 2534 -9599 2587 -9546
rect 2534 -9978 2587 -9925
rect 2713 -9599 2766 -9546
rect 2712 -9979 2765 -9926
rect 3068 -8587 3121 -8534
rect 2980 -8820 3033 -8767
rect 2891 -9978 2944 -9925
rect 3246 -8587 3299 -8534
rect 3158 -8706 3211 -8653
rect 3069 -9978 3122 -9925
rect 3424 -8587 3477 -8534
rect 3336 -8820 3389 -8767
rect 3246 -9978 3299 -9925
rect 3602 -8587 3655 -8534
rect 3513 -8706 3566 -8653
rect 3781 -8587 3834 -8534
rect 3692 -8820 3745 -8767
rect 3869 -8706 3922 -8653
rect 4771 -9367 4824 -9314
rect 4208 -9599 4261 -9546
rect -1827 -10961 -1774 -10908
rect -1470 -10961 -1417 -10908
rect -2004 -11690 -1951 -11637
rect -1915 -11972 -1862 -11919
rect -2005 -12595 -1952 -12542
rect -1649 -11581 -1596 -11528
rect -1738 -11972 -1685 -11919
rect -1559 -11972 -1506 -11919
rect -1649 -12595 -1596 -12542
rect -1114 -10961 -1061 -10908
rect -1293 -11581 -1240 -11528
rect -1381 -11972 -1328 -11919
rect -1203 -11972 -1150 -11919
rect -1294 -12707 -1241 -12654
rect -758 -10961 -705 -10908
rect -937 -11581 -884 -11528
rect -1025 -11972 -972 -11919
rect -848 -11972 -795 -11919
rect -937 -12836 -884 -12783
rect -402 -10961 -349 -10908
rect -46 -10961 7 -10908
rect 309 -10961 362 -10908
rect 665 -10961 718 -10908
rect 931 -10961 984 -10908
rect 1199 -10961 1252 -10908
rect -580 -11690 -527 -11637
rect -670 -11972 -617 -11919
rect -492 -11972 -439 -11919
rect -582 -12706 -529 -12653
rect -224 -11810 -171 -11757
rect -314 -11972 -261 -11919
rect -136 -11972 -83 -11919
rect -224 -12836 -171 -12783
rect 131 -11810 184 -11757
rect 42 -11972 95 -11919
rect 220 -11972 273 -11919
rect 130 -12706 183 -12653
rect -2004 -13598 -1951 -13545
rect -1648 -13725 -1595 -13672
rect -581 -13598 -528 -13545
rect -1291 -13725 -1238 -13672
rect -937 -13725 -884 -13672
rect -225 -13847 -172 -13794
rect 487 -11810 540 -11757
rect 399 -11972 452 -11919
rect 577 -11972 630 -11919
rect 486 -12837 539 -12784
rect 1556 -10961 1609 -10908
rect 1377 -11581 1430 -11528
rect 1288 -11972 1341 -11919
rect 1468 -11972 1521 -11919
rect 1378 -12836 1431 -12783
rect 1913 -10961 1966 -10908
rect 1733 -11581 1786 -11528
rect 1644 -11973 1697 -11920
rect 1823 -11972 1876 -11919
rect 1735 -12707 1788 -12654
rect 2268 -10961 2321 -10908
rect 2623 -10961 2676 -10908
rect 2980 -10961 3033 -10908
rect 3335 -10961 3388 -10908
rect 2089 -11581 2142 -11528
rect 2000 -11972 2053 -11919
rect 2178 -11972 2231 -11919
rect 2088 -12835 2141 -12782
rect 2446 -11690 2499 -11637
rect 2357 -11972 2410 -11919
rect 2534 -11972 2587 -11919
rect 2445 -12706 2498 -12653
rect 2800 -11810 2853 -11757
rect 2713 -11972 2766 -11919
rect 2890 -11972 2943 -11919
rect 2801 -12835 2854 -12782
rect 3157 -11810 3210 -11757
rect 3068 -11972 3121 -11919
rect 3247 -11972 3300 -11919
rect 3158 -12705 3211 -12652
rect 133 -13847 186 -13794
rect 487 -13848 540 -13795
rect 1379 -13725 1432 -13672
rect 1732 -13725 1785 -13672
rect 2091 -13725 2144 -13672
rect 2446 -13598 2499 -13545
rect 2802 -13847 2855 -13794
rect 3692 -10961 3745 -10908
rect 3513 -11810 3566 -11757
rect 3425 -11972 3478 -11919
rect 3603 -11972 3656 -11919
rect 3514 -12595 3567 -12542
rect 3871 -11691 3924 -11638
rect 3781 -11972 3834 -11919
rect 3871 -12595 3924 -12542
rect 3157 -13848 3210 -13795
rect 3870 -13598 3923 -13545
rect 3512 -13847 3565 -13794
rect -2315 -14596 -2262 -14543
rect -2447 -15874 -2394 -15821
rect -2005 -15875 -1952 -15822
rect -1915 -15986 -1862 -15933
rect -3935 -16347 -3883 -16295
rect -5682 -16939 -5629 -16886
rect -6159 -17060 -6106 -17007
rect -5859 -17060 -5806 -17007
rect -5326 -16939 -5273 -16886
rect -4970 -16939 -4917 -16886
rect -5148 -17060 -5095 -17007
rect -5504 -17171 -5451 -17118
rect -4614 -16939 -4561 -16886
rect -4258 -16939 -4205 -16886
rect -4437 -17060 -4384 -17007
rect -1917 -16595 -1864 -16542
rect -1649 -15875 -1596 -15822
rect -1738 -15986 -1685 -15933
rect -1560 -15986 -1507 -15933
rect -1738 -16595 -1685 -16542
rect -1561 -16594 -1508 -16541
rect -1827 -16718 -1774 -16665
rect -1720 -16718 -1548 -16665
rect -1381 -14596 -1328 -14543
rect -1204 -14596 -1151 -14543
rect -1293 -15875 -1240 -15822
rect -1382 -15986 -1329 -15933
rect -1204 -15986 -1151 -15933
rect -1381 -16596 -1328 -16543
rect -1204 -16595 -1151 -16542
rect -1026 -14596 -973 -14543
rect -848 -14596 -795 -14543
rect -847 -14979 -794 -14926
rect -937 -15875 -884 -15822
rect -1025 -15986 -972 -15933
rect -847 -15986 -794 -15933
rect -1026 -16595 -973 -16542
rect -669 -14596 -616 -14543
rect -669 -14979 -616 -14926
rect -491 -14596 -438 -14543
rect -491 -14979 -438 -14926
rect -581 -15875 -528 -15822
rect -670 -15986 -617 -15933
rect -491 -15986 -438 -15933
rect -4792 -17171 -4739 -17118
rect -3935 -17170 -3883 -17118
rect -1471 -16719 -1418 -16666
rect -1114 -16718 -1061 -16665
rect -759 -16717 -706 -16664
rect -314 -14980 -261 -14927
rect -137 -14979 -84 -14926
rect -225 -15875 -172 -15822
rect -313 -15986 -260 -15933
rect -136 -15986 -83 -15933
rect 43 -14979 96 -14926
rect 132 -15874 185 -15821
rect 43 -15986 96 -15933
rect 221 -15986 274 -15933
rect 220 -16595 273 -16542
rect -646 -16718 -471 -16665
rect -403 -16718 -350 -16665
rect -47 -16718 6 -16665
rect 487 -15875 540 -15822
rect 398 -15986 451 -15933
rect 575 -15986 628 -15933
rect 397 -16595 450 -16542
rect 576 -16595 629 -16542
rect 843 -15875 896 -15822
rect 755 -15986 808 -15933
rect 931 -15986 984 -15933
rect 755 -16595 808 -16542
rect 933 -16595 986 -16542
rect 1288 -14596 1341 -14543
rect 1289 -14980 1342 -14927
rect 1201 -15875 1254 -15822
rect 1110 -15986 1163 -15933
rect 1289 -15986 1342 -15933
rect 1111 -16595 1164 -16542
rect 1466 -14596 1519 -14543
rect 1467 -14979 1520 -14926
rect 1644 -14596 1697 -14543
rect 1644 -14979 1697 -14926
rect 1555 -15875 1608 -15822
rect 1466 -15986 1519 -15933
rect 1643 -15986 1696 -15933
rect 1823 -14595 1876 -14542
rect 1822 -14979 1875 -14926
rect 2000 -14596 2053 -14543
rect 1999 -14979 2052 -14926
rect 1910 -15875 1963 -15822
rect 1822 -15986 1875 -15933
rect 2000 -15986 2053 -15933
rect 2178 -14596 2231 -14543
rect 2180 -14979 2233 -14926
rect 2267 -15875 2320 -15822
rect 2179 -15986 2232 -15933
rect 2356 -15986 2409 -15933
rect 2356 -16595 2409 -16542
rect 309 -16719 362 -16666
rect 426 -16718 595 -16665
rect 665 -16718 718 -16665
rect 1021 -16718 1074 -16665
rect 1377 -16718 1430 -16665
rect 1501 -16718 1671 -16665
rect 1735 -16718 1788 -16665
rect 2090 -16717 2143 -16664
rect 2624 -15875 2677 -15822
rect 2534 -15986 2587 -15933
rect 2712 -15986 2765 -15933
rect 2534 -16595 2587 -16542
rect 2713 -16594 2766 -16541
rect 2979 -15875 3032 -15822
rect 2891 -15986 2944 -15933
rect 3068 -15986 3121 -15933
rect 2891 -16595 2944 -16542
rect 3070 -16595 3123 -16542
rect 3246 -14597 3299 -14544
rect 3424 -14596 3477 -14543
rect 3425 -14979 3478 -14926
rect 3335 -15875 3388 -15822
rect 3247 -15986 3300 -15933
rect 3424 -15986 3477 -15933
rect 3249 -16595 3302 -16542
rect 2445 -16718 2498 -16665
rect 2568 -16718 2732 -16665
rect 2801 -16718 2854 -16665
rect 3157 -16717 3210 -16664
rect 3602 -14596 3655 -14543
rect 3603 -14979 3656 -14926
rect 3781 -14596 3834 -14543
rect 3780 -14979 3833 -14926
rect 5184 -7908 5237 -7855
rect 5337 -7903 5390 -7850
rect 5185 -8687 5237 -8635
rect 11054 -8769 11107 -8716
rect 11345 -8769 11398 -8716
rect 11638 -8769 11691 -8716
rect 11932 -8769 11985 -8716
rect 12222 -8769 12275 -8716
rect 6769 -9367 6822 -9314
rect 6679 -9598 6732 -9545
rect 5337 -9978 5390 -9925
rect 6680 -10366 6733 -10313
rect 6947 -9368 7000 -9315
rect 7126 -9368 7179 -9315
rect 6858 -10520 6911 -10467
rect 7303 -9366 7356 -9313
rect 7214 -10519 7267 -10466
rect 7037 -11419 7090 -11366
rect 7482 -9366 7535 -9313
rect 7659 -9368 7712 -9315
rect 7571 -10519 7624 -10466
rect 7393 -11419 7446 -11366
rect 7837 -9367 7890 -9314
rect 8015 -9368 8068 -9315
rect 7927 -10519 7980 -10466
rect 7748 -11420 7801 -11367
rect 8194 -9367 8247 -9314
rect 8371 -9367 8424 -9314
rect 8283 -10520 8336 -10467
rect 8103 -11419 8156 -11366
rect 8549 -9367 8602 -9314
rect 8727 -9368 8780 -9315
rect 8638 -10519 8691 -10466
rect 8461 -11419 8514 -11366
rect 8906 -9367 8959 -9314
rect 11144 -9427 11197 -9374
rect 11436 -9428 11489 -9375
rect 11728 -9428 11781 -9375
rect 12020 -9429 12073 -9376
rect 12312 -9428 12365 -9375
rect 9171 -10367 9224 -10314
rect 8995 -10520 9048 -10467
rect 8817 -11419 8870 -11366
rect 11053 -11727 11106 -11674
rect 11347 -11728 11400 -11675
rect 11638 -11727 11691 -11674
rect 11931 -11727 11984 -11674
rect 12223 -11727 12276 -11674
rect 13022 -11726 13075 -11673
rect 5037 -13349 5090 -13296
rect 5534 -13349 5587 -13296
rect 5031 -13486 5084 -13433
rect 4905 -14598 4958 -14545
rect 4239 -14979 4292 -14926
rect 3692 -15875 3745 -15822
rect 3603 -15986 3656 -15933
rect 3780 -15986 3833 -15933
rect 4238 -15592 4291 -15539
rect 5400 -13598 5453 -13545
rect 5142 -13847 5195 -13794
rect 5143 -14711 5196 -14658
rect 5031 -15593 5084 -15540
rect 4238 -16595 4291 -16542
rect 3514 -16719 3567 -16666
rect 3633 -16718 3804 -16665
rect 3868 -16718 3921 -16665
rect 5534 -13725 5587 -13672
rect 8950 -13486 9003 -13433
rect 9305 -13486 9358 -13433
rect 8772 -13609 8825 -13556
rect 7526 -13725 7579 -13672
rect 7348 -13849 7401 -13796
rect 5833 -13975 5886 -13922
rect 6013 -13975 6066 -13922
rect 6190 -13976 6243 -13923
rect 6369 -13975 6422 -13922
rect 6547 -13976 6600 -13923
rect 6725 -13975 6778 -13922
rect 6902 -13975 6955 -13922
rect 5746 -14598 5799 -14545
rect 5924 -14711 5977 -14658
rect 6101 -14598 6154 -14545
rect 6279 -14711 6332 -14658
rect 6459 -14598 6512 -14545
rect 6813 -14598 6866 -14545
rect 6636 -14711 6689 -14658
rect 6991 -14711 7044 -14658
rect 5745 -15592 5798 -15539
rect 5400 -15706 5453 -15653
rect 5747 -15803 5800 -15750
rect 5923 -15705 5976 -15652
rect 5921 -16001 5974 -15948
rect 6101 -15592 6154 -15539
rect 6101 -15802 6154 -15749
rect 6279 -15705 6332 -15652
rect 6279 -16001 6332 -15948
rect 6458 -15592 6511 -15539
rect 6456 -15803 6509 -15750
rect 7437 -13975 7490 -13922
rect 6993 -14877 7046 -14824
rect 7347 -14877 7400 -14824
rect 6635 -15705 6688 -15652
rect 6713 -15804 6766 -15751
rect 6634 -16001 6687 -15948
rect 6813 -15904 6866 -15851
rect 7080 -14976 7133 -14923
rect 7260 -14977 7313 -14924
rect 7439 -14976 7492 -14923
rect 7882 -13726 7935 -13673
rect 8238 -13724 8291 -13671
rect 7704 -13848 7757 -13795
rect 7615 -13975 7668 -13922
rect 7793 -13976 7846 -13923
rect 8061 -13849 8114 -13796
rect 7970 -13975 8023 -13922
rect 8148 -13975 8201 -13922
rect 8415 -13849 8468 -13796
rect 8326 -13975 8379 -13922
rect 8861 -13975 8914 -13922
rect 9127 -13609 9180 -13556
rect 9038 -13975 9091 -13922
rect 9217 -13975 9270 -13922
rect 9483 -13609 9536 -13556
rect 9394 -13975 9447 -13922
rect 11442 -13725 11495 -13672
rect 11798 -13725 11851 -13672
rect 11264 -13849 11317 -13796
rect 9929 -13976 9982 -13923
rect 10108 -13975 10161 -13922
rect 10284 -13976 10337 -13923
rect 10462 -13976 10515 -13923
rect 10640 -13975 10693 -13922
rect 10819 -13976 10872 -13923
rect 7704 -14878 7757 -14825
rect 8236 -14598 8289 -14545
rect 8060 -14874 8113 -14821
rect 7169 -15803 7222 -15750
rect 7169 -15905 7222 -15852
rect 6994 -16004 7047 -15951
rect 7526 -15802 7579 -15749
rect 7526 -16006 7579 -15953
rect 7882 -15802 7935 -15749
rect 8060 -15904 8113 -15851
rect 8417 -14710 8470 -14657
rect 8327 -14976 8380 -14923
rect 7881 -16005 7934 -15952
rect 8237 -16005 8290 -15952
rect 6548 -16597 6601 -16544
rect 6726 -16597 6779 -16544
rect 6903 -16598 6956 -16545
rect 5399 -16720 5452 -16667
rect 5031 -16835 5084 -16782
rect 7970 -16598 8023 -16545
rect 8149 -16597 8202 -16544
rect 8595 -14598 8648 -14545
rect 8504 -14859 8557 -14806
rect 8505 -14977 8558 -14924
rect 8772 -14711 8825 -14658
rect 8683 -14977 8736 -14924
rect 8950 -14599 9003 -14546
rect 9127 -14712 9180 -14659
rect 9304 -14598 9357 -14545
rect 9661 -14598 9714 -14545
rect 9483 -14711 9536 -14658
rect 9572 -14976 9625 -14923
rect 9837 -14712 9890 -14659
rect 9753 -14859 9806 -14806
rect 9750 -14976 9803 -14923
rect 10016 -14598 10069 -14545
rect 9929 -14976 9982 -14923
rect 10373 -14599 10426 -14546
rect 10196 -14711 10249 -14658
rect 10195 -14875 10248 -14822
rect 10550 -14711 10603 -14658
rect 10552 -14868 10605 -14815
rect 10729 -14598 10782 -14545
rect 10908 -14711 10961 -14658
rect 11087 -14711 11140 -14658
rect 10908 -14866 10961 -14813
rect 11353 -13975 11406 -13922
rect 11620 -13850 11673 -13797
rect 11530 -13975 11583 -13922
rect 11709 -13975 11762 -13922
rect 12152 -13726 12205 -13673
rect 12509 -13725 12562 -13672
rect 11977 -13849 12030 -13796
rect 11886 -13976 11939 -13923
rect 12064 -13975 12117 -13922
rect 12334 -13849 12387 -13796
rect 12242 -13976 12295 -13923
rect 12420 -13975 12473 -13922
rect 11440 -14709 11493 -14656
rect 10819 -14976 10872 -14923
rect 8593 -15905 8646 -15852
rect 9663 -15905 9716 -15852
rect 8771 -16719 8824 -16666
rect 9128 -16719 9181 -16666
rect 10373 -15804 10426 -15751
rect 10194 -15905 10247 -15852
rect 10730 -15803 10783 -15750
rect 11264 -14868 11317 -14815
rect 10996 -14976 11049 -14923
rect 11175 -14976 11228 -14923
rect 11086 -15803 11139 -15750
rect 11619 -15705 11672 -15652
rect 11084 -15905 11137 -15852
rect 11440 -15894 11493 -15841
rect 9484 -16719 9537 -16666
rect 8950 -16835 9003 -16782
rect 9305 -16835 9358 -16782
rect 7347 -16943 7400 -16890
rect 7704 -16943 7757 -16890
rect 8060 -16943 8113 -16890
rect 8416 -16943 8469 -16890
rect 9929 -16597 9982 -16544
rect 9838 -16719 9891 -16666
rect 10107 -16598 10160 -16545
rect 10287 -16598 10340 -16545
rect 10195 -16718 10248 -16665
rect 10550 -16718 10603 -16665
rect 11441 -16005 11494 -15952
rect 11798 -15593 11851 -15540
rect 11797 -16005 11850 -15952
rect 11975 -15705 12028 -15652
rect 12155 -15592 12208 -15539
rect 12154 -16005 12207 -15952
rect 12332 -15705 12385 -15652
rect 12511 -15592 12564 -15539
rect 12511 -16005 12564 -15952
rect 10907 -16718 10960 -16665
rect 10017 -16834 10070 -16781
rect 10374 -16834 10427 -16781
rect 10731 -16832 10784 -16779
rect 11352 -16598 11405 -16545
rect 11530 -16599 11583 -16546
rect 11709 -16598 11762 -16545
rect 11263 -16943 11316 -16890
rect 11620 -16943 11673 -16890
rect 11975 -16942 12028 -16889
rect 12331 -16942 12384 -16889
rect 18337 -13496 18412 -13421
<< metal2 >>
rect -5867 -1910 -5814 -1900
rect -5689 -1910 -5636 -1900
rect -5510 -1910 -5457 -1900
rect -5333 -1910 -5280 -1900
rect -5155 -1910 -5102 -1900
rect -4976 -1910 -4923 -1900
rect -4799 -1910 -4746 -1900
rect -4621 -1910 -4568 -1900
rect -4443 -1910 -4390 -1900
rect -4265 -1910 -4212 -1900
rect -4086 -1910 -4033 -1900
rect -3909 -1910 -3856 -1900
rect -1109 -1910 -1056 -1900
rect -5814 -1963 -5689 -1910
rect -5636 -1963 -5510 -1910
rect -5457 -1963 -5333 -1910
rect -5280 -1963 -5155 -1910
rect -5102 -1963 -4976 -1910
rect -4923 -1963 -4799 -1910
rect -4746 -1963 -4621 -1910
rect -4568 -1963 -4443 -1910
rect -4390 -1963 -4265 -1910
rect -4212 -1963 -4086 -1910
rect -4033 -1963 -3909 -1910
rect -3856 -1963 -1109 -1910
rect -5867 -1973 -5814 -1963
rect -5689 -1973 -5636 -1963
rect -5510 -1973 -5457 -1963
rect -5333 -1973 -5280 -1963
rect -5155 -1973 -5102 -1963
rect -4976 -1973 -4923 -1963
rect -4799 -1973 -4746 -1963
rect -4621 -1973 -4568 -1963
rect -4443 -1973 -4390 -1963
rect -4265 -1973 -4212 -1963
rect -4086 -1973 -4033 -1963
rect -3909 -1973 -3856 -1963
rect -1109 -1973 -1056 -1963
rect 5337 -2205 5390 -2195
rect 6680 -2199 6744 -2189
rect 5390 -2258 6680 -2205
rect 5337 -2268 5390 -2258
rect 6744 -2258 6748 -2205
rect 6680 -2273 6744 -2263
rect -1109 -2425 -1056 -2415
rect -752 -2425 -699 -2415
rect -1056 -2478 -752 -2425
rect -1109 -2488 -1056 -2478
rect -752 -2488 -699 -2478
rect 1919 -2426 1972 -2416
rect 2275 -2426 2328 -2416
rect 3193 -2426 3246 -2417
rect 1972 -2479 2275 -2426
rect 2328 -2427 3246 -2426
rect 2328 -2479 3193 -2427
rect 1919 -2489 1972 -2479
rect 2275 -2489 2328 -2479
rect 3193 -2490 3246 -2480
rect -6498 -2529 -6445 -2519
rect -5777 -2529 -5724 -2520
rect -6445 -2530 -5724 -2529
rect -5066 -2530 -5013 -2520
rect -4354 -2530 -4301 -2520
rect -6445 -2582 -5777 -2530
rect -6498 -2592 -6445 -2582
rect -5724 -2583 -5066 -2530
rect -5013 -2583 -4354 -2530
rect -5777 -2593 -5724 -2583
rect -5066 -2593 -5013 -2583
rect -4354 -2593 -4301 -2583
rect -2624 -2558 -2571 -2548
rect -1285 -2558 -1232 -2548
rect -930 -2558 -877 -2548
rect -2571 -2611 -1285 -2558
rect -1232 -2611 -930 -2558
rect -2624 -2621 -2571 -2611
rect -1285 -2621 -1232 -2611
rect -930 -2621 -877 -2611
rect 2097 -2554 2150 -2544
rect 2453 -2554 2506 -2544
rect 2150 -2607 2453 -2554
rect 2097 -2617 2150 -2607
rect 2453 -2617 2506 -2607
rect -5421 -2668 -5368 -2658
rect -4710 -2668 -4657 -2658
rect -3998 -2668 -3945 -2658
rect -3298 -2668 -3245 -2658
rect -5368 -2721 -4710 -2668
rect -4657 -2721 -3998 -2668
rect -3945 -2721 -3298 -2668
rect -5421 -2731 -5368 -2721
rect -4710 -2731 -4657 -2721
rect -3998 -2731 -3945 -2721
rect -3298 -2731 -3245 -2721
rect -1197 -2665 -1144 -2655
rect -1019 -2665 -966 -2655
rect -841 -2665 -788 -2655
rect -129 -2665 -76 -2655
rect 50 -2665 103 -2655
rect 227 -2665 280 -2655
rect 940 -2665 993 -2655
rect 1117 -2665 1170 -2655
rect 1295 -2665 1348 -2655
rect 2007 -2665 2060 -2655
rect 2186 -2665 2239 -2655
rect 2363 -2665 2416 -2655
rect -1144 -2718 -1019 -2665
rect -966 -2718 -841 -2665
rect -788 -2718 -129 -2665
rect -76 -2718 50 -2665
rect 103 -2718 227 -2665
rect 280 -2718 940 -2665
rect 993 -2718 1117 -2665
rect 1170 -2718 1295 -2665
rect 1348 -2718 2007 -2665
rect 2060 -2718 2186 -2665
rect 2239 -2718 2363 -2665
rect -1197 -2728 -1144 -2718
rect -1019 -2728 -966 -2718
rect -841 -2728 -788 -2718
rect -129 -2728 -76 -2718
rect 50 -2728 103 -2718
rect 227 -2728 280 -2718
rect 940 -2728 993 -2718
rect 1117 -2728 1170 -2718
rect 1295 -2728 1348 -2718
rect 2007 -2728 2060 -2718
rect 2186 -2728 2239 -2718
rect 2363 -2728 2416 -2718
rect -6044 -2780 -5991 -2770
rect -5866 -2780 -5813 -2770
rect -5991 -2833 -5866 -2780
rect -6044 -2843 -5991 -2833
rect -5866 -2843 -5813 -2833
rect -3908 -2780 -3855 -2770
rect -3731 -2780 -3678 -2770
rect -3855 -2833 -3731 -2780
rect -3908 -2843 -3855 -2833
rect -3731 -2843 -3678 -2833
rect -484 -3301 -431 -3291
rect 583 -3301 636 -3291
rect 1654 -3301 1707 -3291
rect -431 -3354 583 -3301
rect 636 -3354 1654 -3301
rect -484 -3364 -431 -3354
rect 583 -3364 636 -3354
rect 1654 -3364 1707 -3354
rect -6625 -3401 -6572 -3391
rect -6134 -3401 -6081 -3391
rect -5066 -3401 -5013 -3391
rect -6572 -3454 -6134 -3401
rect -6081 -3454 -5066 -3401
rect -6625 -3464 -6572 -3454
rect -6134 -3464 -6081 -3454
rect -5066 -3464 -5013 -3454
rect -4710 -3401 -4657 -3391
rect -3642 -3401 -3589 -3391
rect -3131 -3401 -3078 -3391
rect -4657 -3454 -3642 -3401
rect -3589 -3454 -3131 -3401
rect -4710 -3464 -4657 -3454
rect -3642 -3464 -3589 -3454
rect -3131 -3464 -3078 -3454
rect -1645 -3449 -1584 -3439
rect -5777 -3516 -5724 -3506
rect -3998 -3516 -3945 -3506
rect -3298 -3516 -3245 -3506
rect -5724 -3569 -3998 -3516
rect -3945 -3569 -3298 -3516
rect -1108 -3456 -1055 -3446
rect -750 -3456 -697 -3446
rect -396 -3456 -343 -3446
rect -39 -3456 14 -3446
rect 317 -3456 370 -3446
rect -1584 -3509 -1108 -3456
rect -1055 -3509 -750 -3456
rect -697 -3509 -396 -3456
rect -343 -3509 -39 -3456
rect 14 -3509 317 -3456
rect -1645 -3520 -1584 -3510
rect -1108 -3519 -1055 -3509
rect -750 -3519 -697 -3509
rect -396 -3519 -343 -3509
rect -39 -3519 14 -3509
rect 317 -3519 370 -3509
rect 850 -3456 903 -3446
rect 1206 -3456 1259 -3446
rect 1562 -3456 1615 -3446
rect 1919 -3456 1972 -3446
rect 2275 -3456 2328 -3446
rect 3019 -3452 3080 -3442
rect 903 -3509 1206 -3456
rect 1259 -3509 1562 -3456
rect 1615 -3509 1919 -3456
rect 1972 -3509 2275 -3456
rect 2328 -3509 3019 -3456
rect 850 -3519 903 -3509
rect 1206 -3519 1259 -3509
rect 1562 -3519 1615 -3509
rect 1919 -3519 1972 -3509
rect 2275 -3519 2328 -3509
rect 6222 -3451 6286 -3441
rect 3080 -3509 6222 -3456
rect 3019 -3523 3080 -3513
rect 6286 -3509 6297 -3456
rect 6222 -3525 6286 -3515
rect -5777 -3579 -5724 -3569
rect -3998 -3579 -3945 -3569
rect -3298 -3579 -3245 -3569
rect -1286 -3571 -1233 -3561
rect -929 -3571 -876 -3561
rect -573 -3571 -520 -3561
rect -217 -3571 -164 -3561
rect -1702 -3624 -1286 -3571
rect -1233 -3624 -929 -3571
rect -876 -3624 -573 -3571
rect -520 -3624 -217 -3571
rect -6498 -3640 -6445 -3630
rect -5422 -3640 -5369 -3630
rect -4353 -3640 -4300 -3630
rect -1702 -3640 -1649 -3624
rect -1286 -3634 -1233 -3624
rect -929 -3634 -876 -3624
rect -573 -3634 -520 -3624
rect -217 -3634 -164 -3624
rect 1384 -3564 1437 -3554
rect 1741 -3564 1794 -3554
rect 2097 -3564 2150 -3554
rect 2451 -3564 2504 -3554
rect 1437 -3617 1741 -3564
rect 1794 -3617 2097 -3564
rect 2150 -3617 2451 -3564
rect 1384 -3627 1437 -3617
rect 1741 -3627 1794 -3617
rect 2097 -3627 2150 -3617
rect 2451 -3627 2504 -3617
rect -6445 -3693 -5422 -3640
rect -5369 -3693 -4353 -3640
rect -4300 -3693 -1649 -3640
rect -6498 -3703 -6445 -3693
rect -5422 -3703 -5369 -3693
rect -4353 -3703 -4300 -3693
rect -2546 -3928 -2485 -3693
rect -2546 -3999 -2485 -3989
rect -841 -4192 -788 -4182
rect -662 -4192 -609 -4182
rect -483 -4192 -430 -4182
rect -306 -4192 -253 -4182
rect 407 -4192 460 -4182
rect 583 -4192 636 -4182
rect 761 -4192 814 -4182
rect 1474 -4192 1527 -4182
rect 1652 -4192 1705 -4182
rect 1830 -4192 1883 -4182
rect 2008 -4192 2061 -4182
rect -788 -4245 -662 -4192
rect -609 -4245 -483 -4192
rect -430 -4245 -306 -4192
rect -253 -4245 407 -4192
rect 460 -4245 583 -4192
rect 636 -4245 761 -4192
rect 814 -4245 1474 -4192
rect 1527 -4245 1652 -4192
rect 1705 -4245 1830 -4192
rect 1883 -4245 2008 -4192
rect -841 -4255 -788 -4245
rect -662 -4255 -609 -4245
rect -483 -4255 -430 -4245
rect -306 -4255 -253 -4245
rect 407 -4255 460 -4245
rect 583 -4255 636 -4245
rect 761 -4255 814 -4245
rect 1474 -4255 1527 -4245
rect 1652 -4255 1705 -4245
rect 1830 -4255 1883 -4245
rect 2008 -4255 2061 -4245
rect -6498 -4271 -6445 -4261
rect -5778 -4271 -5725 -4261
rect -3998 -4271 -3945 -4261
rect -6445 -4324 -5778 -4271
rect -5725 -4324 -3998 -4271
rect 2538 -4266 2599 -4256
rect 317 -4304 370 -4294
rect 673 -4304 726 -4294
rect -6498 -4334 -6445 -4324
rect -5778 -4334 -5725 -4324
rect -3998 -4334 -3945 -4324
rect -2357 -4357 317 -4304
rect 370 -4357 673 -4304
rect 2538 -4337 2599 -4327
rect -6134 -4390 -6081 -4380
rect -5066 -4390 -5013 -4380
rect -4709 -4390 -4656 -4380
rect -3642 -4390 -3589 -4380
rect -2357 -4390 -2304 -4357
rect 317 -4367 370 -4357
rect 673 -4367 726 -4357
rect -6081 -4443 -5066 -4390
rect -5013 -4443 -4709 -4390
rect -4656 -4443 -3642 -4390
rect -3589 -4443 -2304 -4390
rect -2004 -4412 -1951 -4402
rect 495 -4412 548 -4402
rect 850 -4412 903 -4402
rect -6134 -4453 -6081 -4443
rect -5066 -4453 -5013 -4443
rect -4709 -4453 -4656 -4443
rect -3642 -4453 -3589 -4443
rect -1951 -4465 495 -4412
rect 548 -4465 850 -4412
rect -2004 -4475 -1951 -4465
rect 495 -4475 548 -4465
rect 850 -4475 903 -4465
rect 2746 -4446 2807 -4436
rect -5422 -4506 -5369 -4496
rect -4353 -4506 -4300 -4496
rect -3298 -4506 -3245 -4496
rect -2385 -4505 -2324 -4495
rect -5369 -4559 -4353 -4506
rect -4300 -4559 -3298 -4506
rect -3245 -4559 -2385 -4506
rect -5422 -4569 -5369 -4559
rect -4353 -4569 -4300 -4559
rect -3298 -4569 -3245 -4559
rect 2746 -4517 2807 -4507
rect -2385 -4576 -2324 -4566
rect 3194 -4805 3246 -4795
rect 4771 -4805 4823 -4795
rect 3246 -4857 4771 -4805
rect 3194 -4867 3246 -4857
rect 4771 -4867 4823 -4857
rect 3021 -5002 3082 -4992
rect 5037 -5006 5090 -4996
rect 4985 -5007 5037 -5006
rect 3082 -5059 5037 -5007
rect 3021 -5073 3082 -5063
rect 5037 -5069 5090 -5059
rect -2385 -5093 -2324 -5083
rect -6498 -5141 -6445 -5131
rect -5422 -5141 -5369 -5131
rect -6445 -5187 -5422 -5147
rect -6498 -5204 -6445 -5194
rect -4353 -5141 -4300 -5131
rect -5369 -5188 -4353 -5148
rect -5422 -5204 -5369 -5194
rect -1287 -5097 -1234 -5087
rect -929 -5097 -876 -5087
rect -572 -5097 -519 -5087
rect -218 -5097 -165 -5087
rect -2324 -5150 -1287 -5097
rect -1234 -5150 -929 -5097
rect -876 -5150 -572 -5097
rect -519 -5150 -218 -5097
rect 1385 -5093 1438 -5083
rect 1740 -5093 1793 -5083
rect 2096 -5093 2149 -5083
rect 2453 -5093 2506 -5083
rect -2385 -5164 -2324 -5154
rect -1287 -5160 -1234 -5150
rect -929 -5160 -876 -5150
rect -572 -5160 -519 -5150
rect -218 -5160 -165 -5150
rect 311 -5148 372 -5138
rect -4353 -5204 -4300 -5194
rect -1105 -5213 -1052 -5203
rect -751 -5213 -698 -5203
rect -396 -5213 -343 -5203
rect -41 -5213 12 -5203
rect 1438 -5146 1740 -5093
rect 1793 -5146 2096 -5093
rect 2149 -5146 2453 -5093
rect 1385 -5156 1438 -5146
rect 1740 -5156 1793 -5146
rect 2096 -5156 2149 -5146
rect 2453 -5156 2506 -5146
rect 311 -5213 372 -5209
rect -6134 -5232 -6081 -5222
rect -5066 -5233 -5013 -5223
rect -6081 -5279 -5066 -5239
rect -6134 -5295 -6081 -5285
rect -3130 -5233 -3077 -5223
rect -5013 -5279 -3130 -5239
rect -5066 -5296 -5013 -5286
rect -1876 -5232 -1823 -5222
rect -3077 -5279 -1876 -5239
rect -3130 -5296 -3077 -5286
rect -1052 -5266 -751 -5213
rect -698 -5266 -396 -5213
rect -343 -5266 -41 -5213
rect 12 -5266 316 -5213
rect 369 -5219 372 -5213
rect 846 -5213 903 -5203
rect 1207 -5213 1260 -5203
rect 1563 -5213 1616 -5203
rect 1917 -5213 1970 -5203
rect 2274 -5213 2327 -5203
rect 4905 -5212 4958 -5202
rect -1876 -5295 -1823 -5285
rect -1646 -5278 -1585 -5268
rect -1105 -5276 -1052 -5266
rect -751 -5276 -698 -5266
rect -396 -5276 -343 -5266
rect -41 -5276 12 -5266
rect 316 -5276 369 -5266
rect 846 -5266 850 -5213
rect 903 -5266 1207 -5213
rect 1260 -5266 1563 -5213
rect 1616 -5266 1917 -5213
rect 1970 -5266 2274 -5213
rect 2327 -5265 4905 -5213
rect 5614 -5207 5678 -5197
rect 4958 -5265 5614 -5213
rect 2327 -5266 5614 -5265
rect -6625 -5322 -6572 -5312
rect -4710 -5322 -4657 -5312
rect -6572 -5369 -4710 -5329
rect -6625 -5385 -6572 -5375
rect -3642 -5319 -3589 -5309
rect -4657 -5369 -3642 -5329
rect -4710 -5385 -4657 -5375
rect -2624 -5324 -2571 -5314
rect -3589 -5369 -2624 -5329
rect -3642 -5382 -3589 -5372
rect -1646 -5349 -1585 -5339
rect 846 -5278 907 -5266
rect 1207 -5276 1260 -5266
rect 1563 -5276 1616 -5266
rect 1917 -5276 1970 -5266
rect 2274 -5276 2327 -5266
rect 4905 -5275 4958 -5266
rect 5678 -5266 5685 -5213
rect 5614 -5281 5678 -5271
rect 846 -5349 907 -5339
rect -2624 -5387 -2571 -5377
rect -128 -5380 -75 -5370
rect 50 -5380 103 -5370
rect 228 -5380 281 -5370
rect 940 -5380 993 -5371
rect 1119 -5380 1172 -5370
rect 1296 -5380 1349 -5370
rect -5777 -5415 -5724 -5405
rect -3997 -5415 -3944 -5405
rect -5724 -5462 -3997 -5422
rect -5777 -5478 -5724 -5468
rect -3298 -5416 -3245 -5406
rect -3944 -5462 -3298 -5422
rect -3997 -5478 -3944 -5468
rect -75 -5433 50 -5380
rect 103 -5433 228 -5380
rect 281 -5381 1119 -5380
rect 281 -5433 940 -5381
rect -128 -5443 -75 -5433
rect 50 -5443 103 -5433
rect 228 -5443 281 -5433
rect 993 -5433 1119 -5381
rect 1172 -5433 1296 -5380
rect 940 -5444 993 -5434
rect 1119 -5443 1172 -5433
rect 1296 -5443 1349 -5433
rect -3298 -5479 -3245 -5469
rect 5337 -5527 5390 -5517
rect -5956 -6016 -5903 -6006
rect -5601 -6016 -5548 -6006
rect -5244 -6016 -5191 -6006
rect -4888 -6016 -4835 -6006
rect -4532 -6016 -4479 -6006
rect -4175 -6016 -4122 -6006
rect -3820 -6016 -3767 -6006
rect -5903 -6069 -5601 -6016
rect -5548 -6069 -5244 -6016
rect -5191 -6069 -4888 -6016
rect -4835 -6069 -4532 -6016
rect -4479 -6069 -4175 -6016
rect -4122 -6069 -3820 -6016
rect -5956 -6079 -5903 -6069
rect -5601 -6079 -5548 -6069
rect -5244 -6079 -5191 -6069
rect -4888 -6079 -4835 -6069
rect -4532 -6079 -4479 -6069
rect -4175 -6079 -4122 -6069
rect -3820 -6079 -3767 -6069
rect -2624 -6007 -2571 -5997
rect 2096 -6007 2149 -5997
rect 2452 -6007 2505 -5997
rect -2571 -6060 2096 -6007
rect 2149 -6060 2452 -6007
rect -2624 -6070 -2571 -6060
rect 2096 -6070 2149 -6060
rect 2452 -6070 2505 -6060
rect -5778 -6131 -5725 -6121
rect -5065 -6131 -5012 -6121
rect -4354 -6131 -4301 -6121
rect -3298 -6131 -3245 -6121
rect 1918 -6124 1971 -6114
rect 2275 -6124 2328 -6114
rect -2821 -6125 1918 -6124
rect -5725 -6184 -5065 -6131
rect -5012 -6184 -4354 -6131
rect -4301 -6184 -3298 -6131
rect -5778 -6194 -5725 -6184
rect -5065 -6194 -5012 -6184
rect -4354 -6194 -4301 -6184
rect -3298 -6194 -3245 -6184
rect -2856 -6177 1918 -6125
rect 1971 -6177 2275 -6124
rect -6498 -6248 -6445 -6238
rect -5421 -6248 -5368 -6238
rect -4710 -6248 -4657 -6238
rect -3998 -6247 -3945 -6237
rect -6445 -6301 -5421 -6248
rect -5368 -6301 -4710 -6248
rect -4657 -6300 -3998 -6248
rect -4657 -6301 -3945 -6300
rect -6498 -6311 -6445 -6301
rect -5421 -6311 -5368 -6301
rect -4710 -6311 -4657 -6301
rect -3998 -6310 -3945 -6301
rect -4786 -6378 -4733 -6368
rect -2856 -6401 -2803 -6177
rect 1918 -6187 1971 -6177
rect 2275 -6187 2328 -6177
rect -3874 -6408 -2803 -6401
rect -4733 -6431 -2803 -6408
rect -4786 -6454 -2803 -6431
rect -2702 -6250 -2649 -6249
rect 227 -6250 280 -6240
rect 942 -6250 995 -6240
rect -2702 -6303 227 -6250
rect 280 -6303 942 -6250
rect -4786 -6461 -3820 -6454
rect -3874 -7691 -3821 -6461
rect -2702 -6542 -2649 -6303
rect 227 -6313 280 -6303
rect 942 -6313 995 -6303
rect -1876 -6364 -1823 -6354
rect -1282 -6364 -1229 -6354
rect -1823 -6417 -1282 -6364
rect -1229 -6365 -1177 -6364
rect -928 -6365 -876 -6355
rect 2879 -6365 2931 -6355
rect -1229 -6417 -928 -6365
rect -876 -6417 2879 -6365
rect -1876 -6427 -1823 -6417
rect -1282 -6427 -1229 -6417
rect -928 -6427 -876 -6417
rect 2879 -6427 2931 -6417
rect -1110 -6479 -1057 -6469
rect -752 -6479 -699 -6469
rect -1057 -6532 -752 -6479
rect -1110 -6542 -1057 -6532
rect -752 -6542 -699 -6532
rect -3874 -7743 -3873 -7691
rect -3873 -7753 -3821 -7743
rect -3731 -6595 -2649 -6542
rect -3731 -7785 -3678 -6595
rect -753 -6598 -700 -6588
rect 4772 -6597 4825 -6587
rect -700 -6650 4772 -6598
rect -700 -6651 4825 -6650
rect -753 -6661 -700 -6651
rect 4772 -6660 4825 -6651
rect -2003 -6714 -1950 -6704
rect -1950 -6767 5237 -6714
rect -2003 -6777 -1950 -6767
rect -3545 -6806 -3484 -6796
rect -3545 -6877 -3484 -6867
rect -3679 -7837 -3678 -7785
rect -3541 -7788 -3489 -6877
rect 4770 -6891 4823 -6881
rect -3386 -6979 -3325 -6969
rect 4770 -6996 4823 -6944
rect 4906 -6889 4959 -6879
rect 4906 -6994 4959 -6942
rect -3386 -7050 -3325 -7040
rect -3731 -7847 -3679 -7837
rect -3541 -7850 -3489 -7840
rect -3382 -7933 -3329 -7050
rect 4771 -7844 4823 -6996
rect 4907 -7842 4959 -6994
rect 5038 -6887 5091 -6877
rect 5038 -7840 5091 -6940
rect 4771 -7854 4824 -7844
rect -1382 -7922 -1329 -7912
rect -1203 -7922 -1150 -7913
rect -1025 -7922 -972 -7912
rect -848 -7922 -795 -7912
rect -670 -7922 -617 -7912
rect -490 -7922 -437 -7912
rect 755 -7922 808 -7912
rect 932 -7922 985 -7912
rect 1112 -7922 1165 -7912
rect 1289 -7922 1342 -7913
rect 1467 -7922 1520 -7912
rect 1644 -7922 1697 -7912
rect 2890 -7922 2943 -7912
rect 3069 -7922 3122 -7912
rect 3247 -7922 3300 -7912
rect 3424 -7922 3477 -7912
rect 3603 -7922 3656 -7913
rect 3778 -7922 3831 -7912
rect -1329 -7923 -1025 -7922
rect -1329 -7975 -1203 -7923
rect -1382 -7985 -1329 -7975
rect -1150 -7975 -1025 -7923
rect -972 -7975 -848 -7922
rect -795 -7975 -670 -7922
rect -617 -7975 -490 -7922
rect -437 -7975 755 -7922
rect 808 -7975 932 -7922
rect 985 -7975 1112 -7922
rect 1165 -7923 1467 -7922
rect 1165 -7975 1289 -7923
rect -1203 -7986 -1150 -7976
rect -1025 -7985 -972 -7975
rect -848 -7985 -795 -7975
rect -670 -7985 -617 -7975
rect -490 -7985 -437 -7975
rect 755 -7985 808 -7975
rect 932 -7985 985 -7975
rect 1112 -7985 1165 -7975
rect 1342 -7975 1467 -7923
rect 1520 -7975 1644 -7922
rect 1697 -7975 2890 -7922
rect 2943 -7975 3069 -7922
rect 3122 -7975 3247 -7922
rect 3300 -7975 3424 -7922
rect 3477 -7923 3778 -7922
rect 3477 -7975 3603 -7923
rect 1289 -7986 1342 -7976
rect 1467 -7985 1520 -7975
rect 1644 -7985 1697 -7975
rect 2890 -7985 2943 -7975
rect 3069 -7985 3122 -7975
rect 3247 -7985 3300 -7975
rect 3424 -7985 3477 -7975
rect 3656 -7975 3778 -7923
rect 4208 -7923 4261 -7913
rect 4771 -7917 4824 -7907
rect 4906 -7852 4959 -7842
rect 4906 -7915 4959 -7905
rect 5037 -7850 5091 -7840
rect 5090 -7898 5091 -7850
rect 5184 -7855 5237 -6767
rect 5037 -7913 5090 -7903
rect 5184 -7918 5237 -7908
rect 5337 -7850 5390 -5580
rect 5337 -7913 5390 -7903
rect 17831 -6521 17895 -6511
rect 3831 -7975 4208 -7923
rect 3603 -7986 3656 -7976
rect 3778 -7976 4208 -7975
rect 3778 -7985 3831 -7976
rect 4208 -7986 4261 -7976
rect -3382 -7996 -3329 -7986
rect -1916 -8534 -1863 -8524
rect -1739 -8534 -1686 -8524
rect -1558 -8534 -1505 -8524
rect -1382 -8534 -1329 -8524
rect -1203 -8534 -1150 -8524
rect -1026 -8534 -973 -8524
rect -848 -8534 -795 -8524
rect -670 -8534 -617 -8524
rect -491 -8534 -438 -8524
rect -314 -8534 -261 -8524
rect -136 -8534 -83 -8524
rect 42 -8534 95 -8524
rect 221 -8534 274 -8524
rect 398 -8534 451 -8524
rect 577 -8534 630 -8524
rect 754 -8534 807 -8524
rect 932 -8534 985 -8524
rect 1111 -8534 1164 -8524
rect 1289 -8534 1342 -8524
rect 1466 -8534 1519 -8524
rect 1644 -8534 1697 -8524
rect 1822 -8534 1875 -8524
rect 2000 -8534 2053 -8524
rect 2178 -8534 2231 -8524
rect 2357 -8534 2410 -8524
rect 2534 -8534 2587 -8524
rect 2712 -8534 2765 -8524
rect 2890 -8534 2943 -8524
rect 3068 -8534 3121 -8524
rect 3246 -8534 3299 -8524
rect 3424 -8534 3477 -8524
rect 3602 -8534 3655 -8524
rect 3781 -8534 3834 -8524
rect -1863 -8587 -1739 -8534
rect -1686 -8587 -1558 -8534
rect -1505 -8587 -1382 -8534
rect -1329 -8587 -1203 -8534
rect -1150 -8587 -1026 -8534
rect -973 -8587 -848 -8534
rect -795 -8587 -670 -8534
rect -617 -8587 -491 -8534
rect -438 -8587 -314 -8534
rect -261 -8587 -136 -8534
rect -83 -8587 42 -8534
rect 95 -8587 221 -8534
rect 274 -8587 398 -8534
rect 451 -8587 577 -8534
rect 630 -8587 754 -8534
rect 807 -8587 932 -8534
rect 985 -8587 1111 -8534
rect 1164 -8587 1289 -8534
rect 1342 -8587 1466 -8534
rect 1519 -8587 1644 -8534
rect 1697 -8587 1822 -8534
rect 1875 -8587 2000 -8534
rect 2053 -8587 2178 -8534
rect 2231 -8587 2357 -8534
rect 2410 -8587 2534 -8534
rect 2587 -8587 2712 -8534
rect 2765 -8587 2890 -8534
rect 2943 -8587 3068 -8534
rect 3121 -8587 3246 -8534
rect 3299 -8587 3424 -8534
rect 3477 -8587 3602 -8534
rect 3655 -8587 3781 -8534
rect -1916 -8597 -1863 -8587
rect -1739 -8597 -1686 -8587
rect -1558 -8597 -1505 -8587
rect -1382 -8597 -1329 -8587
rect -1203 -8597 -1150 -8587
rect -1026 -8597 -973 -8587
rect -848 -8597 -795 -8587
rect -670 -8597 -617 -8587
rect -491 -8597 -438 -8587
rect -314 -8597 -261 -8587
rect -136 -8597 -83 -8587
rect 42 -8597 95 -8587
rect 221 -8597 274 -8587
rect 398 -8597 451 -8587
rect 577 -8597 630 -8587
rect 754 -8597 807 -8587
rect 932 -8597 985 -8587
rect 1111 -8597 1164 -8587
rect 1289 -8597 1342 -8587
rect 1466 -8597 1519 -8587
rect 1644 -8597 1697 -8587
rect 1822 -8597 1875 -8587
rect 2000 -8597 2053 -8587
rect 2178 -8597 2231 -8587
rect 2357 -8597 2410 -8587
rect 2534 -8597 2587 -8587
rect 2712 -8597 2765 -8587
rect 2890 -8597 2943 -8587
rect 3068 -8597 3121 -8587
rect 3246 -8597 3299 -8587
rect 3424 -8597 3477 -8587
rect 3602 -8597 3655 -8587
rect 3781 -8597 3834 -8587
rect 5185 -8633 5237 -8625
rect 5185 -8635 10564 -8633
rect -1826 -8653 -1773 -8643
rect -1470 -8653 -1417 -8643
rect -1115 -8653 -1062 -8643
rect -758 -8653 -705 -8643
rect -402 -8653 -349 -8643
rect -47 -8653 6 -8643
rect 310 -8653 363 -8643
rect 666 -8653 719 -8643
rect 1022 -8653 1075 -8643
rect 1377 -8653 1430 -8643
rect 1733 -8653 1786 -8643
rect 2090 -8653 2143 -8643
rect 2446 -8653 2499 -8643
rect 2802 -8653 2855 -8643
rect 3158 -8653 3211 -8643
rect 3513 -8653 3566 -8643
rect 3869 -8653 3922 -8643
rect -1773 -8706 -1470 -8653
rect -1417 -8706 -1115 -8653
rect -1062 -8706 -758 -8653
rect -705 -8706 -402 -8653
rect -349 -8706 -47 -8653
rect 6 -8706 310 -8653
rect 363 -8706 666 -8653
rect 719 -8706 1022 -8653
rect 1075 -8706 1377 -8653
rect 1430 -8706 1733 -8653
rect 1786 -8706 2090 -8653
rect 2143 -8706 2446 -8653
rect 2499 -8706 2802 -8653
rect 2855 -8706 3158 -8653
rect 3211 -8706 3513 -8653
rect 3566 -8706 3869 -8653
rect 5237 -8685 10564 -8635
rect 5185 -8697 5237 -8687
rect -1826 -8716 -1773 -8706
rect -1470 -8716 -1417 -8706
rect -1115 -8716 -1062 -8706
rect -758 -8716 -705 -8706
rect -402 -8716 -349 -8706
rect -47 -8716 6 -8706
rect 310 -8716 363 -8706
rect 666 -8716 719 -8706
rect 1022 -8716 1075 -8706
rect 1377 -8716 1430 -8706
rect 1733 -8716 1786 -8706
rect 2090 -8716 2143 -8706
rect 2446 -8716 2499 -8706
rect 2802 -8716 2855 -8706
rect 3158 -8716 3211 -8706
rect 3513 -8716 3566 -8706
rect 3869 -8716 3922 -8706
rect 10512 -8716 10564 -8685
rect 11054 -8716 11107 -8706
rect 11345 -8716 11398 -8706
rect 11638 -8716 11691 -8706
rect 11932 -8716 11985 -8706
rect 12222 -8716 12275 -8706
rect 17831 -8716 17895 -6585
rect -2447 -8767 -2394 -8757
rect -2005 -8767 -1952 -8757
rect -1648 -8767 -1595 -8757
rect -1293 -8767 -1240 -8757
rect -936 -8767 -883 -8757
rect -580 -8766 -527 -8756
rect -2394 -8820 -2005 -8767
rect -1952 -8820 -1648 -8767
rect -1595 -8820 -1293 -8767
rect -1240 -8820 -936 -8767
rect -883 -8819 -580 -8767
rect -225 -8767 -172 -8757
rect 132 -8767 185 -8758
rect 489 -8766 542 -8756
rect -527 -8819 -225 -8767
rect -883 -8820 -225 -8819
rect -172 -8768 489 -8767
rect -172 -8820 132 -8768
rect -2447 -8830 -2394 -8820
rect -2005 -8830 -1952 -8820
rect -1648 -8830 -1595 -8820
rect -1293 -8830 -1240 -8820
rect -936 -8830 -883 -8820
rect -580 -8829 -527 -8820
rect -225 -8830 -172 -8820
rect 185 -8819 489 -8768
rect 843 -8766 896 -8756
rect 542 -8819 843 -8767
rect 1201 -8767 1254 -8757
rect 1556 -8767 1609 -8757
rect 1911 -8767 1964 -8757
rect 2267 -8767 2320 -8757
rect 2624 -8767 2677 -8757
rect 2980 -8767 3033 -8757
rect 3336 -8767 3389 -8757
rect 3692 -8767 3745 -8757
rect 896 -8819 1201 -8767
rect 185 -8820 1201 -8819
rect 1254 -8820 1556 -8767
rect 1609 -8820 1911 -8767
rect 1964 -8820 2267 -8767
rect 2320 -8820 2624 -8767
rect 2677 -8820 2980 -8767
rect 3033 -8820 3336 -8767
rect 3389 -8820 3692 -8767
rect 10512 -8768 11054 -8716
rect 10584 -8769 11054 -8768
rect 11107 -8769 11345 -8716
rect 11398 -8769 11638 -8716
rect 11691 -8769 11932 -8716
rect 11985 -8769 12222 -8716
rect 12275 -8769 17895 -8716
rect 11054 -8779 11107 -8769
rect 11345 -8779 11398 -8769
rect 11638 -8779 11691 -8769
rect 11932 -8779 11985 -8769
rect 12222 -8779 12275 -8769
rect 132 -8831 185 -8821
rect 489 -8829 542 -8820
rect 843 -8829 896 -8820
rect 1201 -8830 1254 -8820
rect 1556 -8830 1609 -8820
rect 1911 -8830 1964 -8820
rect 2267 -8830 2320 -8820
rect 2624 -8830 2677 -8820
rect 2980 -8830 3033 -8820
rect 3336 -8830 3389 -8820
rect 3692 -8830 3745 -8820
rect 4771 -9314 4824 -9304
rect 6769 -9314 6822 -9304
rect 6947 -9314 7000 -9305
rect 7126 -9314 7179 -9305
rect 7303 -9313 7356 -9303
rect 4824 -9367 6769 -9314
rect 6822 -9315 7303 -9314
rect 6822 -9367 6947 -9315
rect 4771 -9377 4824 -9367
rect 6769 -9377 6822 -9367
rect 7000 -9367 7126 -9315
rect 6947 -9378 7000 -9368
rect 7179 -9366 7303 -9315
rect 7482 -9313 7535 -9303
rect 7356 -9366 7482 -9314
rect 7659 -9314 7712 -9305
rect 7837 -9314 7890 -9304
rect 8015 -9314 8068 -9305
rect 8194 -9314 8247 -9304
rect 8371 -9314 8424 -9304
rect 8549 -9314 8602 -9304
rect 8727 -9314 8780 -9305
rect 8906 -9314 8959 -9304
rect 7535 -9315 7837 -9314
rect 7535 -9366 7659 -9315
rect 7179 -9367 7659 -9366
rect 7126 -9378 7179 -9368
rect 7303 -9376 7356 -9367
rect 7482 -9376 7535 -9367
rect 7712 -9367 7837 -9315
rect 7890 -9315 8194 -9314
rect 7890 -9367 8015 -9315
rect 7659 -9378 7712 -9368
rect 7837 -9377 7890 -9367
rect 8068 -9367 8194 -9315
rect 8247 -9367 8371 -9314
rect 8424 -9367 8549 -9314
rect 8602 -9315 8906 -9314
rect 8602 -9367 8727 -9315
rect 8015 -9378 8068 -9368
rect 8194 -9377 8247 -9367
rect 8371 -9377 8424 -9367
rect 8549 -9377 8602 -9367
rect 8780 -9367 8906 -9315
rect 8727 -9378 8780 -9368
rect 8906 -9377 8959 -9367
rect 11144 -9374 11197 -9364
rect 11436 -9375 11489 -9365
rect 11728 -9375 11781 -9365
rect 12020 -9375 12073 -9366
rect 12312 -9375 12365 -9365
rect 11197 -9427 11436 -9375
rect 11144 -9428 11436 -9427
rect 11489 -9428 11728 -9375
rect 11781 -9376 12312 -9375
rect 11781 -9428 12020 -9376
rect 11144 -9437 11197 -9428
rect 11436 -9438 11489 -9428
rect 11728 -9438 11781 -9428
rect 12073 -9428 12312 -9376
rect 12020 -9439 12073 -9429
rect 12312 -9438 12365 -9428
rect -1916 -9546 -1863 -9536
rect -1738 -9546 -1685 -9536
rect -1558 -9546 -1505 -9536
rect -312 -9546 -259 -9536
rect -136 -9545 -83 -9535
rect -1863 -9599 -1738 -9546
rect -1685 -9599 -1558 -9546
rect -1505 -9599 -312 -9546
rect -259 -9598 -136 -9546
rect 42 -9546 95 -9536
rect 222 -9545 275 -9535
rect -83 -9598 42 -9546
rect -259 -9599 42 -9598
rect 95 -9598 222 -9546
rect 399 -9546 452 -9536
rect 577 -9546 630 -9536
rect 2178 -9546 2231 -9537
rect 2357 -9546 2410 -9536
rect 2534 -9546 2587 -9536
rect 2713 -9546 2766 -9536
rect 4208 -9546 4261 -9536
rect 6679 -9545 6732 -9535
rect 275 -9598 399 -9546
rect 95 -9599 399 -9598
rect 452 -9599 577 -9546
rect 630 -9547 2357 -9546
rect 630 -9599 2178 -9547
rect -1916 -9609 -1863 -9599
rect -1738 -9609 -1685 -9599
rect -1558 -9609 -1505 -9599
rect -312 -9609 -259 -9599
rect -136 -9608 -83 -9599
rect 42 -9609 95 -9599
rect 222 -9608 275 -9599
rect 399 -9609 452 -9599
rect 577 -9609 630 -9599
rect 2231 -9599 2357 -9547
rect 2410 -9599 2534 -9546
rect 2587 -9599 2713 -9546
rect 2766 -9599 4208 -9546
rect 4261 -9598 6679 -9546
rect 4261 -9599 6732 -9598
rect 2178 -9610 2231 -9600
rect 2357 -9609 2410 -9599
rect 2534 -9609 2587 -9599
rect 2713 -9609 2766 -9599
rect 4208 -9609 4261 -9599
rect 6679 -9608 6732 -9599
rect -2315 -9925 -2262 -9915
rect -1916 -9925 -1863 -9915
rect -1738 -9925 -1685 -9916
rect -1560 -9925 -1507 -9915
rect -1382 -9924 -1329 -9914
rect -2262 -9978 -1916 -9925
rect -1863 -9926 -1560 -9925
rect -1863 -9978 -1738 -9926
rect -2315 -9988 -2262 -9978
rect -1916 -9988 -1863 -9978
rect -1685 -9978 -1560 -9926
rect -1507 -9977 -1382 -9925
rect -314 -9925 -261 -9915
rect -136 -9925 -83 -9916
rect 43 -9925 96 -9915
rect 220 -9925 273 -9915
rect 398 -9925 451 -9915
rect 576 -9925 629 -9915
rect 2356 -9925 2409 -9915
rect 2534 -9925 2587 -9915
rect 2712 -9925 2765 -9916
rect 2891 -9925 2944 -9915
rect 3069 -9925 3122 -9915
rect 3246 -9925 3299 -9915
rect 5337 -9925 5390 -9915
rect -1329 -9977 -314 -9925
rect -1507 -9978 -314 -9977
rect -261 -9926 43 -9925
rect -261 -9978 -136 -9926
rect -1738 -9989 -1685 -9979
rect -1560 -9988 -1507 -9978
rect -1382 -9987 -1329 -9978
rect -314 -9988 -261 -9978
rect -83 -9978 43 -9926
rect 96 -9978 220 -9925
rect 273 -9978 398 -9925
rect 451 -9978 576 -9925
rect 629 -9978 2356 -9925
rect 2409 -9978 2534 -9925
rect 2587 -9926 2891 -9925
rect 2587 -9978 2712 -9926
rect -136 -9989 -83 -9979
rect 43 -9988 96 -9978
rect 220 -9988 273 -9978
rect 398 -9988 451 -9978
rect 576 -9988 629 -9978
rect 2356 -9988 2409 -9978
rect 2534 -9988 2587 -9978
rect 2765 -9978 2891 -9926
rect 2944 -9978 3069 -9925
rect 3122 -9978 3246 -9925
rect 3299 -9978 5337 -9925
rect 2712 -9989 2765 -9979
rect 2891 -9988 2944 -9978
rect 3069 -9988 3122 -9978
rect 3246 -9988 3299 -9978
rect 5337 -9988 5390 -9978
rect 6680 -10313 6733 -10303
rect 9171 -10313 9224 -10304
rect 6733 -10314 9224 -10313
rect 6733 -10366 9171 -10314
rect 6680 -10376 6733 -10366
rect 9171 -10377 9224 -10367
rect 6858 -10466 6911 -10457
rect 7214 -10466 7267 -10456
rect 7571 -10466 7624 -10456
rect 7927 -10466 7980 -10456
rect 8283 -10466 8336 -10457
rect 8638 -10466 8691 -10456
rect 8995 -10466 9048 -10457
rect 6858 -10467 7214 -10466
rect 6911 -10519 7214 -10467
rect 7267 -10519 7571 -10466
rect 7624 -10519 7927 -10466
rect 7980 -10467 8638 -10466
rect 7980 -10519 8283 -10467
rect 6858 -10530 6911 -10520
rect 7214 -10529 7267 -10519
rect 7571 -10529 7624 -10519
rect 7927 -10529 7980 -10519
rect 8336 -10519 8638 -10467
rect 8691 -10467 9048 -10466
rect 8691 -10519 8995 -10467
rect 8283 -10530 8336 -10520
rect 8638 -10529 8691 -10519
rect 8995 -10530 9048 -10520
rect -1827 -10908 -1774 -10898
rect -1470 -10908 -1417 -10898
rect -1114 -10908 -1061 -10898
rect -758 -10908 -705 -10898
rect -402 -10908 -349 -10898
rect -46 -10908 7 -10898
rect 309 -10908 362 -10898
rect 665 -10908 718 -10898
rect 931 -10908 984 -10898
rect 1199 -10908 1252 -10898
rect 1556 -10908 1609 -10898
rect 1913 -10908 1966 -10898
rect 2268 -10908 2321 -10898
rect 2623 -10908 2676 -10898
rect 2980 -10908 3033 -10898
rect 3335 -10908 3388 -10898
rect 3692 -10908 3745 -10898
rect -1774 -10961 -1470 -10908
rect -1417 -10961 -1114 -10908
rect -1061 -10961 -758 -10908
rect -705 -10961 -402 -10908
rect -349 -10961 -46 -10908
rect 7 -10961 309 -10908
rect 362 -10961 665 -10908
rect 718 -10961 931 -10908
rect 984 -10961 1199 -10908
rect 1252 -10961 1556 -10908
rect 1609 -10961 1913 -10908
rect 1966 -10961 2268 -10908
rect 2321 -10961 2623 -10908
rect 2676 -10961 2980 -10908
rect 3033 -10961 3335 -10908
rect 3388 -10961 3692 -10908
rect -1827 -10971 -1774 -10961
rect -1470 -10971 -1417 -10961
rect -1114 -10971 -1061 -10961
rect -758 -10971 -705 -10961
rect -402 -10971 -349 -10961
rect -46 -10971 7 -10961
rect 309 -10971 362 -10961
rect 665 -10971 718 -10961
rect 931 -10971 984 -10961
rect 1199 -10971 1252 -10961
rect 1556 -10971 1609 -10961
rect 1913 -10971 1966 -10961
rect 2268 -10971 2321 -10961
rect 2623 -10971 2676 -10961
rect 2980 -10971 3033 -10961
rect 3335 -10971 3388 -10961
rect 3692 -10971 3745 -10961
rect 7037 -11366 7090 -11356
rect 7393 -11366 7446 -11356
rect 7748 -11366 7801 -11357
rect 8103 -11366 8156 -11356
rect 8461 -11366 8514 -11356
rect 8817 -11366 8870 -11356
rect 7090 -11419 7393 -11366
rect 7446 -11367 8103 -11366
rect 7446 -11419 7748 -11367
rect 7037 -11429 7090 -11419
rect 7393 -11429 7446 -11419
rect 7801 -11419 8103 -11367
rect 8156 -11419 8461 -11366
rect 8514 -11419 8817 -11366
rect 7748 -11430 7801 -11420
rect 8103 -11429 8156 -11419
rect 8461 -11429 8514 -11419
rect 8817 -11429 8870 -11419
rect -1649 -11528 -1596 -11518
rect -1293 -11528 -1240 -11518
rect -937 -11528 -884 -11518
rect 1377 -11528 1430 -11518
rect 1733 -11528 1786 -11518
rect 2089 -11528 2142 -11518
rect -1596 -11581 -1293 -11528
rect -1240 -11581 -937 -11528
rect -884 -11581 1377 -11528
rect 1430 -11581 1733 -11528
rect 1786 -11581 2089 -11528
rect -1649 -11591 -1596 -11581
rect -1293 -11591 -1240 -11581
rect -937 -11591 -884 -11581
rect 1377 -11591 1430 -11581
rect 1733 -11591 1786 -11581
rect 2089 -11591 2142 -11581
rect -2004 -11637 -1951 -11627
rect -580 -11637 -527 -11627
rect 2446 -11637 2499 -11627
rect 3871 -11637 3924 -11628
rect -1951 -11690 -580 -11637
rect -527 -11690 2446 -11637
rect 2499 -11638 3924 -11637
rect 2499 -11690 3871 -11638
rect -2004 -11700 -1951 -11690
rect -580 -11700 -527 -11690
rect 2446 -11700 2499 -11690
rect 3871 -11701 3924 -11691
rect 11053 -11674 11106 -11664
rect 11347 -11674 11400 -11665
rect 11638 -11674 11691 -11664
rect 11931 -11674 11984 -11664
rect 12223 -11674 12276 -11664
rect 13022 -11673 13075 -11663
rect 11106 -11675 11638 -11674
rect 11106 -11727 11347 -11675
rect 11053 -11737 11106 -11727
rect 11400 -11727 11638 -11675
rect 11691 -11727 11931 -11674
rect 11984 -11727 12223 -11674
rect 12276 -11726 13022 -11674
rect 12276 -11727 13075 -11726
rect 11347 -11738 11400 -11728
rect 11638 -11737 11691 -11727
rect 11931 -11737 11984 -11727
rect 12223 -11737 12276 -11727
rect 13022 -11736 13075 -11727
rect -224 -11757 -171 -11747
rect 131 -11757 184 -11747
rect 487 -11757 540 -11747
rect 2800 -11757 2853 -11747
rect 3157 -11757 3210 -11747
rect 3513 -11757 3566 -11747
rect -171 -11810 131 -11757
rect 184 -11810 487 -11757
rect 540 -11810 2800 -11757
rect 2853 -11810 3157 -11757
rect 3210 -11810 3513 -11757
rect -224 -11820 -171 -11810
rect 131 -11820 184 -11810
rect 487 -11820 540 -11810
rect 2800 -11820 2853 -11810
rect 3157 -11820 3210 -11810
rect 3513 -11820 3566 -11810
rect -1915 -11919 -1862 -11909
rect -1738 -11919 -1685 -11909
rect -1559 -11919 -1506 -11909
rect -1381 -11919 -1328 -11909
rect -1203 -11919 -1150 -11909
rect -1025 -11919 -972 -11909
rect -848 -11919 -795 -11909
rect -670 -11919 -617 -11909
rect -492 -11919 -439 -11909
rect -314 -11919 -261 -11909
rect -136 -11919 -83 -11909
rect 42 -11919 95 -11909
rect 220 -11919 273 -11909
rect 399 -11919 452 -11909
rect 577 -11919 630 -11909
rect 1288 -11919 1341 -11909
rect 1468 -11919 1521 -11909
rect 1644 -11919 1697 -11910
rect 1823 -11919 1876 -11909
rect 2000 -11919 2053 -11909
rect 2178 -11919 2231 -11909
rect 2357 -11919 2410 -11909
rect 2534 -11919 2587 -11909
rect 2713 -11919 2766 -11909
rect 2890 -11919 2943 -11909
rect 3068 -11919 3121 -11909
rect 3247 -11919 3300 -11909
rect 3425 -11919 3478 -11909
rect 3603 -11919 3656 -11909
rect 3781 -11919 3834 -11909
rect -1862 -11972 -1738 -11919
rect -1685 -11972 -1559 -11919
rect -1506 -11972 -1381 -11919
rect -1328 -11972 -1203 -11919
rect -1150 -11972 -1025 -11919
rect -972 -11972 -848 -11919
rect -795 -11972 -670 -11919
rect -617 -11972 -492 -11919
rect -439 -11972 -314 -11919
rect -261 -11972 -136 -11919
rect -83 -11972 42 -11919
rect 95 -11972 220 -11919
rect 273 -11972 399 -11919
rect 452 -11972 577 -11919
rect 630 -11972 1288 -11919
rect 1341 -11972 1468 -11919
rect 1521 -11920 1823 -11919
rect 1521 -11972 1644 -11920
rect -1915 -11982 -1862 -11972
rect -1738 -11982 -1685 -11972
rect -1559 -11982 -1506 -11972
rect -1381 -11982 -1328 -11972
rect -1203 -11982 -1150 -11972
rect -1025 -11982 -972 -11972
rect -848 -11982 -795 -11972
rect -670 -11982 -617 -11972
rect -492 -11982 -439 -11972
rect -314 -11982 -261 -11972
rect -136 -11982 -83 -11972
rect 42 -11982 95 -11972
rect 220 -11982 273 -11972
rect 399 -11982 452 -11972
rect 577 -11982 630 -11972
rect 1288 -11982 1341 -11972
rect 1468 -11982 1521 -11972
rect 1697 -11972 1823 -11920
rect 1876 -11972 2000 -11919
rect 2053 -11972 2178 -11919
rect 2231 -11972 2357 -11919
rect 2410 -11972 2534 -11919
rect 2587 -11972 2713 -11919
rect 2766 -11972 2890 -11919
rect 2943 -11972 3068 -11919
rect 3121 -11972 3247 -11919
rect 3300 -11972 3425 -11919
rect 3478 -11972 3603 -11919
rect 3656 -11972 3781 -11919
rect 1644 -11983 1697 -11973
rect 1823 -11982 1876 -11972
rect 2000 -11982 2053 -11972
rect 2178 -11982 2231 -11972
rect 2357 -11982 2410 -11972
rect 2534 -11982 2587 -11972
rect 2713 -11982 2766 -11972
rect 2890 -11982 2943 -11972
rect 3068 -11982 3121 -11972
rect 3247 -11982 3300 -11972
rect 3425 -11982 3478 -11972
rect 3603 -11982 3656 -11972
rect 3781 -11982 3834 -11972
rect -5502 -12271 -5449 -12261
rect -5000 -12271 -4947 -12262
rect -4502 -12271 -4449 -12261
rect -5449 -12272 -4502 -12271
rect -5449 -12324 -5000 -12272
rect -5502 -12334 -5449 -12324
rect -4947 -12324 -4502 -12272
rect -2447 -12272 -2394 -12262
rect -4449 -12324 -2447 -12272
rect -5000 -12335 -4947 -12325
rect -4502 -12325 -2447 -12324
rect -4502 -12334 -4449 -12325
rect -2447 -12335 -2394 -12325
rect -5376 -12388 -5323 -12378
rect -5127 -12388 -5074 -12378
rect -4377 -12388 -4324 -12378
rect -3928 -12388 -3875 -12379
rect -5323 -12441 -5127 -12388
rect -5074 -12441 -4377 -12388
rect -4324 -12389 -3875 -12388
rect -4324 -12441 -3928 -12389
rect -5376 -12451 -5323 -12441
rect -5127 -12451 -5074 -12441
rect -4377 -12451 -4324 -12441
rect -3928 -12452 -3875 -12442
rect -6077 -12512 -6024 -12502
rect -5626 -12512 -5573 -12502
rect -4877 -12512 -4824 -12502
rect -4627 -12512 -4574 -12502
rect -6024 -12565 -5626 -12512
rect -5573 -12565 -4877 -12512
rect -4824 -12565 -4627 -12512
rect -6077 -12575 -6024 -12565
rect -5626 -12575 -5573 -12565
rect -4877 -12575 -4824 -12565
rect -4627 -12575 -4574 -12565
rect -2005 -12542 -1952 -12532
rect -1649 -12542 -1596 -12532
rect 3514 -12542 3567 -12532
rect 3871 -12542 3924 -12532
rect -1952 -12595 -1649 -12542
rect -1596 -12544 -1284 -12542
rect -1250 -12544 3514 -12542
rect -1596 -12595 3514 -12544
rect 3567 -12595 3871 -12542
rect -2005 -12605 -1952 -12595
rect -1649 -12605 -1596 -12595
rect 3514 -12605 3567 -12595
rect 3871 -12605 3924 -12595
rect -1294 -12653 -1241 -12644
rect -582 -12653 -529 -12643
rect 130 -12653 183 -12643
rect 1735 -12653 1788 -12644
rect 2445 -12653 2498 -12643
rect 3158 -12652 3211 -12642
rect -1294 -12654 -582 -12653
rect -1241 -12706 -582 -12654
rect -529 -12706 130 -12653
rect 183 -12654 2445 -12653
rect 183 -12706 1735 -12654
rect -1294 -12717 -1241 -12707
rect -582 -12716 -529 -12706
rect 130 -12716 183 -12706
rect 1788 -12706 2445 -12654
rect 2498 -12705 3158 -12653
rect 2498 -12706 3211 -12705
rect 1735 -12717 1788 -12707
rect 2445 -12716 2498 -12706
rect 3158 -12715 3211 -12706
rect -937 -12783 -884 -12773
rect -224 -12783 -171 -12773
rect 486 -12783 539 -12774
rect 1378 -12783 1431 -12773
rect 2088 -12782 2141 -12772
rect -884 -12836 -224 -12783
rect -171 -12784 1378 -12783
rect -171 -12836 486 -12784
rect -937 -12846 -884 -12836
rect -224 -12846 -171 -12836
rect 539 -12836 1378 -12784
rect 1431 -12835 2088 -12783
rect 2801 -12782 2854 -12772
rect 2141 -12835 2801 -12783
rect 1431 -12836 2854 -12835
rect 486 -12847 539 -12837
rect 1378 -12846 1431 -12836
rect 2088 -12845 2141 -12836
rect 2801 -12845 2854 -12836
rect -6223 -13062 -6170 -13052
rect -5751 -13062 -5698 -13052
rect -4752 -13062 -4699 -13052
rect -6170 -13115 -5751 -13062
rect -5698 -13115 -4752 -13062
rect -6223 -13125 -6170 -13115
rect -5751 -13125 -5698 -13115
rect -4752 -13125 -4699 -13115
rect -5251 -13189 -5198 -13179
rect -4251 -13189 -4198 -13179
rect -3788 -13189 -3735 -13179
rect -3542 -13189 -3489 -13179
rect -5198 -13242 -4251 -13189
rect -4198 -13242 -3788 -13189
rect -3735 -13242 -3542 -13189
rect -5251 -13252 -5198 -13242
rect -4251 -13252 -4198 -13242
rect -3788 -13252 -3735 -13242
rect -3542 -13252 -3489 -13242
rect 5037 -13296 5090 -13286
rect 5534 -13296 5587 -13286
rect 5090 -13349 5534 -13296
rect 5037 -13359 5090 -13349
rect 5534 -13359 5587 -13349
rect 18337 -13421 18412 -13411
rect 5031 -13433 5084 -13423
rect 8950 -13433 9003 -13423
rect 9305 -13433 9358 -13423
rect 5084 -13486 8950 -13433
rect 9003 -13486 9305 -13433
rect 9358 -13486 18337 -13433
rect 5031 -13496 5084 -13486
rect 8950 -13496 9003 -13486
rect 9305 -13496 9358 -13486
rect 18412 -13486 18422 -13433
rect 18337 -13506 18412 -13496
rect -2004 -13545 -1951 -13535
rect -581 -13545 -528 -13535
rect 2446 -13545 2499 -13535
rect 3870 -13545 3923 -13535
rect 5400 -13545 5453 -13535
rect -1951 -13598 -581 -13545
rect -528 -13598 2446 -13545
rect 2499 -13598 3870 -13545
rect 3923 -13598 5400 -13545
rect 5453 -13556 8828 -13545
rect 9127 -13556 9180 -13546
rect 9483 -13556 9536 -13546
rect 5453 -13598 8772 -13556
rect -2004 -13608 -1951 -13598
rect -581 -13608 -528 -13598
rect 2446 -13608 2499 -13598
rect 3870 -13608 3923 -13598
rect 5400 -13608 5453 -13598
rect 8825 -13609 9127 -13556
rect 9180 -13609 9483 -13556
rect 8772 -13619 8825 -13609
rect 9127 -13619 9180 -13609
rect 9483 -13619 9536 -13609
rect -1648 -13672 -1595 -13662
rect -1291 -13672 -1238 -13662
rect -937 -13672 -884 -13662
rect 1379 -13672 1432 -13662
rect 1732 -13672 1785 -13662
rect 2091 -13672 2144 -13662
rect 5534 -13672 5587 -13662
rect 7526 -13672 7579 -13662
rect 7882 -13672 7935 -13663
rect 8238 -13671 8291 -13661
rect -1595 -13725 -1291 -13672
rect -1238 -13725 -937 -13672
rect -884 -13725 1379 -13672
rect 1432 -13725 1732 -13672
rect 1785 -13725 2091 -13672
rect 2144 -13725 5323 -13672
rect -1648 -13735 -1595 -13725
rect -1291 -13735 -1238 -13725
rect -937 -13735 -884 -13725
rect 1379 -13735 1432 -13725
rect 1732 -13735 1785 -13725
rect 2091 -13735 2144 -13725
rect -6077 -13745 -6024 -13735
rect -5376 -13745 -5323 -13735
rect -5126 -13745 -5073 -13735
rect -4376 -13745 -4323 -13735
rect -6024 -13798 -5376 -13745
rect -5323 -13798 -5126 -13745
rect -5073 -13798 -4376 -13745
rect -6077 -13808 -6024 -13798
rect -5376 -13808 -5323 -13798
rect -5126 -13808 -5073 -13798
rect -4376 -13808 -4323 -13798
rect -225 -13794 -172 -13784
rect 133 -13794 186 -13784
rect 487 -13794 540 -13785
rect 2802 -13794 2855 -13784
rect 3157 -13794 3210 -13785
rect 3512 -13794 3565 -13784
rect 5142 -13794 5195 -13784
rect -6426 -13852 -6373 -13842
rect -5626 -13852 -5573 -13842
rect -4877 -13852 -4824 -13842
rect -4627 -13852 -4574 -13842
rect -3928 -13852 -3875 -13842
rect -6373 -13905 -5626 -13852
rect -5573 -13905 -4877 -13852
rect -4824 -13905 -4627 -13852
rect -4574 -13905 -3928 -13852
rect -172 -13847 133 -13794
rect 186 -13795 2802 -13794
rect 186 -13847 487 -13795
rect -225 -13857 -172 -13847
rect 133 -13857 186 -13847
rect 540 -13847 2802 -13795
rect 2855 -13795 3512 -13794
rect 2855 -13847 3157 -13795
rect 487 -13858 540 -13848
rect 2802 -13857 2855 -13847
rect 3210 -13847 3512 -13795
rect 3565 -13847 5142 -13794
rect 3157 -13858 3210 -13848
rect 3512 -13857 3565 -13847
rect 5142 -13857 5195 -13847
rect 5270 -13796 5323 -13725
rect 5587 -13725 7526 -13672
rect 7579 -13673 8238 -13672
rect 7579 -13725 7882 -13673
rect 5534 -13735 5587 -13725
rect 7526 -13735 7579 -13725
rect 7935 -13724 8238 -13673
rect 11442 -13672 11495 -13662
rect 11798 -13672 11851 -13662
rect 12152 -13672 12205 -13663
rect 12509 -13672 12562 -13662
rect 8291 -13724 11442 -13672
rect 7935 -13725 11442 -13724
rect 11495 -13725 11798 -13672
rect 11851 -13673 12509 -13672
rect 11851 -13725 12152 -13673
rect 7882 -13736 7935 -13726
rect 8238 -13734 8291 -13725
rect 11442 -13735 11495 -13725
rect 11798 -13735 11851 -13725
rect 12205 -13725 12509 -13673
rect 12152 -13736 12205 -13726
rect 12509 -13735 12562 -13725
rect 7348 -13796 7401 -13786
rect 7704 -13795 7757 -13785
rect 5270 -13849 7348 -13796
rect 7401 -13848 7704 -13796
rect 8061 -13796 8114 -13786
rect 8415 -13796 8468 -13786
rect 11264 -13796 11317 -13786
rect 11620 -13796 11673 -13787
rect 11977 -13796 12030 -13786
rect 12334 -13796 12387 -13786
rect 7757 -13848 8061 -13796
rect 7401 -13849 8061 -13848
rect 8114 -13849 8415 -13796
rect 8468 -13849 11264 -13796
rect 11317 -13797 11977 -13796
rect 11317 -13849 11620 -13797
rect 7348 -13859 7401 -13849
rect 7704 -13858 7757 -13849
rect 8061 -13859 8114 -13849
rect 8415 -13859 8468 -13849
rect 11264 -13859 11317 -13849
rect 11673 -13849 11977 -13797
rect 12030 -13849 12334 -13796
rect 11620 -13860 11673 -13850
rect 11977 -13859 12030 -13849
rect 12334 -13859 12387 -13849
rect -6426 -13915 -6373 -13905
rect -5626 -13915 -5573 -13905
rect -4877 -13915 -4824 -13905
rect -4627 -13915 -4574 -13905
rect -3928 -13915 -3875 -13905
rect 5833 -13922 5886 -13912
rect 6013 -13922 6066 -13912
rect 6190 -13922 6243 -13913
rect 6369 -13922 6422 -13912
rect 6547 -13922 6600 -13913
rect 6725 -13922 6778 -13912
rect 6902 -13922 6955 -13912
rect 7437 -13922 7490 -13912
rect 7615 -13922 7668 -13912
rect 7793 -13922 7846 -13913
rect 7970 -13922 8023 -13912
rect 8148 -13922 8201 -13912
rect 8326 -13922 8379 -13912
rect 8861 -13922 8914 -13912
rect 9038 -13922 9091 -13912
rect 9217 -13922 9270 -13912
rect 9394 -13922 9447 -13912
rect 9929 -13922 9982 -13913
rect 10108 -13922 10161 -13912
rect 10284 -13922 10337 -13913
rect 10462 -13922 10515 -13913
rect 10640 -13922 10693 -13912
rect 10819 -13922 10872 -13913
rect 11353 -13922 11406 -13912
rect 11530 -13922 11583 -13912
rect 11709 -13922 11762 -13912
rect 11886 -13922 11939 -13913
rect 12064 -13922 12117 -13912
rect 12242 -13922 12295 -13913
rect 12420 -13922 12473 -13912
rect -5730 -13957 -5677 -13947
rect -4752 -13957 -4699 -13947
rect -3788 -13957 -3735 -13947
rect -5677 -14010 -4752 -13957
rect -4699 -14010 -3788 -13957
rect 5886 -13975 6013 -13922
rect 6066 -13923 6369 -13922
rect 6066 -13975 6190 -13923
rect 5833 -13985 5886 -13975
rect 6013 -13985 6066 -13975
rect 6243 -13975 6369 -13923
rect 6422 -13923 6725 -13922
rect 6422 -13975 6547 -13923
rect 6190 -13986 6243 -13976
rect 6369 -13985 6422 -13975
rect 6600 -13975 6725 -13923
rect 6778 -13975 6902 -13922
rect 6955 -13975 7437 -13922
rect 7490 -13975 7615 -13922
rect 7668 -13923 7970 -13922
rect 7668 -13975 7793 -13923
rect 6547 -13986 6600 -13976
rect 6725 -13985 6778 -13975
rect 6902 -13985 6955 -13975
rect 7437 -13985 7490 -13975
rect 7615 -13985 7668 -13975
rect 7846 -13975 7970 -13923
rect 8023 -13975 8148 -13922
rect 8201 -13975 8326 -13922
rect 8379 -13975 8861 -13922
rect 8914 -13975 9038 -13922
rect 9091 -13975 9217 -13922
rect 9270 -13975 9394 -13922
rect 9447 -13923 10108 -13922
rect 9447 -13975 9929 -13923
rect 7793 -13986 7846 -13976
rect 7970 -13985 8023 -13975
rect 8148 -13985 8201 -13975
rect 8326 -13985 8379 -13975
rect 8861 -13985 8914 -13975
rect 9038 -13985 9091 -13975
rect 9217 -13985 9270 -13975
rect 9394 -13985 9447 -13975
rect 9982 -13975 10108 -13923
rect 10161 -13923 10640 -13922
rect 10161 -13975 10284 -13923
rect 9929 -13986 9982 -13976
rect 10108 -13985 10161 -13975
rect 10337 -13975 10462 -13923
rect 10284 -13986 10337 -13976
rect 10515 -13975 10640 -13923
rect 10693 -13923 11353 -13922
rect 10693 -13975 10819 -13923
rect 10462 -13986 10515 -13976
rect 10640 -13985 10693 -13975
rect 10872 -13975 11353 -13923
rect 11406 -13975 11530 -13922
rect 11583 -13975 11709 -13922
rect 11762 -13923 12064 -13922
rect 11762 -13975 11886 -13923
rect 10819 -13986 10872 -13976
rect 11353 -13985 11406 -13975
rect 11530 -13985 11583 -13975
rect 11709 -13985 11762 -13975
rect 11939 -13975 12064 -13923
rect 12117 -13923 12420 -13922
rect 12117 -13975 12242 -13923
rect 11886 -13986 11939 -13976
rect 12064 -13985 12117 -13975
rect 12295 -13975 12420 -13923
rect 12242 -13986 12295 -13976
rect 12420 -13985 12473 -13975
rect -5730 -14020 -5677 -14010
rect -4752 -14020 -4699 -14010
rect -3788 -14020 -3735 -14010
rect -6223 -14055 -6170 -14045
rect -5250 -14055 -5197 -14045
rect -4250 -14055 -4197 -14045
rect -3382 -14055 -3329 -14045
rect -6170 -14108 -5250 -14055
rect -5197 -14108 -4250 -14055
rect -4197 -14108 -3382 -14055
rect -6223 -14118 -6170 -14108
rect -5250 -14118 -5197 -14108
rect -4250 -14118 -4197 -14108
rect -3382 -14118 -3329 -14108
rect -2315 -14543 -2262 -14533
rect -1381 -14543 -1328 -14533
rect -1204 -14543 -1151 -14533
rect -1026 -14543 -973 -14533
rect -848 -14543 -795 -14533
rect -669 -14543 -616 -14533
rect -491 -14543 -438 -14533
rect 1288 -14543 1341 -14533
rect 1466 -14543 1519 -14533
rect 1644 -14543 1697 -14533
rect 1823 -14542 1876 -14532
rect -2262 -14596 -1381 -14543
rect -1328 -14596 -1204 -14543
rect -1151 -14596 -1026 -14543
rect -973 -14596 -848 -14543
rect -795 -14596 -669 -14543
rect -616 -14596 -491 -14543
rect -438 -14596 1288 -14543
rect 1341 -14596 1466 -14543
rect 1519 -14596 1644 -14543
rect 1697 -14595 1823 -14543
rect 2000 -14543 2053 -14533
rect 2178 -14543 2231 -14533
rect 3246 -14543 3299 -14534
rect 3424 -14543 3477 -14533
rect 3602 -14543 3655 -14533
rect 3781 -14543 3834 -14533
rect 1876 -14595 2000 -14543
rect 1697 -14596 2000 -14595
rect 2053 -14596 2178 -14543
rect 2231 -14544 3424 -14543
rect 2231 -14596 3246 -14544
rect -2315 -14606 -2262 -14596
rect -1381 -14606 -1328 -14596
rect -1204 -14606 -1151 -14596
rect -1026 -14606 -973 -14596
rect -848 -14606 -795 -14596
rect -669 -14606 -616 -14596
rect -491 -14606 -438 -14596
rect 1288 -14606 1341 -14596
rect 1466 -14606 1519 -14596
rect 1644 -14606 1697 -14596
rect 1823 -14605 1876 -14596
rect 2000 -14606 2053 -14596
rect 2178 -14606 2231 -14596
rect 3299 -14596 3424 -14544
rect 3477 -14596 3602 -14543
rect 3655 -14596 3781 -14543
rect 3246 -14607 3299 -14597
rect 3424 -14606 3477 -14596
rect 3602 -14606 3655 -14596
rect 3781 -14606 3834 -14596
rect 4905 -14545 4958 -14535
rect 5746 -14545 5799 -14535
rect 6101 -14545 6154 -14535
rect 6459 -14545 6512 -14535
rect 6813 -14545 6866 -14535
rect 8236 -14545 8289 -14535
rect 8595 -14545 8648 -14535
rect 8950 -14545 9003 -14536
rect 9304 -14545 9357 -14535
rect 9661 -14545 9714 -14535
rect 10016 -14545 10069 -14535
rect 10373 -14545 10426 -14536
rect 10729 -14545 10782 -14535
rect 4958 -14598 5746 -14545
rect 5799 -14598 6101 -14545
rect 6154 -14598 6459 -14545
rect 6512 -14598 6813 -14545
rect 6866 -14598 8236 -14545
rect 8289 -14598 8595 -14545
rect 8648 -14546 9304 -14545
rect 8648 -14598 8950 -14546
rect 4905 -14608 4958 -14598
rect 5746 -14608 5799 -14598
rect 6101 -14608 6154 -14598
rect 6459 -14608 6512 -14598
rect 6813 -14608 6866 -14598
rect 8236 -14608 8289 -14598
rect 8595 -14608 8648 -14598
rect 9003 -14598 9304 -14546
rect 9357 -14598 9661 -14545
rect 9714 -14598 10016 -14545
rect 10069 -14546 10729 -14545
rect 10069 -14598 10373 -14546
rect 8950 -14609 9003 -14599
rect 9304 -14608 9357 -14598
rect 9661 -14608 9714 -14598
rect 10016 -14608 10069 -14598
rect 10426 -14598 10729 -14546
rect 10373 -14609 10426 -14599
rect 10729 -14608 10782 -14598
rect 5143 -14658 5196 -14648
rect 5924 -14658 5977 -14648
rect 6279 -14658 6332 -14648
rect 6636 -14658 6689 -14648
rect 6991 -14658 7044 -14648
rect 8417 -14657 8470 -14647
rect 5196 -14711 5924 -14658
rect 5977 -14711 6279 -14658
rect 6332 -14711 6636 -14658
rect 6689 -14711 6991 -14658
rect 7044 -14710 8417 -14658
rect 8772 -14658 8825 -14648
rect 9127 -14658 9180 -14649
rect 9483 -14658 9536 -14648
rect 9837 -14658 9890 -14649
rect 10196 -14658 10249 -14648
rect 10550 -14658 10603 -14648
rect 10908 -14658 10961 -14648
rect 8470 -14710 8772 -14658
rect 7044 -14711 8772 -14710
rect 8825 -14659 9483 -14658
rect 8825 -14711 9127 -14659
rect 5143 -14721 5196 -14711
rect 5924 -14721 5977 -14711
rect 6279 -14721 6332 -14711
rect 6636 -14721 6689 -14711
rect 6991 -14721 7044 -14711
rect 8417 -14720 8470 -14711
rect 8772 -14721 8825 -14711
rect 9180 -14711 9483 -14659
rect 9536 -14659 10196 -14658
rect 9536 -14711 9837 -14659
rect 9127 -14722 9180 -14712
rect 9483 -14721 9536 -14711
rect 9890 -14711 10196 -14659
rect 10249 -14711 10550 -14658
rect 10603 -14711 10908 -14658
rect 9837 -14722 9890 -14712
rect 10196 -14721 10249 -14711
rect 10550 -14721 10603 -14711
rect 10908 -14721 10961 -14711
rect 11087 -14656 11140 -14648
rect 11440 -14656 11493 -14646
rect 11087 -14658 11440 -14656
rect 11140 -14708 11440 -14658
rect 11140 -14709 11192 -14708
rect 11087 -14721 11140 -14711
rect 11440 -14719 11493 -14709
rect -6159 -14795 -6106 -14785
rect -5860 -14795 -5807 -14785
rect -5147 -14795 -5094 -14785
rect -4436 -14795 -4383 -14785
rect -6106 -14848 -5860 -14795
rect -5807 -14848 -5147 -14795
rect -5094 -14848 -4436 -14795
rect 8504 -14806 8557 -14796
rect -6159 -14858 -6106 -14848
rect -5860 -14858 -5807 -14848
rect -5147 -14858 -5094 -14848
rect -4436 -14858 -4383 -14848
rect 6993 -14824 7046 -14814
rect 7347 -14824 7400 -14814
rect 7704 -14824 7757 -14815
rect 7046 -14877 7347 -14824
rect 7400 -14825 7757 -14824
rect 7400 -14877 7704 -14825
rect 6993 -14887 7046 -14877
rect 7347 -14887 7400 -14877
rect 7704 -14888 7757 -14878
rect 8060 -14821 8113 -14811
rect 8113 -14859 8504 -14821
rect 9753 -14806 9806 -14796
rect 8557 -14859 9753 -14821
rect 10195 -14821 10248 -14812
rect 9806 -14822 10248 -14821
rect 9806 -14859 10195 -14822
rect 8113 -14874 10195 -14859
rect 8060 -14884 8113 -14874
rect 10195 -14885 10248 -14875
rect 10552 -14814 10605 -14805
rect 10908 -14813 10961 -14803
rect 10552 -14815 10908 -14814
rect 10605 -14866 10908 -14815
rect 10961 -14814 11013 -14813
rect 11264 -14814 11317 -14805
rect 10961 -14815 11317 -14814
rect 10961 -14866 11264 -14815
rect 10552 -14878 10605 -14868
rect 10908 -14876 10961 -14866
rect 11264 -14878 11317 -14868
rect -5504 -14901 -5451 -14891
rect -4791 -14901 -4738 -14891
rect -3936 -14901 -3883 -14891
rect -5451 -14954 -4791 -14901
rect -4738 -14954 -3936 -14901
rect -5504 -14964 -5451 -14954
rect -4791 -14964 -4738 -14954
rect -3936 -14964 -3883 -14954
rect -847 -14926 -794 -14916
rect -669 -14926 -616 -14916
rect -491 -14926 -438 -14916
rect -314 -14926 -261 -14917
rect -137 -14926 -84 -14916
rect 43 -14926 96 -14916
rect 1289 -14926 1342 -14917
rect 1467 -14926 1520 -14916
rect 1644 -14926 1697 -14916
rect 1822 -14926 1875 -14916
rect 1999 -14926 2052 -14916
rect 2180 -14926 2233 -14916
rect 3425 -14926 3478 -14916
rect 3603 -14926 3656 -14916
rect 3780 -14926 3833 -14916
rect 4239 -14926 4292 -14916
rect -794 -14979 -669 -14926
rect -616 -14979 -491 -14926
rect -438 -14927 -137 -14926
rect -438 -14979 -314 -14927
rect -847 -14989 -794 -14979
rect -669 -14989 -616 -14979
rect -491 -14989 -438 -14979
rect -261 -14979 -137 -14927
rect -84 -14979 43 -14926
rect 96 -14927 1467 -14926
rect 96 -14979 1289 -14927
rect -314 -14990 -261 -14980
rect -137 -14989 -84 -14979
rect 43 -14989 96 -14979
rect 1342 -14979 1467 -14927
rect 1520 -14979 1644 -14926
rect 1697 -14979 1822 -14926
rect 1875 -14979 1999 -14926
rect 2052 -14979 2180 -14926
rect 2233 -14979 3425 -14926
rect 3478 -14979 3603 -14926
rect 3656 -14979 3780 -14926
rect 3833 -14979 4239 -14926
rect 1289 -14990 1342 -14980
rect 1467 -14989 1520 -14979
rect 1644 -14989 1697 -14979
rect 1822 -14989 1875 -14979
rect 1999 -14989 2052 -14979
rect 2180 -14989 2233 -14979
rect 3425 -14989 3478 -14979
rect 3603 -14989 3656 -14979
rect 3780 -14989 3833 -14979
rect 4239 -14989 4292 -14979
rect 7080 -14923 7133 -14913
rect 7260 -14923 7313 -14914
rect 7439 -14923 7492 -14913
rect 8327 -14923 8380 -14913
rect 8505 -14923 8558 -14914
rect 8683 -14923 8736 -14914
rect 9572 -14923 9625 -14913
rect 9750 -14923 9803 -14913
rect 9929 -14923 9982 -14913
rect 10819 -14923 10872 -14913
rect 10996 -14923 11049 -14913
rect 11175 -14923 11228 -14913
rect 7133 -14924 7439 -14923
rect 7133 -14976 7260 -14924
rect 7080 -14986 7133 -14976
rect 7313 -14976 7439 -14924
rect 7492 -14976 8327 -14923
rect 8380 -14924 9572 -14923
rect 8380 -14976 8505 -14924
rect 7260 -14987 7313 -14977
rect 7439 -14986 7492 -14976
rect 8327 -14986 8380 -14976
rect 8558 -14976 8683 -14924
rect 8505 -14987 8558 -14977
rect 8736 -14976 9572 -14924
rect 9625 -14976 9750 -14923
rect 9803 -14976 9929 -14923
rect 9982 -14976 10819 -14923
rect 10872 -14976 10996 -14923
rect 11049 -14976 11175 -14923
rect 8683 -14987 8736 -14977
rect 9572 -14986 9625 -14976
rect 9750 -14986 9803 -14976
rect 9929 -14986 9982 -14976
rect 10819 -14986 10872 -14976
rect 10996 -14986 11049 -14976
rect 11175 -14986 11228 -14976
rect -6159 -15481 -6106 -15472
rect -5504 -15481 -5451 -15471
rect -4792 -15481 -4739 -15471
rect -6159 -15482 -5504 -15481
rect -6106 -15534 -5504 -15482
rect -5451 -15534 -4792 -15481
rect -6159 -15545 -6106 -15535
rect -5504 -15544 -5451 -15534
rect -4792 -15544 -4739 -15534
rect 4238 -15539 4291 -15529
rect 5031 -15539 5084 -15530
rect 5745 -15539 5798 -15529
rect 6101 -15539 6154 -15529
rect 6458 -15539 6511 -15529
rect 11798 -15539 11851 -15530
rect 12155 -15539 12208 -15529
rect 12511 -15539 12564 -15529
rect -5860 -15588 -5807 -15578
rect -5148 -15589 -5095 -15579
rect -4435 -15589 -4383 -15579
rect -3935 -15589 -3883 -15579
rect -5807 -15641 -5148 -15589
rect -5860 -15651 -5807 -15641
rect -5095 -15641 -4435 -15589
rect -4383 -15641 -3935 -15589
rect 4291 -15540 5745 -15539
rect 4291 -15592 5031 -15540
rect 4238 -15602 4291 -15592
rect 5084 -15592 5745 -15540
rect 5798 -15592 6101 -15539
rect 6154 -15592 6458 -15539
rect 6511 -15540 12155 -15539
rect 6511 -15592 11798 -15540
rect 5031 -15603 5084 -15593
rect 5745 -15602 5798 -15592
rect 6101 -15602 6154 -15592
rect 6458 -15602 6511 -15592
rect 11851 -15592 12155 -15540
rect 12208 -15592 12511 -15539
rect 11798 -15603 11851 -15593
rect 12155 -15602 12208 -15592
rect 12511 -15602 12564 -15592
rect -5148 -15652 -5095 -15642
rect -4435 -15651 -4383 -15641
rect -3935 -15651 -3883 -15641
rect 5400 -15652 5453 -15643
rect 5923 -15652 5976 -15642
rect 6279 -15652 6332 -15642
rect 6635 -15652 6688 -15642
rect 11619 -15652 11672 -15642
rect 11975 -15652 12028 -15642
rect 12332 -15652 12385 -15642
rect 5400 -15653 5923 -15652
rect 5453 -15705 5923 -15653
rect 5976 -15705 6279 -15652
rect 6332 -15705 6635 -15652
rect 6688 -15705 11619 -15652
rect 11672 -15705 11975 -15652
rect 12028 -15705 12332 -15652
rect 5400 -15716 5453 -15706
rect 5923 -15715 5976 -15705
rect 6279 -15715 6332 -15705
rect 6635 -15715 6688 -15705
rect 11619 -15715 11672 -15705
rect 11975 -15715 12028 -15705
rect 12332 -15715 12385 -15705
rect 5747 -15750 5800 -15740
rect 6101 -15749 6154 -15739
rect 5800 -15802 6101 -15750
rect 6456 -15750 6509 -15740
rect 6713 -15750 6766 -15741
rect 7169 -15750 7222 -15740
rect 7526 -15749 7579 -15739
rect 6154 -15802 6456 -15750
rect 5800 -15803 6456 -15802
rect 6509 -15751 7169 -15750
rect 6509 -15803 6713 -15751
rect -2447 -15821 -2394 -15811
rect -2005 -15821 -1952 -15812
rect -2394 -15822 -1952 -15821
rect -1649 -15822 -1596 -15812
rect -1293 -15822 -1240 -15812
rect -937 -15822 -884 -15812
rect -581 -15822 -528 -15812
rect -225 -15822 -172 -15812
rect 132 -15821 185 -15811
rect -2394 -15874 -2005 -15822
rect -2447 -15884 -2394 -15874
rect -1952 -15875 -1649 -15822
rect -1596 -15875 -1293 -15822
rect -1240 -15875 -937 -15822
rect -884 -15875 -581 -15822
rect -528 -15875 -225 -15822
rect -172 -15874 132 -15822
rect 487 -15822 540 -15812
rect 843 -15822 896 -15812
rect 1201 -15822 1254 -15812
rect 1555 -15822 1608 -15812
rect 1910 -15822 1963 -15812
rect 2267 -15822 2320 -15812
rect 2624 -15822 2677 -15812
rect 2979 -15822 3032 -15812
rect 3335 -15822 3388 -15812
rect 3692 -15822 3745 -15812
rect 5747 -15813 5800 -15803
rect 6101 -15812 6154 -15803
rect 6456 -15813 6509 -15803
rect 6766 -15803 7169 -15751
rect 7222 -15802 7526 -15750
rect 7882 -15749 7935 -15739
rect 7579 -15802 7882 -15750
rect 10373 -15750 10426 -15741
rect 10730 -15750 10783 -15740
rect 11086 -15750 11139 -15740
rect 7935 -15751 10730 -15750
rect 7935 -15802 10373 -15751
rect 7222 -15803 10373 -15802
rect 6713 -15814 6766 -15804
rect 7169 -15813 7222 -15803
rect 7526 -15812 7579 -15803
rect 7882 -15812 7935 -15803
rect 10426 -15803 10730 -15751
rect 10783 -15803 11086 -15750
rect 10373 -15814 10426 -15804
rect 10730 -15813 10783 -15803
rect 11086 -15813 11139 -15803
rect 185 -15874 487 -15822
rect -172 -15875 487 -15874
rect 540 -15875 843 -15822
rect 896 -15875 1201 -15822
rect 1254 -15875 1555 -15822
rect 1608 -15875 1910 -15822
rect 1963 -15875 2267 -15822
rect 2320 -15875 2624 -15822
rect 2677 -15875 2979 -15822
rect 3032 -15875 3335 -15822
rect 3388 -15875 3692 -15822
rect 11440 -15841 11493 -15831
rect -2005 -15885 -1952 -15875
rect -1649 -15885 -1596 -15875
rect -1293 -15885 -1240 -15875
rect -937 -15885 -884 -15875
rect -581 -15885 -528 -15875
rect -225 -15885 -172 -15875
rect 132 -15884 185 -15875
rect 487 -15885 540 -15875
rect 843 -15885 896 -15875
rect 1201 -15885 1254 -15875
rect 1555 -15885 1608 -15875
rect 1910 -15885 1963 -15875
rect 2267 -15885 2320 -15875
rect 2624 -15885 2677 -15875
rect 2979 -15885 3032 -15875
rect 3335 -15885 3388 -15875
rect 3692 -15885 3745 -15875
rect 6813 -15851 6866 -15841
rect 7169 -15851 7222 -15842
rect 8060 -15851 8113 -15841
rect 8593 -15851 8646 -15842
rect 9663 -15851 9716 -15842
rect 10194 -15851 10247 -15842
rect 11084 -15851 11137 -15842
rect 6866 -15852 8060 -15851
rect 6866 -15904 7169 -15852
rect 6813 -15914 6866 -15904
rect 7222 -15904 8060 -15852
rect 8113 -15852 11440 -15851
rect 8113 -15904 8593 -15852
rect 7169 -15915 7222 -15905
rect 8060 -15914 8113 -15904
rect 8646 -15904 9663 -15852
rect 8593 -15915 8646 -15905
rect 9716 -15904 10194 -15852
rect 9663 -15915 9716 -15905
rect 10247 -15904 11084 -15852
rect 10194 -15915 10247 -15905
rect 11137 -15894 11440 -15852
rect 11137 -15904 11493 -15894
rect 11084 -15915 11137 -15905
rect -1915 -15933 -1862 -15923
rect -1738 -15933 -1685 -15923
rect -1560 -15933 -1507 -15923
rect -1382 -15933 -1329 -15923
rect -1204 -15933 -1151 -15923
rect -1025 -15933 -972 -15923
rect -847 -15933 -794 -15923
rect -670 -15933 -617 -15923
rect -491 -15933 -438 -15923
rect -313 -15933 -260 -15923
rect -136 -15933 -83 -15923
rect 43 -15933 96 -15923
rect 221 -15933 274 -15923
rect 398 -15933 451 -15923
rect 575 -15933 628 -15923
rect 755 -15933 808 -15923
rect 931 -15933 984 -15923
rect 1110 -15933 1163 -15923
rect 1289 -15933 1342 -15923
rect 1466 -15933 1519 -15923
rect 1643 -15933 1696 -15923
rect 1822 -15933 1875 -15923
rect 2000 -15933 2053 -15923
rect 2179 -15933 2232 -15923
rect 2356 -15933 2409 -15923
rect 2534 -15933 2587 -15923
rect 2712 -15933 2765 -15923
rect 2891 -15933 2944 -15923
rect 3068 -15933 3121 -15923
rect 3247 -15933 3300 -15923
rect 3424 -15933 3477 -15923
rect 3603 -15933 3656 -15923
rect 3780 -15933 3833 -15923
rect -1862 -15986 -1738 -15933
rect -1685 -15986 -1560 -15933
rect -1507 -15986 -1382 -15933
rect -1329 -15986 -1204 -15933
rect -1151 -15986 -1025 -15933
rect -972 -15986 -847 -15933
rect -794 -15986 -670 -15933
rect -617 -15986 -491 -15933
rect -438 -15986 -313 -15933
rect -260 -15986 -136 -15933
rect -83 -15986 43 -15933
rect 96 -15986 221 -15933
rect 274 -15986 398 -15933
rect 451 -15986 575 -15933
rect 628 -15986 755 -15933
rect 808 -15986 931 -15933
rect 984 -15986 1110 -15933
rect 1163 -15986 1289 -15933
rect 1342 -15986 1466 -15933
rect 1519 -15986 1643 -15933
rect 1696 -15986 1822 -15933
rect 1875 -15986 2000 -15933
rect 2053 -15986 2179 -15933
rect 2232 -15986 2356 -15933
rect 2409 -15986 2534 -15933
rect 2587 -15986 2712 -15933
rect 2765 -15986 2891 -15933
rect 2944 -15986 3068 -15933
rect 3121 -15986 3247 -15933
rect 3300 -15986 3424 -15933
rect 3477 -15986 3603 -15933
rect 3656 -15986 3780 -15933
rect -1915 -15996 -1862 -15986
rect -1738 -15996 -1685 -15986
rect -1560 -15996 -1507 -15986
rect -1382 -15996 -1329 -15986
rect -1204 -15996 -1151 -15986
rect -1025 -15996 -972 -15986
rect -847 -15996 -794 -15986
rect -670 -15996 -617 -15986
rect -491 -15996 -438 -15986
rect -313 -15996 -260 -15986
rect -136 -15996 -83 -15986
rect 43 -15996 96 -15986
rect 221 -15996 274 -15986
rect 398 -15996 451 -15986
rect 575 -15996 628 -15986
rect 755 -15996 808 -15986
rect 931 -15996 984 -15986
rect 1110 -15996 1163 -15986
rect 1289 -15996 1342 -15986
rect 1466 -15996 1519 -15986
rect 1643 -15996 1696 -15986
rect 1822 -15996 1875 -15986
rect 2000 -15996 2053 -15986
rect 2179 -15996 2232 -15986
rect 2356 -15996 2409 -15986
rect 2534 -15996 2587 -15986
rect 2712 -15996 2765 -15986
rect 2891 -15996 2944 -15986
rect 3068 -15996 3121 -15986
rect 3247 -15996 3300 -15986
rect 3424 -15996 3477 -15986
rect 3603 -15996 3656 -15986
rect 3780 -15996 3833 -15986
rect 5921 -15947 5974 -15938
rect 6279 -15947 6332 -15938
rect 6634 -15947 6687 -15938
rect 6994 -15947 7047 -15941
rect 5921 -15948 7047 -15947
rect 5974 -16000 6279 -15948
rect 5921 -16011 5974 -16001
rect 6332 -16000 6634 -15948
rect 6279 -16011 6332 -16001
rect 6687 -15951 7047 -15948
rect 6687 -16000 6994 -15951
rect 6634 -16011 6687 -16001
rect 6994 -16014 7047 -16004
rect 7526 -15952 7579 -15943
rect 7881 -15952 7934 -15942
rect 8237 -15952 8290 -15942
rect 11441 -15952 11494 -15942
rect 11797 -15952 11850 -15942
rect 12154 -15952 12207 -15942
rect 12511 -15952 12564 -15942
rect 7526 -15953 7881 -15952
rect 7579 -16005 7881 -15953
rect 7934 -16005 8237 -15952
rect 8290 -16005 11441 -15952
rect 11494 -16005 11797 -15952
rect 11850 -16005 12154 -15952
rect 12207 -16005 12511 -15952
rect 7526 -16016 7579 -16006
rect 7881 -16015 7934 -16005
rect 8237 -16015 8290 -16005
rect 11441 -16015 11494 -16005
rect 11797 -16015 11850 -16005
rect 12154 -16015 12207 -16005
rect 12511 -16015 12564 -16005
rect -6159 -16193 -6106 -16183
rect -5504 -16193 -5451 -16183
rect -4792 -16193 -4739 -16183
rect -6106 -16246 -5504 -16193
rect -5451 -16246 -4792 -16193
rect -6159 -16256 -6106 -16246
rect -5504 -16256 -5451 -16246
rect -4792 -16256 -4739 -16246
rect -5860 -16294 -5807 -16284
rect -5148 -16294 -5095 -16284
rect -4436 -16294 -4383 -16284
rect -3935 -16294 -3883 -16285
rect -5807 -16347 -5148 -16294
rect -5095 -16346 -4436 -16294
rect -5860 -16357 -5807 -16347
rect -5148 -16357 -5095 -16347
rect -4383 -16295 -3883 -16294
rect -4383 -16346 -3935 -16295
rect -4436 -16357 -4383 -16347
rect -3935 -16357 -3883 -16347
rect -1917 -16542 -1864 -16532
rect -1738 -16542 -1685 -16532
rect -1561 -16541 -1508 -16531
rect -1864 -16595 -1738 -16542
rect -1685 -16594 -1561 -16542
rect -1381 -16542 -1328 -16533
rect -1204 -16542 -1151 -16532
rect -1026 -16542 -973 -16532
rect 220 -16542 273 -16532
rect 397 -16542 450 -16532
rect 576 -16542 629 -16532
rect 755 -16542 808 -16532
rect 933 -16542 986 -16532
rect 1111 -16542 1164 -16532
rect 2356 -16542 2409 -16532
rect 2534 -16542 2587 -16532
rect 2713 -16541 2766 -16531
rect -1508 -16543 -1204 -16542
rect -1508 -16594 -1381 -16543
rect -1685 -16595 -1381 -16594
rect -1917 -16605 -1864 -16595
rect -1738 -16605 -1685 -16595
rect -1561 -16604 -1508 -16595
rect -1328 -16595 -1204 -16543
rect -1151 -16595 -1026 -16542
rect -973 -16595 220 -16542
rect 273 -16595 397 -16542
rect 450 -16595 576 -16542
rect 629 -16595 755 -16542
rect 808 -16595 933 -16542
rect 986 -16595 1111 -16542
rect 1164 -16595 2356 -16542
rect 2409 -16595 2534 -16542
rect 2587 -16594 2713 -16542
rect 2891 -16542 2944 -16532
rect 3070 -16542 3123 -16532
rect 3249 -16542 3302 -16532
rect 4238 -16542 4291 -16532
rect 2766 -16594 2891 -16542
rect 2587 -16595 2891 -16594
rect 2944 -16595 3070 -16542
rect 3123 -16595 3249 -16542
rect 3302 -16595 4238 -16542
rect -1381 -16606 -1328 -16596
rect -1204 -16605 -1151 -16595
rect -1026 -16605 -973 -16595
rect 220 -16605 273 -16595
rect 397 -16605 450 -16595
rect 576 -16605 629 -16595
rect 755 -16605 808 -16595
rect 933 -16605 986 -16595
rect 1111 -16605 1164 -16595
rect 2356 -16605 2409 -16595
rect 2534 -16605 2587 -16595
rect 2713 -16604 2766 -16595
rect 2891 -16605 2944 -16595
rect 3070 -16605 3123 -16595
rect 3249 -16605 3302 -16595
rect 4238 -16605 4291 -16595
rect 6548 -16544 6601 -16534
rect 6726 -16544 6779 -16534
rect 6601 -16597 6726 -16545
rect 6903 -16545 6956 -16535
rect 7970 -16545 8023 -16535
rect 8149 -16544 8202 -16534
rect 6779 -16597 6903 -16545
rect 6548 -16598 6903 -16597
rect 6956 -16598 7970 -16545
rect 8023 -16597 8149 -16545
rect 9929 -16544 9982 -16534
rect 8202 -16597 9929 -16545
rect 10107 -16545 10160 -16535
rect 10287 -16545 10340 -16535
rect 11352 -16545 11405 -16535
rect 11530 -16545 11583 -16536
rect 11709 -16545 11762 -16535
rect 9982 -16597 10107 -16545
rect 8023 -16598 10107 -16597
rect 10160 -16598 10287 -16545
rect 10340 -16598 11352 -16545
rect 11405 -16546 11709 -16545
rect 11405 -16598 11530 -16546
rect 6548 -16607 6601 -16598
rect 6726 -16607 6779 -16598
rect 6903 -16608 6956 -16598
rect 7970 -16608 8023 -16598
rect 8149 -16607 8202 -16598
rect 9929 -16607 9982 -16598
rect 10107 -16608 10160 -16598
rect 10287 -16608 10340 -16598
rect 11352 -16608 11405 -16598
rect 11583 -16598 11709 -16546
rect 11530 -16609 11583 -16599
rect 11709 -16608 11762 -16598
rect -1827 -16665 -1774 -16655
rect -1720 -16665 -1548 -16655
rect -1471 -16665 -1418 -16656
rect -1114 -16665 -1061 -16655
rect -759 -16664 -706 -16654
rect -1774 -16718 -1720 -16665
rect -1548 -16666 -1114 -16665
rect -1548 -16718 -1471 -16666
rect -1827 -16728 -1774 -16718
rect -1720 -16728 -1548 -16718
rect -1418 -16718 -1114 -16666
rect -1061 -16717 -759 -16665
rect -646 -16665 -471 -16655
rect -403 -16665 -350 -16655
rect -47 -16665 6 -16655
rect 309 -16665 362 -16656
rect 426 -16665 595 -16655
rect 665 -16665 718 -16655
rect 1021 -16665 1074 -16655
rect 1377 -16665 1430 -16655
rect 1501 -16665 1671 -16655
rect 1735 -16665 1788 -16655
rect 2090 -16664 2143 -16654
rect -706 -16717 -646 -16665
rect -1061 -16718 -646 -16717
rect -471 -16718 -403 -16665
rect -350 -16718 -47 -16665
rect 6 -16666 426 -16665
rect 6 -16718 309 -16666
rect -1471 -16729 -1418 -16719
rect -1114 -16728 -1061 -16718
rect -759 -16727 -706 -16718
rect -646 -16728 -471 -16718
rect -403 -16728 -350 -16718
rect -47 -16728 6 -16718
rect 362 -16718 426 -16666
rect 595 -16718 665 -16665
rect 718 -16718 1021 -16665
rect 1074 -16718 1377 -16665
rect 1430 -16718 1501 -16665
rect 1671 -16718 1735 -16665
rect 1788 -16717 2090 -16665
rect 2445 -16665 2498 -16655
rect 2568 -16665 2732 -16655
rect 2801 -16665 2854 -16655
rect 3157 -16664 3210 -16654
rect 2143 -16717 2445 -16665
rect 1788 -16718 2445 -16717
rect 2498 -16718 2568 -16665
rect 2732 -16718 2801 -16665
rect 2854 -16717 3157 -16665
rect 3514 -16665 3567 -16656
rect 3633 -16665 3804 -16655
rect 3868 -16665 3921 -16655
rect 3210 -16666 3633 -16665
rect 3210 -16717 3514 -16666
rect 2854 -16718 3514 -16717
rect 309 -16729 362 -16719
rect 426 -16728 595 -16718
rect 665 -16728 718 -16718
rect 1021 -16728 1074 -16718
rect 1377 -16728 1430 -16718
rect 1501 -16728 1671 -16718
rect 1735 -16728 1788 -16718
rect 2090 -16727 2143 -16718
rect 2445 -16728 2498 -16718
rect 2568 -16728 2732 -16718
rect 2801 -16728 2854 -16718
rect 3157 -16727 3210 -16718
rect 3567 -16718 3633 -16666
rect 3804 -16718 3868 -16665
rect 3514 -16729 3567 -16719
rect 3633 -16728 3804 -16718
rect 3868 -16728 3921 -16718
rect 5399 -16666 5452 -16657
rect 8771 -16666 8824 -16656
rect 9128 -16666 9181 -16656
rect 9484 -16666 9537 -16656
rect 5399 -16667 8771 -16666
rect 5452 -16719 8771 -16667
rect 8824 -16719 9128 -16666
rect 9181 -16719 9484 -16666
rect 5399 -16730 5452 -16720
rect 8771 -16729 8824 -16719
rect 9128 -16729 9181 -16719
rect 9484 -16729 9537 -16719
rect 9838 -16665 9891 -16656
rect 10195 -16665 10248 -16655
rect 10550 -16665 10603 -16655
rect 10907 -16665 10960 -16655
rect 9838 -16666 10195 -16665
rect 9891 -16718 10195 -16666
rect 10248 -16718 10550 -16665
rect 10603 -16718 10907 -16665
rect 9838 -16729 9891 -16719
rect 10195 -16728 10248 -16718
rect 10550 -16728 10603 -16718
rect 10907 -16728 10960 -16718
rect 5031 -16782 5084 -16772
rect 8950 -16782 9003 -16772
rect 9305 -16782 9358 -16772
rect 5084 -16835 8950 -16782
rect 9003 -16835 9305 -16782
rect 5031 -16845 5084 -16835
rect 8950 -16845 9003 -16835
rect 9305 -16845 9358 -16835
rect 10017 -16780 10070 -16771
rect 10374 -16780 10427 -16771
rect 10731 -16779 10784 -16769
rect 10017 -16781 10731 -16780
rect 10070 -16833 10374 -16781
rect 10017 -16844 10070 -16834
rect 10427 -16832 10731 -16781
rect 10427 -16833 10784 -16832
rect 10374 -16844 10427 -16834
rect 10731 -16842 10784 -16833
rect -5682 -16886 -5629 -16876
rect -5326 -16886 -5273 -16876
rect -4970 -16886 -4917 -16876
rect -4614 -16886 -4561 -16876
rect -4258 -16886 -4205 -16876
rect -5629 -16939 -5326 -16886
rect -5273 -16939 -4970 -16886
rect -4917 -16939 -4614 -16886
rect -4561 -16939 -4258 -16886
rect -5682 -16949 -5629 -16939
rect -5326 -16949 -5273 -16939
rect -4970 -16949 -4917 -16939
rect -4614 -16949 -4561 -16939
rect -4258 -16949 -4205 -16939
rect 7347 -16890 7400 -16880
rect 7704 -16890 7757 -16880
rect 8060 -16890 8113 -16880
rect 8416 -16890 8469 -16880
rect 11263 -16890 11316 -16880
rect 11620 -16890 11673 -16880
rect 11975 -16889 12028 -16879
rect 7400 -16943 7704 -16890
rect 7757 -16943 8060 -16890
rect 8113 -16943 8416 -16890
rect 8469 -16943 11263 -16890
rect 11316 -16943 11620 -16890
rect 11673 -16942 11975 -16890
rect 12331 -16889 12384 -16879
rect 12028 -16942 12331 -16890
rect 11673 -16943 12384 -16942
rect 7347 -16953 7400 -16943
rect 7704 -16953 7757 -16943
rect 8060 -16953 8113 -16943
rect 8416 -16953 8469 -16943
rect 11263 -16953 11316 -16943
rect 11620 -16953 11673 -16943
rect 11975 -16952 12028 -16943
rect 12331 -16952 12384 -16943
rect -6159 -17007 -6106 -16997
rect -5859 -17007 -5806 -16997
rect -5148 -17007 -5095 -16997
rect -4437 -17007 -4384 -16997
rect -6106 -17060 -5859 -17007
rect -5806 -17060 -5148 -17007
rect -5095 -17060 -4437 -17007
rect -6159 -17070 -6106 -17060
rect -5859 -17070 -5806 -17060
rect -5148 -17070 -5095 -17060
rect -4437 -17070 -4384 -17060
rect -5504 -17118 -5451 -17108
rect -4792 -17118 -4739 -17108
rect -3935 -17118 -3883 -17108
rect -5451 -17170 -4792 -17118
rect -5504 -17181 -5451 -17171
rect -4739 -17170 -3935 -17118
rect -4792 -17181 -4739 -17171
rect -3935 -17180 -3883 -17170
<< via2 >>
rect 3019 -3513 3080 -3452
rect -2546 -3989 -2485 -3928
rect 2538 -4327 2599 -4266
rect -2385 -4566 -2324 -4505
rect 2746 -4507 2807 -4446
rect 3021 -5063 3082 -5002
rect -2385 -5154 -2324 -5093
rect 311 -5209 372 -5148
rect -1646 -5339 -1585 -5278
rect 846 -5339 907 -5278
rect -3545 -6867 -3484 -6806
rect -3386 -7040 -3325 -6979
<< metal3 >>
rect 6451 929 6515 2665
rect 6704 121 6768 1857
rect 17697 122 17761 1858
rect 17950 929 18014 2665
rect 3009 -3452 3090 -3447
rect 3009 -3513 3019 -3452
rect 3080 -3513 3090 -3452
rect 3009 -3518 3090 -3513
rect -2556 -3928 -2475 -3923
rect -2556 -3989 -2546 -3928
rect -2485 -3989 -2475 -3928
rect -2556 -3994 -2475 -3989
rect -2546 -4266 -2485 -3994
rect 2528 -4266 2609 -4261
rect -2546 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect -2546 -6637 -2485 -4327
rect 2528 -4332 2609 -4327
rect 2736 -4446 2817 -4441
rect -2385 -4500 2746 -4446
rect -2395 -4505 2746 -4500
rect -2395 -4566 -2385 -4505
rect -2324 -4507 2746 -4505
rect 2807 -4507 2817 -4446
rect -2324 -4566 -2314 -4507
rect 2736 -4512 2817 -4507
rect -2395 -4571 -2314 -4566
rect -2385 -5088 -2324 -4571
rect 3021 -4997 3082 -3518
rect 3011 -5002 3092 -4997
rect 3011 -5063 3021 -5002
rect 3082 -5063 3092 -5002
rect 3011 -5068 3092 -5063
rect -2395 -5093 -2314 -5088
rect -2395 -5154 -2385 -5093
rect -2324 -5154 -2314 -5093
rect -2395 -5159 -2314 -5154
rect 301 -5147 382 -5143
rect 3021 -5147 3082 -5068
rect 301 -5148 3082 -5147
rect -3545 -6698 -2485 -6637
rect -3545 -6801 -3484 -6698
rect -2385 -6786 -2324 -5159
rect 301 -5209 311 -5148
rect 372 -5208 3082 -5148
rect 372 -5209 382 -5208
rect 301 -5214 382 -5209
rect -1656 -5278 -1575 -5273
rect 836 -5278 917 -5273
rect -1656 -5339 -1646 -5278
rect -1585 -5339 846 -5278
rect 907 -5339 917 -5278
rect -1656 -5344 -1575 -5339
rect 836 -5344 917 -5339
rect 6451 -6271 6515 -4535
rect 6704 -5279 6768 -3543
rect -3555 -6806 -3474 -6801
rect -3555 -6867 -3545 -6806
rect -3484 -6867 -3474 -6806
rect -3555 -6872 -3474 -6867
rect -3386 -6847 -2324 -6786
rect -3386 -6974 -3325 -6847
rect -3396 -6979 -3315 -6974
rect -3396 -7040 -3386 -6979
rect -3325 -7040 -3315 -6979
rect -3396 -7045 -3315 -7040
rect 17697 -7078 17761 -5342
rect 17950 -6271 18014 -4535
use sc_cmfb  sc_cmfb_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/sc_cmfb
timestamp 1654517900
transform 1 0 9102 0 1 -5469
box -3494 -1840 9310 8360
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_0
timestamp 1654517900
transform 1 0 7953 0 1 -9022
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_1
timestamp 1654517900
transform 1 0 7953 0 1 -9922
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_2
timestamp 1654517900
transform 1 0 7953 0 1 -10822
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_AA  sky130_fd_pr__nfet_01v8_AA_3
timestamp 1654517900
transform 1 0 7953 0 1 -11722
box -1453 -228 1453 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_0
timestamp 1654517900
transform 1 0 -5032 0 1 -14522
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_1
timestamp 1654517900
transform 1 0 -5032 0 1 -15222
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_2
timestamp 1654517900
transform 1 0 -5032 0 1 -15922
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_BB  sky130_fd_pr__nfet_01v8_BB_3
timestamp 1654517900
transform 1 0 -5032 0 1 -16622
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_4
timestamp 1654517900
transform 1 0 959 0 1 -15260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_5
timestamp 1654517900
transform 1 0 959 0 1 -14260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_6
timestamp 1654517900
transform 1 0 959 0 1 -13260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_7
timestamp 1654517900
transform 1 0 959 0 1 -12260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_8
timestamp 1654517900
transform 1 0 959 0 1 -11260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_9
timestamp 1654517900
transform 1 0 959 0 1 -10260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_10
timestamp 1654517900
transform 1 0 959 0 1 -9260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_11
timestamp 1654517900
transform 1 0 959 0 1 -8260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_CC  sky130_fd_pr__nfet_01v8_CC_12
timestamp 1654517900
transform 1 0 959 0 1 -16260
box -3144 -228 3144 228
use sky130_fd_pr__nfet_01v8_DD  sky130_fd_pr__nfet_01v8_DD_0
timestamp 1654517900
transform 1 0 9154 0 1 -14260
box -3589 -228 3589 228
use sky130_fd_pr__nfet_01v8_DD  sky130_fd_pr__nfet_01v8_DD_1
timestamp 1654517900
transform 1 0 9154 0 1 -15260
box -3589 -228 3589 228
use sky130_fd_pr__nfet_01v8_DD  sky130_fd_pr__nfet_01v8_DD_2
timestamp 1654517900
transform 1 0 9154 0 1 -16260
box -3589 -228 3589 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_0
timestamp 1654517900
transform 1 0 11754 0 1 -9052
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_1
timestamp 1654517900
transform 1 0 11754 0 1 -9822
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_2
timestamp 1654517900
transform 1 0 11754 0 1 -10592
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_EE  sky130_fd_pr__nfet_01v8_EE_3
timestamp 1654517900
transform 1 0 11754 0 1 -11362
box -994 -228 994 228
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_0
timestamp 1654517900
transform 1 0 -5850 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_1
timestamp 1654517900
transform 1 0 -5850 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_2
timestamp 1654517900
transform 1 0 -5600 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_3
timestamp 1654517900
transform 1 0 -5350 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_4
timestamp 1654517900
transform 1 0 -5100 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_5
timestamp 1654517900
transform 1 0 -4850 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_6
timestamp 1654517900
transform 1 0 -4600 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_7
timestamp 1654517900
transform 1 0 -4350 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_8
timestamp 1654517900
transform 1 0 -4100 0 1 -13500
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_9
timestamp 1654517900
transform 1 0 -5600 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_10
timestamp 1654517900
transform 1 0 -5350 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_11
timestamp 1654517900
transform 1 0 -5100 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_12
timestamp 1654517900
transform 1 0 -4850 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_13
timestamp 1654517900
transform 1 0 -4600 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_14
timestamp 1654517900
transform 1 0 -4350 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_FF  sky130_fd_pr__nfet_01v8_lvt_FF_15
timestamp 1654517900
transform 1 0 -4100 0 1 -12820
box -78 -208 78 208
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_0
timestamp 1654517900
transform 1 0 -4810 0 1 -8002
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_1
timestamp 1654517900
transform 1 0 -4810 0 1 -8552
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_2
timestamp 1654517900
transform 1 0 -4810 0 1 -9102
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_3
timestamp 1654517900
transform 1 0 -4810 0 1 -9652
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_4
timestamp 1654517900
transform 1 0 -4810 0 1 -10202
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_5
timestamp 1654517900
transform 1 0 -4810 0 1 -10752
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_6
timestamp 1654517900
transform 1 0 -4810 0 1 -11302
box -830 -228 830 228
use sky130_fd_pr__nfet_01v8_lvt_GG  sky130_fd_pr__nfet_01v8_lvt_GG_7
timestamp 1654517900
transform 1 0 -4810 0 1 -11852
box -830 -228 830 228
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_0
timestamp 1654517900
transform 1 0 610 0 1 -3012
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_1
timestamp 1654517900
transform 1 0 610 0 1 -3912
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_2
timestamp 1654517900
transform 1 0 610 0 1 -4812
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_HH  sky130_fd_pr__pfet_01v8_HH_3
timestamp 1654517900
transform 1 0 610 0 1 -5712
box -2112 -240 2112 240
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_0
timestamp 1654517900
transform 1 0 -4861 0 1 -2260
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_1
timestamp 1654517900
transform 1 0 -4861 0 1 -3130
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_2
timestamp 1654517900
transform 1 0 -4861 0 1 -4000
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_3
timestamp 1654517900
transform 1 0 -4861 0 1 -4870
box -1489 -241 1489 241
use sky130_fd_pr__pfet_01v8_lvt_II  sky130_fd_pr__pfet_01v8_lvt_II_4
timestamp 1654517900
transform 1 0 -4861 0 1 -5740
box -1489 -241 1489 241
<< labels >>
flabel metal2 3147 -3484 3147 -3484 1 FreeSans 1200 0 0 0 on
port 8 n
flabel metal2 3431 -5243 3431 -5243 1 FreeSans 1200 0 0 0 op
port 7 n
flabel metal2 5049 -9956 5049 -9956 1 FreeSans 1200 0 0 0 cmc
port 15 n
flabel metal1 4262 -15741 4262 -15741 1 FreeSans 1200 0 0 0 bias_a
port 11 n
flabel metal1 6929 -13167 6929 -13167 1 FreeSans 1200 0 0 0 bias_d
port 14 n
flabel metal1 -7420 -1403 -7420 -1403 1 FreeSans 1200 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 -6957 -14245 -6957 -14245 1 FreeSans 1200 0 0 0 i_bias
port 9 n
flabel metal1 -3636 -12323 -3636 -12323 1 FreeSans 1200 0 0 0 bias_c
port 13 n
flabel metal1 -6950 -12541 -6950 -12541 1 FreeSans 1200 0 0 0 ip
port 1 n
flabel metal1 -6952 -13880 -6952 -13880 1 FreeSans 1200 0 0 0 in
port 2 n
flabel metal1 -4277 -7715 -4277 -7715 1 FreeSans 1200 0 0 0 bias_b
port 12 n
flabel metal1 7057 2874 7057 2874 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 7057 1707 7057 1707 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 7058 -83 7058 -83 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 7058 -739 7058 -739 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 7058 -1885 7058 -1885 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 7058 -2537 7058 -2537 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 7051 -4329 7051 -4329 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 7054 -5489 7054 -5489 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 7054 -7288 7054 -7288 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16056 -7290 16056 -7290 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16057 -6136 16057 -6136 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 16055 -5482 16055 -5482 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16057 -2529 16057 -2529 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 16055 -1886 16055 -1886 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16057 -86 16057 -86 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16057 1070 16057 1070 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 16057 1716 16057 1716 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16057 2870 16057 2870 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal3 6479 2585 6479 2585 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal3 6738 1807 6738 1807 1 FreeSans 400 0 0 0 p2
port 5 n
flabel metal3 6486 -6211 6486 -6211 1 FreeSans 400 0 0 0 p1_b
port 4 n
flabel metal3 6735 -5207 6735 -5207 1 FreeSans 400 0 0 0 p1
port 3 n
flabel metal3 17730 1821 17730 1821 1 FreeSans 400 0 0 0 p2
port 5 n
flabel metal3 17980 2631 17980 2631 1 FreeSans 400 0 0 0 p2_b
port 6 n
flabel metal3 17727 -7023 17727 -7023 1 FreeSans 400 0 0 0 p1
port 3 n
flabel metal3 17984 -6236 17984 -6236 1 FreeSans 400 0 0 0 p1_b
port 4 n
flabel metal2 17862 -8732 17862 -8732 1 FreeSans 800 0 0 0 cm
port 10 n
flabel metal1 7058 1058 7058 1058 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 7058 -3672 7058 -3672 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 7058 -6144 7058 -6144 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 16056 -4338 16056 -4338 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 16056 -3678 16056 -3678 1 FreeSans 400 0 0 0 VSS
port 17 n power bidirectional
flabel metal1 16056 -738 16056 -738 1 FreeSans 400 0 0 0 VDD
port 16 n power bidirectional
flabel metal1 1056 -17349 1056 -17349 1 FreeSans 1600 0 0 0 VSS
port 17 n power bidirectional
<< end >>
