magic
tech sky130A
magscale 1 2
timestamp 1655456512
<< error_p >>
rect -4124 181 -4066 187
rect -3704 181 -3646 187
rect -3284 181 -3226 187
rect -2864 181 -2806 187
rect -2444 181 -2386 187
rect -2024 181 -1966 187
rect -1604 181 -1546 187
rect -1184 181 -1126 187
rect -764 181 -706 187
rect -344 181 -286 187
rect 76 181 134 187
rect 496 181 554 187
rect 916 181 974 187
rect 1336 181 1394 187
rect 1756 181 1814 187
rect 2176 181 2234 187
rect 2596 181 2654 187
rect 3016 181 3074 187
rect 3436 181 3494 187
rect 3856 181 3914 187
rect -4124 147 -4112 181
rect -3704 147 -3692 181
rect -3284 147 -3272 181
rect -2864 147 -2852 181
rect -2444 147 -2432 181
rect -2024 147 -2012 181
rect -1604 147 -1592 181
rect -1184 147 -1172 181
rect -764 147 -752 181
rect -344 147 -332 181
rect 76 147 88 181
rect 496 147 508 181
rect 916 147 928 181
rect 1336 147 1348 181
rect 1756 147 1768 181
rect 2176 147 2188 181
rect 2596 147 2608 181
rect 3016 147 3028 181
rect 3436 147 3448 181
rect 3856 147 3868 181
rect -4124 141 -4066 147
rect -3704 141 -3646 147
rect -3284 141 -3226 147
rect -2864 141 -2806 147
rect -2444 141 -2386 147
rect -2024 141 -1966 147
rect -1604 141 -1546 147
rect -1184 141 -1126 147
rect -764 141 -706 147
rect -344 141 -286 147
rect 76 141 134 147
rect 496 141 554 147
rect 916 141 974 147
rect 1336 141 1394 147
rect 1756 141 1814 147
rect 2176 141 2234 147
rect 2596 141 2654 147
rect 3016 141 3074 147
rect 3436 141 3494 147
rect 3856 141 3914 147
rect -3914 -147 -3856 -141
rect -3494 -147 -3436 -141
rect -3074 -147 -3016 -141
rect -2654 -147 -2596 -141
rect -2234 -147 -2176 -141
rect -1814 -147 -1756 -141
rect -1394 -147 -1336 -141
rect -974 -147 -916 -141
rect -554 -147 -496 -141
rect -134 -147 -76 -141
rect 286 -147 344 -141
rect 706 -147 764 -141
rect 1126 -147 1184 -141
rect 1546 -147 1604 -141
rect 1966 -147 2024 -141
rect 2386 -147 2444 -141
rect 2806 -147 2864 -141
rect 3226 -147 3284 -141
rect 3646 -147 3704 -141
rect 4066 -147 4124 -141
rect -3914 -181 -3902 -147
rect -3494 -181 -3482 -147
rect -3074 -181 -3062 -147
rect -2654 -181 -2642 -147
rect -2234 -181 -2222 -147
rect -1814 -181 -1802 -147
rect -1394 -181 -1382 -147
rect -974 -181 -962 -147
rect -554 -181 -542 -147
rect -134 -181 -122 -147
rect 286 -181 298 -147
rect 706 -181 718 -147
rect 1126 -181 1138 -147
rect 1546 -181 1558 -147
rect 1966 -181 1978 -147
rect 2386 -181 2398 -147
rect 2806 -181 2818 -147
rect 3226 -181 3238 -147
rect 3646 -181 3658 -147
rect 4066 -181 4078 -147
rect -3914 -187 -3856 -181
rect -3494 -187 -3436 -181
rect -3074 -187 -3016 -181
rect -2654 -187 -2596 -181
rect -2234 -187 -2176 -181
rect -1814 -187 -1756 -181
rect -1394 -187 -1336 -181
rect -974 -187 -916 -181
rect -554 -187 -496 -181
rect -134 -187 -76 -181
rect 286 -187 344 -181
rect 706 -187 764 -181
rect 1126 -187 1184 -181
rect 1546 -187 1604 -181
rect 1966 -187 2024 -181
rect 2386 -187 2444 -181
rect 2806 -187 2864 -181
rect 3226 -187 3284 -181
rect 3646 -187 3704 -181
rect 4066 -187 4124 -181
rect -4122 -351 -4064 -345
rect -3702 -351 -3644 -345
rect -3282 -351 -3224 -345
rect -2862 -351 -2804 -345
rect -2442 -351 -2384 -345
rect -2022 -351 -1964 -345
rect -1602 -351 -1544 -345
rect -1182 -351 -1124 -345
rect -762 -351 -704 -345
rect -342 -351 -284 -345
rect 78 -351 136 -345
rect 498 -351 556 -345
rect 918 -351 976 -345
rect 1338 -351 1396 -345
rect 1758 -351 1816 -345
rect 2178 -351 2236 -345
rect 2598 -351 2656 -345
rect 3018 -351 3076 -345
rect 3438 -351 3496 -345
rect 3858 -351 3916 -345
rect -4122 -385 -4110 -351
rect -3702 -385 -3690 -351
rect -3282 -385 -3270 -351
rect -2862 -385 -2850 -351
rect -2442 -385 -2430 -351
rect -2022 -385 -2010 -351
rect -1602 -385 -1590 -351
rect -1182 -385 -1170 -351
rect -762 -385 -750 -351
rect -342 -385 -330 -351
rect 78 -385 90 -351
rect 498 -385 510 -351
rect 918 -385 930 -351
rect 1338 -385 1350 -351
rect 1758 -385 1770 -351
rect 2178 -385 2190 -351
rect 2598 -385 2610 -351
rect 3018 -385 3030 -351
rect 3438 -385 3450 -351
rect 3858 -385 3870 -351
rect -4122 -391 -4064 -385
rect -3702 -391 -3644 -385
rect -3282 -391 -3224 -385
rect -2862 -391 -2804 -385
rect -2442 -391 -2384 -385
rect -2022 -391 -1964 -385
rect -1602 -391 -1544 -385
rect -1182 -391 -1124 -385
rect -762 -391 -704 -385
rect -342 -391 -284 -385
rect 78 -391 136 -385
rect 498 -391 556 -385
rect 918 -391 976 -385
rect 1338 -391 1396 -385
rect 1758 -391 1816 -385
rect 2178 -391 2236 -385
rect 2598 -391 2656 -385
rect 3018 -391 3076 -385
rect 3438 -391 3496 -385
rect 3858 -391 3916 -385
rect -3912 -680 -3854 -674
rect -3492 -680 -3434 -674
rect -3072 -680 -3014 -674
rect -2652 -680 -2594 -674
rect -2232 -680 -2174 -674
rect -1812 -680 -1754 -674
rect -1392 -680 -1334 -674
rect -972 -680 -914 -674
rect -552 -680 -494 -674
rect -132 -680 -74 -674
rect 288 -680 346 -674
rect 708 -680 766 -674
rect 1128 -680 1186 -674
rect 1548 -680 1606 -674
rect 1968 -680 2026 -674
rect 2388 -680 2446 -674
rect 2808 -680 2866 -674
rect 3228 -680 3286 -674
rect 3648 -680 3706 -674
rect 4068 -680 4126 -674
rect -3912 -714 -3900 -680
rect -3492 -714 -3480 -680
rect -3072 -714 -3060 -680
rect -2652 -714 -2640 -680
rect -2232 -714 -2220 -680
rect -1812 -714 -1800 -680
rect -1392 -714 -1380 -680
rect -972 -714 -960 -680
rect -552 -714 -540 -680
rect -132 -714 -120 -680
rect 288 -714 300 -680
rect 708 -714 720 -680
rect 1128 -714 1140 -680
rect 1548 -714 1560 -680
rect 1968 -714 1980 -680
rect 2388 -714 2400 -680
rect 2808 -714 2820 -680
rect 3228 -714 3240 -680
rect 3648 -714 3660 -680
rect 4068 -714 4080 -680
rect -3912 -720 -3854 -714
rect -3492 -720 -3434 -714
rect -3072 -720 -3014 -714
rect -2652 -720 -2594 -714
rect -2232 -720 -2174 -714
rect -1812 -720 -1754 -714
rect -1392 -720 -1334 -714
rect -972 -720 -914 -714
rect -552 -720 -494 -714
rect -132 -720 -74 -714
rect 288 -720 346 -714
rect 708 -720 766 -714
rect 1128 -720 1186 -714
rect 1548 -720 1606 -714
rect 1968 -720 2026 -714
rect 2388 -720 2446 -714
rect 2808 -720 2866 -714
rect 3228 -720 3286 -714
rect 3648 -720 3706 -714
rect 4068 -720 4126 -714
<< nwell >>
rect -4520 -852 4520 319
<< pmos >>
rect -4320 -100 -4290 100
rect -4110 -100 -4080 100
rect -3900 -100 -3870 100
rect -3690 -100 -3660 100
rect -3480 -100 -3450 100
rect -3270 -100 -3240 100
rect -3060 -100 -3030 100
rect -2850 -100 -2820 100
rect -2640 -100 -2610 100
rect -2430 -100 -2400 100
rect -2220 -100 -2190 100
rect -2010 -100 -1980 100
rect -1800 -100 -1770 100
rect -1590 -100 -1560 100
rect -1380 -100 -1350 100
rect -1170 -100 -1140 100
rect -960 -100 -930 100
rect -750 -100 -720 100
rect -540 -100 -510 100
rect -330 -100 -300 100
rect -120 -100 -90 100
rect 90 -100 120 100
rect 300 -100 330 100
rect 510 -100 540 100
rect 720 -100 750 100
rect 930 -100 960 100
rect 1140 -100 1170 100
rect 1350 -100 1380 100
rect 1560 -100 1590 100
rect 1770 -100 1800 100
rect 1980 -100 2010 100
rect 2190 -100 2220 100
rect 2400 -100 2430 100
rect 2610 -100 2640 100
rect 2820 -100 2850 100
rect 3030 -100 3060 100
rect 3240 -100 3270 100
rect 3450 -100 3480 100
rect 3660 -100 3690 100
rect 3870 -100 3900 100
rect 4080 -100 4110 100
rect 4290 -100 4320 100
rect -4318 -633 -4288 -433
rect -4108 -633 -4078 -433
rect -3898 -633 -3868 -433
rect -3688 -633 -3658 -433
rect -3478 -633 -3448 -433
rect -3268 -633 -3238 -433
rect -3058 -633 -3028 -433
rect -2848 -633 -2818 -433
rect -2638 -633 -2608 -433
rect -2428 -633 -2398 -433
rect -2218 -633 -2188 -433
rect -2008 -633 -1978 -433
rect -1798 -633 -1768 -433
rect -1588 -633 -1558 -433
rect -1378 -633 -1348 -433
rect -1168 -633 -1138 -433
rect -958 -633 -928 -433
rect -748 -633 -718 -433
rect -538 -633 -508 -433
rect -328 -633 -298 -433
rect -118 -633 -88 -433
rect 92 -633 122 -433
rect 302 -633 332 -433
rect 512 -633 542 -433
rect 722 -633 752 -433
rect 932 -633 962 -433
rect 1142 -633 1172 -433
rect 1352 -633 1382 -433
rect 1562 -633 1592 -433
rect 1772 -633 1802 -433
rect 1982 -633 2012 -433
rect 2192 -633 2222 -433
rect 2402 -633 2432 -433
rect 2612 -633 2642 -433
rect 2822 -633 2852 -433
rect 3032 -633 3062 -433
rect 3242 -633 3272 -433
rect 3452 -633 3482 -433
rect 3662 -633 3692 -433
rect 3872 -633 3902 -433
rect 4082 -633 4112 -433
rect 4292 -633 4322 -433
<< pdiff >>
rect -4382 88 -4320 100
rect -4382 -88 -4370 88
rect -4336 -88 -4320 88
rect -4382 -100 -4320 -88
rect -4290 88 -4228 100
rect -4290 -88 -4274 88
rect -4240 -88 -4228 88
rect -4290 -100 -4228 -88
rect -4172 88 -4110 100
rect -4172 -88 -4160 88
rect -4126 -88 -4110 88
rect -4172 -100 -4110 -88
rect -4080 88 -4018 100
rect -4080 -88 -4064 88
rect -4030 -88 -4018 88
rect -4080 -100 -4018 -88
rect -3962 88 -3900 100
rect -3962 -88 -3950 88
rect -3916 -88 -3900 88
rect -3962 -100 -3900 -88
rect -3870 88 -3808 100
rect -3870 -88 -3854 88
rect -3820 -88 -3808 88
rect -3870 -100 -3808 -88
rect -3752 88 -3690 100
rect -3752 -88 -3740 88
rect -3706 -88 -3690 88
rect -3752 -100 -3690 -88
rect -3660 88 -3598 100
rect -3660 -88 -3644 88
rect -3610 -88 -3598 88
rect -3660 -100 -3598 -88
rect -3542 88 -3480 100
rect -3542 -88 -3530 88
rect -3496 -88 -3480 88
rect -3542 -100 -3480 -88
rect -3450 88 -3388 100
rect -3450 -88 -3434 88
rect -3400 -88 -3388 88
rect -3450 -100 -3388 -88
rect -3332 88 -3270 100
rect -3332 -88 -3320 88
rect -3286 -88 -3270 88
rect -3332 -100 -3270 -88
rect -3240 88 -3178 100
rect -3240 -88 -3224 88
rect -3190 -88 -3178 88
rect -3240 -100 -3178 -88
rect -3122 88 -3060 100
rect -3122 -88 -3110 88
rect -3076 -88 -3060 88
rect -3122 -100 -3060 -88
rect -3030 88 -2968 100
rect -3030 -88 -3014 88
rect -2980 -88 -2968 88
rect -3030 -100 -2968 -88
rect -2912 88 -2850 100
rect -2912 -88 -2900 88
rect -2866 -88 -2850 88
rect -2912 -100 -2850 -88
rect -2820 88 -2758 100
rect -2820 -88 -2804 88
rect -2770 -88 -2758 88
rect -2820 -100 -2758 -88
rect -2702 88 -2640 100
rect -2702 -88 -2690 88
rect -2656 -88 -2640 88
rect -2702 -100 -2640 -88
rect -2610 88 -2548 100
rect -2610 -88 -2594 88
rect -2560 -88 -2548 88
rect -2610 -100 -2548 -88
rect -2492 88 -2430 100
rect -2492 -88 -2480 88
rect -2446 -88 -2430 88
rect -2492 -100 -2430 -88
rect -2400 88 -2338 100
rect -2400 -88 -2384 88
rect -2350 -88 -2338 88
rect -2400 -100 -2338 -88
rect -2282 88 -2220 100
rect -2282 -88 -2270 88
rect -2236 -88 -2220 88
rect -2282 -100 -2220 -88
rect -2190 88 -2128 100
rect -2190 -88 -2174 88
rect -2140 -88 -2128 88
rect -2190 -100 -2128 -88
rect -2072 88 -2010 100
rect -2072 -88 -2060 88
rect -2026 -88 -2010 88
rect -2072 -100 -2010 -88
rect -1980 88 -1918 100
rect -1980 -88 -1964 88
rect -1930 -88 -1918 88
rect -1980 -100 -1918 -88
rect -1862 88 -1800 100
rect -1862 -88 -1850 88
rect -1816 -88 -1800 88
rect -1862 -100 -1800 -88
rect -1770 88 -1708 100
rect -1770 -88 -1754 88
rect -1720 -88 -1708 88
rect -1770 -100 -1708 -88
rect -1652 88 -1590 100
rect -1652 -88 -1640 88
rect -1606 -88 -1590 88
rect -1652 -100 -1590 -88
rect -1560 88 -1498 100
rect -1560 -88 -1544 88
rect -1510 -88 -1498 88
rect -1560 -100 -1498 -88
rect -1442 88 -1380 100
rect -1442 -88 -1430 88
rect -1396 -88 -1380 88
rect -1442 -100 -1380 -88
rect -1350 88 -1288 100
rect -1350 -88 -1334 88
rect -1300 -88 -1288 88
rect -1350 -100 -1288 -88
rect -1232 88 -1170 100
rect -1232 -88 -1220 88
rect -1186 -88 -1170 88
rect -1232 -100 -1170 -88
rect -1140 88 -1078 100
rect -1140 -88 -1124 88
rect -1090 -88 -1078 88
rect -1140 -100 -1078 -88
rect -1022 88 -960 100
rect -1022 -88 -1010 88
rect -976 -88 -960 88
rect -1022 -100 -960 -88
rect -930 88 -868 100
rect -930 -88 -914 88
rect -880 -88 -868 88
rect -930 -100 -868 -88
rect -812 88 -750 100
rect -812 -88 -800 88
rect -766 -88 -750 88
rect -812 -100 -750 -88
rect -720 88 -658 100
rect -720 -88 -704 88
rect -670 -88 -658 88
rect -720 -100 -658 -88
rect -602 88 -540 100
rect -602 -88 -590 88
rect -556 -88 -540 88
rect -602 -100 -540 -88
rect -510 88 -448 100
rect -510 -88 -494 88
rect -460 -88 -448 88
rect -510 -100 -448 -88
rect -392 88 -330 100
rect -392 -88 -380 88
rect -346 -88 -330 88
rect -392 -100 -330 -88
rect -300 88 -238 100
rect -300 -88 -284 88
rect -250 -88 -238 88
rect -300 -100 -238 -88
rect -182 88 -120 100
rect -182 -88 -170 88
rect -136 -88 -120 88
rect -182 -100 -120 -88
rect -90 88 -28 100
rect -90 -88 -74 88
rect -40 -88 -28 88
rect -90 -100 -28 -88
rect 28 88 90 100
rect 28 -88 40 88
rect 74 -88 90 88
rect 28 -100 90 -88
rect 120 88 182 100
rect 120 -88 136 88
rect 170 -88 182 88
rect 120 -100 182 -88
rect 238 88 300 100
rect 238 -88 250 88
rect 284 -88 300 88
rect 238 -100 300 -88
rect 330 88 392 100
rect 330 -88 346 88
rect 380 -88 392 88
rect 330 -100 392 -88
rect 448 88 510 100
rect 448 -88 460 88
rect 494 -88 510 88
rect 448 -100 510 -88
rect 540 88 602 100
rect 540 -88 556 88
rect 590 -88 602 88
rect 540 -100 602 -88
rect 658 88 720 100
rect 658 -88 670 88
rect 704 -88 720 88
rect 658 -100 720 -88
rect 750 88 812 100
rect 750 -88 766 88
rect 800 -88 812 88
rect 750 -100 812 -88
rect 868 88 930 100
rect 868 -88 880 88
rect 914 -88 930 88
rect 868 -100 930 -88
rect 960 88 1022 100
rect 960 -88 976 88
rect 1010 -88 1022 88
rect 960 -100 1022 -88
rect 1078 88 1140 100
rect 1078 -88 1090 88
rect 1124 -88 1140 88
rect 1078 -100 1140 -88
rect 1170 88 1232 100
rect 1170 -88 1186 88
rect 1220 -88 1232 88
rect 1170 -100 1232 -88
rect 1288 88 1350 100
rect 1288 -88 1300 88
rect 1334 -88 1350 88
rect 1288 -100 1350 -88
rect 1380 88 1442 100
rect 1380 -88 1396 88
rect 1430 -88 1442 88
rect 1380 -100 1442 -88
rect 1498 88 1560 100
rect 1498 -88 1510 88
rect 1544 -88 1560 88
rect 1498 -100 1560 -88
rect 1590 88 1652 100
rect 1590 -88 1606 88
rect 1640 -88 1652 88
rect 1590 -100 1652 -88
rect 1708 88 1770 100
rect 1708 -88 1720 88
rect 1754 -88 1770 88
rect 1708 -100 1770 -88
rect 1800 88 1862 100
rect 1800 -88 1816 88
rect 1850 -88 1862 88
rect 1800 -100 1862 -88
rect 1918 88 1980 100
rect 1918 -88 1930 88
rect 1964 -88 1980 88
rect 1918 -100 1980 -88
rect 2010 88 2072 100
rect 2010 -88 2026 88
rect 2060 -88 2072 88
rect 2010 -100 2072 -88
rect 2128 88 2190 100
rect 2128 -88 2140 88
rect 2174 -88 2190 88
rect 2128 -100 2190 -88
rect 2220 88 2282 100
rect 2220 -88 2236 88
rect 2270 -88 2282 88
rect 2220 -100 2282 -88
rect 2338 88 2400 100
rect 2338 -88 2350 88
rect 2384 -88 2400 88
rect 2338 -100 2400 -88
rect 2430 88 2492 100
rect 2430 -88 2446 88
rect 2480 -88 2492 88
rect 2430 -100 2492 -88
rect 2548 88 2610 100
rect 2548 -88 2560 88
rect 2594 -88 2610 88
rect 2548 -100 2610 -88
rect 2640 88 2702 100
rect 2640 -88 2656 88
rect 2690 -88 2702 88
rect 2640 -100 2702 -88
rect 2758 88 2820 100
rect 2758 -88 2770 88
rect 2804 -88 2820 88
rect 2758 -100 2820 -88
rect 2850 88 2912 100
rect 2850 -88 2866 88
rect 2900 -88 2912 88
rect 2850 -100 2912 -88
rect 2968 88 3030 100
rect 2968 -88 2980 88
rect 3014 -88 3030 88
rect 2968 -100 3030 -88
rect 3060 88 3122 100
rect 3060 -88 3076 88
rect 3110 -88 3122 88
rect 3060 -100 3122 -88
rect 3178 88 3240 100
rect 3178 -88 3190 88
rect 3224 -88 3240 88
rect 3178 -100 3240 -88
rect 3270 88 3332 100
rect 3270 -88 3286 88
rect 3320 -88 3332 88
rect 3270 -100 3332 -88
rect 3388 88 3450 100
rect 3388 -88 3400 88
rect 3434 -88 3450 88
rect 3388 -100 3450 -88
rect 3480 88 3542 100
rect 3480 -88 3496 88
rect 3530 -88 3542 88
rect 3480 -100 3542 -88
rect 3598 88 3660 100
rect 3598 -88 3610 88
rect 3644 -88 3660 88
rect 3598 -100 3660 -88
rect 3690 88 3752 100
rect 3690 -88 3706 88
rect 3740 -88 3752 88
rect 3690 -100 3752 -88
rect 3808 88 3870 100
rect 3808 -88 3820 88
rect 3854 -88 3870 88
rect 3808 -100 3870 -88
rect 3900 88 3962 100
rect 3900 -88 3916 88
rect 3950 -88 3962 88
rect 3900 -100 3962 -88
rect 4018 88 4080 100
rect 4018 -88 4030 88
rect 4064 -88 4080 88
rect 4018 -100 4080 -88
rect 4110 88 4172 100
rect 4110 -88 4126 88
rect 4160 -88 4172 88
rect 4110 -100 4172 -88
rect 4228 88 4290 100
rect 4228 -88 4240 88
rect 4274 -88 4290 88
rect 4228 -100 4290 -88
rect 4320 88 4382 100
rect 4320 -88 4336 88
rect 4370 -88 4382 88
rect 4320 -100 4382 -88
rect -4380 -445 -4318 -433
rect -4380 -621 -4368 -445
rect -4334 -621 -4318 -445
rect -4380 -633 -4318 -621
rect -4288 -445 -4226 -433
rect -4288 -621 -4272 -445
rect -4238 -621 -4226 -445
rect -4288 -633 -4226 -621
rect -4170 -445 -4108 -433
rect -4170 -621 -4158 -445
rect -4124 -621 -4108 -445
rect -4170 -633 -4108 -621
rect -4078 -445 -4016 -433
rect -4078 -621 -4062 -445
rect -4028 -621 -4016 -445
rect -4078 -633 -4016 -621
rect -3960 -445 -3898 -433
rect -3960 -621 -3948 -445
rect -3914 -621 -3898 -445
rect -3960 -633 -3898 -621
rect -3868 -445 -3806 -433
rect -3868 -621 -3852 -445
rect -3818 -621 -3806 -445
rect -3868 -633 -3806 -621
rect -3750 -445 -3688 -433
rect -3750 -621 -3738 -445
rect -3704 -621 -3688 -445
rect -3750 -633 -3688 -621
rect -3658 -445 -3596 -433
rect -3658 -621 -3642 -445
rect -3608 -621 -3596 -445
rect -3658 -633 -3596 -621
rect -3540 -445 -3478 -433
rect -3540 -621 -3528 -445
rect -3494 -621 -3478 -445
rect -3540 -633 -3478 -621
rect -3448 -445 -3386 -433
rect -3448 -621 -3432 -445
rect -3398 -621 -3386 -445
rect -3448 -633 -3386 -621
rect -3330 -445 -3268 -433
rect -3330 -621 -3318 -445
rect -3284 -621 -3268 -445
rect -3330 -633 -3268 -621
rect -3238 -445 -3176 -433
rect -3238 -621 -3222 -445
rect -3188 -621 -3176 -445
rect -3238 -633 -3176 -621
rect -3120 -445 -3058 -433
rect -3120 -621 -3108 -445
rect -3074 -621 -3058 -445
rect -3120 -633 -3058 -621
rect -3028 -445 -2966 -433
rect -3028 -621 -3012 -445
rect -2978 -621 -2966 -445
rect -3028 -633 -2966 -621
rect -2910 -445 -2848 -433
rect -2910 -621 -2898 -445
rect -2864 -621 -2848 -445
rect -2910 -633 -2848 -621
rect -2818 -445 -2756 -433
rect -2818 -621 -2802 -445
rect -2768 -621 -2756 -445
rect -2818 -633 -2756 -621
rect -2700 -445 -2638 -433
rect -2700 -621 -2688 -445
rect -2654 -621 -2638 -445
rect -2700 -633 -2638 -621
rect -2608 -445 -2546 -433
rect -2608 -621 -2592 -445
rect -2558 -621 -2546 -445
rect -2608 -633 -2546 -621
rect -2490 -445 -2428 -433
rect -2490 -621 -2478 -445
rect -2444 -621 -2428 -445
rect -2490 -633 -2428 -621
rect -2398 -445 -2336 -433
rect -2398 -621 -2382 -445
rect -2348 -621 -2336 -445
rect -2398 -633 -2336 -621
rect -2280 -445 -2218 -433
rect -2280 -621 -2268 -445
rect -2234 -621 -2218 -445
rect -2280 -633 -2218 -621
rect -2188 -445 -2126 -433
rect -2188 -621 -2172 -445
rect -2138 -621 -2126 -445
rect -2188 -633 -2126 -621
rect -2070 -445 -2008 -433
rect -2070 -621 -2058 -445
rect -2024 -621 -2008 -445
rect -2070 -633 -2008 -621
rect -1978 -445 -1916 -433
rect -1978 -621 -1962 -445
rect -1928 -621 -1916 -445
rect -1978 -633 -1916 -621
rect -1860 -445 -1798 -433
rect -1860 -621 -1848 -445
rect -1814 -621 -1798 -445
rect -1860 -633 -1798 -621
rect -1768 -445 -1706 -433
rect -1768 -621 -1752 -445
rect -1718 -621 -1706 -445
rect -1768 -633 -1706 -621
rect -1650 -445 -1588 -433
rect -1650 -621 -1638 -445
rect -1604 -621 -1588 -445
rect -1650 -633 -1588 -621
rect -1558 -445 -1496 -433
rect -1558 -621 -1542 -445
rect -1508 -621 -1496 -445
rect -1558 -633 -1496 -621
rect -1440 -445 -1378 -433
rect -1440 -621 -1428 -445
rect -1394 -621 -1378 -445
rect -1440 -633 -1378 -621
rect -1348 -445 -1286 -433
rect -1348 -621 -1332 -445
rect -1298 -621 -1286 -445
rect -1348 -633 -1286 -621
rect -1230 -445 -1168 -433
rect -1230 -621 -1218 -445
rect -1184 -621 -1168 -445
rect -1230 -633 -1168 -621
rect -1138 -445 -1076 -433
rect -1138 -621 -1122 -445
rect -1088 -621 -1076 -445
rect -1138 -633 -1076 -621
rect -1020 -445 -958 -433
rect -1020 -621 -1008 -445
rect -974 -621 -958 -445
rect -1020 -633 -958 -621
rect -928 -445 -866 -433
rect -928 -621 -912 -445
rect -878 -621 -866 -445
rect -928 -633 -866 -621
rect -810 -445 -748 -433
rect -810 -621 -798 -445
rect -764 -621 -748 -445
rect -810 -633 -748 -621
rect -718 -445 -656 -433
rect -718 -621 -702 -445
rect -668 -621 -656 -445
rect -718 -633 -656 -621
rect -600 -445 -538 -433
rect -600 -621 -588 -445
rect -554 -621 -538 -445
rect -600 -633 -538 -621
rect -508 -445 -446 -433
rect -508 -621 -492 -445
rect -458 -621 -446 -445
rect -508 -633 -446 -621
rect -390 -445 -328 -433
rect -390 -621 -378 -445
rect -344 -621 -328 -445
rect -390 -633 -328 -621
rect -298 -445 -236 -433
rect -298 -621 -282 -445
rect -248 -621 -236 -445
rect -298 -633 -236 -621
rect -180 -445 -118 -433
rect -180 -621 -168 -445
rect -134 -621 -118 -445
rect -180 -633 -118 -621
rect -88 -445 -26 -433
rect -88 -621 -72 -445
rect -38 -621 -26 -445
rect -88 -633 -26 -621
rect 30 -445 92 -433
rect 30 -621 42 -445
rect 76 -621 92 -445
rect 30 -633 92 -621
rect 122 -445 184 -433
rect 122 -621 138 -445
rect 172 -621 184 -445
rect 122 -633 184 -621
rect 240 -445 302 -433
rect 240 -621 252 -445
rect 286 -621 302 -445
rect 240 -633 302 -621
rect 332 -445 394 -433
rect 332 -621 348 -445
rect 382 -621 394 -445
rect 332 -633 394 -621
rect 450 -445 512 -433
rect 450 -621 462 -445
rect 496 -621 512 -445
rect 450 -633 512 -621
rect 542 -445 604 -433
rect 542 -621 558 -445
rect 592 -621 604 -445
rect 542 -633 604 -621
rect 660 -445 722 -433
rect 660 -621 672 -445
rect 706 -621 722 -445
rect 660 -633 722 -621
rect 752 -445 814 -433
rect 752 -621 768 -445
rect 802 -621 814 -445
rect 752 -633 814 -621
rect 870 -445 932 -433
rect 870 -621 882 -445
rect 916 -621 932 -445
rect 870 -633 932 -621
rect 962 -445 1024 -433
rect 962 -621 978 -445
rect 1012 -621 1024 -445
rect 962 -633 1024 -621
rect 1080 -445 1142 -433
rect 1080 -621 1092 -445
rect 1126 -621 1142 -445
rect 1080 -633 1142 -621
rect 1172 -445 1234 -433
rect 1172 -621 1188 -445
rect 1222 -621 1234 -445
rect 1172 -633 1234 -621
rect 1290 -445 1352 -433
rect 1290 -621 1302 -445
rect 1336 -621 1352 -445
rect 1290 -633 1352 -621
rect 1382 -445 1444 -433
rect 1382 -621 1398 -445
rect 1432 -621 1444 -445
rect 1382 -633 1444 -621
rect 1500 -445 1562 -433
rect 1500 -621 1512 -445
rect 1546 -621 1562 -445
rect 1500 -633 1562 -621
rect 1592 -445 1654 -433
rect 1592 -621 1608 -445
rect 1642 -621 1654 -445
rect 1592 -633 1654 -621
rect 1710 -445 1772 -433
rect 1710 -621 1722 -445
rect 1756 -621 1772 -445
rect 1710 -633 1772 -621
rect 1802 -445 1864 -433
rect 1802 -621 1818 -445
rect 1852 -621 1864 -445
rect 1802 -633 1864 -621
rect 1920 -445 1982 -433
rect 1920 -621 1932 -445
rect 1966 -621 1982 -445
rect 1920 -633 1982 -621
rect 2012 -445 2074 -433
rect 2012 -621 2028 -445
rect 2062 -621 2074 -445
rect 2012 -633 2074 -621
rect 2130 -445 2192 -433
rect 2130 -621 2142 -445
rect 2176 -621 2192 -445
rect 2130 -633 2192 -621
rect 2222 -445 2284 -433
rect 2222 -621 2238 -445
rect 2272 -621 2284 -445
rect 2222 -633 2284 -621
rect 2340 -445 2402 -433
rect 2340 -621 2352 -445
rect 2386 -621 2402 -445
rect 2340 -633 2402 -621
rect 2432 -445 2494 -433
rect 2432 -621 2448 -445
rect 2482 -621 2494 -445
rect 2432 -633 2494 -621
rect 2550 -445 2612 -433
rect 2550 -621 2562 -445
rect 2596 -621 2612 -445
rect 2550 -633 2612 -621
rect 2642 -445 2704 -433
rect 2642 -621 2658 -445
rect 2692 -621 2704 -445
rect 2642 -633 2704 -621
rect 2760 -445 2822 -433
rect 2760 -621 2772 -445
rect 2806 -621 2822 -445
rect 2760 -633 2822 -621
rect 2852 -445 2914 -433
rect 2852 -621 2868 -445
rect 2902 -621 2914 -445
rect 2852 -633 2914 -621
rect 2970 -445 3032 -433
rect 2970 -621 2982 -445
rect 3016 -621 3032 -445
rect 2970 -633 3032 -621
rect 3062 -445 3124 -433
rect 3062 -621 3078 -445
rect 3112 -621 3124 -445
rect 3062 -633 3124 -621
rect 3180 -445 3242 -433
rect 3180 -621 3192 -445
rect 3226 -621 3242 -445
rect 3180 -633 3242 -621
rect 3272 -445 3334 -433
rect 3272 -621 3288 -445
rect 3322 -621 3334 -445
rect 3272 -633 3334 -621
rect 3390 -445 3452 -433
rect 3390 -621 3402 -445
rect 3436 -621 3452 -445
rect 3390 -633 3452 -621
rect 3482 -445 3544 -433
rect 3482 -621 3498 -445
rect 3532 -621 3544 -445
rect 3482 -633 3544 -621
rect 3600 -445 3662 -433
rect 3600 -621 3612 -445
rect 3646 -621 3662 -445
rect 3600 -633 3662 -621
rect 3692 -445 3754 -433
rect 3692 -621 3708 -445
rect 3742 -621 3754 -445
rect 3692 -633 3754 -621
rect 3810 -445 3872 -433
rect 3810 -621 3822 -445
rect 3856 -621 3872 -445
rect 3810 -633 3872 -621
rect 3902 -445 3964 -433
rect 3902 -621 3918 -445
rect 3952 -621 3964 -445
rect 3902 -633 3964 -621
rect 4020 -445 4082 -433
rect 4020 -621 4032 -445
rect 4066 -621 4082 -445
rect 4020 -633 4082 -621
rect 4112 -445 4174 -433
rect 4112 -621 4128 -445
rect 4162 -621 4174 -445
rect 4112 -633 4174 -621
rect 4230 -445 4292 -433
rect 4230 -621 4242 -445
rect 4276 -621 4292 -445
rect 4230 -633 4292 -621
rect 4322 -445 4384 -433
rect 4322 -621 4338 -445
rect 4372 -621 4384 -445
rect 4322 -633 4384 -621
<< pdiffc >>
rect -4370 -88 -4336 88
rect -4274 -88 -4240 88
rect -4160 -88 -4126 88
rect -4064 -88 -4030 88
rect -3950 -88 -3916 88
rect -3854 -88 -3820 88
rect -3740 -88 -3706 88
rect -3644 -88 -3610 88
rect -3530 -88 -3496 88
rect -3434 -88 -3400 88
rect -3320 -88 -3286 88
rect -3224 -88 -3190 88
rect -3110 -88 -3076 88
rect -3014 -88 -2980 88
rect -2900 -88 -2866 88
rect -2804 -88 -2770 88
rect -2690 -88 -2656 88
rect -2594 -88 -2560 88
rect -2480 -88 -2446 88
rect -2384 -88 -2350 88
rect -2270 -88 -2236 88
rect -2174 -88 -2140 88
rect -2060 -88 -2026 88
rect -1964 -88 -1930 88
rect -1850 -88 -1816 88
rect -1754 -88 -1720 88
rect -1640 -88 -1606 88
rect -1544 -88 -1510 88
rect -1430 -88 -1396 88
rect -1334 -88 -1300 88
rect -1220 -88 -1186 88
rect -1124 -88 -1090 88
rect -1010 -88 -976 88
rect -914 -88 -880 88
rect -800 -88 -766 88
rect -704 -88 -670 88
rect -590 -88 -556 88
rect -494 -88 -460 88
rect -380 -88 -346 88
rect -284 -88 -250 88
rect -170 -88 -136 88
rect -74 -88 -40 88
rect 40 -88 74 88
rect 136 -88 170 88
rect 250 -88 284 88
rect 346 -88 380 88
rect 460 -88 494 88
rect 556 -88 590 88
rect 670 -88 704 88
rect 766 -88 800 88
rect 880 -88 914 88
rect 976 -88 1010 88
rect 1090 -88 1124 88
rect 1186 -88 1220 88
rect 1300 -88 1334 88
rect 1396 -88 1430 88
rect 1510 -88 1544 88
rect 1606 -88 1640 88
rect 1720 -88 1754 88
rect 1816 -88 1850 88
rect 1930 -88 1964 88
rect 2026 -88 2060 88
rect 2140 -88 2174 88
rect 2236 -88 2270 88
rect 2350 -88 2384 88
rect 2446 -88 2480 88
rect 2560 -88 2594 88
rect 2656 -88 2690 88
rect 2770 -88 2804 88
rect 2866 -88 2900 88
rect 2980 -88 3014 88
rect 3076 -88 3110 88
rect 3190 -88 3224 88
rect 3286 -88 3320 88
rect 3400 -88 3434 88
rect 3496 -88 3530 88
rect 3610 -88 3644 88
rect 3706 -88 3740 88
rect 3820 -88 3854 88
rect 3916 -88 3950 88
rect 4030 -88 4064 88
rect 4126 -88 4160 88
rect 4240 -88 4274 88
rect 4336 -88 4370 88
rect -4368 -621 -4334 -445
rect -4272 -621 -4238 -445
rect -4158 -621 -4124 -445
rect -4062 -621 -4028 -445
rect -3948 -621 -3914 -445
rect -3852 -621 -3818 -445
rect -3738 -621 -3704 -445
rect -3642 -621 -3608 -445
rect -3528 -621 -3494 -445
rect -3432 -621 -3398 -445
rect -3318 -621 -3284 -445
rect -3222 -621 -3188 -445
rect -3108 -621 -3074 -445
rect -3012 -621 -2978 -445
rect -2898 -621 -2864 -445
rect -2802 -621 -2768 -445
rect -2688 -621 -2654 -445
rect -2592 -621 -2558 -445
rect -2478 -621 -2444 -445
rect -2382 -621 -2348 -445
rect -2268 -621 -2234 -445
rect -2172 -621 -2138 -445
rect -2058 -621 -2024 -445
rect -1962 -621 -1928 -445
rect -1848 -621 -1814 -445
rect -1752 -621 -1718 -445
rect -1638 -621 -1604 -445
rect -1542 -621 -1508 -445
rect -1428 -621 -1394 -445
rect -1332 -621 -1298 -445
rect -1218 -621 -1184 -445
rect -1122 -621 -1088 -445
rect -1008 -621 -974 -445
rect -912 -621 -878 -445
rect -798 -621 -764 -445
rect -702 -621 -668 -445
rect -588 -621 -554 -445
rect -492 -621 -458 -445
rect -378 -621 -344 -445
rect -282 -621 -248 -445
rect -168 -621 -134 -445
rect -72 -621 -38 -445
rect 42 -621 76 -445
rect 138 -621 172 -445
rect 252 -621 286 -445
rect 348 -621 382 -445
rect 462 -621 496 -445
rect 558 -621 592 -445
rect 672 -621 706 -445
rect 768 -621 802 -445
rect 882 -621 916 -445
rect 978 -621 1012 -445
rect 1092 -621 1126 -445
rect 1188 -621 1222 -445
rect 1302 -621 1336 -445
rect 1398 -621 1432 -445
rect 1512 -621 1546 -445
rect 1608 -621 1642 -445
rect 1722 -621 1756 -445
rect 1818 -621 1852 -445
rect 1932 -621 1966 -445
rect 2028 -621 2062 -445
rect 2142 -621 2176 -445
rect 2238 -621 2272 -445
rect 2352 -621 2386 -445
rect 2448 -621 2482 -445
rect 2562 -621 2596 -445
rect 2658 -621 2692 -445
rect 2772 -621 2806 -445
rect 2868 -621 2902 -445
rect 2982 -621 3016 -445
rect 3078 -621 3112 -445
rect 3192 -621 3226 -445
rect 3288 -621 3322 -445
rect 3402 -621 3436 -445
rect 3498 -621 3532 -445
rect 3612 -621 3646 -445
rect 3708 -621 3742 -445
rect 3822 -621 3856 -445
rect 3918 -621 3952 -445
rect 4032 -621 4066 -445
rect 4128 -621 4162 -445
rect 4242 -621 4276 -445
rect 4338 -621 4372 -445
<< nsubdiff >>
rect -4484 249 -4388 283
rect 4388 249 4484 283
rect -4484 187 -4450 249
rect 4450 187 4484 249
rect -4484 -345 -4450 -187
rect 4450 -345 4484 -187
rect -4484 -782 -4450 -720
rect 4450 -782 4484 -720
rect -4484 -816 -4388 -782
rect 4388 -816 4484 -782
<< nsubdiffcont >>
rect -4388 249 4388 283
rect -4484 -187 -4450 187
rect 4450 -187 4484 187
rect -4484 -720 -4450 -345
rect 4450 -720 4484 -345
rect -4388 -816 4388 -782
<< poly >>
rect -4128 181 -4062 197
rect -4128 147 -4112 181
rect -4078 147 -4062 181
rect -4128 131 -4062 147
rect -3708 181 -3642 197
rect -3708 147 -3692 181
rect -3658 147 -3642 181
rect -3708 131 -3642 147
rect -3288 181 -3222 197
rect -3288 147 -3272 181
rect -3238 147 -3222 181
rect -3288 131 -3222 147
rect -2868 181 -2802 197
rect -2868 147 -2852 181
rect -2818 147 -2802 181
rect -2868 131 -2802 147
rect -2448 181 -2382 197
rect -2448 147 -2432 181
rect -2398 147 -2382 181
rect -2448 131 -2382 147
rect -2028 181 -1962 197
rect -2028 147 -2012 181
rect -1978 147 -1962 181
rect -2028 131 -1962 147
rect -1608 181 -1542 197
rect -1608 147 -1592 181
rect -1558 147 -1542 181
rect -1608 131 -1542 147
rect -1188 181 -1122 197
rect -1188 147 -1172 181
rect -1138 147 -1122 181
rect -1188 131 -1122 147
rect -768 181 -702 197
rect -768 147 -752 181
rect -718 147 -702 181
rect -768 131 -702 147
rect -348 181 -282 197
rect -348 147 -332 181
rect -298 147 -282 181
rect -348 131 -282 147
rect 72 181 138 197
rect 72 147 88 181
rect 122 147 138 181
rect 72 131 138 147
rect 492 181 558 197
rect 492 147 508 181
rect 542 147 558 181
rect 492 131 558 147
rect 912 181 978 197
rect 912 147 928 181
rect 962 147 978 181
rect 912 131 978 147
rect 1332 181 1398 197
rect 1332 147 1348 181
rect 1382 147 1398 181
rect 1332 131 1398 147
rect 1752 181 1818 197
rect 1752 147 1768 181
rect 1802 147 1818 181
rect 1752 131 1818 147
rect 2172 181 2238 197
rect 2172 147 2188 181
rect 2222 147 2238 181
rect 2172 131 2238 147
rect 2592 181 2658 197
rect 2592 147 2608 181
rect 2642 147 2658 181
rect 2592 131 2658 147
rect 3012 181 3078 197
rect 3012 147 3028 181
rect 3062 147 3078 181
rect 3012 131 3078 147
rect 3432 181 3498 197
rect 3432 147 3448 181
rect 3482 147 3498 181
rect 3432 131 3498 147
rect 3852 181 3918 197
rect 3852 147 3868 181
rect 3902 147 3918 181
rect 3852 131 3918 147
rect 4272 181 4338 197
rect 4272 147 4288 181
rect 4322 147 4338 181
rect 4272 131 4338 147
rect -4320 100 -4290 127
rect -4110 100 -4080 131
rect -3900 100 -3870 127
rect -3690 100 -3660 131
rect -3480 100 -3450 127
rect -3270 100 -3240 131
rect -3060 100 -3030 127
rect -2850 100 -2820 131
rect -2640 100 -2610 127
rect -2430 100 -2400 131
rect -2220 100 -2190 127
rect -2010 100 -1980 131
rect -1800 100 -1770 127
rect -1590 100 -1560 131
rect -1380 100 -1350 127
rect -1170 100 -1140 131
rect -960 100 -930 127
rect -750 100 -720 131
rect -540 100 -510 127
rect -330 100 -300 131
rect -120 100 -90 127
rect 90 100 120 131
rect 300 100 330 127
rect 510 100 540 131
rect 720 100 750 127
rect 930 100 960 131
rect 1140 100 1170 127
rect 1350 100 1380 131
rect 1560 100 1590 127
rect 1770 100 1800 131
rect 1980 100 2010 127
rect 2190 100 2220 131
rect 2400 100 2430 127
rect 2610 100 2640 131
rect 2820 100 2850 127
rect 3030 100 3060 131
rect 3240 100 3270 127
rect 3450 100 3480 131
rect 3660 100 3690 127
rect 3870 100 3900 131
rect 4080 100 4110 127
rect 4290 100 4320 131
rect -4320 -131 -4290 -100
rect -4110 -127 -4080 -100
rect -3900 -131 -3870 -100
rect -3690 -127 -3660 -100
rect -3480 -131 -3450 -100
rect -3270 -127 -3240 -100
rect -3060 -131 -3030 -100
rect -2850 -127 -2820 -100
rect -2640 -131 -2610 -100
rect -2430 -127 -2400 -100
rect -2220 -131 -2190 -100
rect -2010 -127 -1980 -100
rect -1800 -131 -1770 -100
rect -1590 -127 -1560 -100
rect -1380 -131 -1350 -100
rect -1170 -127 -1140 -100
rect -960 -131 -930 -100
rect -750 -127 -720 -100
rect -540 -131 -510 -100
rect -330 -127 -300 -100
rect -120 -131 -90 -100
rect 90 -127 120 -100
rect 300 -131 330 -100
rect 510 -127 540 -100
rect 720 -131 750 -100
rect 930 -127 960 -100
rect 1140 -131 1170 -100
rect 1350 -127 1380 -100
rect 1560 -131 1590 -100
rect 1770 -127 1800 -100
rect 1980 -131 2010 -100
rect 2190 -127 2220 -100
rect 2400 -131 2430 -100
rect 2610 -127 2640 -100
rect 2820 -131 2850 -100
rect 3030 -127 3060 -100
rect 3240 -131 3270 -100
rect 3450 -127 3480 -100
rect 3660 -131 3690 -100
rect 3870 -127 3900 -100
rect 4080 -131 4110 -100
rect 4290 -127 4320 -100
rect -4338 -147 -4272 -131
rect -4338 -181 -4322 -147
rect -4288 -181 -4272 -147
rect -4338 -197 -4272 -181
rect -3918 -147 -3852 -131
rect -3918 -181 -3902 -147
rect -3868 -181 -3852 -147
rect -3918 -197 -3852 -181
rect -3498 -147 -3432 -131
rect -3498 -181 -3482 -147
rect -3448 -181 -3432 -147
rect -3498 -197 -3432 -181
rect -3078 -147 -3012 -131
rect -3078 -181 -3062 -147
rect -3028 -181 -3012 -147
rect -3078 -197 -3012 -181
rect -2658 -147 -2592 -131
rect -2658 -181 -2642 -147
rect -2608 -181 -2592 -147
rect -2658 -197 -2592 -181
rect -2238 -147 -2172 -131
rect -2238 -181 -2222 -147
rect -2188 -181 -2172 -147
rect -2238 -197 -2172 -181
rect -1818 -147 -1752 -131
rect -1818 -181 -1802 -147
rect -1768 -181 -1752 -147
rect -1818 -197 -1752 -181
rect -1398 -147 -1332 -131
rect -1398 -181 -1382 -147
rect -1348 -181 -1332 -147
rect -1398 -197 -1332 -181
rect -978 -147 -912 -131
rect -978 -181 -962 -147
rect -928 -181 -912 -147
rect -978 -197 -912 -181
rect -558 -147 -492 -131
rect -558 -181 -542 -147
rect -508 -181 -492 -147
rect -558 -197 -492 -181
rect -138 -147 -72 -131
rect -138 -181 -122 -147
rect -88 -181 -72 -147
rect -138 -197 -72 -181
rect 282 -147 348 -131
rect 282 -181 298 -147
rect 332 -181 348 -147
rect 282 -197 348 -181
rect 702 -147 768 -131
rect 702 -181 718 -147
rect 752 -181 768 -147
rect 702 -197 768 -181
rect 1122 -147 1188 -131
rect 1122 -181 1138 -147
rect 1172 -181 1188 -147
rect 1122 -197 1188 -181
rect 1542 -147 1608 -131
rect 1542 -181 1558 -147
rect 1592 -181 1608 -147
rect 1542 -197 1608 -181
rect 1962 -147 2028 -131
rect 1962 -181 1978 -147
rect 2012 -181 2028 -147
rect 1962 -197 2028 -181
rect 2382 -147 2448 -131
rect 2382 -181 2398 -147
rect 2432 -181 2448 -147
rect 2382 -197 2448 -181
rect 2802 -147 2868 -131
rect 2802 -181 2818 -147
rect 2852 -181 2868 -147
rect 2802 -197 2868 -181
rect 3222 -147 3288 -131
rect 3222 -181 3238 -147
rect 3272 -181 3288 -147
rect 3222 -197 3288 -181
rect 3642 -147 3708 -131
rect 3642 -181 3658 -147
rect 3692 -181 3708 -147
rect 3642 -197 3708 -181
rect 4062 -147 4128 -131
rect 4062 -181 4078 -147
rect 4112 -181 4128 -147
rect 4062 -197 4128 -181
rect -4126 -351 -4060 -335
rect -4126 -385 -4110 -351
rect -4076 -385 -4060 -351
rect -4126 -401 -4060 -385
rect -3706 -351 -3640 -335
rect -3706 -385 -3690 -351
rect -3656 -385 -3640 -351
rect -3706 -401 -3640 -385
rect -3286 -351 -3220 -335
rect -3286 -385 -3270 -351
rect -3236 -385 -3220 -351
rect -3286 -401 -3220 -385
rect -2866 -351 -2800 -335
rect -2866 -385 -2850 -351
rect -2816 -385 -2800 -351
rect -2866 -401 -2800 -385
rect -2446 -351 -2380 -335
rect -2446 -385 -2430 -351
rect -2396 -385 -2380 -351
rect -2446 -401 -2380 -385
rect -2026 -351 -1960 -335
rect -2026 -385 -2010 -351
rect -1976 -385 -1960 -351
rect -2026 -401 -1960 -385
rect -1606 -351 -1540 -335
rect -1606 -385 -1590 -351
rect -1556 -385 -1540 -351
rect -1606 -401 -1540 -385
rect -1186 -351 -1120 -335
rect -1186 -385 -1170 -351
rect -1136 -385 -1120 -351
rect -1186 -401 -1120 -385
rect -766 -351 -700 -335
rect -766 -385 -750 -351
rect -716 -385 -700 -351
rect -766 -401 -700 -385
rect -346 -351 -280 -335
rect -346 -385 -330 -351
rect -296 -385 -280 -351
rect -346 -401 -280 -385
rect 74 -351 140 -335
rect 74 -385 90 -351
rect 124 -385 140 -351
rect 74 -401 140 -385
rect 494 -351 560 -335
rect 494 -385 510 -351
rect 544 -385 560 -351
rect 494 -401 560 -385
rect 914 -351 980 -335
rect 914 -385 930 -351
rect 964 -385 980 -351
rect 914 -401 980 -385
rect 1334 -351 1400 -335
rect 1334 -385 1350 -351
rect 1384 -385 1400 -351
rect 1334 -401 1400 -385
rect 1754 -351 1820 -335
rect 1754 -385 1770 -351
rect 1804 -385 1820 -351
rect 1754 -401 1820 -385
rect 2174 -351 2240 -335
rect 2174 -385 2190 -351
rect 2224 -385 2240 -351
rect 2174 -401 2240 -385
rect 2594 -351 2660 -335
rect 2594 -385 2610 -351
rect 2644 -385 2660 -351
rect 2594 -401 2660 -385
rect 3014 -351 3080 -335
rect 3014 -385 3030 -351
rect 3064 -385 3080 -351
rect 3014 -401 3080 -385
rect 3434 -351 3500 -335
rect 3434 -385 3450 -351
rect 3484 -385 3500 -351
rect 3434 -401 3500 -385
rect 3854 -351 3920 -335
rect 3854 -385 3870 -351
rect 3904 -385 3920 -351
rect 3854 -401 3920 -385
rect 4274 -351 4340 -335
rect 4274 -385 4290 -351
rect 4324 -385 4340 -351
rect 4274 -401 4340 -385
rect -4318 -433 -4288 -407
rect -4108 -433 -4078 -401
rect -3898 -433 -3868 -407
rect -3688 -433 -3658 -401
rect -3478 -433 -3448 -407
rect -3268 -433 -3238 -401
rect -3058 -433 -3028 -407
rect -2848 -433 -2818 -401
rect -2638 -433 -2608 -407
rect -2428 -433 -2398 -401
rect -2218 -433 -2188 -407
rect -2008 -433 -1978 -401
rect -1798 -433 -1768 -407
rect -1588 -433 -1558 -401
rect -1378 -433 -1348 -407
rect -1168 -433 -1138 -401
rect -958 -433 -928 -407
rect -748 -433 -718 -401
rect -538 -433 -508 -407
rect -328 -433 -298 -401
rect -118 -433 -88 -407
rect 92 -433 122 -401
rect 302 -433 332 -407
rect 512 -433 542 -401
rect 722 -433 752 -407
rect 932 -433 962 -401
rect 1142 -433 1172 -407
rect 1352 -433 1382 -401
rect 1562 -433 1592 -407
rect 1772 -433 1802 -401
rect 1982 -433 2012 -407
rect 2192 -433 2222 -401
rect 2402 -433 2432 -407
rect 2612 -433 2642 -401
rect 2822 -433 2852 -407
rect 3032 -433 3062 -401
rect 3242 -433 3272 -407
rect 3452 -433 3482 -401
rect 3662 -433 3692 -407
rect 3872 -433 3902 -401
rect 4082 -433 4112 -407
rect 4292 -433 4322 -401
rect -4318 -664 -4288 -633
rect -4108 -660 -4078 -633
rect -3898 -664 -3868 -633
rect -3688 -660 -3658 -633
rect -3478 -664 -3448 -633
rect -3268 -660 -3238 -633
rect -3058 -664 -3028 -633
rect -2848 -660 -2818 -633
rect -2638 -664 -2608 -633
rect -2428 -660 -2398 -633
rect -2218 -664 -2188 -633
rect -2008 -660 -1978 -633
rect -1798 -664 -1768 -633
rect -1588 -660 -1558 -633
rect -1378 -664 -1348 -633
rect -1168 -660 -1138 -633
rect -958 -664 -928 -633
rect -748 -660 -718 -633
rect -538 -664 -508 -633
rect -328 -660 -298 -633
rect -118 -664 -88 -633
rect 92 -660 122 -633
rect 302 -664 332 -633
rect 512 -660 542 -633
rect 722 -664 752 -633
rect 932 -660 962 -633
rect 1142 -664 1172 -633
rect 1352 -660 1382 -633
rect 1562 -664 1592 -633
rect 1772 -660 1802 -633
rect 1982 -664 2012 -633
rect 2192 -660 2222 -633
rect 2402 -664 2432 -633
rect 2612 -660 2642 -633
rect 2822 -664 2852 -633
rect 3032 -660 3062 -633
rect 3242 -664 3272 -633
rect 3452 -660 3482 -633
rect 3662 -664 3692 -633
rect 3872 -660 3902 -633
rect 4082 -664 4112 -633
rect 4292 -660 4322 -633
rect -4336 -680 -4270 -664
rect -4336 -714 -4320 -680
rect -4286 -714 -4270 -680
rect -4336 -730 -4270 -714
rect -3916 -680 -3850 -664
rect -3916 -714 -3900 -680
rect -3866 -714 -3850 -680
rect -3916 -730 -3850 -714
rect -3496 -680 -3430 -664
rect -3496 -714 -3480 -680
rect -3446 -714 -3430 -680
rect -3496 -730 -3430 -714
rect -3076 -680 -3010 -664
rect -3076 -714 -3060 -680
rect -3026 -714 -3010 -680
rect -3076 -730 -3010 -714
rect -2656 -680 -2590 -664
rect -2656 -714 -2640 -680
rect -2606 -714 -2590 -680
rect -2656 -730 -2590 -714
rect -2236 -680 -2170 -664
rect -2236 -714 -2220 -680
rect -2186 -714 -2170 -680
rect -2236 -730 -2170 -714
rect -1816 -680 -1750 -664
rect -1816 -714 -1800 -680
rect -1766 -714 -1750 -680
rect -1816 -730 -1750 -714
rect -1396 -680 -1330 -664
rect -1396 -714 -1380 -680
rect -1346 -714 -1330 -680
rect -1396 -730 -1330 -714
rect -976 -680 -910 -664
rect -976 -714 -960 -680
rect -926 -714 -910 -680
rect -976 -730 -910 -714
rect -556 -680 -490 -664
rect -556 -714 -540 -680
rect -506 -714 -490 -680
rect -556 -730 -490 -714
rect -136 -680 -70 -664
rect -136 -714 -120 -680
rect -86 -714 -70 -680
rect -136 -730 -70 -714
rect 284 -680 350 -664
rect 284 -714 300 -680
rect 334 -714 350 -680
rect 284 -730 350 -714
rect 704 -680 770 -664
rect 704 -714 720 -680
rect 754 -714 770 -680
rect 704 -730 770 -714
rect 1124 -680 1190 -664
rect 1124 -714 1140 -680
rect 1174 -714 1190 -680
rect 1124 -730 1190 -714
rect 1544 -680 1610 -664
rect 1544 -714 1560 -680
rect 1594 -714 1610 -680
rect 1544 -730 1610 -714
rect 1964 -680 2030 -664
rect 1964 -714 1980 -680
rect 2014 -714 2030 -680
rect 1964 -730 2030 -714
rect 2384 -680 2450 -664
rect 2384 -714 2400 -680
rect 2434 -714 2450 -680
rect 2384 -730 2450 -714
rect 2804 -680 2870 -664
rect 2804 -714 2820 -680
rect 2854 -714 2870 -680
rect 2804 -730 2870 -714
rect 3224 -680 3290 -664
rect 3224 -714 3240 -680
rect 3274 -714 3290 -680
rect 3224 -730 3290 -714
rect 3644 -680 3710 -664
rect 3644 -714 3660 -680
rect 3694 -714 3710 -680
rect 3644 -730 3710 -714
rect 4064 -680 4130 -664
rect 4064 -714 4080 -680
rect 4114 -714 4130 -680
rect 4064 -730 4130 -714
<< polycont >>
rect -4112 147 -4078 181
rect -3692 147 -3658 181
rect -3272 147 -3238 181
rect -2852 147 -2818 181
rect -2432 147 -2398 181
rect -2012 147 -1978 181
rect -1592 147 -1558 181
rect -1172 147 -1138 181
rect -752 147 -718 181
rect -332 147 -298 181
rect 88 147 122 181
rect 508 147 542 181
rect 928 147 962 181
rect 1348 147 1382 181
rect 1768 147 1802 181
rect 2188 147 2222 181
rect 2608 147 2642 181
rect 3028 147 3062 181
rect 3448 147 3482 181
rect 3868 147 3902 181
rect 4288 147 4322 181
rect -4322 -181 -4288 -147
rect -3902 -181 -3868 -147
rect -3482 -181 -3448 -147
rect -3062 -181 -3028 -147
rect -2642 -181 -2608 -147
rect -2222 -181 -2188 -147
rect -1802 -181 -1768 -147
rect -1382 -181 -1348 -147
rect -962 -181 -928 -147
rect -542 -181 -508 -147
rect -122 -181 -88 -147
rect 298 -181 332 -147
rect 718 -181 752 -147
rect 1138 -181 1172 -147
rect 1558 -181 1592 -147
rect 1978 -181 2012 -147
rect 2398 -181 2432 -147
rect 2818 -181 2852 -147
rect 3238 -181 3272 -147
rect 3658 -181 3692 -147
rect 4078 -181 4112 -147
rect -4110 -385 -4076 -351
rect -3690 -385 -3656 -351
rect -3270 -385 -3236 -351
rect -2850 -385 -2816 -351
rect -2430 -385 -2396 -351
rect -2010 -385 -1976 -351
rect -1590 -385 -1556 -351
rect -1170 -385 -1136 -351
rect -750 -385 -716 -351
rect -330 -385 -296 -351
rect 90 -385 124 -351
rect 510 -385 544 -351
rect 930 -385 964 -351
rect 1350 -385 1384 -351
rect 1770 -385 1804 -351
rect 2190 -385 2224 -351
rect 2610 -385 2644 -351
rect 3030 -385 3064 -351
rect 3450 -385 3484 -351
rect 3870 -385 3904 -351
rect 4290 -385 4324 -351
rect -4320 -714 -4286 -680
rect -3900 -714 -3866 -680
rect -3480 -714 -3446 -680
rect -3060 -714 -3026 -680
rect -2640 -714 -2606 -680
rect -2220 -714 -2186 -680
rect -1800 -714 -1766 -680
rect -1380 -714 -1346 -680
rect -960 -714 -926 -680
rect -540 -714 -506 -680
rect -120 -714 -86 -680
rect 300 -714 334 -680
rect 720 -714 754 -680
rect 1140 -714 1174 -680
rect 1560 -714 1594 -680
rect 1980 -714 2014 -680
rect 2400 -714 2434 -680
rect 2820 -714 2854 -680
rect 3240 -714 3274 -680
rect 3660 -714 3694 -680
rect 4080 -714 4114 -680
<< locali >>
rect -4484 249 -4388 283
rect 4388 249 4484 283
rect -4484 187 -4450 249
rect 4450 187 4484 249
rect -4128 147 -4112 181
rect -4078 147 -4062 181
rect -3708 147 -3692 181
rect -3658 147 -3642 181
rect -3288 147 -3272 181
rect -3238 147 -3222 181
rect -2868 147 -2852 181
rect -2818 147 -2802 181
rect -2448 147 -2432 181
rect -2398 147 -2382 181
rect -2028 147 -2012 181
rect -1978 147 -1962 181
rect -1608 147 -1592 181
rect -1558 147 -1542 181
rect -1188 147 -1172 181
rect -1138 147 -1122 181
rect -768 147 -752 181
rect -718 147 -702 181
rect -348 147 -332 181
rect -298 147 -282 181
rect 72 147 88 181
rect 122 147 138 181
rect 492 147 508 181
rect 542 147 558 181
rect 912 147 928 181
rect 962 147 978 181
rect 1332 147 1348 181
rect 1382 147 1398 181
rect 1752 147 1768 181
rect 1802 147 1818 181
rect 2172 147 2188 181
rect 2222 147 2238 181
rect 2592 147 2608 181
rect 2642 147 2658 181
rect 3012 147 3028 181
rect 3062 147 3078 181
rect 3432 147 3448 181
rect 3482 147 3498 181
rect 3852 147 3868 181
rect 3902 147 3918 181
rect 4240 147 4288 181
rect 4322 147 4450 181
rect -4370 88 -4336 104
rect -4370 -147 -4336 -88
rect -4274 88 -4240 104
rect -4274 -147 -4240 -88
rect -4160 88 -4126 104
rect -4160 -104 -4126 -88
rect -4064 88 -4030 104
rect -4064 -104 -4030 -88
rect -3950 88 -3916 104
rect -3950 -104 -3916 -88
rect -3854 88 -3820 104
rect -3854 -104 -3820 -88
rect -3740 88 -3706 104
rect -3740 -104 -3706 -88
rect -3644 88 -3610 104
rect -3644 -104 -3610 -88
rect -3530 88 -3496 104
rect -3530 -104 -3496 -88
rect -3434 88 -3400 104
rect -3434 -104 -3400 -88
rect -3320 88 -3286 104
rect -3320 -104 -3286 -88
rect -3224 88 -3190 104
rect -3224 -104 -3190 -88
rect -3110 88 -3076 104
rect -3110 -104 -3076 -88
rect -3014 88 -2980 104
rect -3014 -104 -2980 -88
rect -2900 88 -2866 104
rect -2900 -104 -2866 -88
rect -2804 88 -2770 104
rect -2804 -104 -2770 -88
rect -2690 88 -2656 104
rect -2690 -104 -2656 -88
rect -2594 88 -2560 104
rect -2594 -104 -2560 -88
rect -2480 88 -2446 104
rect -2480 -104 -2446 -88
rect -2384 88 -2350 104
rect -2384 -104 -2350 -88
rect -2270 88 -2236 104
rect -2270 -104 -2236 -88
rect -2174 88 -2140 104
rect -2174 -104 -2140 -88
rect -2060 88 -2026 104
rect -2060 -104 -2026 -88
rect -1964 88 -1930 104
rect -1964 -104 -1930 -88
rect -1850 88 -1816 104
rect -1850 -104 -1816 -88
rect -1754 88 -1720 104
rect -1754 -104 -1720 -88
rect -1640 88 -1606 104
rect -1640 -104 -1606 -88
rect -1544 88 -1510 104
rect -1544 -104 -1510 -88
rect -1430 88 -1396 104
rect -1430 -104 -1396 -88
rect -1334 88 -1300 104
rect -1334 -104 -1300 -88
rect -1220 88 -1186 104
rect -1220 -104 -1186 -88
rect -1124 88 -1090 104
rect -1124 -104 -1090 -88
rect -1010 88 -976 104
rect -1010 -104 -976 -88
rect -914 88 -880 104
rect -914 -104 -880 -88
rect -800 88 -766 104
rect -800 -104 -766 -88
rect -704 88 -670 104
rect -704 -104 -670 -88
rect -590 88 -556 104
rect -590 -104 -556 -88
rect -494 88 -460 104
rect -494 -104 -460 -88
rect -380 88 -346 104
rect -380 -104 -346 -88
rect -284 88 -250 104
rect -284 -104 -250 -88
rect -170 88 -136 104
rect -170 -104 -136 -88
rect -74 88 -40 104
rect -74 -104 -40 -88
rect 40 88 74 104
rect 40 -104 74 -88
rect 136 88 170 104
rect 136 -104 170 -88
rect 250 88 284 104
rect 250 -104 284 -88
rect 346 88 380 104
rect 346 -104 380 -88
rect 460 88 494 104
rect 460 -104 494 -88
rect 556 88 590 104
rect 556 -104 590 -88
rect 670 88 704 104
rect 670 -104 704 -88
rect 766 88 800 104
rect 766 -104 800 -88
rect 880 88 914 104
rect 880 -104 914 -88
rect 976 88 1010 104
rect 976 -104 1010 -88
rect 1090 88 1124 104
rect 1090 -104 1124 -88
rect 1186 88 1220 104
rect 1186 -104 1220 -88
rect 1300 88 1334 104
rect 1300 -104 1334 -88
rect 1396 88 1430 104
rect 1396 -104 1430 -88
rect 1510 88 1544 104
rect 1510 -104 1544 -88
rect 1606 88 1640 104
rect 1606 -104 1640 -88
rect 1720 88 1754 104
rect 1720 -104 1754 -88
rect 1816 88 1850 104
rect 1816 -104 1850 -88
rect 1930 88 1964 104
rect 1930 -104 1964 -88
rect 2026 88 2060 104
rect 2026 -104 2060 -88
rect 2140 88 2174 104
rect 2140 -104 2174 -88
rect 2236 88 2270 104
rect 2236 -104 2270 -88
rect 2350 88 2384 104
rect 2350 -104 2384 -88
rect 2446 88 2480 104
rect 2446 -104 2480 -88
rect 2560 88 2594 104
rect 2560 -104 2594 -88
rect 2656 88 2690 104
rect 2656 -104 2690 -88
rect 2770 88 2804 104
rect 2770 -104 2804 -88
rect 2866 88 2900 104
rect 2866 -104 2900 -88
rect 2980 88 3014 104
rect 2980 -104 3014 -88
rect 3076 88 3110 104
rect 3076 -104 3110 -88
rect 3190 88 3224 104
rect 3190 -104 3224 -88
rect 3286 88 3320 104
rect 3286 -104 3320 -88
rect 3400 88 3434 104
rect 3400 -104 3434 -88
rect 3496 88 3530 104
rect 3496 -104 3530 -88
rect 3610 88 3644 104
rect 3610 -104 3644 -88
rect 3706 88 3740 104
rect 3706 -104 3740 -88
rect 3820 88 3854 104
rect 3820 -104 3854 -88
rect 3916 88 3950 104
rect 3916 -104 3950 -88
rect 4030 88 4064 104
rect 4030 -104 4064 -88
rect 4126 88 4160 104
rect 4126 -104 4160 -88
rect 4240 88 4274 147
rect 4240 -104 4274 -88
rect 4336 88 4370 147
rect 4336 -104 4370 -88
rect -4450 -181 -4322 -147
rect -4288 -181 -4240 -147
rect -3918 -181 -3902 -147
rect -3868 -181 -3852 -147
rect -3498 -181 -3482 -147
rect -3448 -181 -3432 -147
rect -3078 -181 -3062 -147
rect -3028 -181 -3012 -147
rect -2658 -181 -2642 -147
rect -2608 -181 -2592 -147
rect -2238 -181 -2222 -147
rect -2188 -181 -2172 -147
rect -1818 -181 -1802 -147
rect -1768 -181 -1752 -147
rect -1398 -181 -1382 -147
rect -1348 -181 -1332 -147
rect -978 -181 -962 -147
rect -928 -181 -912 -147
rect -558 -181 -542 -147
rect -508 -181 -492 -147
rect -138 -181 -122 -147
rect -88 -181 -72 -147
rect 282 -181 298 -147
rect 332 -181 348 -147
rect 702 -181 718 -147
rect 752 -181 768 -147
rect 1122 -181 1138 -147
rect 1172 -181 1188 -147
rect 1542 -181 1558 -147
rect 1592 -181 1608 -147
rect 1962 -181 1978 -147
rect 2012 -181 2028 -147
rect 2382 -181 2398 -147
rect 2432 -181 2448 -147
rect 2802 -181 2818 -147
rect 2852 -181 2868 -147
rect 3222 -181 3238 -147
rect 3272 -181 3288 -147
rect 3642 -181 3658 -147
rect 3692 -181 3708 -147
rect 4062 -181 4078 -147
rect 4112 -181 4128 -147
rect -4484 -345 -4450 -187
rect 4450 -345 4484 -187
rect -4126 -385 -4110 -351
rect -4076 -385 -4060 -351
rect -3706 -385 -3690 -351
rect -3656 -385 -3640 -351
rect -3286 -385 -3270 -351
rect -3236 -385 -3220 -351
rect -2866 -385 -2850 -351
rect -2816 -385 -2800 -351
rect -2446 -385 -2430 -351
rect -2396 -385 -2380 -351
rect -2026 -385 -2010 -351
rect -1976 -385 -1960 -351
rect -1606 -385 -1590 -351
rect -1556 -385 -1540 -351
rect -1186 -385 -1170 -351
rect -1136 -385 -1120 -351
rect -766 -385 -750 -351
rect -716 -385 -700 -351
rect -346 -385 -330 -351
rect -296 -385 -280 -351
rect 74 -385 90 -351
rect 124 -385 140 -351
rect 494 -385 510 -351
rect 544 -385 560 -351
rect 914 -385 930 -351
rect 964 -385 980 -351
rect 1334 -385 1350 -351
rect 1384 -385 1400 -351
rect 1754 -385 1770 -351
rect 1804 -385 1820 -351
rect 2174 -385 2190 -351
rect 2224 -385 2240 -351
rect 2594 -385 2610 -351
rect 2644 -385 2660 -351
rect 3014 -385 3030 -351
rect 3064 -385 3080 -351
rect 3434 -385 3450 -351
rect 3484 -385 3500 -351
rect 3854 -385 3870 -351
rect 3904 -385 3920 -351
rect 4242 -385 4290 -351
rect 4324 -385 4450 -351
rect -4368 -445 -4334 -429
rect -4368 -680 -4334 -621
rect -4272 -445 -4238 -429
rect -4272 -680 -4238 -621
rect -4158 -445 -4124 -429
rect -4158 -637 -4124 -621
rect -4062 -445 -4028 -429
rect -4062 -637 -4028 -621
rect -3948 -445 -3914 -429
rect -3948 -637 -3914 -621
rect -3852 -445 -3818 -429
rect -3852 -637 -3818 -621
rect -3738 -445 -3704 -429
rect -3738 -637 -3704 -621
rect -3642 -445 -3608 -429
rect -3642 -637 -3608 -621
rect -3528 -445 -3494 -429
rect -3528 -637 -3494 -621
rect -3432 -445 -3398 -429
rect -3432 -637 -3398 -621
rect -3318 -445 -3284 -429
rect -3318 -637 -3284 -621
rect -3222 -445 -3188 -429
rect -3222 -637 -3188 -621
rect -3108 -445 -3074 -429
rect -3108 -637 -3074 -621
rect -3012 -445 -2978 -429
rect -3012 -637 -2978 -621
rect -2898 -445 -2864 -429
rect -2898 -637 -2864 -621
rect -2802 -445 -2768 -429
rect -2802 -637 -2768 -621
rect -2688 -445 -2654 -429
rect -2688 -637 -2654 -621
rect -2592 -445 -2558 -429
rect -2592 -637 -2558 -621
rect -2478 -445 -2444 -429
rect -2478 -637 -2444 -621
rect -2382 -445 -2348 -429
rect -2382 -637 -2348 -621
rect -2268 -445 -2234 -429
rect -2268 -637 -2234 -621
rect -2172 -445 -2138 -429
rect -2172 -637 -2138 -621
rect -2058 -445 -2024 -429
rect -2058 -637 -2024 -621
rect -1962 -445 -1928 -429
rect -1962 -637 -1928 -621
rect -1848 -445 -1814 -429
rect -1848 -637 -1814 -621
rect -1752 -445 -1718 -429
rect -1752 -637 -1718 -621
rect -1638 -445 -1604 -429
rect -1638 -637 -1604 -621
rect -1542 -445 -1508 -429
rect -1542 -637 -1508 -621
rect -1428 -445 -1394 -429
rect -1428 -637 -1394 -621
rect -1332 -445 -1298 -429
rect -1332 -637 -1298 -621
rect -1218 -445 -1184 -429
rect -1218 -637 -1184 -621
rect -1122 -445 -1088 -429
rect -1122 -637 -1088 -621
rect -1008 -445 -974 -429
rect -1008 -637 -974 -621
rect -912 -445 -878 -429
rect -912 -637 -878 -621
rect -798 -445 -764 -429
rect -798 -637 -764 -621
rect -702 -445 -668 -429
rect -702 -637 -668 -621
rect -588 -445 -554 -429
rect -588 -637 -554 -621
rect -492 -445 -458 -429
rect -492 -637 -458 -621
rect -378 -445 -344 -429
rect -378 -637 -344 -621
rect -282 -445 -248 -429
rect -282 -637 -248 -621
rect -168 -445 -134 -429
rect -168 -637 -134 -621
rect -72 -445 -38 -429
rect -72 -637 -38 -621
rect 42 -445 76 -429
rect 42 -637 76 -621
rect 138 -445 172 -429
rect 138 -637 172 -621
rect 252 -445 286 -429
rect 252 -637 286 -621
rect 348 -445 382 -429
rect 348 -637 382 -621
rect 462 -445 496 -429
rect 462 -637 496 -621
rect 558 -445 592 -429
rect 558 -637 592 -621
rect 672 -445 706 -429
rect 672 -637 706 -621
rect 768 -445 802 -429
rect 768 -637 802 -621
rect 882 -445 916 -429
rect 882 -637 916 -621
rect 978 -445 1012 -429
rect 978 -637 1012 -621
rect 1092 -445 1126 -429
rect 1092 -637 1126 -621
rect 1188 -445 1222 -429
rect 1188 -637 1222 -621
rect 1302 -445 1336 -429
rect 1302 -637 1336 -621
rect 1398 -445 1432 -429
rect 1398 -637 1432 -621
rect 1512 -445 1546 -429
rect 1512 -637 1546 -621
rect 1608 -445 1642 -429
rect 1608 -637 1642 -621
rect 1722 -445 1756 -429
rect 1722 -637 1756 -621
rect 1818 -445 1852 -429
rect 1818 -637 1852 -621
rect 1932 -445 1966 -429
rect 1932 -637 1966 -621
rect 2028 -445 2062 -429
rect 2028 -637 2062 -621
rect 2142 -445 2176 -429
rect 2142 -637 2176 -621
rect 2238 -445 2272 -429
rect 2238 -637 2272 -621
rect 2352 -445 2386 -429
rect 2352 -637 2386 -621
rect 2448 -445 2482 -429
rect 2448 -637 2482 -621
rect 2562 -445 2596 -429
rect 2562 -637 2596 -621
rect 2658 -445 2692 -429
rect 2658 -637 2692 -621
rect 2772 -445 2806 -429
rect 2772 -637 2806 -621
rect 2868 -445 2902 -429
rect 2868 -637 2902 -621
rect 2982 -445 3016 -429
rect 2982 -637 3016 -621
rect 3078 -445 3112 -429
rect 3078 -637 3112 -621
rect 3192 -445 3226 -429
rect 3192 -637 3226 -621
rect 3288 -445 3322 -429
rect 3288 -637 3322 -621
rect 3402 -445 3436 -429
rect 3402 -637 3436 -621
rect 3498 -445 3532 -429
rect 3498 -637 3532 -621
rect 3612 -445 3646 -429
rect 3612 -637 3646 -621
rect 3708 -445 3742 -429
rect 3708 -637 3742 -621
rect 3822 -445 3856 -429
rect 3822 -637 3856 -621
rect 3918 -445 3952 -429
rect 3918 -637 3952 -621
rect 4032 -445 4066 -429
rect 4032 -637 4066 -621
rect 4128 -445 4162 -429
rect 4128 -637 4162 -621
rect 4242 -445 4276 -385
rect 4242 -637 4276 -621
rect 4338 -445 4372 -385
rect 4338 -637 4372 -621
rect -4450 -714 -4320 -680
rect -4286 -714 -4238 -680
rect -3916 -714 -3900 -680
rect -3866 -714 -3850 -680
rect -3496 -714 -3480 -680
rect -3446 -714 -3430 -680
rect -3076 -714 -3060 -680
rect -3026 -714 -3010 -680
rect -2656 -714 -2640 -680
rect -2606 -714 -2590 -680
rect -2236 -714 -2220 -680
rect -2186 -714 -2170 -680
rect -1816 -714 -1800 -680
rect -1766 -714 -1750 -680
rect -1396 -714 -1380 -680
rect -1346 -714 -1330 -680
rect -976 -714 -960 -680
rect -926 -714 -910 -680
rect -556 -714 -540 -680
rect -506 -714 -490 -680
rect -136 -714 -120 -680
rect -86 -714 -70 -680
rect 284 -714 300 -680
rect 334 -714 350 -680
rect 704 -714 720 -680
rect 754 -714 770 -680
rect 1124 -714 1140 -680
rect 1174 -714 1190 -680
rect 1544 -714 1560 -680
rect 1594 -714 1610 -680
rect 1964 -714 1980 -680
rect 2014 -714 2030 -680
rect 2384 -714 2400 -680
rect 2434 -714 2450 -680
rect 2804 -714 2820 -680
rect 2854 -714 2870 -680
rect 3224 -714 3240 -680
rect 3274 -714 3290 -680
rect 3644 -714 3660 -680
rect 3694 -714 3710 -680
rect 4064 -714 4080 -680
rect 4114 -714 4130 -680
rect -4484 -782 -4450 -720
rect 4450 -782 4484 -720
rect -4484 -816 -4388 -782
rect 4388 -816 4484 -782
<< viali >>
rect -4112 147 -4078 181
rect -3692 147 -3658 181
rect -3272 147 -3238 181
rect -2852 147 -2818 181
rect -2432 147 -2398 181
rect -2012 147 -1978 181
rect -1592 147 -1558 181
rect -1172 147 -1138 181
rect -752 147 -718 181
rect -332 147 -298 181
rect 88 147 122 181
rect 508 147 542 181
rect 928 147 962 181
rect 1348 147 1382 181
rect 1768 147 1802 181
rect 2188 147 2222 181
rect 2608 147 2642 181
rect 3028 147 3062 181
rect 3448 147 3482 181
rect 3868 147 3902 181
rect -3902 -181 -3868 -147
rect -3482 -181 -3448 -147
rect -3062 -181 -3028 -147
rect -2642 -181 -2608 -147
rect -2222 -181 -2188 -147
rect -1802 -181 -1768 -147
rect -1382 -181 -1348 -147
rect -962 -181 -928 -147
rect -542 -181 -508 -147
rect -122 -181 -88 -147
rect 298 -181 332 -147
rect 718 -181 752 -147
rect 1138 -181 1172 -147
rect 1558 -181 1592 -147
rect 1978 -181 2012 -147
rect 2398 -181 2432 -147
rect 2818 -181 2852 -147
rect 3238 -181 3272 -147
rect 3658 -181 3692 -147
rect 4078 -181 4112 -147
rect -4110 -385 -4076 -351
rect -3690 -385 -3656 -351
rect -3270 -385 -3236 -351
rect -2850 -385 -2816 -351
rect -2430 -385 -2396 -351
rect -2010 -385 -1976 -351
rect -1590 -385 -1556 -351
rect -1170 -385 -1136 -351
rect -750 -385 -716 -351
rect -330 -385 -296 -351
rect 90 -385 124 -351
rect 510 -385 544 -351
rect 930 -385 964 -351
rect 1350 -385 1384 -351
rect 1770 -385 1804 -351
rect 2190 -385 2224 -351
rect 2610 -385 2644 -351
rect 3030 -385 3064 -351
rect 3450 -385 3484 -351
rect 3870 -385 3904 -351
rect -3900 -714 -3866 -680
rect -3480 -714 -3446 -680
rect -3060 -714 -3026 -680
rect -2640 -714 -2606 -680
rect -2220 -714 -2186 -680
rect -1800 -714 -1766 -680
rect -1380 -714 -1346 -680
rect -960 -714 -926 -680
rect -540 -714 -506 -680
rect -120 -714 -86 -680
rect 300 -714 334 -680
rect 720 -714 754 -680
rect 1140 -714 1174 -680
rect 1560 -714 1594 -680
rect 1980 -714 2014 -680
rect 2400 -714 2434 -680
rect 2820 -714 2854 -680
rect 3240 -714 3274 -680
rect 3660 -714 3694 -680
rect 4080 -714 4114 -680
<< metal1 >>
rect -4124 181 -4066 187
rect -4124 147 -4112 181
rect -4078 147 -4066 181
rect -4124 141 -4066 147
rect -3704 181 -3646 187
rect -3704 147 -3692 181
rect -3658 147 -3646 181
rect -3704 141 -3646 147
rect -3284 181 -3226 187
rect -3284 147 -3272 181
rect -3238 147 -3226 181
rect -3284 141 -3226 147
rect -2864 181 -2806 187
rect -2864 147 -2852 181
rect -2818 147 -2806 181
rect -2864 141 -2806 147
rect -2444 181 -2386 187
rect -2444 147 -2432 181
rect -2398 147 -2386 181
rect -2444 141 -2386 147
rect -2024 181 -1966 187
rect -2024 147 -2012 181
rect -1978 147 -1966 181
rect -2024 141 -1966 147
rect -1604 181 -1546 187
rect -1604 147 -1592 181
rect -1558 147 -1546 181
rect -1604 141 -1546 147
rect -1184 181 -1126 187
rect -1184 147 -1172 181
rect -1138 147 -1126 181
rect -1184 141 -1126 147
rect -764 181 -706 187
rect -764 147 -752 181
rect -718 147 -706 181
rect -764 141 -706 147
rect -344 181 -286 187
rect -344 147 -332 181
rect -298 147 -286 181
rect -344 141 -286 147
rect 76 181 134 187
rect 76 147 88 181
rect 122 147 134 181
rect 76 141 134 147
rect 496 181 554 187
rect 496 147 508 181
rect 542 147 554 181
rect 496 141 554 147
rect 916 181 974 187
rect 916 147 928 181
rect 962 147 974 181
rect 916 141 974 147
rect 1336 181 1394 187
rect 1336 147 1348 181
rect 1382 147 1394 181
rect 1336 141 1394 147
rect 1756 181 1814 187
rect 1756 147 1768 181
rect 1802 147 1814 181
rect 1756 141 1814 147
rect 2176 181 2234 187
rect 2176 147 2188 181
rect 2222 147 2234 181
rect 2176 141 2234 147
rect 2596 181 2654 187
rect 2596 147 2608 181
rect 2642 147 2654 181
rect 2596 141 2654 147
rect 3016 181 3074 187
rect 3016 147 3028 181
rect 3062 147 3074 181
rect 3016 141 3074 147
rect 3436 181 3494 187
rect 3436 147 3448 181
rect 3482 147 3494 181
rect 3436 141 3494 147
rect 3856 181 3914 187
rect 3856 147 3868 181
rect 3902 147 3914 181
rect 3856 141 3914 147
rect -3914 -147 -3856 -141
rect -3914 -181 -3902 -147
rect -3868 -181 -3856 -147
rect -3914 -187 -3856 -181
rect -3494 -147 -3436 -141
rect -3494 -181 -3482 -147
rect -3448 -181 -3436 -147
rect -3494 -187 -3436 -181
rect -3074 -147 -3016 -141
rect -3074 -181 -3062 -147
rect -3028 -181 -3016 -147
rect -3074 -187 -3016 -181
rect -2654 -147 -2596 -141
rect -2654 -181 -2642 -147
rect -2608 -181 -2596 -147
rect -2654 -187 -2596 -181
rect -2234 -147 -2176 -141
rect -2234 -181 -2222 -147
rect -2188 -181 -2176 -147
rect -2234 -187 -2176 -181
rect -1814 -147 -1756 -141
rect -1814 -181 -1802 -147
rect -1768 -181 -1756 -147
rect -1814 -187 -1756 -181
rect -1394 -147 -1336 -141
rect -1394 -181 -1382 -147
rect -1348 -181 -1336 -147
rect -1394 -187 -1336 -181
rect -974 -147 -916 -141
rect -974 -181 -962 -147
rect -928 -181 -916 -147
rect -974 -187 -916 -181
rect -554 -147 -496 -141
rect -554 -181 -542 -147
rect -508 -181 -496 -147
rect -554 -187 -496 -181
rect -134 -147 -76 -141
rect -134 -181 -122 -147
rect -88 -181 -76 -147
rect -134 -187 -76 -181
rect 286 -147 344 -141
rect 286 -181 298 -147
rect 332 -181 344 -147
rect 286 -187 344 -181
rect 706 -147 764 -141
rect 706 -181 718 -147
rect 752 -181 764 -147
rect 706 -187 764 -181
rect 1126 -147 1184 -141
rect 1126 -181 1138 -147
rect 1172 -181 1184 -147
rect 1126 -187 1184 -181
rect 1546 -147 1604 -141
rect 1546 -181 1558 -147
rect 1592 -181 1604 -147
rect 1546 -187 1604 -181
rect 1966 -147 2024 -141
rect 1966 -181 1978 -147
rect 2012 -181 2024 -147
rect 1966 -187 2024 -181
rect 2386 -147 2444 -141
rect 2386 -181 2398 -147
rect 2432 -181 2444 -147
rect 2386 -187 2444 -181
rect 2806 -147 2864 -141
rect 2806 -181 2818 -147
rect 2852 -181 2864 -147
rect 2806 -187 2864 -181
rect 3226 -147 3284 -141
rect 3226 -181 3238 -147
rect 3272 -181 3284 -147
rect 3226 -187 3284 -181
rect 3646 -147 3704 -141
rect 3646 -181 3658 -147
rect 3692 -181 3704 -147
rect 3646 -187 3704 -181
rect 4066 -147 4124 -141
rect 4066 -181 4078 -147
rect 4112 -181 4124 -147
rect 4066 -187 4124 -181
rect -4122 -351 -4064 -345
rect -4122 -385 -4110 -351
rect -4076 -385 -4064 -351
rect -4122 -391 -4064 -385
rect -3702 -351 -3644 -345
rect -3702 -385 -3690 -351
rect -3656 -385 -3644 -351
rect -3702 -391 -3644 -385
rect -3282 -351 -3224 -345
rect -3282 -385 -3270 -351
rect -3236 -385 -3224 -351
rect -3282 -391 -3224 -385
rect -2862 -351 -2804 -345
rect -2862 -385 -2850 -351
rect -2816 -385 -2804 -351
rect -2862 -391 -2804 -385
rect -2442 -351 -2384 -345
rect -2442 -385 -2430 -351
rect -2396 -385 -2384 -351
rect -2442 -391 -2384 -385
rect -2022 -351 -1964 -345
rect -2022 -385 -2010 -351
rect -1976 -385 -1964 -351
rect -2022 -391 -1964 -385
rect -1602 -351 -1544 -345
rect -1602 -385 -1590 -351
rect -1556 -385 -1544 -351
rect -1602 -391 -1544 -385
rect -1182 -351 -1124 -345
rect -1182 -385 -1170 -351
rect -1136 -385 -1124 -351
rect -1182 -391 -1124 -385
rect -762 -351 -704 -345
rect -762 -385 -750 -351
rect -716 -385 -704 -351
rect -762 -391 -704 -385
rect -342 -351 -284 -345
rect -342 -385 -330 -351
rect -296 -385 -284 -351
rect -342 -391 -284 -385
rect 78 -351 136 -345
rect 78 -385 90 -351
rect 124 -385 136 -351
rect 78 -391 136 -385
rect 498 -351 556 -345
rect 498 -385 510 -351
rect 544 -385 556 -351
rect 498 -391 556 -385
rect 918 -351 976 -345
rect 918 -385 930 -351
rect 964 -385 976 -351
rect 918 -391 976 -385
rect 1338 -351 1396 -345
rect 1338 -385 1350 -351
rect 1384 -385 1396 -351
rect 1338 -391 1396 -385
rect 1758 -351 1816 -345
rect 1758 -385 1770 -351
rect 1804 -385 1816 -351
rect 1758 -391 1816 -385
rect 2178 -351 2236 -345
rect 2178 -385 2190 -351
rect 2224 -385 2236 -351
rect 2178 -391 2236 -385
rect 2598 -351 2656 -345
rect 2598 -385 2610 -351
rect 2644 -385 2656 -351
rect 2598 -391 2656 -385
rect 3018 -351 3076 -345
rect 3018 -385 3030 -351
rect 3064 -385 3076 -351
rect 3018 -391 3076 -385
rect 3438 -351 3496 -345
rect 3438 -385 3450 -351
rect 3484 -385 3496 -351
rect 3438 -391 3496 -385
rect 3858 -351 3916 -345
rect 3858 -385 3870 -351
rect 3904 -385 3916 -351
rect 3858 -391 3916 -385
rect -3912 -680 -3854 -674
rect -3912 -714 -3900 -680
rect -3866 -714 -3854 -680
rect -3912 -720 -3854 -714
rect -3492 -680 -3434 -674
rect -3492 -714 -3480 -680
rect -3446 -714 -3434 -680
rect -3492 -720 -3434 -714
rect -3072 -680 -3014 -674
rect -3072 -714 -3060 -680
rect -3026 -714 -3014 -680
rect -3072 -720 -3014 -714
rect -2652 -680 -2594 -674
rect -2652 -714 -2640 -680
rect -2606 -714 -2594 -680
rect -2652 -720 -2594 -714
rect -2232 -680 -2174 -674
rect -2232 -714 -2220 -680
rect -2186 -714 -2174 -680
rect -2232 -720 -2174 -714
rect -1812 -680 -1754 -674
rect -1812 -714 -1800 -680
rect -1766 -714 -1754 -680
rect -1812 -720 -1754 -714
rect -1392 -680 -1334 -674
rect -1392 -714 -1380 -680
rect -1346 -714 -1334 -680
rect -1392 -720 -1334 -714
rect -972 -680 -914 -674
rect -972 -714 -960 -680
rect -926 -714 -914 -680
rect -972 -720 -914 -714
rect -552 -680 -494 -674
rect -552 -714 -540 -680
rect -506 -714 -494 -680
rect -552 -720 -494 -714
rect -132 -680 -74 -674
rect -132 -714 -120 -680
rect -86 -714 -74 -680
rect -132 -720 -74 -714
rect 288 -680 346 -674
rect 288 -714 300 -680
rect 334 -714 346 -680
rect 288 -720 346 -714
rect 708 -680 766 -674
rect 708 -714 720 -680
rect 754 -714 766 -680
rect 708 -720 766 -714
rect 1128 -680 1186 -674
rect 1128 -714 1140 -680
rect 1174 -714 1186 -680
rect 1128 -720 1186 -714
rect 1548 -680 1606 -674
rect 1548 -714 1560 -680
rect 1594 -714 1606 -680
rect 1548 -720 1606 -714
rect 1968 -680 2026 -674
rect 1968 -714 1980 -680
rect 2014 -714 2026 -680
rect 1968 -720 2026 -714
rect 2388 -680 2446 -674
rect 2388 -714 2400 -680
rect 2434 -714 2446 -680
rect 2388 -720 2446 -714
rect 2808 -680 2866 -674
rect 2808 -714 2820 -680
rect 2854 -714 2866 -680
rect 2808 -720 2866 -714
rect 3228 -680 3286 -674
rect 3228 -714 3240 -680
rect 3274 -714 3286 -680
rect 3228 -720 3286 -714
rect 3648 -680 3706 -674
rect 3648 -714 3660 -680
rect 3694 -714 3706 -680
rect 3648 -720 3706 -714
rect 4068 -680 4126 -674
rect 4068 -714 4080 -680
rect 4114 -714 4126 -680
rect 4068 -720 4126 -714
<< properties >>
string FIXED_BBOX -4466 -266 4466 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 42 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
