magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< metal3 >>
rect -1310 -1260 1210 1260
<< mimcap >>
rect -1210 1120 1110 1160
rect -1210 -1120 -1170 1120
rect 1070 -1120 1110 1120
rect -1210 -1160 1110 -1120
<< mimcapcontact >>
rect -1170 -1120 1070 1120
<< metal4 >>
rect -1171 1120 1071 1121
rect -1171 -1120 -1170 1120
rect 1070 -1120 1071 1120
rect -1171 -1121 1071 -1120
<< properties >>
string FIXED_BBOX -1310 -1260 1210 1260
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 11.6 l 11.6 val 277.936 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
