* NGSPICE file created from clock.ext - technology: sky130A

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X a_110_47# VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VPB A 0.23fF
C1 VPB VPWR 0.78fF
C2 VPB X 0.03fF
C3 A VPWR 0.07fF
C4 A X 0.00fF
C5 A VGND 0.10fF
C6 VPWR X 2.96fF
C7 a_110_47# VPB 0.81fF
C8 VPWR VGND 0.28fF
C9 a_110_47# A 0.51fF
C10 X VGND 1.95fF
C11 a_110_47# VPWR 0.98fF
C12 a_110_47# X 2.36fF
C13 a_110_47# VGND 0.78fF
C14 VGND VNB 1.05fF
C15 X VNB 0.10fF
C16 VPWR VNB 0.39fF
C17 A VNB 0.43fF
C18 VPB VNB 1.85fF
C19 a_110_47# VNB 1.28fF
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
C0 VPB VGND 0.25fF
C1 VGND VPWR 0.82fF
C2 VPB VPWR 0.27fF
C3 VPWR VNB 0.41fF
C4 VGND VNB 0.37fF
C5 VPB VNB 0.43fF
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
C0 VGND VPWR 3.03fF
C1 VGND VPB 0.87fF
C2 VPB VPWR 0.47fF
C3 VPWR VNB 1.33fF
C4 VGND VNB 0.77fF
C5 VPB VNB 1.14fF
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VPWR X VNB VPB a_283_47# a_390_47#
+ a_27_47#
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=6.517e+11p ps=5.37e+06u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=4.027e+11p pd=3.97e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
C0 a_283_47# VGND 0.14fF
C1 a_283_47# A 0.02fF
C2 a_27_47# X 0.02fF
C3 a_27_47# VPB 0.16fF
C4 VPB X 0.05fF
C5 a_283_47# VPWR 0.17fF
C6 a_27_47# a_390_47# 0.05fF
C7 a_390_47# X 0.12fF
C8 a_27_47# VGND 0.24fF
C9 a_27_47# A 0.29fF
C10 a_390_47# VPB 0.06fF
C11 X VGND 0.14fF
C12 A X 0.00fF
C13 VPB A 0.06fF
C14 a_390_47# VGND 0.14fF
C15 a_27_47# VPWR 0.31fF
C16 a_390_47# A 0.01fF
C17 A VGND 0.02fF
C18 VPWR X 0.19fF
C19 VPB VPWR 0.32fF
C20 a_390_47# VPWR 0.16fF
C21 VPWR VGND 0.11fF
C22 A VPWR 0.02fF
C23 a_283_47# a_27_47# 0.18fF
C24 a_283_47# X 0.04fF
C25 a_283_47# VPB 0.12fF
C26 a_283_47# a_390_47# 0.44fF
C27 VGND VNB 0.43fF
C28 X VNB 0.05fF
C29 VPWR VNB 0.16fF
C30 A VNB 0.13fF
C31 VPB VNB 0.78fF
C32 a_390_47# VNB 0.10fF
C33 a_283_47# VNB 0.18fF
C34 a_27_47# VNB 0.18fF
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 Y A 0.88fF
C1 VGND VPWR 0.10fF
C2 VGND Y 0.56fF
C3 VGND A 0.13fF
C4 VPWR VPB 0.34fF
C5 VPB Y 0.05fF
C6 VPWR Y 1.13fF
C7 VPB A 0.21fF
C8 VPWR A 0.13fF
C9 VGND VNB 0.40fF
C10 Y VNB 0.10fF
C11 VPWR VNB 0.14fF
C12 A VNB 0.47fF
C13 VPB VNB 0.69fF
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB a_27_47#
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 a_27_47# VGND 0.77fF
C1 a_27_47# A 0.10fF
C2 VGND A 0.08fF
C3 a_27_47# B 0.33fF
C4 B VGND 0.10fF
C5 B A 0.16fF
C6 Y VPB 0.02fF
C7 Y VPWR 1.44fF
C8 Y a_27_47# 0.41fF
C9 Y VGND 0.13fF
C10 Y A 0.35fF
C11 Y B 0.30fF
C12 VPB VPWR 0.43fF
C13 VPB A 0.18fF
C14 VPB B 0.21fF
C15 a_27_47# VPWR 0.07fF
C16 VGND VPWR 0.12fF
C17 A VPWR 0.09fF
C18 B VPWR 0.12fF
C19 VGND VNB 0.48fF
C20 Y VNB 0.01fF
C21 VPWR VNB 0.18fF
C22 A VNB 0.26fF
C23 B VNB 0.30fF
C24 VPB VNB 0.87fF
C25 a_27_47# VNB 0.06fF
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
C0 VGND VPB 0.16fF
C1 VPWR VPB 0.24fF
C2 VPWR VGND 0.54fF
C3 VPWR VNB 0.28fF
C4 VGND VNB 0.31fF
C5 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
C0 VGND VPB 0.55fF
C1 VPWR VPB 0.37fF
C2 VPWR VGND 1.92fF
C3 VPWR VNB 0.86fF
C4 VGND VNB 0.56fF
C5 VPB VNB 0.78fF
.ends

.subckt sky130_fd_sc_hd__dfxbp_1 CLK D VGND VPWR Q Q_N a_975_413# a_891_413# VNB VPB
+ a_466_413# a_592_47# a_1059_315# a_193_47# a_561_413# a_634_159# a_381_47# a_1017_47#
+ a_1490_369# a_27_47#
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=9.432e+11p ps=1.006e+07u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.32905e+12p pd=1.228e+07u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X6 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1059_315# a_1490_369# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X17 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23 Q_N a_1490_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q_N a_1490_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 VPWR a_1059_315# a_1490_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
C0 a_193_47# a_891_413# 0.38fF
C1 a_891_413# VPB 0.08fF
C2 a_634_159# CLK 0.01fF
C3 a_381_47# VGND 0.09fF
C4 VPWR Q_N 0.25fF
C5 VGND Q 0.14fF
C6 a_1059_315# a_1490_369# 0.18fF
C7 a_466_413# a_1059_315# 0.05fF
C8 a_27_47# CLK 0.33fF
C9 a_466_413# a_1490_369# 0.02fF
C10 a_891_413# CLK 0.01fF
C11 a_634_159# D 0.04fF
C12 a_193_47# a_1059_315# 0.13fF
C13 a_1059_315# VPB 0.24fF
C14 a_381_47# Q 0.01fF
C15 VGND Q_N 0.11fF
C16 a_193_47# a_1490_369# 0.03fF
C17 a_1490_369# VPB 0.06fF
C18 a_193_47# a_466_413# 0.20fF
C19 a_466_413# VPB 0.08fF
C20 a_27_47# D 0.17fF
C21 a_891_413# D 0.01fF
C22 a_193_47# VPB 0.21fF
C23 a_634_159# VPWR 0.21fF
C24 a_1059_315# CLK 0.01fF
C25 a_381_47# Q_N 0.01fF
C26 Q Q_N 0.05fF
C27 a_592_47# VGND 0.00fF
C28 a_1490_369# CLK 0.00fF
C29 a_466_413# CLK 0.01fF
C30 a_27_47# VPWR 0.60fF
C31 a_891_413# VPWR 0.20fF
C32 a_193_47# CLK 0.06fF
C33 a_634_159# VGND 0.18fF
C34 VPB CLK 0.14fF
C35 a_1059_315# D 0.02fF
C36 a_1490_369# D 0.01fF
C37 a_1017_47# VGND 0.00fF
C38 a_466_413# D 0.03fF
C39 a_27_47# VGND 0.30fF
C40 a_381_47# a_634_159# 0.03fF
C41 a_975_413# VPWR 0.01fF
C42 a_891_413# VGND 0.18fF
C43 a_634_159# Q 0.02fF
C44 a_193_47# D 0.30fF
C45 VPB D 0.13fF
C46 a_1059_315# VPWR 0.37fF
C47 a_1490_369# VPWR 0.29fF
C48 a_466_413# VPWR 0.31fF
C49 a_381_47# a_27_47# 0.16fF
C50 a_27_47# Q 0.03fF
C51 a_381_47# a_891_413# 0.02fF
C52 a_891_413# Q 0.04fF
C53 a_634_159# Q_N 0.01fF
C54 a_193_47# VPWR 0.37fF
C55 CLK D 0.04fF
C56 VPB VPWR 0.73fF
C57 a_1059_315# VGND 0.22fF
C58 a_1490_369# VGND 0.12fF
C59 a_466_413# VGND 0.15fF
C60 a_27_47# Q_N 0.02fF
C61 a_466_413# a_561_413# 0.01fF
C62 a_891_413# Q_N 0.02fF
C63 a_193_47# VGND 0.24fF
C64 a_381_47# a_1059_315# 0.01fF
C65 CLK VPWR 0.03fF
C66 a_1059_315# Q 0.19fF
C67 a_381_47# a_1490_369# 0.01fF
C68 a_1490_369# Q 0.31fF
C69 a_381_47# a_466_413# 0.09fF
C70 a_466_413# Q 0.02fF
C71 a_381_47# a_193_47# 0.22fF
C72 a_193_47# Q 0.03fF
C73 a_381_47# VPB 0.03fF
C74 CLK VGND 0.04fF
C75 VPB Q 0.02fF
C76 D VPWR 0.03fF
C77 a_1059_315# Q_N 0.03fF
C78 a_1490_369# Q_N 0.14fF
C79 a_27_47# a_634_159# 0.29fF
C80 a_466_413# Q_N 0.01fF
C81 a_634_159# a_891_413# 0.10fF
C82 a_193_47# Q_N 0.02fF
C83 a_381_47# CLK 0.01fF
C84 CLK Q 0.00fF
C85 D VGND 0.05fF
C86 VPB Q_N 0.05fF
C87 a_891_413# a_1017_47# 0.01fF
C88 a_27_47# a_891_413# 0.09fF
C89 a_466_413# a_592_47# 0.01fF
C90 a_634_159# a_1059_315# 0.06fF
C91 a_381_47# D 0.21fF
C92 CLK Q_N 0.00fF
C93 VPWR VGND 0.26fF
C94 D Q 0.00fF
C95 a_634_159# a_1490_369# 0.02fF
C96 a_634_159# a_466_413# 0.36fF
C97 a_561_413# VPWR 0.01fF
C98 a_27_47# a_1059_315# 0.14fF
C99 a_27_47# a_1490_369# 0.03fF
C100 a_891_413# a_975_413# 0.02fF
C101 a_27_47# a_466_413# 0.51fF
C102 a_634_159# a_193_47# 0.21fF
C103 a_634_159# VPB 0.08fF
C104 a_1059_315# a_891_413# 0.44fF
C105 a_381_47# VPWR 0.13fF
C106 VPWR Q 0.24fF
C107 D Q_N 0.00fF
C108 a_1490_369# a_891_413# 0.04fF
C109 a_466_413# a_891_413# 0.04fF
C110 a_27_47# a_193_47# 1.69fF
C111 a_27_47# VPB 0.30fF
C112 Q_N VNB 0.05fF
C113 Q VNB 0.01fF
C114 VGND VNB 0.95fF
C115 VPWR VNB 0.37fF
C116 D VNB 0.12fF
C117 CLK VNB 0.18fF
C118 VPB VNB 1.76fF
C119 a_381_47# VNB 0.03fF
C120 a_1490_369# VNB 0.09fF
C121 a_891_413# VNB 0.12fF
C122 a_1059_315# VNB 0.24fF
C123 a_466_413# VNB 0.11fF
C124 a_634_159# VNB 0.12fF
C125 a_193_47# VNB 0.21fF
C126 a_27_47# VNB 0.31fF
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VGND B 0.06fF
C1 VGND a_113_47# 0.01fF
C2 A VPB 0.06fF
C3 VPWR A 0.05fF
C4 VPWR VPB 0.24fF
C5 VGND A 0.02fF
C6 VGND VPWR 0.05fF
C7 Y B 0.05fF
C8 Y a_113_47# 0.01fF
C9 Y A 0.11fF
C10 Y VPB 0.02fF
C11 Y VPWR 0.40fF
C12 Y VGND 0.21fF
C13 A B 0.07fF
C14 VPB B 0.06fF
C15 VPWR B 0.06fF
C16 VGND VNB 0.23fF
C17 Y VNB 0.05fF
C18 VPWR VNB 0.06fF
C19 A VNB 0.10fF
C20 B VNB 0.10fF
C21 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 A Y 0.26fF
C1 VPB A 0.14fF
C2 VPB Y 0.00fF
C3 VPWR VGND 0.04fF
C4 A VGND 0.05fF
C5 Y VGND 0.17fF
C6 A VPWR 0.04fF
C7 Y VPWR 0.35fF
C8 VPB VPWR 0.23fF
C9 VGND VNB 0.23fF
C10 Y VNB 0.04fF
C11 VPWR VNB 0.06fF
C12 A VNB 0.24fF
C13 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB a_505_21# a_439_47# a_218_47#
+ a_76_199# a_218_374#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 a_76_199# X 0.18fF
C1 a_505_21# VPWR 0.12fF
C2 VPB a_505_21# 0.09fF
C3 X VPWR 0.23fF
C4 A0 S 0.09fF
C5 a_76_199# VPWR 0.15fF
C6 VPB X 0.06fF
C7 VPB a_76_199# 0.08fF
C8 A0 VGND 0.08fF
C9 VPB VPWR 0.44fF
C10 a_505_21# S 0.26fF
C11 A0 A1 0.41fF
C12 X S 0.08fF
C13 a_76_199# S 0.54fF
C14 a_218_47# VGND 0.01fF
C15 a_505_21# VGND 0.16fF
C16 a_535_374# S 0.01fF
C17 X VGND 0.09fF
C18 VPWR S 0.64fF
C19 a_76_199# VGND 0.24fF
C20 VPB S 0.24fF
C21 a_505_21# A1 0.16fF
C22 a_439_47# VGND 0.01fF
C23 X A1 0.04fF
C24 VPWR VGND 0.12fF
C25 a_76_199# A1 0.41fF
C26 a_439_47# A1 0.00fF
C27 VPWR A1 0.04fF
C28 a_76_199# a_218_374# 0.00fF
C29 VPB A1 0.06fF
C30 S VGND 0.07fF
C31 S A1 0.25fF
C32 a_505_21# A0 0.08fF
C33 a_218_374# S 0.01fF
C34 A0 X 0.02fF
C35 VGND A1 0.12fF
C36 a_76_199# A0 0.14fF
C37 a_439_47# A0 0.01fF
C38 A0 VPWR 0.01fF
C39 VPB A0 0.08fF
C40 a_505_21# X 0.02fF
C41 a_218_47# a_76_199# 0.01fF
C42 a_76_199# a_505_21# 0.04fF
C43 VGND VNB 0.48fF
C44 A1 VNB 0.09fF
C45 A0 VNB 0.08fF
C46 S VNB 0.17fF
C47 VPWR VNB 0.18fF
C48 X VNB 0.06fF
C49 VPB VNB 0.87fF
C50 a_505_21# VNB 0.15fF
C51 a_76_199# VNB 0.11fF
.ends

.subckt clock clk p2d_b p2d p2_b p2 p1d_b p1d p1_b p1 Ad_b Ad A_b A Bd_b Bd B_b B
+ VDD VSS
Xsky130_fd_sc_hd__clkbuf_16_11 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD p1d_b sky130_fd_sc_hd__clkbuf_16_11/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_226 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_204 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_12 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD p2d_b sky130_fd_sc_hd__clkbuf_16_12/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_13 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD p2d sky130_fd_sc_hd__clkbuf_16_13/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_217 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_0 sky130_fd_sc_hd__clkinv_1_0/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_14 sky130_fd_sc_hd__clkinv_4_10/Y VSS VDD p2_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_10 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_4_10/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_1 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_15 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD p2 sky130_fd_sc_hd__clkbuf_16_15/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_11 sky130_fd_sc_hd__nand2_4_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_2 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_3 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS VDD sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/A
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_4 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_2 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__nand2_4_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__nand2_4_2/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_190 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_5 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_180 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_4_3 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__nand2_4_3/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_6 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_7/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_7 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_193 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_8 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_9/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_4_4/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_172 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_183 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_9 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_9/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_5/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_195 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_140 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_162 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_6 sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/A
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_190 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_196 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_90 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_7 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_191 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_180 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_181/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_186 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_80 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_81/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_91 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_8 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__clkinv_4_8/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_192 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_181 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_170 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_165 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_198 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_70 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_81 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_92 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_9 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__clkinv_4_9/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_193 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_182 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_183/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_171 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_160 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_111 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_166 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_188 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_60 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_71 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_82 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_83/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_93 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_0 p2 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__mux2_1_0/S
+ sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__dfxbp_1_0/a_975_413# sky130_fd_sc_hd__dfxbp_1_0/a_891_413#
+ VSS VDD sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_592_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__dfxbp_1_0/a_1017_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_194 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_183 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_172 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_150 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_161 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_178 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_189 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_50 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_61 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_62/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_72 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_83 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_94 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_1 clk sky130_fd_sc_hd__dfxbp_1_1/D VSS VDD sky130_fd_sc_hd__nand2_1_1/A
+ sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__dfxbp_1_1/a_975_413# sky130_fd_sc_hd__dfxbp_1_1/a_891_413#
+ VSS VDD sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_592_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# sky130_fd_sc_hd__dfxbp_1_1/a_1017_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_195 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_184 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_185/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_173 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_151 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_140 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_162 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_157 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_168 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_179 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_40 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_51 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_62 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_73 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_84 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_85/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_95 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_130 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_141 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_196 sky130_fd_sc_hd__clkinv_1_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_185 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_174 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_152 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_163 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_165/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_158 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_41 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_30 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_52 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_63 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_64/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_74 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_85 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_96 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_197 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_186 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_175 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_164 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_166/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_120 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_131 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_142 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_153 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD B sky130_fd_sc_hd__clkbuf_16_0/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_159 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_42 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_20 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_21/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_31 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_53 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_64 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_75 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_86 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_97 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_1/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_198 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_187 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_176 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_165 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_165/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_110 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_121 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_132 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_133/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_154 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_143 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD Bd sky130_fd_sc_hd__clkbuf_16_1/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_10 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_41/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_21 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_43 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_43/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_54 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_32 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_40/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_65 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_66/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_76 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_98 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_87 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_199 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_3/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_188 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_177 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_155 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_166 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_111 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_100 sky130_fd_sc_hd__clkinv_1_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_122 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD
+ sky130_fd_sc_hd__nand2_1_4/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_133 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_144 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD B_b sky130_fd_sc_hd__clkbuf_16_2/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_22 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_23/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_44 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_11 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_46/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_55 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_33 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_66 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_77 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_99 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_88 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_189 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_178 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_179/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_167 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_112 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_101 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_123 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_134 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_135/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_156 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_145 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD Bd_b sky130_fd_sc_hd__clkbuf_16_3/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_23 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_12 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_45 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_45/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_56 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_34 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_67 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_78 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_79/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_89 sky130_fd_sc_hd__clkinv_1_1/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_157 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_102 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_113 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_114/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_124 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_135 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_146 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_179 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_168 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_4 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD Ad_b sky130_fd_sc_hd__clkbuf_16_4/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_24 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_13 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_46 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_57 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_35 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_68 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_0/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_79 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_169 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_2/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_103 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_2/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_114 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_125 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_136 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_137/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_147 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_158 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_5 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD Ad sky130_fd_sc_hd__clkbuf_16_5/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_14 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_25 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_26/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_47 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_58 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_36 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_69 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_104 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_115 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_126 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_137 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_148 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_159 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_160/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_6 sky130_fd_sc_hd__clkinv_4_4/Y VSS VDD A_b sky130_fd_sc_hd__clkbuf_16_6/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_15 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_48 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_26 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_37 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_59 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_60/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_105 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_116 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_127 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_138 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_139/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_149 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_7 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD A sky130_fd_sc_hd__clkbuf_16_7/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_16 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_49 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_1/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_27 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_28/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_38 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_250 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_106 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_117 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_119/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_128 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_139 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_8 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD p1 sky130_fd_sc_hd__clkbuf_16_8/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_17 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_28 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_39 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_107 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_118 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_120/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_129 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_9 sky130_fd_sc_hd__clkinv_4_7/Y VSS VDD p1_b sky130_fd_sc_hd__clkbuf_16_9/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_1_0/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_18 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_19/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_29 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_30/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_108 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_119 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_119/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__nand2_1_2/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_19 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_1_1/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_109 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_110/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_1_3/A clk VSS VDD sky130_fd_sc_hd__nand2_4_3/A
+ VSS VDD sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_254 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_232 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_210 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/B
+ VSS VDD sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1_4/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_211 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_200 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux2_1_0 Ad_b Bd_b sky130_fd_sc_hd__mux2_1_0/S VSS VDD sky130_fd_sc_hd__mux2_1_0/X
+ VSS VDD sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/a_439_47#
+ sky130_fd_sc_hd__mux2_1_0/a_218_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374#
+ sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_234 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_246 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_224 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_10 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD p1d sky130_fd_sc_hd__clkbuf_16_10/a_110_47#
+ VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_6 clk VSS VDD sky130_fd_sc_hd__nand2_1_2/A VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_247 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_225 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
C0 p2 Bd_b 0.56fF
C1 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.01fF
C2 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.08fF
C3 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.02fF
C4 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C5 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C6 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.01fF
C7 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C8 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.01fF
C9 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.02fF
C10 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.01fF
C11 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C12 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# VDD 0.48fF
C13 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.01fF
C14 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C15 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C16 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C17 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C18 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.08fF
C19 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.04fF
C20 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.01fF
C21 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C22 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.04fF
C23 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.04fF
C24 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# VDD 0.16fF
C25 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.03fF
C26 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C27 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C28 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.00fF
C29 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.02fF
C30 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.00fF
C31 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C32 B B_b 0.47fF
C33 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.14fF
C34 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.09fF
C35 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C36 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.00fF
C37 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C38 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C39 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.01fF
C40 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.01fF
C41 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.01fF
C42 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.01fF
C43 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__dfxbp_1_0/a_1017_47# -0.00fF
C44 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_1_1/A 0.06fF
C45 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_1/A 0.47fF
C46 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C47 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C48 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C49 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.08fF
C50 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.04fF
C51 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.16fF
C52 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# VDD 0.15fF
C53 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.09fF
C54 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.04fF
C55 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.04fF
C56 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C57 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C58 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.02fF
C59 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_2/B 0.23fF
C60 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.02fF
C61 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C62 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C63 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# VDD 0.11fF
C64 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C65 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.01fF
C66 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C67 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C68 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C69 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C70 Ad sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.15fF
C71 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# A_b 0.15fF
C72 VDD sky130_fd_sc_hd__clkinv_4_5/Y 4.36fF
C73 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.00fF
C74 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.04fF
C75 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.04fF
C76 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.01fF
C77 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C78 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C79 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C80 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.01fF
C81 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.00fF
C82 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.00fF
C83 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.00fF
C84 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.01fF
C85 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C86 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C87 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.11fF
C88 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.01fF
C89 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.01fF
C90 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C91 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VDD 0.59fF
C92 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C93 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C94 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C95 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C96 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C97 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C98 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C99 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C100 sky130_fd_sc_hd__nand2_4_0/B VDD 0.55fF
C101 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.01fF
C102 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.02fF
C103 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C104 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C105 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.03fF
C106 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C107 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.02fF
C108 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.02fF
C109 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C110 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.11fF
C111 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C112 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C113 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C114 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C115 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C116 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C117 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C118 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.11fF
C119 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C120 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.03fF
C121 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C122 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C123 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.00fF
C124 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.01fF
C125 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.03fF
C126 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.01fF
C127 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.02fF
C128 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.02fF
C129 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C130 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C131 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C132 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.09fF
C133 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.01fF
C134 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C135 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.02fF
C136 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C137 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.11fF
C138 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.04fF
C139 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C140 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C141 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C142 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C143 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C144 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C145 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C146 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C147 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# VDD 0.15fF
C148 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.03fF
C149 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C150 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C151 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C152 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C153 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__mux2_1_0/X 0.05fF
C154 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.16fF
C155 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C156 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.04fF
C157 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C158 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C159 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C160 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.12fF
C161 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.00fF
C162 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C163 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.01fF
C164 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C165 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C166 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C167 p2d_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.07fF
C168 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2_b 0.06fF
C169 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.02fF
C170 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.02fF
C171 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C172 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C173 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# VDD 0.14fF
C174 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.09fF
C175 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.01fF
C176 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# VDD 0.10fF
C177 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C178 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C179 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C180 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VDD 0.14fF
C181 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C182 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C183 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C184 VDD p1_b 1.24fF
C185 sky130_fd_sc_hd__mux2_1_0/a_505_21# Bd_b 0.04fF
C186 sky130_fd_sc_hd__clkinv_4_4/Y A_b 0.03fF
C187 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C188 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C189 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C190 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C191 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C192 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 1.69fF
C193 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# VDD 0.14fF
C194 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C195 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C196 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# VDD 0.16fF
C197 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C198 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.01fF
C199 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C200 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.01fF
C201 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.02fF
C202 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.01fF
C203 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C204 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# 0.05fF
C205 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.69fF
C206 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VDD 0.48fF
C207 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C208 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# VDD 0.30fF
C209 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.01fF
C210 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.02fF
C211 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C212 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C213 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C214 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.02fF
C215 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C216 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.05fF
C217 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.03fF
C218 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C219 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.84fF
C220 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C221 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.06fF
C222 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.02fF
C223 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.01fF
C224 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C225 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.05fF
C226 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.11fF
C227 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.04fF
C228 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.00fF
C229 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.00fF
C230 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C231 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C232 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.08fF
C233 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.00fF
C234 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.09fF
C235 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.05fF
C236 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C237 Ad_b Bd_b 4.81fF
C238 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C239 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C240 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.01fF
C241 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C242 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C243 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.00fF
C244 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.84fF
C245 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.00fF
C246 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.00fF
C247 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C248 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C249 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C250 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C251 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C252 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.02fF
C253 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C254 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.01fF
C255 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C256 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.01fF
C257 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C258 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C259 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C260 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.01fF
C261 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.03fF
C262 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C263 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C264 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.00fF
C265 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C266 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C267 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.02fF
C268 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# 0.10fF
C269 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.09fF
C270 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C271 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.00fF
C272 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.00fF
C273 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.11fF
C274 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C275 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.33fF
C276 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.11fF
C277 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C278 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.01fF
C279 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.00fF
C280 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C281 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.02fF
C282 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C283 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C284 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.01fF
C285 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.02fF
C286 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# 0.12fF
C287 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C288 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.01fF
C289 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.03fF
C290 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__nand2_4_0/Y 0.09fF
C291 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.02fF
C292 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C293 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.02fF
C294 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.01fF
C295 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.02fF
C296 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.55fF
C297 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkinv_4_5/Y 0.85fF
C298 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C299 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C300 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C301 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A 0.73fF
C302 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.00fF
C303 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C304 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.01fF
C305 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.00fF
C306 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.00fF
C307 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C308 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C309 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.02fF
C310 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C311 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# VDD 0.12fF
C312 sky130_fd_sc_hd__nand2_1_1/A clk 0.06fF
C313 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.04fF
C314 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.04fF
C315 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C316 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# -0.33fF
C317 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.03fF
C318 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.00fF
C319 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.09fF
C320 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.00fF
C321 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A VDD 0.52fF
C322 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C323 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VDD 6.26fF
C324 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.00fF
C325 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.00fF
C326 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.01fF
C327 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C328 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C329 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C330 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C331 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.01fF
C332 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C333 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C334 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.00fF
C335 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C336 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.08fF
C337 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C338 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# 0.15fF
C339 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.01fF
C340 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.01fF
C341 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.05fF
C342 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C343 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# -0.08fF
C344 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.00fF
C345 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.04fF
C346 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.04fF
C347 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.03fF
C348 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.01fF
C349 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C350 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.01fF
C351 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.29fF
C352 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C353 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.00fF
C354 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C355 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.17fF
C356 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C357 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C358 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.06fF
C359 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C360 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C361 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.02fF
C362 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# VDD 0.14fF
C363 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.00fF
C364 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.00fF
C365 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.00fF
C366 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.00fF
C367 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkinv_4_7/A 0.85fF
C368 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.33fF
C369 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C370 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C371 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C372 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.11fF
C373 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.40fF
C374 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Bd_b 0.03fF
C375 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.08fF
C376 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C377 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.57fF
C378 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.02fF
C379 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.01fF
C380 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.08fF
C381 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.04fF
C382 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C383 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.02fF
C384 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.01fF
C385 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# VDD 0.17fF
C386 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C387 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C388 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VDD 0.52fF
C389 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# VDD 0.15fF
C390 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.00fF
C391 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C392 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.08fF
C393 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C394 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C395 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# VDD 0.14fF
C396 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.04fF
C397 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0.04fF
C398 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.04fF
C399 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.04fF
C400 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A VDD 0.56fF
C401 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.05fF
C402 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.05fF
C403 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VDD 0.67fF
C404 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.00fF
C405 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.02fF
C406 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# VDD 0.13fF
C407 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.02fF
C408 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C409 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C410 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C411 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.09fF
C412 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C413 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.02fF
C414 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.69fF
C415 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C416 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C417 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.08fF
C418 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.02fF
C419 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# VDD 0.12fF
C420 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.00fF
C421 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.00fF
C422 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C423 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.03fF
C424 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.09fF
C425 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.00fF
C426 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.00fF
C427 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.00fF
C428 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.08fF
C429 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.67fF
C430 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# VDD 0.29fF
C431 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C432 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C433 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C434 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C435 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C436 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C437 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.15fF
C438 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.02fF
C439 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.02fF
C440 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C441 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C442 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C443 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C444 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C445 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C446 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C447 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.02fF
C448 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.17fF
C449 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C450 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.02fF
C451 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.08fF
C452 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A -0.02fF
C453 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.04fF
C454 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.04fF
C455 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C456 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.30fF
C457 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C458 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.02fF
C459 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C460 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C461 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# 0.01fF
C462 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C463 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.33fF
C464 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# 0.02fF
C465 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# 0.01fF
C466 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C467 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C468 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C469 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C470 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# VDD 0.15fF
C471 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C472 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.03fF
C473 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C474 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.00fF
C475 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.00fF
C476 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C477 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C478 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# VDD 0.13fF
C479 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.02fF
C480 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.02fF
C481 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C482 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# VDD 0.14fF
C483 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# VDD 0.15fF
C484 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VDD 0.52fF
C485 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C486 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.04fF
C487 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.04fF
C488 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.01fF
C489 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.06fF
C490 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# VDD 0.25fF
C491 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# VDD 0.11fF
C492 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C493 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C494 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C495 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C496 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.05fF
C497 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C498 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.00fF
C499 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Ad_b 0.04fF
C500 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C501 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.00fF
C502 VDD sky130_fd_sc_hd__nand2_4_0/A 16.63fF
C503 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.02fF
C504 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.02fF
C505 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C506 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.11fF
C507 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C508 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C509 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C510 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C511 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.01fF
C512 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C513 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.02fF
C514 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VDD 0.69fF
C515 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C516 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C517 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.03fF
C518 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C519 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.02fF
C520 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.14fF
C521 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.51fF
C522 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C523 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C524 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C525 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C526 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C527 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.16fF
C528 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# 0.05fF
C529 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.06fF
C530 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.01fF
C531 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C532 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# 0.00fF
C533 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# 0.00fF
C534 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C535 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C536 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C537 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.00fF
C538 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C539 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.08fF
C540 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.01fF
C541 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.73fF
C542 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.01fF
C543 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# 0.02fF
C544 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# 0.01fF
C545 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# 0.01fF
C546 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C547 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.06fF
C548 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.05fF
C549 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.02fF
C550 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.11fF
C551 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.00fF
C552 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.00fF
C553 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.07fF
C554 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.02fF
C555 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.02fF
C556 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.02fF
C557 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C558 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.06fF
C559 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C560 p2d_b VDD 0.79fF
C561 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.02fF
C562 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.02fF
C563 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.00fF
C564 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.06fF
C565 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.03fF
C566 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VDD 0.14fF
C567 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.08fF
C568 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C569 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.06fF
C570 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.03fF
C571 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C572 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C573 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C574 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.06fF
C575 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C576 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.34fF
C577 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C578 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C579 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C580 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C581 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C582 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C583 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C584 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.02fF
C585 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C586 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C587 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.10fF
C588 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C589 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.01fF
C590 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C591 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_1/Y 0.08fF
C592 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VDD 0.59fF
C593 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# VDD 0.14fF
C594 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C595 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C596 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C597 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C598 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C599 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C600 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C601 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.43fF
C602 Ad A 0.19fF
C603 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# VDD 0.17fF
C604 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.01fF
C605 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.05fF
C606 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.03fF
C607 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C608 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C609 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.08fF
C610 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.00fF
C611 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.03fF
C612 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C613 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.03fF
C614 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__nand2_1_2/B 0.02fF
C615 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C616 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C617 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.03fF
C618 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.05fF
C619 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.05fF
C620 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C621 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C622 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C623 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.01fF
C624 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.03fF
C625 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C626 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.03fF
C627 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.01fF
C628 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.04fF
C629 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.59fF
C630 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.05fF
C631 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C632 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C633 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.00fF
C634 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C635 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C636 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C637 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C638 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.01fF
C639 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.01fF
C640 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C641 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C642 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.00fF
C643 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.01fF
C644 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/B 0.04fF
C645 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C646 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C647 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C648 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C649 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.01fF
C650 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.01fF
C651 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C652 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C653 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C654 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C655 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.06fF
C656 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C657 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.01fF
C658 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.01fF
C659 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C660 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C661 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.03fF
C662 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.01fF
C663 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C664 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.01fF
C665 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.05fF
C666 p1 sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C667 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.06fF
C668 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C669 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.03fF
C670 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.00fF
C671 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.00fF
C672 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C673 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C674 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.03fF
C675 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C676 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C677 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.08fF
C678 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C679 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C680 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C681 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C682 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C683 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C684 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C685 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C686 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C687 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.03fF
C688 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C689 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C690 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.02fF
C691 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.02fF
C692 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.02fF
C693 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C694 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C695 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C696 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.02fF
C697 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C698 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.01fF
C699 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C700 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.09fF
C701 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C702 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.01fF
C703 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# VDD 0.44fF
C704 VDD sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.67fF
C705 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C706 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VDD 0.14fF
C707 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C708 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C709 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C710 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.00fF
C711 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.01fF
C712 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.03fF
C713 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C714 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.02fF
C715 sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C716 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.01fF
C717 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C718 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.06fF
C719 sky130_fd_sc_hd__dfxbp_1_0/Q_N Ad_b 0.01fF
C720 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.01fF
C721 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C722 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C723 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C724 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.01fF
C725 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C726 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.02fF
C727 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.02fF
C728 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.00fF
C729 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C730 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.09fF
C731 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.09fF
C732 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C733 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C734 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C735 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.01fF
C736 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.33fF
C737 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__clkinv_4_5/Y 0.03fF
C738 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C739 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.04fF
C740 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C741 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C742 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C743 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.00fF
C744 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.00fF
C745 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.00fF
C746 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.11fF
C747 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.05fF
C748 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.00fF
C749 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.00fF
C750 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# 0.00fF
C751 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C752 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.04fF
C753 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.04fF
C754 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C755 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C756 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C757 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C758 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.00fF
C759 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.00fF
C760 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C761 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C762 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C763 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.01fF
C764 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.01fF
C765 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_4/B 0.04fF
C766 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.15fF
C767 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.01fF
C768 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.03fF
C769 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C770 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C771 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C772 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C773 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C774 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.01fF
C775 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C776 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C777 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C778 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.02fF
C779 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C780 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.03fF
C781 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.55fF
C782 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C783 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C784 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.02fF
C785 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.02fF
C786 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.01fF
C787 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.01fF
C788 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VDD 0.58fF
C789 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.05fF
C790 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.08fF
C791 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C792 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C793 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C794 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C795 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C796 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.02fF
C797 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.00fF
C798 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C799 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.03fF
C800 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C801 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.60fF
C802 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C803 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C804 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C805 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C806 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C807 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C808 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.04fF
C809 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.04fF
C810 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.02fF
C811 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C812 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.00fF
C813 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C814 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C815 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C816 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C817 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.09fF
C818 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.02fF
C819 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.07fF
C820 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_3/Y 0.03fF
C821 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C822 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.00fF
C823 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C824 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.01fF
C825 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.04fF
C826 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.04fF
C827 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.00fF
C828 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.02fF
C829 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C830 p2d_b sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.14fF
C831 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2d 0.12fF
C832 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C833 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C834 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C835 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C836 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C837 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C838 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkinv_1_0/Y 0.00fF
C839 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C840 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# VDD 0.16fF
C841 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C842 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.01fF
C843 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C844 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.00fF
C845 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.01fF
C846 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.02fF
C847 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.03fF
C848 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C849 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.12fF
C850 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.07fF
C851 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.01fF
C852 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C853 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C854 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C855 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C856 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.01fF
C857 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C858 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.17fF
C859 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C860 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C861 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C862 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.04fF
C863 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C864 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.14fF
C865 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.14fF
C866 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# VDD 0.14fF
C867 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.00fF
C868 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.00fF
C869 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C870 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.03fF
C871 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.06fF
C872 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C873 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C874 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.01fF
C875 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.02fF
C876 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.01fF
C877 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C878 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.34fF
C879 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C880 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.05fF
C881 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.16fF
C882 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# VDD 0.11fF
C883 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C884 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.01fF
C885 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C886 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.00fF
C887 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.03fF
C888 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# VDD 0.30fF
C889 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.00fF
C890 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C891 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.01fF
C892 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C893 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.01fF
C894 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C895 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C896 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.02fF
C897 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.04fF
C898 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.00fF
C899 sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C900 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.03fF
C901 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C902 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.02fF
C903 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.00fF
C904 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.01fF
C905 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C906 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C907 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.01fF
C908 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.05fF
C909 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C910 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C911 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.04fF
C912 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C913 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.02fF
C914 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C915 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.02fF
C916 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.08fF
C917 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.01fF
C918 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.01fF
C919 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.01fF
C920 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.01fF
C921 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.04fF
C922 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.04fF
C923 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C924 sky130_fd_sc_hd__nand2_4_2/Y VDD 5.23fF
C925 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.00fF
C926 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.00fF
C927 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.01fF
C928 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.02fF
C929 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B 0.12fF
C930 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C931 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.04fF
C932 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.04fF
C933 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Bd_b 0.02fF
C934 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C935 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C936 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.06fF
C937 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C938 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C939 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.04fF
C940 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.04fF
C941 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C942 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.01fF
C943 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.01fF
C944 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.01fF
C945 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.02fF
C946 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C947 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C948 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C949 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C950 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.00fF
C951 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VDD 0.51fF
C952 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.02fF
C953 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_27_47# 0.08fF
C954 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C955 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.02fF
C956 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.01fF
C957 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.00fF
C958 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C959 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.02fF
C960 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C961 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.00fF
C962 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C963 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C964 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C965 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.01fF
C966 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.00fF
C967 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_3/A 0.49fF
C968 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.01fF
C969 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C970 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C971 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.10fF
C972 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C973 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.01fF
C974 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.01fF
C975 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.00fF
C976 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.02fF
C977 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C978 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C979 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.01fF
C980 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C981 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.01fF
C982 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.11fF
C983 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VDD 0.29fF
C984 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.02fF
C985 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.02fF
C986 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VDD 0.27fF
C987 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C988 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.01fF
C989 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.00fF
C990 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.02fF
C991 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.01fF
C992 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.00fF
C993 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C994 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C995 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C996 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C997 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C998 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.00fF
C999 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.02fF
C1000 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.02fF
C1001 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.11fF
C1002 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C1003 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C1004 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C1005 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C1006 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.03fF
C1007 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# VDD 0.13fF
C1008 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.57fF
C1009 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.04fF
C1010 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.05fF
C1011 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.06fF
C1012 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.03fF
C1013 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C1014 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# 0.04fF
C1015 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C1016 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.01fF
C1017 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.01fF
C1018 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C1019 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C1020 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_4/B 0.12fF
C1021 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C1022 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# VDD 0.18fF
C1023 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.09fF
C1024 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C1025 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C1026 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C1027 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.06fF
C1028 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C1029 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C1030 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C1031 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C1032 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.00fF
C1033 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C1034 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# 0.01fF
C1035 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C1036 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.03fF
C1037 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.09fF
C1038 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C1039 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C1040 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C1041 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C1042 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.01fF
C1043 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C1044 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.01fF
C1045 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C1046 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C1047 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C1048 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.02fF
C1049 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C1050 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.02fF
C1051 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C1052 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C1053 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C1054 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.00fF
C1055 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.00fF
C1056 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.03fF
C1057 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C1058 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1059 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.02fF
C1060 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C1061 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C1062 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.03fF
C1063 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.02fF
C1064 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.02fF
C1065 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C1066 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C1067 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C1068 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.00fF
C1069 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.02fF
C1070 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C1071 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.02fF
C1072 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.02fF
C1073 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C1074 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C1075 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# VDD 0.20fF
C1076 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.01fF
C1077 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.00fF
C1078 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C1079 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.02fF
C1080 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.04fF
C1081 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.04fF
C1082 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C1083 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C1084 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C1085 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# VDD 0.15fF
C1086 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C1087 VDD sky130_fd_sc_hd__mux2_1_0/X 0.62fF
C1088 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C1089 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# VDD 0.34fF
C1090 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# VDD 0.31fF
C1091 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C1092 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.02fF
C1093 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C1094 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C1095 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C1096 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.01fF
C1097 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C1098 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C1099 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C1100 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.02fF
C1101 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.02fF
C1102 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_1_1/A 0.10fF
C1103 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C1104 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C1105 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C1106 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.05fF
C1107 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.05fF
C1108 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.04fF
C1109 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.14fF
C1110 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1111 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C1112 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C1113 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C1114 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# 0.04fF
C1115 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C1116 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_2/A 0.05fF
C1117 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.84fF
C1118 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.00fF
C1119 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C1120 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C1121 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.02fF
C1122 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.01fF
C1123 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.37fF
C1124 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkinv_4_5/Y 0.08fF
C1125 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C1126 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# VDD 0.13fF
C1127 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C1128 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C1129 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.02fF
C1130 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.02fF
C1131 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C1132 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_1/B 0.00fF
C1133 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__nand2_4_0/Y 0.20fF
C1134 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C1135 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.02fF
C1136 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C1137 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.01fF
C1138 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C1139 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C1140 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C1141 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Ad_b 0.02fF
C1142 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.01fF
C1143 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.02fF
C1144 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C1145 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C1146 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.02fF
C1147 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C1148 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.00fF
C1149 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.00fF
C1150 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C1151 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.06fF
C1152 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.02fF
C1153 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.04fF
C1154 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C1155 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.03fF
C1156 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C1157 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.04fF
C1158 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C1159 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1160 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C1161 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C1162 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C1163 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.00fF
C1164 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C1165 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.02fF
C1166 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.01fF
C1167 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.00fF
C1168 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C1169 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.03fF
C1170 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkinv_4_5/Y 0.85fF
C1171 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C1172 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C1173 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.02fF
C1174 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_1_1/Y 0.12fF
C1175 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.02fF
C1176 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VDD 0.73fF
C1177 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C1178 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C1179 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VDD 0.73fF
C1180 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C1181 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C1182 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.00fF
C1183 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.00fF
C1184 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# p2_b 0.12fF
C1185 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C1186 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C1187 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.09fF
C1188 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_47# -0.00fF
C1189 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C1190 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.03fF
C1191 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.05fF
C1192 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.06fF
C1193 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C1194 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C1195 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C1196 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C1197 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C1198 p2 sky130_fd_sc_hd__clkinv_4_9/Y 0.04fF
C1199 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C1200 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C1201 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_1_2/A 0.00fF
C1202 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.12fF
C1203 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.00fF
C1204 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.00fF
C1205 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C1206 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C1207 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.01fF
C1208 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C1209 Ad Ad_b 0.60fF
C1210 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1211 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.00fF
C1212 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C1213 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1214 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.05fF
C1215 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C1216 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.03fF
C1217 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C1218 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.03fF
C1219 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.06fF
C1220 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C1221 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C1222 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C1223 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.07fF
C1224 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.03fF
C1225 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C1226 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C1227 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.03fF
C1228 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.06fF
C1229 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C1230 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.04fF
C1231 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.04fF
C1232 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C1233 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.02fF
C1234 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C1235 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C1236 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.01fF
C1237 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C1238 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.03fF
C1239 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C1240 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C1241 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C1242 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C1243 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C1244 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C1245 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C1246 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C1247 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C1248 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C1249 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C1250 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# VDD 0.12fF
C1251 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.03fF
C1252 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# VDD 0.12fF
C1253 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C1254 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C1255 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C1256 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.02fF
C1257 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.02fF
C1258 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C1259 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C1260 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.02fF
C1261 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C1262 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.00fF
C1263 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C1264 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C1265 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# VDD 0.15fF
C1266 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# VDD 0.20fF
C1267 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.01fF
C1268 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C1269 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.55fF
C1270 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.00fF
C1271 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.02fF
C1272 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.01fF
C1273 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C1274 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C1275 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.07fF
C1276 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.05fF
C1277 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.05fF
C1278 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.00fF
C1279 sky130_fd_sc_hd__dfxbp_1_1/D clk 0.04fF
C1280 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VDD 0.52fF
C1281 VDD clk 1.78fF
C1282 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.01fF
C1283 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C1284 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.00fF
C1285 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C1286 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.01fF
C1287 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C1288 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# VDD 0.33fF
C1289 A sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C1290 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.00fF
C1291 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.02fF
C1292 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C1293 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_0/Y 0.03fF
C1294 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.05fF
C1295 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.09fF
C1296 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C1297 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.02fF
C1298 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C1299 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.13fF
C1300 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C1301 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.03fF
C1302 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.01fF
C1303 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.03fF
C1304 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_4_5/Y 1.26fF
C1305 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.01fF
C1306 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.01fF
C1307 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C1308 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C1309 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C1310 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.08fF
C1311 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_8/Y 0.04fF
C1312 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C1313 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.04fF
C1314 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C1315 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C1316 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C1317 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C1318 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.02fF
C1319 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C1320 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.00fF
C1321 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.02fF
C1322 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C1323 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.01fF
C1324 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C1325 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.01fF
C1326 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.02fF
C1327 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C1328 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C1329 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.09fF
C1330 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.08fF
C1331 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.01fF
C1332 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.02fF
C1333 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.00fF
C1334 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C1335 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# 0.07fF
C1336 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.11fF
C1337 sky130_fd_sc_hd__clkinv_4_1/Y VDD 0.49fF
C1338 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.02fF
C1339 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.00fF
C1340 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.00fF
C1341 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.00fF
C1342 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.05fF
C1343 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.07fF
C1344 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.04fF
C1345 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C1346 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.01fF
C1347 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C1348 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C1349 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# VDD 0.35fF
C1350 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C1351 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.10fF
C1352 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# 0.07fF
C1353 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# 0.09fF
C1354 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.00fF
C1355 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.00fF
C1356 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.00fF
C1357 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# VDD 0.54fF
C1358 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.73fF
C1359 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.02fF
C1360 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.04fF
C1361 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.04fF
C1362 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.06fF
C1363 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.09fF
C1364 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.08fF
C1365 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C1366 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C1367 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.04fF
C1368 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.84fF
C1369 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.02fF
C1370 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C1371 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.11fF
C1372 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# 0.01fF
C1373 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C1374 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.01fF
C1375 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.01fF
C1376 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.01fF
C1377 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C1378 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C1379 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# 0.07fF
C1380 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.03fF
C1381 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.01fF
C1382 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.03fF
C1383 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C1384 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.01fF
C1385 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C1386 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.01fF
C1387 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.03fF
C1388 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.00fF
C1389 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.04fF
C1390 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.03fF
C1391 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C1392 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.09fF
C1393 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C1394 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C1395 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C1396 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.03fF
C1397 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.00fF
C1398 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C1399 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C1400 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C1401 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C1402 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C1403 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.01fF
C1404 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C1405 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.03fF
C1406 Ad_b sky130_fd_sc_hd__clkinv_4_9/Y 0.03fF
C1407 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.03fF
C1408 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.04fF
C1409 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C1410 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C1411 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.01fF
C1412 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C1413 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.05fF
C1414 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.00fF
C1415 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C1416 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.10fF
C1417 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C1418 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C1419 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.02fF
C1420 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.02fF
C1421 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.00fF
C1422 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C1423 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.00fF
C1424 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.03fF
C1425 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C1426 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.12fF
C1427 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VDD 0.68fF
C1428 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.00fF
C1429 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.00fF
C1430 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C1431 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C1432 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C1433 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C1434 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C1435 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.02fF
C1436 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.00fF
C1437 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C1438 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# VDD 0.13fF
C1439 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C1440 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.00fF
C1441 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.14fF
C1442 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C1443 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C1444 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.86fF
C1445 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C1446 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C1447 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.06fF
C1448 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C1449 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C1450 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.02fF
C1451 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.01fF
C1452 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.00fF
C1453 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.05fF
C1454 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.12fF
C1455 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.02fF
C1456 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.02fF
C1457 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# 0.06fF
C1458 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# VDD 0.14fF
C1459 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C1460 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C1461 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.00fF
C1462 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.00fF
C1463 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.00fF
C1464 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.09fF
C1465 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.01fF
C1466 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C1467 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C1468 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C1469 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0.01fF
C1470 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.02fF
C1471 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.01fF
C1472 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.01fF
C1473 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.01fF
C1474 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C1475 p1d_b p1 0.08fF
C1476 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.02fF
C1477 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# VDD 0.13fF
C1478 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.04fF
C1479 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.09fF
C1480 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_3/A 0.21fF
C1481 sky130_fd_sc_hd__nand2_4_1/Y VDD 5.73fF
C1482 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.04fF
C1483 VDD sky130_fd_sc_hd__nand2_1_2/B 1.61fF
C1484 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C1485 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.03fF
C1486 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C1487 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.01fF
C1488 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.01fF
C1489 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.02fF
C1490 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C1491 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.02fF
C1492 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C1493 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C1494 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C1495 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C1496 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.02fF
C1497 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C1498 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C1499 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.02fF
C1500 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# VDD 0.12fF
C1501 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C1502 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_1_0/B 0.00fF
C1503 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A 0.62fF
C1504 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C1505 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C1506 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.00fF
C1507 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.00fF
C1508 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.00fF
C1509 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C1510 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# VDD 0.14fF
C1511 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C1512 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C1513 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C1514 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C1515 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C1516 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C1517 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.02fF
C1518 VDD sky130_fd_sc_hd__nand2_4_2/B 0.50fF
C1519 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# VDD 0.29fF
C1520 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C1521 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C1522 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C1523 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.08fF
C1524 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.01fF
C1525 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C1526 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.14fF
C1527 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_1/A 0.18fF
C1528 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C1529 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# 0.00fF
C1530 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C1531 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.16fF
C1532 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.00fF
C1533 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C1534 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.01fF
C1535 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.02fF
C1536 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C1537 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C1538 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.02fF
C1539 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C1540 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.00fF
C1541 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.17fF
C1542 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C1543 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C1544 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C1545 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C1546 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C1547 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# 0.02fF
C1548 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# 0.01fF
C1549 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# 0.00fF
C1550 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C1551 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C1552 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C1553 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C1554 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C1555 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C1556 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.01fF
C1557 p2 sky130_fd_sc_hd__clkinv_4_5/Y 0.16fF
C1558 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.05fF
C1559 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C1560 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C1561 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__nand2_4_3/Y 0.19fF
C1562 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C1563 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.01fF
C1564 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C1565 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# VDD 0.12fF
C1566 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# VDD 0.12fF
C1567 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.06fF
C1568 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C1569 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C1570 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C1571 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C1572 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.01fF
C1573 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.07fF
C1574 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# VDD 0.09fF
C1575 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# VDD 0.09fF
C1576 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.04fF
C1577 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C1578 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C1579 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C1580 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C1581 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C1582 p2_b VDD 0.77fF
C1583 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C1584 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C1585 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.01fF
C1586 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.04fF
C1587 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Bd_b 0.05fF
C1588 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# VDD 0.31fF
C1589 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C1590 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C1591 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C1592 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.02fF
C1593 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C1594 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C1595 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C1596 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C1597 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C1598 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.02fF
C1599 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C1600 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# Bd_b 0.12fF
C1601 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.00fF
C1602 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C1603 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.11fF
C1604 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.05fF
C1605 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.02fF
C1606 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.02fF
C1607 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1608 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C1609 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C1610 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C1611 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.12fF
C1612 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C1613 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C1614 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.03fF
C1615 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C1616 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C1617 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# 0.00fF
C1618 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# 0.00fF
C1619 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# 0.00fF
C1620 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C1621 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C1622 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.00fF
C1623 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.01fF
C1624 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.21fF
C1625 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# 0.02fF
C1626 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# 0.02fF
C1627 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C1628 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.06fF
C1629 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.02fF
C1630 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.02fF
C1631 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C1632 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.09fF
C1633 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.00fF
C1634 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C1635 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.02fF
C1636 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.00fF
C1637 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C1638 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C1639 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C1640 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.01fF
C1641 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.02fF
C1642 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C1643 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__nand2_1_0/A 0.10fF
C1644 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C1645 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C1646 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C1647 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C1648 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C1649 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.03fF
C1650 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C1651 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.02fF
C1652 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.06fF
C1653 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C1654 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C1655 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.03fF
C1656 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.11fF
C1657 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.06fF
C1658 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C1659 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C1660 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C1661 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.02fF
C1662 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.01fF
C1663 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.00fF
C1664 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C1665 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.03fF
C1666 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C1667 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C1668 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.01fF
C1669 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.02fF
C1670 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C1671 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C1672 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.03fF
C1673 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C1674 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C1675 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C1676 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C1677 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C1678 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C1679 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C1680 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C1681 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.16fF
C1682 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.03fF
C1683 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.03fF
C1684 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.06fF
C1685 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.08fF
C1686 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C1687 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# VDD 0.14fF
C1688 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1689 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.00fF
C1690 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.08fF
C1691 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C1692 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.03fF
C1693 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.00fF
C1694 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C1695 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.02fF
C1696 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C1697 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C1698 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C1699 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C1700 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C1701 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C1702 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.01fF
C1703 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.02fF
C1704 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.05fF
C1705 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.05fF
C1706 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C1707 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.05fF
C1708 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.00fF
C1709 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.02fF
C1710 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C1711 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/A 0.46fF
C1712 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.08fF
C1713 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C1714 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.01fF
C1715 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C1716 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.01fF
C1717 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C1718 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C1719 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.00fF
C1720 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.00fF
C1721 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C1722 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C1723 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VDD 0.52fF
C1724 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C1725 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C1726 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.04fF
C1727 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.06fF
C1728 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.01fF
C1729 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.01fF
C1730 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C1731 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C1732 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C1733 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.01fF
C1734 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.03fF
C1735 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.01fF
C1736 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C1737 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C1738 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C1739 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C1740 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C1741 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C1742 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# 0.00fF
C1743 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C1744 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.02fF
C1745 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.02fF
C1746 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.02fF
C1747 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C1748 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C1749 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.02fF
C1750 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.00fF
C1751 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.00fF
C1752 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C1753 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C1754 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.02fF
C1755 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.00fF
C1756 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.03fF
C1757 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C1758 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C1759 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.02fF
C1760 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C1761 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C1762 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C1763 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.01fF
C1764 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.02fF
C1765 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.04fF
C1766 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.04fF
C1767 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C1768 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C1769 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.01fF
C1770 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# VDD 0.17fF
C1771 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C1772 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C1773 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.03fF
C1774 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.11fF
C1775 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C1776 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C1777 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C1778 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C1779 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C1780 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C1781 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.03fF
C1782 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# VDD 0.30fF
C1783 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C1784 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1785 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.02fF
C1786 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C1787 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C1788 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.03fF
C1789 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C1790 sky130_fd_sc_hd__dfxbp_1_0/Q_N Bd_b 0.01fF
C1791 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C1792 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.00fF
C1793 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.02fF
C1794 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.02fF
C1795 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C1796 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C1797 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C1798 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C1799 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C1800 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.09fF
C1801 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.08fF
C1802 Ad_b sky130_fd_sc_hd__clkinv_4_5/Y 0.31fF
C1803 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.02fF
C1804 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.17fF
C1805 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# p2_b 0.15fF
C1806 p2d sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.15fF
C1807 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C1808 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.00fF
C1809 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.00fF
C1810 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C1811 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.04fF
C1812 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.04fF
C1813 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.07fF
C1814 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.04fF
C1815 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.04fF
C1816 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.02fF
C1817 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.01fF
C1818 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.08fF
C1819 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.00fF
C1820 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.00fF
C1821 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.01fF
C1822 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.01fF
C1823 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C1824 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C1825 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C1826 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C1827 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C1828 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# B 0.02fF
C1829 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.08fF
C1830 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C1831 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C1832 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C1833 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C1834 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C1835 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C1836 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C1837 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# VDD 0.44fF
C1838 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C1839 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.04fF
C1840 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.04fF
C1841 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.07fF
C1842 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.08fF
C1843 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.01fF
C1844 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.59fF
C1845 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C1846 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C1847 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.02fF
C1848 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C1849 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.02fF
C1850 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C1851 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.04fF
C1852 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.04fF
C1853 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C1854 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.01fF
C1855 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C1856 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C1857 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C1858 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.02fF
C1859 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.02fF
C1860 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.04fF
C1861 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.04fF
C1862 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.01fF
C1863 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C1864 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C1865 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.02fF
C1866 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.02fF
C1867 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.01fF
C1868 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C1869 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C1870 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C1871 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C1872 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C1873 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C1874 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C1875 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C1876 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.05fF
C1877 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C1878 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C1879 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C1880 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C1881 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VDD 0.53fF
C1882 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.06fF
C1883 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.05fF
C1884 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C1885 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C1886 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C1887 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C1888 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.00fF
C1889 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VDD 0.53fF
C1890 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.05fF
C1891 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.05fF
C1892 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C1893 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C1894 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# 0.00fF
C1895 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# 0.00fF
C1896 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C1897 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.01fF
C1898 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.01fF
C1899 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.01fF
C1900 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.02fF
C1901 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.03fF
C1902 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C1903 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C1904 sky130_fd_sc_hd__clkinv_1_2/Y sky130_fd_sc_hd__clkinv_4_7/A 0.36fF
C1905 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VDD 0.35fF
C1906 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C1907 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.01fF
C1908 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.22fF
C1909 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# 0.01fF
C1910 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# 0.01fF
C1911 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.06fF
C1912 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C1913 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.03fF
C1914 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.03fF
C1915 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C1916 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.04fF
C1917 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.04fF
C1918 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# VDD 0.13fF
C1919 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.05fF
C1920 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.03fF
C1921 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.01fF
C1922 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.03fF
C1923 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.11fF
C1924 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C1925 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C1926 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.00fF
C1927 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C1928 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C1929 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.00fF
C1930 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.00fF
C1931 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# 0.00fF
C1932 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.00fF
C1933 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C1934 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C1935 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C1936 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.03fF
C1937 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C1938 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.03fF
C1939 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.84fF
C1940 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.00fF
C1941 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.27fF
C1942 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C1943 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C1944 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C1945 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.02fF
C1946 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.01fF
C1947 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.04fF
C1948 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.04fF
C1949 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C1950 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.14fF
C1951 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# A 0.02fF
C1952 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.04fF
C1953 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C1954 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C1955 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C1956 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.02fF
C1957 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/B 0.04fF
C1958 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C1959 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.02fF
C1960 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.02fF
C1961 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.17fF
C1962 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C1963 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.03fF
C1964 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# VDD 0.14fF
C1965 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.84fF
C1966 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.13fF
C1967 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.04fF
C1968 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.04fF
C1969 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.06fF
C1970 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C1971 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C1972 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C1973 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.04fF
C1974 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.01fF
C1975 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.24fF
C1976 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# VDD 0.18fF
C1977 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.06fF
C1978 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C1979 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C1980 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# VDD 0.33fF
C1981 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.04fF
C1982 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.04fF
C1983 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.02fF
C1984 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.01fF
C1985 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1986 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.01fF
C1987 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C1988 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C1989 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C1990 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C1991 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.02fF
C1992 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C1993 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C1994 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C1995 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.02fF
C1996 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C1997 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C1998 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# VDD 0.31fF
C1999 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.03fF
C2000 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# VDD 0.28fF
C2001 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/A 0.03fF
C2002 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C2003 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C2004 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.00fF
C2005 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C2006 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# 0.00fF
C2007 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C2008 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.31fF
C2009 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C2010 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkinv_4_5/Y 0.85fF
C2011 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# 0.11fF
C2012 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.01fF
C2013 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# 0.01fF
C2014 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.08fF
C2015 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.00fF
C2016 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C2017 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.02fF
C2018 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.01fF
C2019 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.01fF
C2020 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.01fF
C2021 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.02fF
C2022 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.02fF
C2023 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C2024 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.02fF
C2025 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.04fF
C2026 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C2027 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.02fF
C2028 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VDD 0.68fF
C2029 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/B 0.11fF
C2030 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C2031 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C2032 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C2033 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C2034 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.09fF
C2035 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.00fF
C2036 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.03fF
C2037 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C2038 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C2039 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C2040 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C2041 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.06fF
C2042 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C2043 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.01fF
C2044 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.12fF
C2045 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.01fF
C2046 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C2047 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.01fF
C2048 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.01fF
C2049 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.03fF
C2050 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VDD 0.35fF
C2051 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.01fF
C2052 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C2053 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C2054 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C2055 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.13fF
C2056 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.02fF
C2057 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.02fF
C2058 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.03fF
C2059 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C2060 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C2061 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C2062 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C2063 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.02fF
C2064 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.00fF
C2065 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.12fF
C2066 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.12fF
C2067 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C2068 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.01fF
C2069 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C2070 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C2071 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C2072 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C2073 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C2074 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C2075 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C2076 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C2077 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.14fF
C2078 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.04fF
C2079 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C2080 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C2081 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C2082 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C2083 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.04fF
C2084 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.04fF
C2085 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VDD 6.88fF
C2086 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.01fF
C2087 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C2088 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.02fF
C2089 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0.00fF
C2090 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.02fF
C2091 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C2092 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C2093 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.03fF
C2094 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C2095 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C2096 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C2097 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C2098 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C2099 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.01fF
C2100 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.01fF
C2101 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.03fF
C2102 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.00fF
C2103 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C2104 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C2105 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C2106 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VDD 0.63fF
C2107 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C2108 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.00fF
C2109 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C2110 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C2111 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C2112 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.03fF
C2113 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C2114 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C2115 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C2116 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C2117 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.01fF
C2118 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.05fF
C2119 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.04fF
C2120 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.03fF
C2121 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.02fF
C2122 VDD sky130_fd_sc_hd__clkinv_1_1/Y 0.40fF
C2123 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# VDD 0.14fF
C2124 VDD sky130_fd_sc_hd__clkinv_1_0/Y 0.26fF
C2125 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.03fF
C2126 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.31fF
C2127 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C2128 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C2129 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C2130 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# VDD 0.30fF
C2131 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C2132 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C2133 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C2134 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.01fF
C2135 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C2136 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C2137 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C2138 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.02fF
C2139 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C2140 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C2141 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C2142 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# VDD 0.31fF
C2143 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.03fF
C2144 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.03fF
C2145 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.06fF
C2146 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C2147 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C2148 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.02fF
C2149 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C2150 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.00fF
C2151 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C2152 VDD sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.30fF
C2153 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.02fF
C2154 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C2155 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.06fF
C2156 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C2157 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C2158 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.00fF
C2159 p2d_b p2 0.09fF
C2160 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C2161 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.01fF
C2162 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C2163 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C2164 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C2165 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C2166 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C2167 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.00fF
C2168 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C2169 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.01fF
C2170 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C2171 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C2172 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C2173 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# VDD 0.14fF
C2174 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.00fF
C2175 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.00fF
C2176 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.04fF
C2177 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C2178 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.01fF
C2179 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C2180 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.00fF
C2181 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.00fF
C2182 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C2183 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.04fF
C2184 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.02fF
C2185 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C2186 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C2187 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C2188 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C2189 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# VDD 0.17fF
C2190 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C2191 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# VDD 0.20fF
C2192 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.01fF
C2193 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.03fF
C2194 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C2195 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C2196 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C2197 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C2198 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.02fF
C2199 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.07fF
C2200 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C2201 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C2202 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C2203 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C2204 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C2205 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# VDD 0.28fF
C2206 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C2207 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# VDD 0.25fF
C2208 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C2209 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C2210 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C2211 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C2212 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.04fF
C2213 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C2214 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C2215 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C2216 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C2217 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# 0.09fF
C2218 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.05fF
C2219 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C2220 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C2221 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.02fF
C2222 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.00fF
C2223 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.01fF
C2224 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C2225 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_1_0/A 0.01fF
C2226 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C2227 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C2228 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C2229 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C2230 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.00fF
C2231 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C2232 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C2233 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C2234 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C2235 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C2236 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.02fF
C2237 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.02fF
C2238 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C2239 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C2240 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# VDD 0.25fF
C2241 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.00fF
C2242 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.00fF
C2243 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Bd_b 0.03fF
C2244 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C2245 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C2246 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.00fF
C2247 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.00fF
C2248 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.00fF
C2249 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.00fF
C2250 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.00fF
C2251 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.01fF
C2252 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.02fF
C2253 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.02fF
C2254 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C2255 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.00fF
C2256 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C2257 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C2258 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C2259 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C2260 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C2261 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C2262 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.01fF
C2263 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.03fF
C2264 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.03fF
C2265 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C2266 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C2267 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C2268 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.01fF
C2269 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C2270 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.00fF
C2271 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.01fF
C2272 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.01fF
C2273 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C2274 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C2275 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.01fF
C2276 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.02fF
C2277 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C2278 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.00fF
C2279 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.02fF
C2280 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C2281 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.06fF
C2282 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C2283 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C2284 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C2285 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C2286 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.11fF
C2287 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C2288 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C2289 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.00fF
C2290 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C2291 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C2292 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A VDD 0.57fF
C2293 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VDD 6.52fF
C2294 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.04fF
C2295 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VDD 0.53fF
C2296 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.00fF
C2297 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C2298 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C2299 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.05fF
C2300 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.02fF
C2301 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C2302 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_1_4/B 0.11fF
C2303 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# VDD 0.29fF
C2304 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C2305 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VDD 0.22fF
C2306 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.04fF
C2307 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C2308 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.01fF
C2309 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.07fF
C2310 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.08fF
C2311 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C2312 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.01fF
C2313 p2d VDD 1.53fF
C2314 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.01fF
C2315 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.10fF
C2316 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.04fF
C2317 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.04fF
C2318 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C2319 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C2320 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.01fF
C2321 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C2322 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C2323 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.08fF
C2324 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C2325 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C2326 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.01fF
C2327 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.09fF
C2328 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.02fF
C2329 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.01fF
C2330 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C2331 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C2332 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C2333 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.06fF
C2334 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.06fF
C2335 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.01fF
C2336 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1_b 0.06fF
C2337 p1d_b sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.06fF
C2338 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C2339 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C2340 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C2341 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C2342 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.14fF
C2343 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C2344 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C2345 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C2346 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.03fF
C2347 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.02fF
C2348 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.02fF
C2349 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C2350 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C2351 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C2352 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C2353 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.01fF
C2354 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.02fF
C2355 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.04fF
C2356 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.04fF
C2357 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# VDD 0.14fF
C2358 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.08fF
C2359 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# VDD 0.15fF
C2360 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.01fF
C2361 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.01fF
C2362 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.03fF
C2363 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.01fF
C2364 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.01fF
C2365 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# VDD 0.33fF
C2366 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.01fF
C2367 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.00fF
C2368 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C2369 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C2370 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C2371 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C2372 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C2373 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# VDD 0.17fF
C2374 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C2375 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.00fF
C2376 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.00fF
C2377 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.01fF
C2378 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C2379 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# VDD 0.24fF
C2380 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C2381 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.03fF
C2382 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C2383 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.03fF
C2384 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C2385 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VDD 0.53fF
C2386 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C2387 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C2388 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C2389 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C2390 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.02fF
C2391 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C2392 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.05fF
C2393 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.04fF
C2394 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.09fF
C2395 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.05fF
C2396 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C2397 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C2398 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C2399 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C2400 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C2401 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C2402 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.02fF
C2403 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C2404 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.01fF
C2405 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C2406 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C2407 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.00fF
C2408 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.02fF
C2409 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C2410 B_b Bd_b 0.20fF
C2411 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.09fF
C2412 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.01fF
C2413 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C2414 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.11fF
C2415 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# 0.07fF
C2416 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.04fF
C2417 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.08fF
C2418 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.00fF
C2419 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.00fF
C2420 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C2421 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C2422 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.04fF
C2423 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.01fF
C2424 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# VDD 0.20fF
C2425 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.11fF
C2426 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.03fF
C2427 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C2428 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C2429 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VDD 0.54fF
C2430 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# 0.06fF
C2431 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.00fF
C2432 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.02fF
C2433 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VDD 0.33fF
C2434 VDD sky130_fd_sc_hd__nand2_1_3/A 4.52fF
C2435 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.05fF
C2436 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.02fF
C2437 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# 0.01fF
C2438 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C2439 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.00fF
C2440 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.02fF
C2441 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.05fF
C2442 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.00fF
C2443 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C2444 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C2445 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.01fF
C2446 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.01fF
C2447 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.01fF
C2448 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C2449 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# VDD 0.32fF
C2450 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.01fF
C2451 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.00fF
C2452 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C2453 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.03fF
C2454 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.01fF
C2455 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.02fF
C2456 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.02fF
C2457 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C2458 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# 0.06fF
C2459 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.00fF
C2460 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C2461 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.01fF
C2462 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.01fF
C2463 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.07fF
C2464 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C2465 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C2466 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C2467 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C2468 p2 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.02fF
C2469 sky130_fd_sc_hd__clkinv_1_3/A VDD 4.38fF
C2470 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.04fF
C2471 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.01fF
C2472 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# p2d 0.02fF
C2473 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Ad_b 0.12fF
C2474 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.04fF
C2475 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C2476 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.01fF
C2477 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C2478 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C2479 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.09fF
C2480 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C2481 Bd_b sky130_fd_sc_hd__clkinv_4_9/Y 0.00fF
C2482 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C2483 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VDD 0.74fF
C2484 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C2485 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C2486 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C2487 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.00fF
C2488 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.04fF
C2489 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C2490 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.01fF
C2491 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.04fF
C2492 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.04fF
C2493 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.00fF
C2494 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.00fF
C2495 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.00fF
C2496 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C2497 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C2498 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.01fF
C2499 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C2500 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.01fF
C2501 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C2502 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C2503 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C2504 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.14fF
C2505 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VDD 0.34fF
C2506 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C2507 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C2508 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.57fF
C2509 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.07fF
C2510 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C2511 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C2512 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.01fF
C2513 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.01fF
C2514 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C2515 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C2516 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.07fF
C2517 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# 0.01fF
C2518 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C2519 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.06fF
C2520 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C2521 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.07fF
C2522 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.02fF
C2523 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C2524 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C2525 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C2526 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.05fF
C2527 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.02fF
C2528 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.02fF
C2529 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C2530 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.02fF
C2531 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# 0.09fF
C2532 VDD sky130_fd_sc_hd__nand2_1_2/A -0.72fF
C2533 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.02fF
C2534 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.02fF
C2535 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.00fF
C2536 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C2537 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.03fF
C2538 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C2539 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.02fF
C2540 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C2541 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.04fF
C2542 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C2543 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.00fF
C2544 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C2545 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.02fF
C2546 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.07fF
C2547 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.02fF
C2548 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.04fF
C2549 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C2550 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C2551 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.04fF
C2552 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.09fF
C2553 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.04fF
C2554 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.04fF
C2555 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C2556 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.00fF
C2557 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VDD 0.52fF
C2558 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.03fF
C2559 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.00fF
C2560 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.00fF
C2561 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C2562 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2563 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# VDD 0.12fF
C2564 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C2565 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.01fF
C2566 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.00fF
C2567 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C2568 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C2569 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C2570 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C2571 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C2572 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C2573 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.02fF
C2574 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# VDD 0.15fF
C2575 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0.09fF
C2576 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C2577 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# 0.01fF
C2578 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C2579 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C2580 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C2581 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C2582 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.03fF
C2583 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# VDD 0.23fF
C2584 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C2585 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.15fF
C2586 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C2587 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C2588 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.02fF
C2589 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.02fF
C2590 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C2591 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C2592 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.14fF
C2593 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C2594 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C2595 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C2596 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# 0.01fF
C2597 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# 0.01fF
C2598 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C2599 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C2600 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C2601 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.00fF
C2602 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C2603 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.00fF
C2604 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C2605 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C2606 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkinv_4_1/A 0.08fF
C2607 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C2608 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C2609 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C2610 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C2611 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C2612 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.01fF
C2613 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.07fF
C2614 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C2615 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.02fF
C2616 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.02fF
C2617 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C2618 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.08fF
C2619 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C2620 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# VDD 0.12fF
C2621 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C2622 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C2623 VDD A_b 0.82fF
C2624 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.03fF
C2625 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C2626 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C2627 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.01fF
C2628 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C2629 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# VDD 0.18fF
C2630 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.08fF
C2631 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__nand2_4_2/A 2.12fF
C2632 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C2633 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.01fF
C2634 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C2635 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.09fF
C2636 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C2637 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C2638 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C2639 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C2640 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.06fF
C2641 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C2642 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.01fF
C2643 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.00fF
C2644 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C2645 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C2646 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# VDD 0.33fF
C2647 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C2648 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C2649 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.03fF
C2650 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.02fF
C2651 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.03fF
C2652 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.03fF
C2653 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.04fF
C2654 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.04fF
C2655 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C2656 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkinv_4_5/Y 0.87fF
C2657 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C2658 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# B_b 0.15fF
C2659 Bd sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.15fF
C2660 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C2661 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# 0.02fF
C2662 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C2663 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C2664 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.02fF
C2665 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# 0.00fF
C2666 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# 0.00fF
C2667 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C2668 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.01fF
C2669 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.03fF
C2670 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.11fF
C2671 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.05fF
C2672 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.05fF
C2673 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.14fF
C2674 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.03fF
C2675 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# VDD 0.30fF
C2676 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.06fF
C2677 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.08fF
C2678 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.01fF
C2679 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C2680 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.04fF
C2681 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.04fF
C2682 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C2683 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# Ad_b 0.06fF
C2684 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkinv_4_3/Y 0.04fF
C2685 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C2686 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C2687 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C2688 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_3/A 0.47fF
C2689 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C2690 p1d_b sky130_fd_sc_hd__clkbuf_16_12/a_110_47# 0.02fF
C2691 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p2d_b 0.02fF
C2692 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.04fF
C2693 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.08fF
C2694 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.04fF
C2695 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C2696 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C2697 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.01fF
C2698 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.03fF
C2699 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.31fF
C2700 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.09fF
C2701 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C2702 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.02fF
C2703 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.02fF
C2704 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.06fF
C2705 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.02fF
C2706 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C2707 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C2708 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.11fF
C2709 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C2710 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C2711 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.02fF
C2712 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C2713 p1 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.12fF
C2714 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1_b 0.12fF
C2715 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/A 0.62fF
C2716 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.04fF
C2717 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.04fF
C2718 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C2719 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C2720 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2721 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C2722 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C2723 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C2724 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.02fF
C2725 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.02fF
C2726 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.02fF
C2727 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C2728 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.01fF
C2729 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.03fF
C2730 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C2731 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.01fF
C2732 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C2733 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C2734 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2735 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2736 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C2737 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C2738 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C2739 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C2740 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C2741 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C2742 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.00fF
C2743 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C2744 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.03fF
C2745 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C2746 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.03fF
C2747 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.13fF
C2748 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.00fF
C2749 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C2750 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.00fF
C2751 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C2752 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C2753 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C2754 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.03fF
C2755 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2756 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.02fF
C2757 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y -0.01fF
C2758 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2759 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C2760 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C2761 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.00fF
C2762 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C2763 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C2764 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.02fF
C2765 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C2766 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.02fF
C2767 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.02fF
C2768 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C2769 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C2770 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C2771 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C2772 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C2773 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C2774 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.01fF
C2775 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.02fF
C2776 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C2777 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C2778 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C2779 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C2780 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.01fF
C2781 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.02fF
C2782 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.06fF
C2783 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C2784 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C2785 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.00fF
C2786 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C2787 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.03fF
C2788 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C2789 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# -0.08fF
C2790 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.03fF
C2791 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C2792 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C2793 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.02fF
C2794 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C2795 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.00fF
C2796 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C2797 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.04fF
C2798 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.10fF
C2799 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.03fF
C2800 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C2801 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C2802 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C2803 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C2804 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C2805 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C2806 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.03fF
C2807 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.01fF
C2808 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.03fF
C2809 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C2810 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C2811 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.01fF
C2812 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.01fF
C2813 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VDD 0.51fF
C2814 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__nand2_4_3/Y 0.04fF
C2815 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C2816 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C2817 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C2818 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C2819 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.03fF
C2820 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.09fF
C2821 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.02fF
C2822 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C2823 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C2824 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkinv_1_2/Y 0.06fF
C2825 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.08fF
C2826 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.06fF
C2827 sky130_fd_sc_hd__mux2_1_0/X Ad_b 0.00fF
C2828 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C2829 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C2830 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.00fF
C2831 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C2832 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C2833 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C2834 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C2835 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.03fF
C2836 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.05fF
C2837 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# VDD 0.14fF
C2838 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C2839 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C2840 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2841 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C2842 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2843 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.08fF
C2844 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C2845 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C2846 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.02fF
C2847 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C2848 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C2849 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C2850 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.01fF
C2851 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.03fF
C2852 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.70fF
C2853 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C2854 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C2855 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C2856 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C2857 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C2858 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C2859 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# VDD 0.16fF
C2860 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.03fF
C2861 sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.11fF
C2862 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.02fF
C2863 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# 0.00fF
C2864 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C2865 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C2866 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C2867 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C2868 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C2869 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.01fF
C2870 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.09fF
C2871 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C2872 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C2873 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.02fF
C2874 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C2875 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C2876 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.05fF
C2877 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.05fF
C2878 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.03fF
C2879 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C2880 Bd_b sky130_fd_sc_hd__clkinv_4_5/Y 0.46fF
C2881 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.14fF
C2882 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.09fF
C2883 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C2884 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.00fF
C2885 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C2886 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C2887 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C2888 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C2889 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C2890 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.01fF
C2891 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.01fF
C2892 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C2893 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.01fF
C2894 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C2895 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C2896 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.00fF
C2897 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.02fF
C2898 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.02fF
C2899 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C2900 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C2901 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C2902 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C2903 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C2904 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C2905 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.01fF
C2906 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C2907 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C2908 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.09fF
C2909 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C2910 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# VDD 0.16fF
C2911 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.01fF
C2912 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C2913 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C2914 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C2915 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.02fF
C2916 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.01fF
C2917 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C2918 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C2919 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.04fF
C2920 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.04fF
C2921 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# 0.04fF
C2922 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# 0.04fF
C2923 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.09fF
C2924 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# VDD 0.32fF
C2925 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C2926 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.03fF
C2927 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C2928 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.02fF
C2929 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C2930 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.51fF
C2931 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C2932 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C2933 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.01fF
C2934 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.02fF
C2935 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C2936 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.01fF
C2937 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C2938 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C2939 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C2940 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkinv_4_1/A 1.80fF
C2941 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.02fF
C2942 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.02fF
C2943 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.01fF
C2944 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.03fF
C2945 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.02fF
C2946 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.02fF
C2947 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C2948 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.03fF
C2949 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C2950 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.15fF
C2951 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C2952 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.04fF
C2953 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.01fF
C2954 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.02fF
C2955 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C2956 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.08fF
C2957 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.16fF
C2958 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_2/B 0.07fF
C2959 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A VDD 0.56fF
C2960 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.04fF
C2961 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.05fF
C2962 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C2963 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C2964 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.06fF
C2965 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.03fF
C2966 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C2967 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C2968 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C2969 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C2970 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C2971 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C2972 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.04fF
C2973 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.10fF
C2974 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C2975 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C2976 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C2977 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.02fF
C2978 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.02fF
C2979 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C2980 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C2981 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C2982 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# 0.00fF
C2983 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# 0.00fF
C2984 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# 0.00fF
C2985 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.01fF
C2986 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.06fF
C2987 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C2988 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VDD 0.21fF
C2989 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.01fF
C2990 sky130_fd_sc_hd__clkinv_4_8/Y VDD 1.51fF
C2991 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.41fF
C2992 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.00fF
C2993 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.00fF
C2994 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C2995 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C2996 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C2997 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C2998 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.06fF
C2999 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C3000 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.01fF
C3001 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.01fF
C3002 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C3003 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.06fF
C3004 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C3005 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C3006 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.00fF
C3007 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.04fF
C3008 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C3009 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C3010 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C3011 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.02fF
C3012 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# 0.02fF
C3013 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C3014 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.04fF
C3015 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.00fF
C3016 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C3017 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C3018 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.04fF
C3019 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.01fF
C3020 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.11fF
C3021 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C3022 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C3023 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C3024 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.03fF
C3025 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C3026 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.01fF
C3027 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.00fF
C3028 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.00fF
C3029 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.33fF
C3030 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.02fF
C3031 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C3032 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C3033 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.00fF
C3034 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.30fF
C3035 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.14fF
C3036 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkinv_4_1/A 0.12fF
C3037 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.03fF
C3038 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.03fF
C3039 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.09fF
C3040 p2 sky130_fd_sc_hd__nand2_4_1/Y 0.00fF
C3041 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C3042 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C3043 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C3044 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C3045 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3046 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C3047 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C3048 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C3049 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C3050 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C3051 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C3052 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C3053 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C3054 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.00fF
C3055 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.00fF
C3056 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.12fF
C3057 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.01fF
C3058 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.03fF
C3059 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C3060 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.00fF
C3061 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# VDD 0.14fF
C3062 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.04fF
C3063 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.04fF
C3064 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.03fF
C3065 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.14fF
C3066 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.01fF
C3067 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.02fF
C3068 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.00fF
C3069 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# VDD 0.15fF
C3070 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C3071 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C3072 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C3073 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C3074 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C3075 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C3076 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C3077 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C3078 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C3079 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C3080 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.02fF
C3081 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C3082 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.00fF
C3083 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# VDD 0.14fF
C3084 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.03fF
C3085 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C3086 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# VDD 0.15fF
C3087 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/A 0.01fF
C3088 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# VDD 0.28fF
C3089 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.04fF
C3090 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.00fF
C3091 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C3092 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.03fF
C3093 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# VDD 0.20fF
C3094 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.01fF
C3095 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.01fF
C3096 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C3097 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C3098 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C3099 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C3100 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.02fF
C3101 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C3102 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.00fF
C3103 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.02fF
C3104 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.02fF
C3105 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# 0.00fF
C3106 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__nand2_4_2/Y 0.04fF
C3107 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.02fF
C3108 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.02fF
C3109 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.01fF
C3110 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.84fF
C3111 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C3112 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C3113 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C3114 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C3115 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.02fF
C3116 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.01fF
C3117 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C3118 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C3119 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C3120 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C3121 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C3122 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C3123 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C3124 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.07fF
C3125 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C3126 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C3127 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_4/Y 0.04fF
C3128 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.03fF
C3129 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.08fF
C3130 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VDD 0.07fF
C3131 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.01fF
C3132 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C3133 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C3134 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C3135 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__nand2_4_0/Y 0.16fF
C3136 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.07fF
C3137 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C3138 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_3/A 0.25fF
C3139 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C3140 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3141 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C3142 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C3143 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C3144 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C3145 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.00fF
C3146 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.10fF
C3147 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C3148 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C3149 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C3150 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C3151 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C3152 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C3153 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C3154 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C3155 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C3156 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C3157 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C3158 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C3159 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.04fF
C3160 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.01fF
C3161 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.00fF
C3162 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C3163 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C3164 p2_b p2 0.47fF
C3165 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C3166 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.04fF
C3167 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.04fF
C3168 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A VDD 0.58fF
C3169 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C3170 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.01fF
C3171 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.01fF
C3172 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.04fF
C3173 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.03fF
C3174 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C3175 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.09fF
C3176 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# 0.09fF
C3177 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C3178 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.02fF
C3179 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__nand2_1_1/B 0.03fF
C3180 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C3181 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.01fF
C3182 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C3183 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C3184 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C3185 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C3186 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C3187 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C3188 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C3189 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C3190 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C3191 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.01fF
C3192 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.07fF
C3193 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C3194 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.04fF
C3195 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.04fF
C3196 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VDD 0.53fF
C3197 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.04fF
C3198 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.01fF
C3199 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C3200 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C3201 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.01fF
C3202 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# 0.12fF
C3203 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.05fF
C3204 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# VDD 0.18fF
C3205 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.11fF
C3206 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C3207 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C3208 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.08fF
C3209 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.04fF
C3210 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.06fF
C3211 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.03fF
C3212 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.05fF
C3213 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3214 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C3215 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C3216 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C3217 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C3218 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.00fF
C3219 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.03fF
C3220 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C3221 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.00fF
C3222 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# VDD 0.17fF
C3223 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C3224 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C3225 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C3226 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C3227 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C3228 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.00fF
C3229 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.00fF
C3230 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C3231 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C3232 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C3233 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C3234 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkinv_4_5/Y 0.08fF
C3235 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.09fF
C3236 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C3237 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# VDD 0.23fF
C3238 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.00fF
C3239 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.01fF
C3240 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C3241 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C3242 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C3243 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.01fF
C3244 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C3245 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C3246 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C3247 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.00fF
C3248 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.01fF
C3249 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.02fF
C3250 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C3251 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C3252 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C3253 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.02fF
C3254 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.02fF
C3255 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C3256 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C3257 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C3258 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C3259 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# VDD 0.14fF
C3260 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.06fF
C3261 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# VDD 0.15fF
C3262 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.01fF
C3263 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C3264 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C3265 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C3266 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.01fF
C3267 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C3268 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C3269 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C3270 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.05fF
C3271 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.05fF
C3272 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C3273 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C3274 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C3275 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# VDD 0.12fF
C3276 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C3277 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# VDD 0.15fF
C3278 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C3279 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C3280 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C3281 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C3282 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C3283 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C3284 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C3285 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C3286 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.05fF
C3287 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.05fF
C3288 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C3289 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C3290 p1d_b p1d 0.47fF
C3291 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C3292 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# VDD 0.34fF
C3293 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C3294 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.01fF
C3295 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.01fF
C3296 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.01fF
C3297 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C3298 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.01fF
C3299 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C3300 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.05fF
C3301 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.05fF
C3302 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/A 0.45fF
C3303 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C3304 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.01fF
C3305 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C3306 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C3307 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C3308 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C3309 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.05fF
C3310 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.05fF
C3311 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C3312 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C3313 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.03fF
C3314 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C3315 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C3316 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C3317 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.00fF
C3318 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C3319 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.00fF
C3320 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C3321 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C3322 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.00fF
C3323 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# VDD 0.15fF
C3324 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.50fF
C3325 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.02fF
C3326 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.00fF
C3327 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C3328 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.01fF
C3329 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.01fF
C3330 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.00fF
C3331 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.00fF
C3332 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.00fF
C3333 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.00fF
C3334 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.00fF
C3335 sky130_fd_sc_hd__nand2_4_1/Y Ad_b 0.00fF
C3336 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C3337 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C3338 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C3339 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C3340 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C3341 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C3342 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.01fF
C3343 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.02fF
C3344 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C3345 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.01fF
C3346 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C3347 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.02fF
C3348 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.02fF
C3349 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C3350 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.02fF
C3351 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.05fF
C3352 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.03fF
C3353 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.01fF
C3354 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.06fF
C3355 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C3356 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C3357 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C3358 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.02fF
C3359 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# A_b 0.09fF
C3360 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.01fF
C3361 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.00fF
C3362 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.00fF
C3363 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.05fF
C3364 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.02fF
C3365 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.01fF
C3366 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C3367 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C3368 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C3369 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.00fF
C3370 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C3371 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C3372 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C3373 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.03fF
C3374 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.04fF
C3375 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C3376 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C3377 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C3378 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_1/A 2.16fF
C3379 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C3380 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C3381 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.03fF
C3382 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C3383 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C3384 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# VDD 0.15fF
C3385 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.01fF
C3386 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3387 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3388 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/a_27_47# 0.00fF
C3389 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VDD 0.11fF
C3390 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.08fF
C3391 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.06fF
C3392 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.02fF
C3393 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C3394 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.12fF
C3395 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# A 0.04fF
C3396 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C3397 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.11fF
C3398 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C3399 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C3400 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.02fF
C3401 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.00fF
C3402 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.00fF
C3403 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.31fF
C3404 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_1/Y 0.73fF
C3405 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.01fF
C3406 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C3407 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.02fF
C3408 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.00fF
C3409 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.03fF
C3410 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C3411 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C3412 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C3413 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkinv_4_7/A 0.05fF
C3414 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C3415 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C3416 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.00fF
C3417 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.00fF
C3418 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C3419 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C3420 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C3421 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.01fF
C3422 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.02fF
C3423 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.00fF
C3424 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C3425 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C3426 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C3427 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.11fF
C3428 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.02fF
C3429 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.02fF
C3430 sky130_fd_sc_hd__mux2_1_0/a_439_47# Ad_b 0.02fF
C3431 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C3432 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C3433 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C3434 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C3435 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_1_1/A 0.03fF
C3436 VDD sky130_fd_sc_hd__clkinv_4_7/A 3.99fF
C3437 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C3438 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C3439 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.00fF
C3440 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C3441 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C3442 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C3443 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C3444 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.01fF
C3445 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C3446 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# 0.09fF
C3447 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C3448 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C3449 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.01fF
C3450 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.02fF
C3451 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.01fF
C3452 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C3453 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C3454 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# VDD 0.15fF
C3455 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C3456 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C3457 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.02fF
C3458 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__nand2_1_4/B 0.10fF
C3459 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# VDD 0.14fF
C3460 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# 0.04fF
C3461 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.01fF
C3462 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.03fF
C3463 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.03fF
C3464 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# VDD 0.12fF
C3465 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C3466 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C3467 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.03fF
C3468 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.02fF
C3469 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.05fF
C3470 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.06fF
C3471 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.04fF
C3472 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.04fF
C3473 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.02fF
C3474 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# VDD 0.31fF
C3475 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C3476 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.01fF
C3477 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.09fF
C3478 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C3479 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.00fF
C3480 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.00fF
C3481 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.04fF
C3482 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VDD 0.53fF
C3483 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.03fF
C3484 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.01fF
C3485 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.02fF
C3486 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C3487 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C3488 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C3489 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C3490 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C3491 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C3492 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.29fF
C3493 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.05fF
C3494 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C3495 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C3496 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.08fF
C3497 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C3498 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C3499 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C3500 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.08fF
C3501 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C3502 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C3503 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C3504 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C3505 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C3506 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C3507 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.30fF
C3508 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# VDD 0.15fF
C3509 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C3510 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C3511 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.06fF
C3512 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C3513 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C3514 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C3515 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_1/A 0.10fF
C3516 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# 0.05fF
C3517 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.09fF
C3518 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C3519 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VDD 0.17fF
C3520 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C3521 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C3522 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.03fF
C3523 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.00fF
C3524 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.00fF
C3525 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.01fF
C3526 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.01fF
C3527 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_0/A 0.21fF
C3528 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.00fF
C3529 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C3530 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.00fF
C3531 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# VDD 0.14fF
C3532 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.05fF
C3533 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C3534 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/B 0.02fF
C3535 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.01fF
C3536 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C3537 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C3538 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C3539 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C3540 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.01fF
C3541 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C3542 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# VDD 0.31fF
C3543 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.02fF
C3544 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.05fF
C3545 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.05fF
C3546 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.04fF
C3547 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.05fF
C3548 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.05fF
C3549 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C3550 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C3551 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.01fF
C3552 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C3553 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.01fF
C3554 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C3555 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.01fF
C3556 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.01fF
C3557 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.02fF
C3558 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.04fF
C3559 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.03fF
C3560 p2 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.02fF
C3561 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.03fF
C3562 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C3563 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.03fF
C3564 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.02fF
C3565 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.01fF
C3566 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C3567 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Bd_b 0.14fF
C3568 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C3569 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.01fF
C3570 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.03fF
C3571 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C3572 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C3573 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.04fF
C3574 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C3575 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.00fF
C3576 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C3577 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C3578 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.08fF
C3579 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.02fF
C3580 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.04fF
C3581 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.04fF
C3582 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.00fF
C3583 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.03fF
C3584 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.01fF
C3585 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C3586 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.00fF
C3587 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.00fF
C3588 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C3589 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.01fF
C3590 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C3591 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C3592 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C3593 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.00fF
C3594 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.04fF
C3595 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.04fF
C3596 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C3597 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.08fF
C3598 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.08fF
C3599 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C3600 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C3601 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C3602 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.01fF
C3603 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# VDD 0.23fF
C3604 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.06fF
C3605 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.02fF
C3606 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C3607 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# 0.01fF
C3608 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VDD 0.52fF
C3609 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C3610 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C3611 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.08fF
C3612 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.02fF
C3613 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C3614 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.02fF
C3615 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C3616 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C3617 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.06fF
C3618 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.09fF
C3619 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_4_3/A 0.30fF
C3620 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.05fF
C3621 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.04fF
C3622 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.11fF
C3623 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.01fF
C3624 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.44fF
C3625 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C3626 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C3627 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C3628 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C3629 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C3630 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.02fF
C3631 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C3632 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C3633 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C3634 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C3635 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C3636 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C3637 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C3638 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C3639 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C3640 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X Ad_b 0.02fF
C3641 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkinv_4_1/A 0.11fF
C3642 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.08fF
C3643 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A VDD 0.56fF
C3644 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.01fF
C3645 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.02fF
C3646 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.01fF
C3647 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.01fF
C3648 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C3649 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# 0.01fF
C3650 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C3651 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.04fF
C3652 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.01fF
C3653 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C3654 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C3655 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.00fF
C3656 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.04fF
C3657 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.01fF
C3658 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C3659 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C3660 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C3661 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C3662 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C3663 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C3664 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VDD 0.53fF
C3665 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C3666 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C3667 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.01fF
C3668 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.04fF
C3669 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.04fF
C3670 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C3671 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C3672 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# VDD 0.12fF
C3673 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C3674 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C3675 p1 p1d 0.20fF
C3676 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_3/A 0.13fF
C3677 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# VDD 0.11fF
C3678 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C3679 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.02fF
C3680 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C3681 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.11fF
C3682 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C3683 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.03fF
C3684 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.01fF
C3685 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C3686 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.59fF
C3687 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C3688 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# 0.00fF
C3689 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.04fF
C3690 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# 0.01fF
C3691 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# VDD 0.46fF
C3692 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C3693 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C3694 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C3695 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.01fF
C3696 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.00fF
C3697 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C3698 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.03fF
C3699 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.01fF
C3700 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C3701 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.09fF
C3702 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VDD 0.87fF
C3703 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C3704 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C3705 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C3706 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C3707 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C3708 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 1.68fF
C3709 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.01fF
C3710 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.03fF
C3711 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.01fF
C3712 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C3713 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.01fF
C3714 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C3715 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.04fF
C3716 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.04fF
C3717 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.00fF
C3718 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C3719 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VDD 0.54fF
C3720 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.05fF
C3721 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C3722 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.02fF
C3723 sky130_fd_sc_hd__clkinv_4_7/Y p1_b 0.03fF
C3724 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C3725 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3726 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C3727 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C3728 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C3729 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.03fF
C3730 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# VDD 0.14fF
C3731 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.02fF
C3732 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C3733 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C3734 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.02fF
C3735 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.00fF
C3736 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.00fF
C3737 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3738 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.00fF
C3739 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C3740 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# VDD 0.16fF
C3741 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C3742 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C3743 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C3744 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.07fF
C3745 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.03fF
C3746 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C3747 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C3748 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C3749 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.03fF
C3750 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C3751 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.02fF
C3752 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C3753 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# VDD 0.33fF
C3754 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C3755 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C3756 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.01fF
C3757 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C3758 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.01fF
C3759 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkinv_4_5/Y 1.81fF
C3760 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C3761 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C3762 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C3763 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.32fF
C3764 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.01fF
C3765 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# VDD 0.18fF
C3766 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.01fF
C3767 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B 0.16fF
C3768 p2d p2 0.20fF
C3769 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C3770 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C3771 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C3772 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.07fF
C3773 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C3774 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.02fF
C3775 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# VDD 0.71fF
C3776 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C3777 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# Ad_b 0.07fF
C3778 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# Bd_b 0.05fF
C3779 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C3780 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C3781 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.11fF
C3782 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.01fF
C3783 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.01fF
C3784 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.01fF
C3785 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.08fF
C3786 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.09fF
C3787 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# VDD 0.45fF
C3788 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.03fF
C3789 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A -0.00fF
C3790 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.02fF
C3791 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C3792 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C3793 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Ad_b 0.12fF
C3794 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C3795 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.04fF
C3796 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.04fF
C3797 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C3798 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C3799 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C3800 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.01fF
C3801 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C3802 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.00fF
C3803 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.02fF
C3804 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C3805 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C3806 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C3807 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C3808 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C3809 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C3810 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C3811 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C3812 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C3813 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C3814 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.02fF
C3815 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C3816 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.04fF
C3817 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C3818 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.02fF
C3819 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C3820 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C3821 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C3822 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.01fF
C3823 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C3824 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C3825 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C3826 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.02fF
C3827 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.03fF
C3828 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C3829 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C3830 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VDD 0.35fF
C3831 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C3832 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C3833 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.11fF
C3834 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C3835 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C3836 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C3837 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.02fF
C3838 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C3839 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C3840 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C3841 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C3842 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.00fF
C3843 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C3844 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__nand2_4_2/A 0.80fF
C3845 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C3846 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C3847 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C3848 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C3849 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.01fF
C3850 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.01fF
C3851 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C3852 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C3853 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C3854 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.01fF
C3855 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.09fF
C3856 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C3857 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.10fF
C3858 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.02fF
C3859 A_b A 0.47fF
C3860 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.04fF
C3861 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.00fF
C3862 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C3863 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# Ad_b 0.12fF
C3864 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C3865 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C3866 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.00fF
C3867 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# 0.03fF
C3868 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.01fF
C3869 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.07fF
C3870 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.30fF
C3871 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# 0.10fF
C3872 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C3873 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.00fF
C3874 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.00fF
C3875 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.04fF
C3876 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.06fF
C3877 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C3878 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C3879 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.03fF
C3880 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.01fF
C3881 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.03fF
C3882 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C3883 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.01fF
C3884 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.00fF
C3885 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.00fF
C3886 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C3887 sky130_fd_sc_hd__mux2_1_0/X Bd_b 0.01fF
C3888 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.04fF
C3889 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C3890 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C3891 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C3892 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.02fF
C3893 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C3894 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C3895 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C3896 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C3897 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C3898 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.02fF
C3899 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.02fF
C3900 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C3901 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.02fF
C3902 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.01fF
C3903 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C3904 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C3905 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C3906 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.00fF
C3907 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C3908 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C3909 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C3910 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C3911 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C3912 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# 0.04fF
C3913 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.04fF
C3914 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C3915 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.03fF
C3916 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C3917 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C3918 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C3919 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C3920 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C3921 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# VDD 0.15fF
C3922 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C3923 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.02fF
C3924 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.02fF
C3925 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C3926 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C3927 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C3928 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.10fF
C3929 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.44fF
C3930 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C3931 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C3932 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# p2 0.02fF
C3933 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C3934 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C3935 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.02fF
C3936 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.05fF
C3937 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.05fF
C3938 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.05fF
C3939 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.04fF
C3940 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.04fF
C3941 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.02fF
C3942 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.02fF
C3943 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C3944 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C3945 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C3946 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C3947 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.05fF
C3948 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C3949 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.01fF
C3950 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.02fF
C3951 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C3952 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C3953 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/A 0.47fF
C3954 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# VDD 0.13fF
C3955 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.43fF
C3956 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.04fF
C3957 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.31fF
C3958 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C3959 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.02fF
C3960 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# 0.02fF
C3961 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# 0.01fF
C3962 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# 0.01fF
C3963 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C3964 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C3965 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C3966 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C3967 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C3968 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.09fF
C3969 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# VDD 0.14fF
C3970 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C3971 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C3972 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.03fF
C3973 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.02fF
C3974 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.00fF
C3975 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.01fF
C3976 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.02fF
C3977 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.02fF
C3978 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.01fF
C3979 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C3980 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C3981 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VDD 0.50fF
C3982 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C3983 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.02fF
C3984 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.01fF
C3985 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C3986 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.16fF
C3987 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_2/A 0.00fF
C3988 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Ad_b 0.09fF
C3989 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C3990 sky130_fd_sc_hd__clkinv_1_3/A p2 0.24fF
C3991 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C3992 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C3993 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C3994 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C3995 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C3996 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C3997 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.01fF
C3998 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.06fF
C3999 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4000 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C4001 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4002 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C4003 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.00fF
C4004 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.02fF
C4005 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.02fF
C4006 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VDD -0.81fF
C4007 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.07fF
C4008 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# 0.00fF
C4009 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# 0.00fF
C4010 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.06fF
C4011 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C4012 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C4013 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.05fF
C4014 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.05fF
C4015 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C4016 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.07fF
C4017 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/D -0.03fF
C4018 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# VDD -0.06fF
C4019 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VDD 0.60fF
C4020 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C4021 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# 0.11fF
C4022 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.00fF
C4023 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.01fF
C4024 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C4025 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C4026 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.08fF
C4027 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.02fF
C4028 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.02fF
C4029 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C4030 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C4031 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C4032 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.00fF
C4033 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.00fF
C4034 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C4035 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.09fF
C4036 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.01fF
C4037 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C4038 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.02fF
C4039 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C4040 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.13fF
C4041 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.00fF
C4042 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.02fF
C4043 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.02fF
C4044 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.02fF
C4045 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# 0.01fF
C4046 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.04fF
C4047 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C4048 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.02fF
C4049 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.17fF
C4050 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C4051 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C4052 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.03fF
C4053 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.16fF
C4054 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C4055 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.02fF
C4056 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C4057 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.00fF
C4058 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.00fF
C4059 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C4060 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkinv_4_1/A 0.07fF
C4061 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.84fF
C4062 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.02fF
C4063 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C4064 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/A 0.87fF
C4065 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.21fF
C4066 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C4067 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C4068 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C4069 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4070 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C4071 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C4072 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C4073 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C4074 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C4075 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C4076 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C4077 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.09fF
C4078 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.00fF
C4079 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.00fF
C4080 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.02fF
C4081 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.11fF
C4082 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C4083 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C4084 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.02fF
C4085 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C4086 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C4087 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# VDD 0.15fF
C4088 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C4089 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C4090 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.01fF
C4091 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.01fF
C4092 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.03fF
C4093 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.01fF
C4094 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.01fF
C4095 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/A 1.27fF
C4096 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C4097 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C4098 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C4099 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C4100 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.01fF
C4101 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.02fF
C4102 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# VDD 0.14fF
C4103 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.01fF
C4104 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.04fF
C4105 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# VDD 0.12fF
C4106 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/A 0.01fF
C4107 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C4108 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# VDD 0.16fF
C4109 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C4110 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.08fF
C4111 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C4112 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# 0.09fF
C4113 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.00fF
C4114 Bd sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.12fF
C4115 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# VDD 0.08fF
C4116 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C4117 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# VDD 0.29fF
C4118 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.06fF
C4119 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.03fF
C4120 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# 0.11fF
C4121 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.02fF
C4122 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.01fF
C4123 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C4124 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C4125 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C4126 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.03fF
C4127 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C4128 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.00fF
C4129 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.02fF
C4130 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C4131 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C4132 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# 0.00fF
C4133 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# VDD 0.24fF
C4134 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C4135 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.00fF
C4136 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.00fF
C4137 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.08fF
C4138 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C4139 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C4140 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.01fF
C4141 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A VDD 0.56fF
C4142 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C4143 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C4144 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.05fF
C4145 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.08fF
C4146 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.01fF
C4147 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C4148 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# 0.09fF
C4149 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C4150 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C4151 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C4152 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.06fF
C4153 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C4154 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.01fF
C4155 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.00fF
C4156 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.03fF
C4157 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.03fF
C4158 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C4159 sky130_fd_sc_hd__nand2_4_1/B VDD 0.68fF
C4160 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.02fF
C4161 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.00fF
C4162 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C4163 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.04fF
C4164 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VDD 0.11fF
C4165 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C4166 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4167 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.00fF
C4168 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.07fF
C4169 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C4170 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.11fF
C4171 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C4172 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C4173 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C4174 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.06fF
C4175 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C4176 p1d_b VDD 0.80fF
C4177 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C4178 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C4179 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.02fF
C4180 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VDD 0.58fF
C4181 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C4182 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C4183 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkinv_4_10/Y 0.08fF
C4184 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C4185 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C4186 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C4187 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C4188 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# 0.07fF
C4189 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.01fF
C4190 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.00fF
C4191 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C4192 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C4193 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C4194 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C4195 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.01fF
C4196 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C4197 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C4198 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C4199 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.00fF
C4200 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.01fF
C4201 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.01fF
C4202 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.02fF
C4203 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# Bd_b 0.02fF
C4204 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C4205 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.03fF
C4206 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.09fF
C4207 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VDD 0.31fF
C4208 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C4209 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C4210 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C4211 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C4212 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C4213 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.01fF
C4214 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.03fF
C4215 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X -0.00fF
C4216 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.01fF
C4217 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C4218 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.02fF
C4219 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.01fF
C4220 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C4221 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C4222 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# 0.07fF
C4223 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C4224 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.03fF
C4225 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C4226 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C4227 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VDD 0.51fF
C4228 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C4229 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# VDD 0.14fF
C4230 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C4231 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.03fF
C4232 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.01fF
C4233 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.03fF
C4234 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C4235 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C4236 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.09fF
C4237 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C4238 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C4239 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C4240 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C4241 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.11fF
C4242 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C4243 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C4244 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VDD 0.31fF
C4245 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.02fF
C4246 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C4247 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4248 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C4249 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.01fF
C4250 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# VDD 0.14fF
C4251 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.04fF
C4252 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C4253 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/A 0.01fF
C4254 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.00fF
C4255 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.00fF
C4256 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.00fF
C4257 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C4258 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C4259 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.01fF
C4260 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C4261 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.11fF
C4262 sky130_fd_sc_hd__clkinv_1_3/A Ad_b 0.25fF
C4263 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C4264 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# VDD 0.14fF
C4265 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.01fF
C4266 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.06fF
C4267 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.03fF
C4268 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C4269 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.09fF
C4270 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C4271 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C4272 sky130_fd_sc_hd__nand2_4_3/Y VDD 5.51fF
C4273 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.03fF
C4274 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# VDD 0.29fF
C4275 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C4276 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.04fF
C4277 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C4278 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C4279 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C4280 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.01fF
C4281 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C4282 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.00fF
C4283 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.00fF
C4284 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C4285 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C4286 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.01fF
C4287 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.05fF
C4288 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# VDD 0.12fF
C4289 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C4290 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C4291 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.01fF
C4292 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C4293 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C4294 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C4295 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C4296 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C4297 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C4298 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# VDD 0.12fF
C4299 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C4300 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.00fF
C4301 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C4302 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C4303 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X VDD 0.57fF
C4304 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C4305 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.01fF
C4306 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.01fF
C4307 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C4308 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4309 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# 0.05fF
C4310 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C4311 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# VDD 0.17fF
C4312 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.01fF
C4313 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C4314 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C4315 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.02fF
C4316 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C4317 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C4318 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.04fF
C4319 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.06fF
C4320 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VDD 0.54fF
C4321 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.01fF
C4322 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C4323 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.02fF
C4324 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.04fF
C4325 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.04fF
C4326 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C4327 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# VDD 0.32fF
C4328 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.01fF
C4329 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.09fF
C4330 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C4331 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C4332 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C4333 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C4334 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C4335 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C4336 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C4337 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C4338 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C4339 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.02fF
C4340 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.52fF
C4341 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C4342 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C4343 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.09fF
C4344 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.05fF
C4345 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.05fF
C4346 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# VDD 0.12fF
C4347 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C4348 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.00fF
C4349 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.11fF
C4350 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# 0.09fF
C4351 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C4352 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.00fF
C4353 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.00fF
C4354 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.01fF
C4355 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.03fF
C4356 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.01fF
C4357 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.00fF
C4358 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.00fF
C4359 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C4360 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C4361 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C4362 sky130_fd_sc_hd__nand2_4_1/Y Bd_b 0.22fF
C4363 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C4364 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.02fF
C4365 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C4366 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C4367 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.00fF
C4368 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.02fF
C4369 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C4370 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.00fF
C4371 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C4372 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C4373 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C4374 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C4375 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.03fF
C4376 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C4377 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C4378 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C4379 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.01fF
C4380 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.02fF
C4381 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.01fF
C4382 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.04fF
C4383 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C4384 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.01fF
C4385 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.02fF
C4386 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.00fF
C4387 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.01fF
C4388 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C4389 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.00fF
C4390 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C4391 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C4392 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.01fF
C4393 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkinv_1_0/Y 0.06fF
C4394 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C4395 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C4396 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C4397 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.05fF
C4398 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# 0.05fF
C4399 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C4400 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C4401 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.02fF
C4402 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C4403 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C4404 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# VDD 0.14fF
C4405 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.07fF
C4406 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VDD 0.09fF
C4407 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.07fF
C4408 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VDD 0.34fF
C4409 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C4410 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.13fF
C4411 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C4412 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.03fF
C4413 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.11fF
C4414 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.09fF
C4415 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# 0.07fF
C4416 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C4417 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C4418 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C4419 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.02fF
C4420 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.02fF
C4421 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.32fF
C4422 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C4423 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.14fF
C4424 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C4425 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.01fF
C4426 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C4427 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C4428 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.00fF
C4429 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.01fF
C4430 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.02fF
C4431 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C4432 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.00fF
C4433 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C4434 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C4435 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B 0.69fF
C4436 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.04fF
C4437 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C4438 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.02fF
C4439 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.05fF
C4440 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.06fF
C4441 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C4442 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C4443 A_b Ad_b 0.33fF
C4444 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.01fF
C4445 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.01fF
C4446 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C4447 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C4448 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C4449 sky130_fd_sc_hd__mux2_1_0/a_439_47# Bd_b 0.00fF
C4450 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C4451 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.06fF
C4452 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C4453 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C4454 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.22fF
C4455 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C4456 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C4457 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C4458 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C4459 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.02fF
C4460 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C4461 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C4462 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C4463 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C4464 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.02fF
C4465 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.02fF
C4466 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C4467 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# VDD 0.14fF
C4468 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.03fF
C4469 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C4470 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_1_4/B 0.13fF
C4471 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.08fF
C4472 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.52fF
C4473 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C4474 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VDD 0.49fF
C4475 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C4476 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C4477 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C4478 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C4479 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# VDD 0.11fF
C4480 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_7/Y 0.19fF
C4481 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.03fF
C4482 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C4483 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.04fF
C4484 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C4485 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.04fF
C4486 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.01fF
C4487 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.01fF
C4488 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.01fF
C4489 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C4490 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C4491 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.06fF
C4492 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# VDD 0.16fF
C4493 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.02fF
C4494 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.04fF
C4495 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.04fF
C4496 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.09fF
C4497 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C4498 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C4499 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C4500 p1_b sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.15fF
C4501 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# p1d 0.15fF
C4502 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C4503 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C4504 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.05fF
C4505 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.07fF
C4506 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.01fF
C4507 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C4508 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.01fF
C4509 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkinv_4_3/Y -0.00fF
C4510 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Ad 0.12fF
C4511 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.15fF
C4512 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.03fF
C4513 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C4514 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4515 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C4516 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C4517 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.17fF
C4518 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.03fF
C4519 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.05fF
C4520 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4521 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.03fF
C4522 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.37fF
C4523 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.07fF
C4524 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C4525 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C4526 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C4527 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.06fF
C4528 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C4529 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C4530 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C4531 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.01fF
C4532 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.17fF
C4533 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C4534 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.04fF
C4535 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.01fF
C4536 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C4537 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C4538 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C4539 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C4540 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C4541 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C4542 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.03fF
C4543 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.32fF
C4544 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C4545 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VDD 0.14fF
C4546 VDD sky130_fd_sc_hd__nand2_4_3/A 10.99fF
C4547 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.01fF
C4548 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# 0.11fF
C4549 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.02fF
C4550 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C4551 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C4552 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C4553 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.00fF
C4554 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.00fF
C4555 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.00fF
C4556 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.04fF
C4557 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# VDD 0.14fF
C4558 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C4559 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C4560 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C4561 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C4562 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C4563 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C4564 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# VDD 0.14fF
C4565 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkinv_4_7/A 0.03fF
C4566 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# 0.09fF
C4567 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.02fF
C4568 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.01fF
C4569 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.01fF
C4570 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C4571 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.09fF
C4572 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A VDD 0.52fF
C4573 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.01fF
C4574 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VDD 0.27fF
C4575 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C4576 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.02fF
C4577 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.03fF
C4578 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C4579 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C4580 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C4581 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.06fF
C4582 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.03fF
C4583 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.05fF
C4584 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.00fF
C4585 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C4586 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C4587 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C4588 sky130_fd_sc_hd__clkinv_4_10/Y VDD 0.49fF
C4589 VDD p1 1.45fF
C4590 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.02fF
C4591 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C4592 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.00fF
C4593 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C4594 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.05fF
C4595 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.01fF
C4596 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.03fF
C4597 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.03fF
C4598 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C4599 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C4600 p2d_b sky130_fd_sc_hd__clkinv_4_9/Y 0.03fF
C4601 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C4602 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4603 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.03fF
C4604 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C4605 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C4606 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C4607 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.00fF
C4608 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C4609 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C4610 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C4611 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.02fF
C4612 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.02fF
C4613 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C4614 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C4615 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.04fF
C4616 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C4617 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C4618 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C4619 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.02fF
C4620 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# 0.04fF
C4621 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# 0.04fF
C4622 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C4623 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C4624 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# 0.00fF
C4625 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.03fF
C4626 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C4627 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VDD 0.33fF
C4628 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.01fF
C4629 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# 0.03fF
C4630 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.00fF
C4631 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C4632 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C4633 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.01fF
C4634 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C4635 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C4636 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C4637 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# VDD 0.14fF
C4638 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.02fF
C4639 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C4640 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C4641 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C4642 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# VDD 0.32fF
C4643 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# VDD 0.34fF
C4644 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C4645 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C4646 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C4647 VDD sky130_fd_sc_hd__clkbuf_16_5/a_110_47# -0.06fF
C4648 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C4649 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.03fF
C4650 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# 0.05fF
C4651 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.06fF
C4652 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.03fF
C4653 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C4654 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C4655 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C4656 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C4657 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C4658 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.01fF
C4659 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C4660 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C4661 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C4662 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C4663 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.05fF
C4664 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X Bd_b 0.03fF
C4665 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.01fF
C4666 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C4667 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C4668 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C4669 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.02fF
C4670 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.02fF
C4671 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C4672 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C4673 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.04fF
C4674 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.04fF
C4675 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.04fF
C4676 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C4677 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C4678 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.02fF
C4679 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkinv_1_1/Y 0.06fF
C4680 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.00fF
C4681 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C4682 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.00fF
C4683 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C4684 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C4685 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.01fF
C4686 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C4687 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C4688 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C4689 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C4690 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C4691 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0.04fF
C4692 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C4693 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# 0.01fF
C4694 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# 0.04fF
C4695 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.04fF
C4696 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C4697 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkinv_1_0/Y 0.02fF
C4698 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C4699 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.04fF
C4700 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# VDD 0.10fF
C4701 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4702 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C4703 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VDD 0.68fF
C4704 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.04fF
C4705 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# VDD 0.19fF
C4706 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C4707 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.01fF
C4708 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.06fF
C4709 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C4710 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.00fF
C4711 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# VDD 0.34fF
C4712 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C4713 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C4714 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C4715 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.01fF
C4716 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.03fF
C4717 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C4718 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.02fF
C4719 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C4720 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.02fF
C4721 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C4722 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.00fF
C4723 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C4724 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.03fF
C4725 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C4726 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.01fF
C4727 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C4728 sky130_fd_sc_hd__clkinv_4_3/Y VDD 1.73fF
C4729 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C4730 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C4731 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.07fF
C4732 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C4733 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.09fF
C4734 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C4735 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.06fF
C4736 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.13fF
C4737 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# 0.02fF
C4738 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.00fF
C4739 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C4740 sky130_fd_sc_hd__clkinv_4_4/Y VDD 0.57fF
C4741 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.03fF
C4742 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# VDD 0.13fF
C4743 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.06fF
C4744 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.03fF
C4745 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# VDD 0.22fF
C4746 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.02fF
C4747 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C4748 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C4749 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C4750 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C4751 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.02fF
C4752 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.02fF
C4753 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C4754 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# VDD 0.15fF
C4755 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C4756 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C4757 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C4758 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.00fF
C4759 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# 0.01fF
C4760 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C4761 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# VDD 0.29fF
C4762 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.01fF
C4763 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C4764 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.08fF
C4765 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.06fF
C4766 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__nand2_1_2/B 0.02fF
C4767 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C4768 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C4769 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.04fF
C4770 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.17fF
C4771 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C4772 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.01fF
C4773 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.00fF
C4774 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4775 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C4776 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# VDD 0.30fF
C4777 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# VDD 0.14fF
C4778 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C4779 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C4780 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.29fF
C4781 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C4782 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C4783 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.01fF
C4784 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C4785 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# VDD 0.18fF
C4786 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4787 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# Bd_b 0.06fF
C4788 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.02fF
C4789 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.02fF
C4790 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.04fF
C4791 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.04fF
C4792 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.05fF
C4793 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.04fF
C4794 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.04fF
C4795 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# VDD 0.17fF
C4796 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.04fF
C4797 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.04fF
C4798 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A -0.00fF
C4799 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C4800 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C4801 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C4802 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Bd_b 0.14fF
C4803 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_4_2/A 0.15fF
C4804 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C4805 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.02fF
C4806 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.01fF
C4807 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C4808 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.01fF
C4809 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# VDD 0.21fF
C4810 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.01fF
C4811 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.03fF
C4812 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C4813 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.02fF
C4814 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C4815 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C4816 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.01fF
C4817 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C4818 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C4819 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C4820 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C4821 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C4822 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C4823 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C4824 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C4825 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C4826 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C4827 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C4828 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.00fF
C4829 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.02fF
C4830 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C4831 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.02fF
C4832 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C4833 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_1/Y 0.33fF
C4834 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C4835 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_4/B 0.92fF
C4836 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# 0.03fF
C4837 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C4838 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.03fF
C4839 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C4840 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C4841 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C4842 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.00fF
C4843 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C4844 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C4845 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.08fF
C4846 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.01fF
C4847 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.00fF
C4848 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.03fF
C4849 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C4850 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C4851 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C4852 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.03fF
C4853 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C4854 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.01fF
C4855 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C4856 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.02fF
C4857 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0.02fF
C4858 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C4859 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.01fF
C4860 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C4861 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# 0.01fF
C4862 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VDD 0.29fF
C4863 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.01fF
C4864 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C4865 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.01fF
C4866 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.02fF
C4867 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C4868 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C4869 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.03fF
C4870 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 1.80fF
C4871 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C4872 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C4873 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# Bd_b 0.10fF
C4874 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.01fF
C4875 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C4876 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.18fF
C4877 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.02fF
C4878 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.55fF
C4879 sky130_fd_sc_hd__nand2_4_0/Y Bd 0.00fF
C4880 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.01fF
C4881 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C4882 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.00fF
C4883 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.04fF
C4884 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C4885 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.01fF
C4886 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C4887 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C4888 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C4889 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C4890 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C4891 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C4892 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.01fF
C4893 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.02fF
C4894 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.09fF
C4895 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C4896 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/A 1.15fF
C4897 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.03fF
C4898 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C4899 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.00fF
C4900 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C4901 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C4902 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C4903 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C4904 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.02fF
C4905 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.01fF
C4906 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# 0.01fF
C4907 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# 0.01fF
C4908 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.02fF
C4909 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.00fF
C4910 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.01fF
C4911 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C4912 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C4913 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C4914 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C4915 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C4916 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C4917 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.01fF
C4918 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.03fF
C4919 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C4920 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.00fF
C4921 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C4922 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.05fF
C4923 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C4924 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.00fF
C4925 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C4926 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C4927 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C4928 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C4929 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C4930 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C4931 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.04fF
C4932 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C4933 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.01fF
C4934 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# 0.01fF
C4935 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.01fF
C4936 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.02fF
C4937 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.01fF
C4938 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# 0.01fF
C4939 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.01fF
C4940 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.01fF
C4941 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C4942 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.03fF
C4943 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.02fF
C4944 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.03fF
C4945 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4946 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C4947 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.09fF
C4948 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.05fF
C4949 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# 0.12fF
C4950 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.11fF
C4951 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.11fF
C4952 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.18fF
C4953 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.01fF
C4954 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.01fF
C4955 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# 0.02fF
C4956 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# 0.02fF
C4957 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4958 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.07fF
C4959 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# VDD 0.14fF
C4960 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C4961 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C4962 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.33fF
C4963 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C4964 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C4965 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.35fF
C4966 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.01fF
C4967 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.01fF
C4968 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.09fF
C4969 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.01fF
C4970 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4971 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.09fF
C4972 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C4973 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.00fF
C4974 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C4975 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.10fF
C4976 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VDD 0.21fF
C4977 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C4978 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Bd_b 0.07fF
C4979 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C4980 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.00fF
C4981 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.02fF
C4982 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C4983 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C4984 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C4985 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C4986 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.03fF
C4987 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.09fF
C4988 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C4989 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.40fF
C4990 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C4991 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C4992 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.01fF
C4993 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4994 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C4995 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.07fF
C4996 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VDD 0.74fF
C4997 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.02fF
C4998 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C4999 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C5000 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C5001 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.02fF
C5002 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.06fF
C5003 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.02fF
C5004 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# VDD 0.08fF
C5005 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.07fF
C5006 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.07fF
C5007 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/D 0.02fF
C5008 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.03fF
C5009 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C5010 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.02fF
C5011 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.03fF
C5012 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C5013 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C5014 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.02fF
C5015 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C5016 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.02fF
C5017 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C5018 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C5019 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.01fF
C5020 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C5021 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.00fF
C5022 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.00fF
C5023 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VDD 0.47fF
C5024 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.01fF
C5025 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C5026 sky130_fd_sc_hd__nand2_4_2/a_27_47# VDD 0.04fF
C5027 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C5028 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C5029 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C5030 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# 0.03fF
C5031 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C5032 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C5033 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.14fF
C5034 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.00fF
C5035 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.00fF
C5036 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.03fF
C5037 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.00fF
C5038 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.15fF
C5039 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C5040 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C5041 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.00fF
C5042 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C5043 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C5044 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkinv_4_1/A 0.06fF
C5045 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C5046 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.06fF
C5047 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.07fF
C5048 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.09fF
C5049 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.00fF
C5050 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C5051 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C5052 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5053 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.03fF
C5054 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.00fF
C5055 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.00fF
C5056 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.00fF
C5057 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C5058 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C5059 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.00fF
C5060 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.00fF
C5061 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.04fF
C5062 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.04fF
C5063 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.30fF
C5064 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C5065 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.04fF
C5066 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.04fF
C5067 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.02fF
C5068 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.02fF
C5069 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.03fF
C5070 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C5071 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.01fF
C5072 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C5073 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.01fF
C5074 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C5075 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C5076 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# VDD 0.12fF
C5077 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkinv_1_3/Y 0.06fF
C5078 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.06fF
C5079 Bd VDD 1.53fF
C5080 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C5081 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C5082 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.00fF
C5083 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C5084 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.00fF
C5085 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# VDD 0.09fF
C5086 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# VDD 0.11fF
C5087 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.03fF
C5088 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# 0.00fF
C5089 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.01fF
C5090 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.02fF
C5091 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C5092 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.04fF
C5093 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C5094 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C5095 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C5096 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C5097 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C5098 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# VDD 0.12fF
C5099 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.02fF
C5100 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.08fF
C5101 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# VDD 0.31fF
C5102 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C5103 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.05fF
C5104 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.05fF
C5105 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C5106 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.00fF
C5107 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C5108 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__nand2_4_2/B 0.08fF
C5109 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.01fF
C5110 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C5111 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C5112 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C5113 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C5114 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# VDD 0.30fF
C5115 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/B 0.02fF
C5116 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C5117 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C5118 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.09fF
C5119 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.08fF
C5120 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.01fF
C5121 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.01fF
C5122 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# 0.11fF
C5123 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C5124 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.02fF
C5125 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C5126 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C5127 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VDD 0.59fF
C5128 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.09fF
C5129 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C5130 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.00fF
C5131 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# 0.06fF
C5132 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VDD 0.32fF
C5133 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.02fF
C5134 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.01fF
C5135 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C5136 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C5137 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.00fF
C5138 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.01fF
C5139 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.31fF
C5140 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C5141 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.01fF
C5142 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C5143 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.00fF
C5144 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C5145 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.03fF
C5146 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.16fF
C5147 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.01fF
C5148 sky130_fd_sc_hd__clkinv_4_1/Y B_b 0.03fF
C5149 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C5150 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C5151 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.06fF
C5152 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.00fF
C5153 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.03fF
C5154 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.05fF
C5155 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__mux2_1_0/S 0.11fF
C5156 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# 0.03fF
C5157 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.01fF
C5158 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.02fF
C5159 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# 0.00fF
C5160 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.02fF
C5161 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C5162 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.00fF
C5163 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C5164 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C5165 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C5166 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.03fF
C5167 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.02fF
C5168 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.02fF
C5169 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C5170 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C5171 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C5172 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.01fF
C5173 B sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.12fF
C5174 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# B_b 0.12fF
C5175 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C5176 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.03fF
C5177 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.06fF
C5178 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.09fF
C5179 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C5180 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C5181 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C5182 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.03fF
C5183 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# 0.06fF
C5184 sky130_fd_sc_hd__nand2_4_1/Y Ad 0.00fF
C5185 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.01fF
C5186 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.03fF
C5187 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C5188 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C5189 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.01fF
C5190 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C5191 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C5192 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C5193 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C5194 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.06fF
C5195 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.03fF
C5196 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C5197 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.01fF
C5198 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.01fF
C5199 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.09fF
C5200 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.04fF
C5201 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C5202 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.00fF
C5203 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C5204 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C5205 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C5206 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.00fF
C5207 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.00fF
C5208 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.34fF
C5209 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C5210 sky130_fd_sc_hd__clkinv_1_3/A Bd_b 0.22fF
C5211 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.05fF
C5212 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# VDD 0.11fF
C5213 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.00fF
C5214 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C5215 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.00fF
C5216 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.00fF
C5217 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.03fF
C5218 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C5219 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C5220 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C5221 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# VDD 0.11fF
C5222 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C5223 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.02fF
C5224 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.01fF
C5225 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# VDD 0.31fF
C5226 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/A 0.84fF
C5227 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C5228 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.01fF
C5229 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C5230 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C5231 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C5232 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.02fF
C5233 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C5234 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C5235 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C5236 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.01fF
C5237 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.02fF
C5238 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.09fF
C5239 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.00fF
C5240 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C5241 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C5242 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C5243 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C5244 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C5245 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C5246 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C5247 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C5248 VDD sky130_fd_sc_hd__nand2_1_1/B 1.42fF
C5249 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.02fF
C5250 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.02fF
C5251 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C5252 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C5253 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C5254 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.02fF
C5255 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C5256 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# VDD 0.14fF
C5257 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C5258 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.02fF
C5259 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C5260 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C5261 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C5262 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C5263 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.02fF
C5264 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.00fF
C5265 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C5266 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C5267 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C5268 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C5269 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.02fF
C5270 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.02fF
C5271 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# VDD 0.14fF
C5272 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.02fF
C5273 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C5274 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C5275 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C5276 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.06fF
C5277 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C5278 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C5279 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C5280 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C5281 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C5282 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C5283 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C5284 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C5285 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.02fF
C5286 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# VDD 0.29fF
C5287 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C5288 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.02fF
C5289 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C5290 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C5291 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C5292 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.00fF
C5293 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.00fF
C5294 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C5295 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C5296 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.01fF
C5297 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C5298 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.06fF
C5299 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C5300 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.02fF
C5301 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C5302 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C5303 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C5304 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.03fF
C5305 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C5306 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C5307 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.01fF
C5308 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_1/A 0.87fF
C5309 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C5310 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C5311 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C5312 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C5313 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C5314 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C5315 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.01fF
C5316 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C5317 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.06fF
C5318 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.00fF
C5319 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C5320 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C5321 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.01fF
C5322 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.01fF
C5323 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C5324 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C5325 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.04fF
C5326 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.04fF
C5327 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C5328 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.01fF
C5329 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.01fF
C5330 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.07fF
C5331 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C5332 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C5333 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C5334 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C5335 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.02fF
C5336 VDD sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.46fF
C5337 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# 0.12fF
C5338 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C5339 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.07fF
C5340 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# 0.01fF
C5341 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.01fF
C5342 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.01fF
C5343 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.02fF
C5344 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.00fF
C5345 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C5346 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.01fF
C5347 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C5348 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C5349 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.01fF
C5350 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.02fF
C5351 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.04fF
C5352 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.04fF
C5353 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# 0.11fF
C5354 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.03fF
C5355 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.01fF
C5356 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.00fF
C5357 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C5358 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.11fF
C5359 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C5360 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.11fF
C5361 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C5362 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.08fF
C5363 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VDD 0.17fF
C5364 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.03fF
C5365 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C5366 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VDD -0.76fF
C5367 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C5368 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C5369 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# 0.07fF
C5370 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.16fF
C5371 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.13fF
C5372 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C5373 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C5374 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C5375 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.01fF
C5376 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.01fF
C5377 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.02fF
C5378 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C5379 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.09fF
C5380 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.03fF
C5381 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.00fF
C5382 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C5383 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C5384 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C5385 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.02fF
C5386 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C5387 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.02fF
C5388 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C5389 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.11fF
C5390 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.03fF
C5391 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.01fF
C5392 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C5393 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.02fF
C5394 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.56fF
C5395 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.06fF
C5396 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C5397 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.00fF
C5398 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C5399 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.03fF
C5400 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C5401 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C5402 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C5403 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C5404 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.03fF
C5405 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.02fF
C5406 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C5407 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C5408 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C5409 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C5410 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C5411 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.00fF
C5412 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C5413 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C5414 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C5415 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C5416 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.02fF
C5417 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# 0.05fF
C5418 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C5419 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.09fF
C5420 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C5421 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C5422 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.04fF
C5423 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.04fF
C5424 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.04fF
C5425 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.06fF
C5426 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C5427 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.04fF
C5428 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.01fF
C5429 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C5430 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.03fF
C5431 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.01fF
C5432 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.02fF
C5433 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.02fF
C5434 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C5435 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C5436 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C5437 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.01fF
C5438 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.01fF
C5439 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.01fF
C5440 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.01fF
C5441 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# VDD 0.14fF
C5442 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.03fF
C5443 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C5444 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.02fF
C5445 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C5446 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C5447 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.11fF
C5448 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C5449 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C5450 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.02fF
C5451 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.01fF
C5452 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C5453 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C5454 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.06fF
C5455 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.01fF
C5456 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.02fF
C5457 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C5458 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.14fF
C5459 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.01fF
C5460 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C5461 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C5462 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.19fF
C5463 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C5464 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C5465 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C5466 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C5467 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.70fF
C5468 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.00fF
C5469 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# 0.00fF
C5470 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C5471 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.01fF
C5472 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C5473 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.08fF
C5474 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C5475 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.11fF
C5476 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.00fF
C5477 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C5478 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A Ad_b 0.00fF
C5479 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.06fF
C5480 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C5481 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C5482 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.14fF
C5483 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C5484 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C5485 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C5486 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C5487 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C5488 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C5489 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.01fF
C5490 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.01fF
C5491 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.01fF
C5492 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.07fF
C5493 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.14fF
C5494 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.00fF
C5495 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.00fF
C5496 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C5497 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# 0.01fF
C5498 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C5499 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C5500 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.01fF
C5501 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.09fF
C5502 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.08fF
C5503 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.00fF
C5504 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.00fF
C5505 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C5506 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.00fF
C5507 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C5508 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# 0.01fF
C5509 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VDD 0.52fF
C5510 B Bd 0.20fF
C5511 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.06fF
C5512 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VDD 0.32fF
C5513 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_1_0/Y 0.37fF
C5514 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C5515 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C5516 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.00fF
C5517 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.04fF
C5518 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.04fF
C5519 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# VDD 0.14fF
C5520 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.02fF
C5521 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.02fF
C5522 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C5523 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C5524 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# 0.23fF
C5525 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C5526 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C5527 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C5528 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C5529 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C5530 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C5531 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C5532 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C5533 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VDD 0.53fF
C5534 p2 sky130_fd_sc_hd__nand2_4_1/B 0.04fF
C5535 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C5536 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C5537 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.03fF
C5538 p2 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.00fF
C5539 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C5540 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C5541 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.00fF
C5542 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C5543 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C5544 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C5545 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.04fF
C5546 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C5547 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C5548 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A 1.13fF
C5549 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.10fF
C5550 sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.05fF
C5551 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# 0.02fF
C5552 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.01fF
C5553 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.02fF
C5554 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C5555 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C5556 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C5557 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.03fF
C5558 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.03fF
C5559 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C5560 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C5561 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C5562 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# Ad_b 0.00fF
C5563 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.01fF
C5564 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C5565 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.03fF
C5566 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C5567 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.02fF
C5568 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.03fF
C5569 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C5570 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C5571 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C5572 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C5573 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.02fF
C5574 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.02fF
C5575 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.04fF
C5576 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C5577 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.04fF
C5578 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C5579 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C5580 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# 0.01fF
C5581 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# 0.01fF
C5582 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# 0.01fF
C5583 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.01fF
C5584 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C5585 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.01fF
C5586 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C5587 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.03fF
C5588 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VDD 0.18fF
C5589 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.00fF
C5590 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.00fF
C5591 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C5592 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VDD 0.34fF
C5593 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.02fF
C5594 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.02fF
C5595 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# VDD 0.11fF
C5596 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.01fF
C5597 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C5598 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# VDD 0.14fF
C5599 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# VDD 0.17fF
C5600 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C5601 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.06fF
C5602 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.02fF
C5603 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# VDD 0.30fF
C5604 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.08fF
C5605 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# VDD 0.30fF
C5606 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# VDD 0.32fF
C5607 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C5608 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C5609 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.11fF
C5610 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.06fF
C5611 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C5612 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C5613 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.04fF
C5614 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.04fF
C5615 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C5616 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C5617 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C5618 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.21fF
C5619 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.01fF
C5620 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkinv_1_0/Y 0.02fF
C5621 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.02fF
C5622 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.00fF
C5623 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.00fF
C5624 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C5625 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.04fF
C5626 p2 sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C5627 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# 0.11fF
C5628 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C5629 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C5630 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.11fF
C5631 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C5632 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C5633 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C5634 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.09fF
C5635 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.01fF
C5636 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C5637 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.01fF
C5638 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C5639 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C5640 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C5641 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.00fF
C5642 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.00fF
C5643 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.00fF
C5644 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.02fF
C5645 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C5646 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.00fF
C5647 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C5648 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C5649 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C5650 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C5651 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkinv_1_2/Y 0.02fF
C5652 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C5653 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.00fF
C5654 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.02fF
C5655 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# 0.01fF
C5656 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# 0.01fF
C5657 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.01fF
C5658 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.02fF
C5659 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C5660 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C5661 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C5662 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C5663 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkinv_4_1/A 0.11fF
C5664 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C5665 VDD sky130_fd_sc_hd__clkinv_1_2/Y 0.21fF
C5666 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C5667 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_3/A 0.32fF
C5668 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C5669 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C5670 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C5671 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C5672 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C5673 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# VDD 0.15fF
C5674 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.00fF
C5675 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C5676 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C5677 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C5678 sky130_fd_sc_hd__nand2_1_4/B VDD 2.14fF
C5679 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C5680 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VDD 0.18fF
C5681 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.01fF
C5682 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.03fF
C5683 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.52fF
C5684 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C5685 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.03fF
C5686 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C5687 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C5688 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.02fF
C5689 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C5690 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.13fF
C5691 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.01fF
C5692 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.03fF
C5693 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.02fF
C5694 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C5695 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C5696 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.01fF
C5697 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.01fF
C5698 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C5699 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VDD 0.42fF
C5700 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C5701 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C5702 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C5703 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C5704 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.01fF
C5705 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.05fF
C5706 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.05fF
C5707 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C5708 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C5709 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.04fF
C5710 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C5711 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C5712 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.02fF
C5713 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C5714 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C5715 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.02fF
C5716 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C5717 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C5718 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C5719 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C5720 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# VDD 0.14fF
C5721 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C5722 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# 0.00fF
C5723 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# 0.00fF
C5724 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C5725 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C5726 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C5727 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.00fF
C5728 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.00fF
C5729 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# VDD 0.16fF
C5730 Ad sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.06fF
C5731 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# A 0.06fF
C5732 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C5733 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.00fF
C5734 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.02fF
C5735 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.14fF
C5736 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.73fF
C5737 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# VDD 0.30fF
C5738 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C5739 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.00fF
C5740 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C5741 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# VDD 0.16fF
C5742 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C5743 sky130_fd_sc_hd__nand2_4_1/B Ad_b 0.06fF
C5744 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.16fF
C5745 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VDD 0.52fF
C5746 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C5747 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C5748 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.05fF
C5749 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# VDD 0.13fF
C5750 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C5751 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# VDD 0.23fF
C5752 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C5753 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.00fF
C5754 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C5755 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C5756 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.33fF
C5757 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.08fF
C5758 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.01fF
C5759 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.02fF
C5760 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.01fF
C5761 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.07fF
C5762 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.28fF
C5763 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C5764 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# VDD 0.15fF
C5765 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.01fF
C5766 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.01fF
C5767 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.01fF
C5768 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C5769 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C5770 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C5771 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.02fF
C5772 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.02fF
C5773 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.02fF
C5774 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C5775 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C5776 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5777 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# VDD 0.09fF
C5778 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C5779 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C5780 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C5781 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.02fF
C5782 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C5783 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.00fF
C5784 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C5785 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C5786 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# VDD 0.18fF
C5787 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C5788 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C5789 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.04fF
C5790 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.01fF
C5791 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C5792 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.02fF
C5793 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C5794 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C5795 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C5796 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C5797 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C5798 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.09fF
C5799 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.00fF
C5800 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.00fF
C5801 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C5802 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.01fF
C5803 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C5804 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C5805 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C5806 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C5807 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C5808 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C5809 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.01fF
C5810 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C5811 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C5812 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C5813 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.02fF
C5814 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C5815 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C5816 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VDD 0.16fF
C5817 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C5818 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.03fF
C5819 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C5820 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C5821 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.04fF
C5822 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.05fF
C5823 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C5824 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.01fF
C5825 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C5826 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VDD 0.34fF
C5827 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C5828 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.01fF
C5829 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.04fF
C5830 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.56fF
C5831 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C5832 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C5833 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C5834 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.15fF
C5835 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.03fF
C5836 sky130_fd_sc_hd__nand2_4_3/Y Ad_b 0.00fF
C5837 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.03fF
C5838 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C5839 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.01fF
C5840 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C5841 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C5842 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.01fF
C5843 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C5844 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C5845 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5846 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VDD 6.42fF
C5847 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C5848 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C5849 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.00fF
C5850 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C5851 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.01fF
C5852 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C5853 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.06fF
C5854 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.02fF
C5855 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C5856 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.08fF
C5857 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C5858 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C5859 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C5860 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C5861 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# 0.02fF
C5862 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.02fF
C5863 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.01fF
C5864 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.01fF
C5865 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.01fF
C5866 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.01fF
C5867 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C5868 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C5869 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.01fF
C5870 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C5871 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.02fF
C5872 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.01fF
C5873 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C5874 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C5875 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.01fF
C5876 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.44fF
C5877 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C5878 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.00fF
C5879 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C5880 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C5881 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C5882 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C5883 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.02fF
C5884 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.00fF
C5885 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.00fF
C5886 p2 sky130_fd_sc_hd__nand2_4_3/A 0.34fF
C5887 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.02fF
C5888 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.02fF
C5889 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.02fF
C5890 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C5891 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.06fF
C5892 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.02fF
C5893 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# 0.02fF
C5894 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.31fF
C5895 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C5896 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.06fF
C5897 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.09fF
C5898 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.07fF
C5899 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.14fF
C5900 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C5901 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.01fF
C5902 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.01fF
C5903 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C5904 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.15fF
C5905 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C5906 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C5907 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.00fF
C5908 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.01fF
C5909 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C5910 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C5911 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C5912 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C5913 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.01fF
C5914 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.29fF
C5915 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VDD 0.15fF
C5916 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C5917 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C5918 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C5919 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C5920 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C5921 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C5922 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C5923 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C5924 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.01fF
C5925 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.02fF
C5926 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.04fF
C5927 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.35fF
C5928 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C5929 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C5930 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.03fF
C5931 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.01fF
C5932 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.09fF
C5933 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.00fF
C5934 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C5935 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C5936 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C5937 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C5938 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.02fF
C5939 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.02fF
C5940 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.04fF
C5941 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.03fF
C5942 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C5943 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A sky130_fd_sc_hd__clkinv_1_0/Y 0.00fF
C5944 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.05fF
C5945 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C5946 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C5947 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# VDD 0.19fF
C5948 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/D 0.10fF
C5949 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C5950 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C5951 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C5952 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VDD 0.35fF
C5953 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C5954 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.03fF
C5955 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.02fF
C5956 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C5957 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.00fF
C5958 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C5959 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.00fF
C5960 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VDD 0.52fF
C5961 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C5962 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.00fF
C5963 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C5964 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_1_1/B 0.05fF
C5965 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C5966 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C5967 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.01fF
C5968 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.01fF
C5969 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD 0.23fF
C5970 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C5971 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C5972 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.11fF
C5973 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C5974 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.01fF
C5975 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C5976 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.02fF
C5977 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.01fF
C5978 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C5979 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C5980 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C5981 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C5982 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.00fF
C5983 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.09fF
C5984 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5985 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.01fF
C5986 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.00fF
C5987 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.00fF
C5988 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.05fF
C5989 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C5990 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.00fF
C5991 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.01fF
C5992 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# 0.00fF
C5993 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.11fF
C5994 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.09fF
C5995 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.01fF
C5996 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.16fF
C5997 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.04fF
C5998 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C5999 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C6000 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.01fF
C6001 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.23fF
C6002 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C6003 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C6004 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.01fF
C6005 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C6006 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.01fF
C6007 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VDD 0.42fF
C6008 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C6009 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C6010 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.29fF
C6011 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Ad_b 0.03fF
C6012 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.01fF
C6013 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C6014 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.01fF
C6015 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.01fF
C6016 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C6017 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# 0.05fF
C6018 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C6019 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C6020 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.00fF
C6021 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.03fF
C6022 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C6023 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# VDD 0.13fF
C6024 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C6025 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C6026 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C6027 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkinv_4_5/Y 0.03fF
C6028 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C6029 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# 0.01fF
C6030 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.00fF
C6031 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__nand2_1_2/B 0.03fF
C6032 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C6033 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# VDD 0.19fF
C6034 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C6035 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.00fF
C6036 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# VDD 0.11fF
C6037 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C6038 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C6039 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C6040 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C6041 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.01fF
C6042 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.04fF
C6043 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.04fF
C6044 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C6045 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C6046 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C6047 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C6048 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C6049 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.00fF
C6050 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.00fF
C6051 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.01fF
C6052 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# VDD 0.32fF
C6053 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# VDD 0.17fF
C6054 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# 0.05fF
C6055 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.02fF
C6056 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C6057 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C6058 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.03fF
C6059 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.01fF
C6060 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C6061 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C6062 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C6063 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.03fF
C6064 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.03fF
C6065 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# VDD 0.40fF
C6066 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C6067 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C6068 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkinv_4_5/Y 0.85fF
C6069 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.07fF
C6070 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VDD 0.13fF
C6071 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 1.69fF
C6072 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.01fF
C6073 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.01fF
C6074 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.11fF
C6075 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# VDD 0.12fF
C6076 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C6077 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.02fF
C6078 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1d_b 0.10fF
C6079 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.11fF
C6080 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C6081 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.00fF
C6082 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C6083 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.01fF
C6084 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.02fF
C6085 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.19fF
C6086 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.03fF
C6087 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.01fF
C6088 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# VDD 0.33fF
C6089 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.08fF
C6090 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.00fF
C6091 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.00fF
C6092 p2 sky130_fd_sc_hd__clkinv_4_3/Y 0.03fF
C6093 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.11fF
C6094 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C6095 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.09fF
C6096 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.01fF
C6097 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C6098 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C6099 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C6100 sky130_fd_sc_hd__nand2_4_3/A Ad_b 0.32fF
C6101 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.06fF
C6102 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# 0.01fF
C6103 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.01fF
C6104 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VDD 0.28fF
C6105 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# 0.03fF
C6106 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.02fF
C6107 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.02fF
C6108 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__nand2_4_2/A 0.42fF
C6109 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C6110 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C6111 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.01fF
C6112 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.08fF
C6113 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C6114 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.12fF
C6115 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.09fF
C6116 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C6117 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C6118 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.01fF
C6119 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C6120 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C6121 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.04fF
C6122 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.03fF
C6123 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_561_413# 0.01fF
C6124 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.03fF
C6125 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.01fF
C6126 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.02fF
C6127 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C6128 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C6129 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C6130 VDD p1d 1.51fF
C6131 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C6132 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C6133 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C6134 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C6135 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C6136 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C6137 sky130_fd_sc_hd__nand2_1_1/A VDD 13.45fF
C6138 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.07fF
C6139 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/D 0.91fF
C6140 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.02fF
C6141 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C6142 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C6143 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.01fF
C6144 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C6145 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.07fF
C6146 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.05fF
C6147 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.05fF
C6148 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C6149 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C6150 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VDD 0.34fF
C6151 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.00fF
C6152 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.10fF
C6153 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C6154 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C6155 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.11fF
C6156 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C6157 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.00fF
C6158 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.00fF
C6159 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C6160 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.03fF
C6161 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.05fF
C6162 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C6163 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.01fF
C6164 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C6165 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.02fF
C6166 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.04fF
C6167 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.04fF
C6168 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.37fF
C6169 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# VDD 0.13fF
C6170 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C6171 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.01fF
C6172 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.03fF
C6173 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.01fF
C6174 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C6175 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C6176 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C6177 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C6178 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.04fF
C6179 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# VDD 0.18fF
C6180 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C6181 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C6182 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.09fF
C6183 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C6184 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C6185 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C6186 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C6187 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.02fF
C6188 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.00fF
C6189 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C6190 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.02fF
C6191 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# VDD 0.33fF
C6192 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.06fF
C6193 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.03fF
C6194 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C6195 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C6196 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C6197 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.03fF
C6198 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.03fF
C6199 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C6200 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C6201 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C6202 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C6203 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C6204 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C6205 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.01fF
C6206 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.00fF
C6207 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C6208 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.01fF
C6209 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C6210 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.02fF
C6211 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C6212 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C6213 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C6214 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.02fF
C6215 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.02fF
C6216 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C6217 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C6218 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.06fF
C6219 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# VDD 0.14fF
C6220 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.82fF
C6221 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C6222 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C6223 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C6224 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.00fF
C6225 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C6226 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C6227 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C6228 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C6229 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.04fF
C6230 Ad A_b 0.53fF
C6231 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C6232 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.02fF
C6233 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.51fF
C6234 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.04fF
C6235 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# VDD 0.15fF
C6236 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_4_5/Y 0.45fF
C6237 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.06fF
C6238 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.02fF
C6239 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.02fF
C6240 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# 0.05fF
C6241 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.01fF
C6242 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Ad_b 0.22fF
C6243 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.01fF
C6244 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.02fF
C6245 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C6246 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C6247 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.02fF
C6248 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# VDD 0.17fF
C6249 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C6250 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C6251 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.01fF
C6252 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C6253 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.02fF
C6254 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# VDD 0.35fF
C6255 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C6256 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C6257 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.00fF
C6258 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.00fF
C6259 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C6260 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C6261 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C6262 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C6263 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.09fF
C6264 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.01fF
C6265 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.04fF
C6266 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.04fF
C6267 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C6268 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.00fF
C6269 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.04fF
C6270 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.01fF
C6271 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C6272 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.02fF
C6273 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C6274 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C6275 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C6276 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C6277 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C6278 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C6279 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C6280 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.01fF
C6281 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# 0.02fF
C6282 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.00fF
C6283 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C6284 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.00fF
C6285 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0.07fF
C6286 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.02fF
C6287 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.02fF
C6288 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.37fF
C6289 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.02fF
C6290 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.03fF
C6291 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C6292 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.03fF
C6293 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_9/Y 0.68fF
C6294 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.14fF
C6295 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.01fF
C6296 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.01fF
C6297 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.02fF
C6298 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C6299 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.01fF
C6300 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.02fF
C6301 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.01fF
C6302 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C6303 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C6304 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C6305 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.02fF
C6306 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VDD 0.14fF
C6307 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.07fF
C6308 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C6309 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C6310 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# 0.05fF
C6311 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.02fF
C6312 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C6313 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C6314 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C6315 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C6316 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.14fF
C6317 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C6318 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C6319 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VDD 0.63fF
C6320 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.00fF
C6321 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C6322 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C6323 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.02fF
C6324 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.00fF
C6325 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.01fF
C6326 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C6327 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.00fF
C6328 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.06fF
C6329 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C6330 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C6331 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C6332 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.00fF
C6333 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C6334 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.08fF
C6335 p2d_b p2_b 0.22fF
C6336 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkinv_4_9/Y 0.04fF
C6337 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C6338 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C6339 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.02fF
C6340 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C6341 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.00fF
C6342 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.01fF
C6343 sky130_fd_sc_hd__clkinv_4_3/Y Ad_b 0.07fF
C6344 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.06fF
C6345 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.69fF
C6346 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C6347 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.28fF
C6348 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.03fF
C6349 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.00fF
C6350 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C6351 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C6352 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C6353 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.09fF
C6354 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C6355 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.04fF
C6356 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C6357 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.11fF
C6358 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C6359 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C6360 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C6361 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.00fF
C6362 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C6363 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C6364 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C6365 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# 0.00fF
C6366 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C6367 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.03fF
C6368 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C6369 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C6370 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.01fF
C6371 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C6372 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C6373 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VDD 0.58fF
C6374 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.09fF
C6375 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.00fF
C6376 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.01fF
C6377 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C6378 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C6379 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.01fF
C6380 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C6381 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_1/A 0.03fF
C6382 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.02fF
C6383 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.01fF
C6384 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.02fF
C6385 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C6386 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.02fF
C6387 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.07fF
C6388 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C6389 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# VDD 0.29fF
C6390 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C6391 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.03fF
C6392 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# VDD 0.28fF
C6393 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C6394 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.44fF
C6395 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.00fF
C6396 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.01fF
C6397 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.02fF
C6398 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C6399 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C6400 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.02fF
C6401 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C6402 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C6403 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C6404 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C6405 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C6406 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C6407 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C6408 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C6409 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C6410 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.00fF
C6411 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.02fF
C6412 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.02fF
C6413 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.00fF
C6414 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C6415 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.11fF
C6416 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.02fF
C6417 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.06fF
C6418 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.08fF
C6419 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.33fF
C6420 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.01fF
C6421 sky130_fd_sc_hd__nand2_4_0/a_27_47# VDD 0.04fF
C6422 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.14fF
C6423 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C6424 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C6425 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C6426 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.00fF
C6427 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.03fF
C6428 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C6429 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C6430 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A Bd_b 0.00fF
C6431 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C6432 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.01fF
C6433 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.11fF
C6434 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# 0.01fF
C6435 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C6436 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.02fF
C6437 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C6438 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0.03fF
C6439 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.14fF
C6440 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# VDD 0.32fF
C6441 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.01fF
C6442 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.01fF
C6443 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.02fF
C6444 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C6445 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C6446 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_4/Y -0.43fF
C6447 B sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.02fF
C6448 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VDD -0.76fF
C6449 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.00fF
C6450 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.09fF
C6451 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# 0.01fF
C6452 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C6453 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C6454 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.09fF
C6455 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C6456 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.00fF
C6457 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C6458 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C6459 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C6460 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.01fF
C6461 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C6462 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C6463 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.00fF
C6464 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.00fF
C6465 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C6466 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# 0.05fF
C6467 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C6468 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# 0.05fF
C6469 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C6470 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.09fF
C6471 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.00fF
C6472 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# 0.00fF
C6473 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C6474 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C6475 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C6476 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# 0.01fF
C6477 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C6478 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C6479 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C6480 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.04fF
C6481 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.04fF
C6482 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C6483 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C6484 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.04fF
C6485 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.01fF
C6486 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VDD 0.51fF
C6487 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.00fF
C6488 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.00fF
C6489 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C6490 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C6491 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C6492 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.03fF
C6493 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C6494 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VDD 0.59fF
C6495 p2 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# -0.00fF
C6496 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VDD 0.66fF
C6497 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C6498 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.01fF
C6499 p1d_b sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.02fF
C6500 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1 0.02fF
C6501 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C6502 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.04fF
C6503 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.52fF
C6504 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# 0.02fF
C6505 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.01fF
C6506 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C6507 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.02fF
C6508 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.01fF
C6509 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C6510 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C6511 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C6512 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.23fF
C6513 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C6514 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C6515 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C6516 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# Bd_b 0.00fF
C6517 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/X 0.01fF
C6518 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C6519 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C6520 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C6521 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C6522 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C6523 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C6524 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C6525 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# 0.02fF
C6526 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# 0.02fF
C6527 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C6528 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C6529 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C6530 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.03fF
C6531 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VDD 0.14fF
C6532 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C6533 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VDD 0.17fF
C6534 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.00fF
C6535 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.01fF
C6536 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C6537 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C6538 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C6539 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# 0.04fF
C6540 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# 0.04fF
C6541 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.23fF
C6542 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C6543 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.00fF
C6544 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# VDD 0.14fF
C6545 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# VDD 0.14fF
C6546 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C6547 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.02fF
C6548 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# 0.01fF
C6549 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# VDD 0.16fF
C6550 sky130_fd_sc_hd__nand2_4_3/B VDD 0.58fF
C6551 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# VDD 0.14fF
C6552 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C6553 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# VDD 0.16fF
C6554 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C6555 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C6556 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.01fF
C6557 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# VDD 0.34fF
C6558 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C6559 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C6560 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C6561 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/B 0.14fF
C6562 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.02fF
C6563 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.01fF
C6564 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.01fF
C6565 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.09fF
C6566 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# VDD 0.33fF
C6567 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# VDD 0.29fF
C6568 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.02fF
C6569 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.01fF
C6570 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C6571 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.04fF
C6572 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.04fF
C6573 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.32fF
C6574 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.02fF
C6575 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkinv_4_2/Y 0.03fF
C6576 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C6577 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C6578 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.02fF
C6579 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.02fF
C6580 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C6581 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.02fF
C6582 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VDD 0.22fF
C6583 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.00fF
C6584 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.00fF
C6585 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C6586 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C6587 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.04fF
C6588 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# 0.09fF
C6589 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C6590 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C6591 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C6592 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.04fF
C6593 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.02fF
C6594 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# 0.02fF
C6595 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.02fF
C6596 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.01fF
C6597 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# 0.00fF
C6598 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X VDD 0.69fF
C6599 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.04fF
C6600 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.04fF
C6601 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.04fF
C6602 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.00fF
C6603 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C6604 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkinv_4_1/A 0.06fF
C6605 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C6606 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.02fF
C6607 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.04fF
C6608 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.04fF
C6609 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C6610 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C6611 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VDD 0.42fF
C6612 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.69fF
C6613 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__mux2_1_0/S 0.02fF
C6614 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X VDD 0.51fF
C6615 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.01fF
C6616 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.05fF
C6617 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.05fF
C6618 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.03fF
C6619 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__nand2_4_2/A 0.05fF
C6620 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VDD 0.15fF
C6621 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.02fF
C6622 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.02fF
C6623 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.02fF
C6624 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# 0.02fF
C6625 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.01fF
C6626 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.02fF
C6627 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C6628 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C6629 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.00fF
C6630 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C6631 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.01fF
C6632 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkinv_4_7/A 0.32fF
C6633 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.04fF
C6634 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.04fF
C6635 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.09fF
C6636 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C6637 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.05fF
C6638 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C6639 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C6640 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.02fF
C6641 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.08fF
C6642 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.00fF
C6643 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.00fF
C6644 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C6645 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C6646 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.03fF
C6647 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C6648 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C6649 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C6650 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C6651 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C6652 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/X 0.00fF
C6653 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C6654 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C6655 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C6656 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C6657 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.03fF
C6658 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C6659 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C6660 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C6661 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.02fF
C6662 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# 0.02fF
C6663 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C6664 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C6665 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# VDD 0.15fF
C6666 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C6667 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.01fF
C6668 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C6669 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.02fF
C6670 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.04fF
C6671 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.03fF
C6672 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A VDD 0.57fF
C6673 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# VDD 0.16fF
C6674 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.04fF
C6675 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.04fF
C6676 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C6677 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.01fF
C6678 sky130_fd_sc_hd__nand2_4_1/B Bd_b 0.07fF
C6679 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# VDD 0.12fF
C6680 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C6681 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C6682 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C6683 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C6684 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkinv_1_0/Y 0.77fF
C6685 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.15fF
C6686 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C6687 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.04fF
C6688 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# VDD 0.34fF
C6689 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.06fF
C6690 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# Ad_b 0.01fF
C6691 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C6692 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.00fF
C6693 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# VDD 0.12fF
C6694 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C6695 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C6696 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.02fF
C6697 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.02fF
C6698 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.16fF
C6699 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.02fF
C6700 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.02fF
C6701 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.01fF
C6702 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.01fF
C6703 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C6704 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.00fF
C6705 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C6706 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.00fF
C6707 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C6708 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.07fF
C6709 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.02fF
C6710 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.02fF
C6711 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C6712 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C6713 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# VDD 0.10fF
C6714 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.04fF
C6715 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.04fF
C6716 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.02fF
C6717 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C6718 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.04fF
C6719 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# VDD 0.05fF
C6720 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C6721 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkinv_1_2/Y 0.02fF
C6722 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.01fF
C6723 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.01fF
C6724 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C6725 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C6726 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkinv_4_7/A 1.80fF
C6727 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.02fF
C6728 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.04fF
C6729 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# 0.09fF
C6730 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C6731 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C6732 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# 0.04fF
C6733 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.04fF
C6734 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.02fF
C6735 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C6736 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C6737 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.06fF
C6738 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.03fF
C6739 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.01fF
C6740 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.00fF
C6741 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.00fF
C6742 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C6743 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C6744 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.00fF
C6745 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.13fF
C6746 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.03fF
C6747 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C6748 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.01fF
C6749 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.02fF
C6750 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.02fF
C6751 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C6752 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.00fF
C6753 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.06fF
C6754 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C6755 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C6756 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.01fF
C6757 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C6758 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.04fF
C6759 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.04fF
C6760 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__nand2_4_2/B 0.04fF
C6761 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.04fF
C6762 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.04fF
C6763 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.01fF
C6764 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.02fF
C6765 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C6766 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VDD 0.14fF
C6767 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C6768 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.00fF
C6769 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C6770 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C6771 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C6772 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.01fF
C6773 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.02fF
C6774 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.02fF
C6775 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C6776 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C6777 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C6778 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VDD 0.18fF
C6779 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C6780 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C6781 sky130_fd_sc_hd__nand2_4_0/Y VDD 5.50fF
C6782 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C6783 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C6784 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.34fF
C6785 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C6786 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.02fF
C6787 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C6788 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.09fF
C6789 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C6790 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_1/A 0.31fF
C6791 sky130_fd_sc_hd__nand2_4_3/Y Bd_b 0.00fF
C6792 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# 0.03fF
C6793 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.03fF
C6794 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.01fF
C6795 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.05fF
C6796 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C6797 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C6798 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C6799 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.01fF
C6800 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.02fF
C6801 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C6802 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C6803 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.02fF
C6804 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C6805 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C6806 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.01fF
C6807 sky130_fd_sc_hd__nand2_1_2/B clk 0.04fF
C6808 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C6809 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C6810 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C6811 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C6812 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.00fF
C6813 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.00fF
C6814 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.00fF
C6815 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C6816 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.01fF
C6817 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C6818 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.00fF
C6819 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.02fF
C6820 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C6821 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.01fF
C6822 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.02fF
C6823 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C6824 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C6825 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.00fF
C6826 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.00fF
C6827 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.00fF
C6828 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.00fF
C6829 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C6830 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C6831 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.02fF
C6832 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C6833 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C6834 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C6835 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C6836 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.02fF
C6837 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.00fF
C6838 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C6839 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# 0.00fF
C6840 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.00fF
C6841 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.00fF
C6842 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.02fF
C6843 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.02fF
C6844 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.30fF
C6845 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.04fF
C6846 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.00fF
C6847 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# 0.09fF
C6848 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.01fF
C6849 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.00fF
C6850 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.07fF
C6851 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C6852 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C6853 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.06fF
C6854 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.05fF
C6855 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.02fF
C6856 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C6857 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C6858 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C6859 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C6860 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.06fF
C6861 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C6862 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.05fF
C6863 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C6864 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C6865 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.14fF
C6866 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.03fF
C6867 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.09fF
C6868 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C6869 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C6870 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.01fF
C6871 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C6872 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C6873 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.05fF
C6874 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C6875 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C6876 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.04fF
C6877 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.17fF
C6878 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.02fF
C6879 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C6880 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C6881 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.01fF
C6882 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C6883 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.01fF
C6884 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C6885 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C6886 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.04fF
C6887 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1 -0.03fF
C6888 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C6889 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.02fF
C6890 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C6891 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C6892 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.57fF
C6893 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.02fF
C6894 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C6895 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.08fF
C6896 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C6897 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C6898 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C6899 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C6900 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_4/Y 0.06fF
C6901 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.02fF
C6902 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.02fF
C6903 p2d_b p2d 0.52fF
C6904 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C6905 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C6906 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C6907 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# VDD 0.10fF
C6908 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C6909 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.02fF
C6910 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C6911 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C6912 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C6913 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C6914 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.00fF
C6915 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/D 0.08fF
C6916 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.01fF
C6917 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.04fF
C6918 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.04fF
C6919 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Ad_b 0.03fF
C6920 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.01fF
C6921 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.02fF
C6922 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.02fF
C6923 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A VDD 0.56fF
C6924 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.03fF
C6925 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C6926 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.03fF
C6927 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C6928 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C6929 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.00fF
C6930 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C6931 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C6932 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C6933 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.03fF
C6934 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C6935 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.02fF
C6936 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C6937 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.00fF
C6938 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.00fF
C6939 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C6940 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.00fF
C6941 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C6942 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A VDD 0.57fF
C6943 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C6944 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.00fF
C6945 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C6946 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C6947 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.07fF
C6948 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C6949 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C6950 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C6951 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.03fF
C6952 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C6953 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C6954 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.08fF
C6955 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C6956 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C6957 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.04fF
C6958 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C6959 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C6960 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.01fF
C6961 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_4/B 0.40fF
C6962 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C6963 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.02fF
C6964 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C6965 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.05fF
C6966 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C6967 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C6968 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C6969 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.03fF
C6970 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C6971 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.56fF
C6972 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.08fF
C6973 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# 0.00fF
C6974 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.00fF
C6975 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.01fF
C6976 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.15fF
C6977 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C6978 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.02fF
C6979 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C6980 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.01fF
C6981 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.02fF
C6982 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.02fF
C6983 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.12fF
C6984 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C6985 sky130_fd_sc_hd__dfxbp_1_1/D VDD 0.61fF
C6986 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C6987 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.03fF
C6988 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.02fF
C6989 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C6990 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C6991 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C6992 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.15fF
C6993 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Bd_b 0.03fF
C6994 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C6995 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C6996 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.30fF
C6997 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.01fF
C6998 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# 0.01fF
C6999 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.03fF
C7000 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C7001 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C7002 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C7003 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C7004 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C7005 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C7006 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C7007 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C7008 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C7009 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.07fF
C7010 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C7011 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.02fF
C7012 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# VDD 0.15fF
C7013 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.02fF
C7014 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.01fF
C7015 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.01fF
C7016 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.02fF
C7017 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C7018 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C7019 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C7020 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C7021 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.02fF
C7022 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.03fF
C7023 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C7024 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C7025 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.03fF
C7026 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C7027 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.01fF
C7028 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.02fF
C7029 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.00fF
C7030 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.00fF
C7031 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.00fF
C7032 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C7033 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C7034 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C7035 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# VDD 0.15fF
C7036 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.02fF
C7037 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# VDD 0.14fF
C7038 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.01fF
C7039 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C7040 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.02fF
C7041 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C7042 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C7043 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C7044 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C7045 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C7046 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C7047 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C7048 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.06fF
C7049 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.01fF
C7050 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.02fF
C7051 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# VDD 0.22fF
C7052 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# VDD 0.29fF
C7053 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.03fF
C7054 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.01fF
C7055 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C7056 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C7057 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C7058 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C7059 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.03fF
C7060 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VDD 0.10fF
C7061 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.02fF
C7062 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.00fF
C7063 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.04fF
C7064 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.05fF
C7065 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.01fF
C7066 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C7067 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C7068 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.06fF
C7069 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.06fF
C7070 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.00fF
C7071 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C7072 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C7073 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.01fF
C7074 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.02fF
C7075 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C7076 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.14fF
C7077 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C7078 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.03fF
C7079 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.01fF
C7080 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# VDD 0.19fF
C7081 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.04fF
C7082 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.00fF
C7083 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C7084 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2 0.02fF
C7085 p2d_b sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.03fF
C7086 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C7087 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VDD 0.56fF
C7088 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C7089 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C7090 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C7091 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C7092 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# VDD 0.31fF
C7093 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.01fF
C7094 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C7095 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C7096 sky130_fd_sc_hd__nand2_4_3/A Bd_b 0.27fF
C7097 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.01fF
C7098 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.01fF
C7099 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C7100 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C7101 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.03fF
C7102 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# 0.01fF
C7103 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C7104 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C7105 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C7106 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C7107 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C7108 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.02fF
C7109 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.11fF
C7110 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.05fF
C7111 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.11fF
C7112 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.00fF
C7113 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.00fF
C7114 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C7115 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.01fF
C7116 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C7117 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.00fF
C7118 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.00fF
C7119 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.02fF
C7120 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.01fF
C7121 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C7122 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C7123 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C7124 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C7125 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.01fF
C7126 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C7127 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C7128 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.01fF
C7129 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.09fF
C7130 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.05fF
C7131 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.05fF
C7132 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.00fF
C7133 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X VDD 0.68fF
C7134 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.04fF
C7135 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.04fF
C7136 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.04fF
C7137 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C7138 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.09fF
C7139 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C7140 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.09fF
C7141 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C7142 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.03fF
C7143 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C7144 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C7145 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.02fF
C7146 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.01fF
C7147 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.01fF
C7148 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.02fF
C7149 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C7150 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C7151 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C7152 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.00fF
C7153 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.07fF
C7154 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C7155 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C7156 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C7157 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.03fF
C7158 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C7159 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__nand2_1_1/A 0.03fF
C7160 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.09fF
C7161 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.00fF
C7162 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.04fF
C7163 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C7164 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C7165 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C7166 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C7167 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C7168 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.01fF
C7169 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C7170 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.01fF
C7171 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C7172 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# 0.11fF
C7173 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# VDD 0.15fF
C7174 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.02fF
C7175 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.05fF
C7176 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.05fF
C7177 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C7178 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C7179 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# 0.00fF
C7180 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C7181 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C7182 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C7183 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C7184 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C7185 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# VDD 0.14fF
C7186 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C7187 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__nand2_1_1/A 0.07fF
C7188 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.04fF
C7189 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.04fF
C7190 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C7191 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# VDD 0.24fF
C7192 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.06fF
C7193 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.04fF
C7194 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C7195 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__nand2_1_2/B 0.00fF
C7196 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C7197 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C7198 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C7199 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.01fF
C7200 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.01fF
C7201 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C7202 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.04fF
C7203 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.04fF
C7204 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C7205 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C7206 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C7207 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C7208 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C7209 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.01fF
C7210 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C7211 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clk 0.05fF
C7212 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.04fF
C7213 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.04fF
C7214 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# VDD 0.14fF
C7215 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C7216 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VDD 0.37fF
C7217 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C7218 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C7219 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Bd_b 0.10fF
C7220 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.02fF
C7221 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.00fF
C7222 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.01fF
C7223 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C7224 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C7225 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C7226 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C7227 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.00fF
C7228 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.00fF
C7229 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# VDD 0.17fF
C7230 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C7231 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C7232 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C7233 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C7234 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# VDD 0.30fF
C7235 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkinv_4_5/Y 0.05fF
C7236 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.02fF
C7237 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.01fF
C7238 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# VDD 0.28fF
C7239 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.01fF
C7240 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.01fF
C7241 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.01fF
C7242 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C7243 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C7244 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.00fF
C7245 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.00fF
C7246 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C7247 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_72/X 0.01fF
C7248 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C7249 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C7250 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C7251 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.01fF
C7252 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C7253 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.02fF
C7254 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD 0.25fF
C7255 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C7256 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.10fF
C7257 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C7258 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkinv_4_1/A 0.01fF
C7259 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.07fF
C7260 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0.06fF
C7261 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C7262 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.01fF
C7263 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C7264 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.09fF
C7265 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.02fF
C7266 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.02fF
C7267 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.01fF
C7268 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C7269 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.02fF
C7270 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.00fF
C7271 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C7272 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C7273 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C7274 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.01fF
C7275 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.09fF
C7276 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C7277 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.01fF
C7278 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C7279 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.00fF
C7280 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C7281 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C7282 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C7283 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C7284 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.06fF
C7285 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.02fF
C7286 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.01fF
C7287 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.02fF
C7288 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkinv_1_3/Y 0.02fF
C7289 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C7290 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C7291 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C7292 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C7293 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.06fF
C7294 sky130_fd_sc_hd__nand2_1_4/B Ad_b 0.02fF
C7295 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C7296 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.04fF
C7297 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.04fF
C7298 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VDD 0.59fF
C7299 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.00fF
C7300 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.00fF
C7301 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C7302 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C7303 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C7304 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.07fF
C7305 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C7306 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.01fF
C7307 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C7308 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C7309 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_4_1/A 1.35fF
C7310 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C7311 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.00fF
C7312 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.00fF
C7313 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.00fF
C7314 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.01fF
C7315 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C7316 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C7317 sky130_fd_sc_hd__clkinv_4_3/Y Bd_b 0.18fF
C7318 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.01fF
C7319 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C7320 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C7321 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.06fF
C7322 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.02fF
C7323 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C7324 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.02fF
C7325 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C7326 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.02fF
C7327 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C7328 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C7329 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.02fF
C7330 sky130_fd_sc_hd__clkinv_4_4/Y Bd_b 0.08fF
C7331 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# VDD 0.38fF
C7332 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.02fF
C7333 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C7334 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# Bd_b 0.06fF
C7335 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C7336 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C7337 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.03fF
C7338 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C7339 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.01fF
C7340 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.03fF
C7341 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.00fF
C7342 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C7343 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.07fF
C7344 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# 0.01fF
C7345 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C7346 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.01fF
C7347 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.01fF
C7348 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.02fF
C7349 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.02fF
C7350 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C7351 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C7352 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__mux2_1_0/X 0.05fF
C7353 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C7354 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C7355 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C7356 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.02fF
C7357 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C7358 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.01fF
C7359 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_1_0/B 0.06fF
C7360 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C7361 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.04fF
C7362 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C7363 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X Ad_b 0.02fF
C7364 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C7365 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C7366 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C7367 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C7368 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C7369 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C7370 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.02fF
C7371 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.03fF
C7372 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.03fF
C7373 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C7374 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.08fF
C7375 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# VDD 0.33fF
C7376 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# VDD 0.13fF
C7377 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C7378 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C7379 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.02fF
C7380 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.01fF
C7381 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C7382 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C7383 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C7384 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C7385 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C7386 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.01fF
C7387 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C7388 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.02fF
C7389 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C7390 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C7391 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.02fF
C7392 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.00fF
C7393 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.01fF
C7394 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.03fF
C7395 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C7396 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C7397 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.05fF
C7398 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.14fF
C7399 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.11fF
C7400 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.06fF
C7401 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.09fF
C7402 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C7403 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.07fF
C7404 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C7405 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.31fF
C7406 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.44fF
C7407 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C7408 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C7409 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C7410 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# A_b 0.06fF
C7411 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.09fF
C7412 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# 0.02fF
C7413 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# 0.01fF
C7414 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C7415 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C7416 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C7417 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C7418 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# 0.05fF
C7419 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.04fF
C7420 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# VDD 0.17fF
C7421 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.02fF
C7422 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C7423 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C7424 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C7425 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C7426 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C7427 B VDD 1.54fF
C7428 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.09fF
C7429 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.05fF
C7430 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.01fF
C7431 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C7432 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.06fF
C7433 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C7434 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.06fF
C7435 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C7436 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C7437 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.44fF
C7438 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C7439 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C7440 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.02fF
C7441 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.02fF
C7442 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# 0.03fF
C7443 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C7444 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.66fF
C7445 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.00fF
C7446 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.01fF
C7447 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.08fF
C7448 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# 0.00fF
C7449 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.01fF
C7450 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C7451 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C7452 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A VDD 0.57fF
C7453 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C7454 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C7455 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.00fF
C7456 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C7457 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C7458 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X VDD 0.57fF
C7459 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.04fF
C7460 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.00fF
C7461 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C7462 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C7463 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C7464 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C7465 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C7466 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C7467 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C7468 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C7469 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.00fF
C7470 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.03fF
C7471 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.08fF
C7472 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.07fF
C7473 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.03fF
C7474 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C7475 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.08fF
C7476 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.04fF
C7477 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.00fF
C7478 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# 0.02fF
C7479 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.01fF
C7480 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VDD 0.49fF
C7481 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.01fF
C7482 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.01fF
C7483 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.05fF
C7484 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C7485 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.03fF
C7486 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.01fF
C7487 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C7488 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C7489 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C7490 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# VDD 0.33fF
C7491 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C7492 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C7493 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.31fF
C7494 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.01fF
C7495 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C7496 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C7497 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C7498 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C7499 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C7500 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C7501 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.02fF
C7502 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C7503 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.03fF
C7504 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.11fF
C7505 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VDD 0.14fF
C7506 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C7507 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.01fF
C7508 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/A 0.03fF
C7509 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.01fF
C7510 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.02fF
C7511 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C7512 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.05fF
C7513 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.08fF
C7514 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C7515 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C7516 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C7517 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# 0.01fF
C7518 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# 0.01fF
C7519 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# 0.02fF
C7520 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.02fF
C7521 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.02fF
C7522 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C7523 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.00fF
C7524 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C7525 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.02fF
C7526 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C7527 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.03fF
C7528 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C7529 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.09fF
C7530 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# 0.01fF
C7531 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# 0.02fF
C7532 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD 0.52fF
C7533 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# VDD 0.15fF
C7534 p2 sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C7535 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C7536 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# VDD 0.15fF
C7537 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# VDD 0.14fF
C7538 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C7539 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C7540 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C7541 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# VDD 0.17fF
C7542 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.02fF
C7543 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.02fF
C7544 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.09fF
C7545 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# VDD 0.15fF
C7546 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.03fF
C7547 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.02fF
C7548 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# VDD 0.17fF
C7549 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.00fF
C7550 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C7551 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.01fF
C7552 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.02fF
C7553 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.00fF
C7554 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C7555 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.03fF
C7556 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C7557 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.03fF
C7558 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C7559 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C7560 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C7561 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C7562 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C7563 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.58fF
C7564 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.14fF
C7565 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# VDD 0.30fF
C7566 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.10fF
C7567 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.04fF
C7568 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.04fF
C7569 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C7570 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C7571 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.05fF
C7572 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C7573 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C7574 VDD sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.45fF
C7575 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.31fF
C7576 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.06fF
C7577 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.01fF
C7578 VDD sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.14fF
C7579 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.11fF
C7580 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# 0.10fF
C7581 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C7582 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C7583 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C7584 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.01fF
C7585 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.01fF
C7586 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.02fF
C7587 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C7588 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C7589 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.04fF
C7590 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C7591 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkinv_4_1/A 0.05fF
C7592 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.02fF
C7593 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.01fF
C7594 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.01fF
C7595 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.01fF
C7596 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.06fF
C7597 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C7598 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.02fF
C7599 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.00fF
C7600 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.02fF
C7601 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.01fF
C7602 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.01fF
C7603 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.01fF
C7604 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VDD 0.56fF
C7605 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C7606 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.03fF
C7607 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.41fF
C7608 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.09fF
C7609 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C7610 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C7611 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C7612 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C7613 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/X 0.00fF
C7614 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C7615 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.02fF
C7616 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Ad_b 0.02fF
C7617 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.01fF
C7618 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C7619 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.02fF
C7620 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C7621 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.01fF
C7622 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.02fF
C7623 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# VDD 0.34fF
C7624 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C7625 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C7626 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C7627 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.01fF
C7628 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.03fF
C7629 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.00fF
C7630 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C7631 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C7632 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C7633 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C7634 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.00fF
C7635 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.00fF
C7636 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C7637 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_12/a_110_47# 0.04fF
C7638 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C7639 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C7640 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.02fF
C7641 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.04fF
C7642 VDD sky130_fd_sc_hd__mux2_1_0/S -0.30fF
C7643 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.32fF
C7644 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C7645 VDD sky130_fd_sc_hd__clkinv_4_2/Y 1.52fF
C7646 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# Ad_b 0.02fF
C7647 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.02fF
C7648 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C7649 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.00fF
C7650 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C7651 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.02fF
C7652 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.04fF
C7653 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.03fF
C7654 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C7655 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C7656 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C7657 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.03fF
C7658 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.01fF
C7659 Bd Bd_b 0.47fF
C7660 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C7661 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C7662 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.31fF
C7663 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C7664 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C7665 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C7666 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C7667 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C7668 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C7669 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.01fF
C7670 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.04fF
C7671 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.00fF
C7672 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.00fF
C7673 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.03fF
C7674 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.03fF
C7675 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C7676 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.01fF
C7677 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C7678 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.07fF
C7679 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.01fF
C7680 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.06fF
C7681 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# VDD 0.15fF
C7682 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkinv_4_7/A 0.02fF
C7683 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C7684 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C7685 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.02fF
C7686 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C7687 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.01fF
C7688 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C7689 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C7690 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.01fF
C7691 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.03fF
C7692 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__nand2_1_3/A 0.03fF
C7693 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C7694 sky130_fd_sc_hd__nand2_1_3/A clk 0.02fF
C7695 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C7696 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C7697 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C7698 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C7699 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.00fF
C7700 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C7701 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C7702 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# Ad_b 0.00fF
C7703 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# VDD 0.19fF
C7704 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.00fF
C7705 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C7706 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.00fF
C7707 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.09fF
C7708 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.00fF
C7709 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.00fF
C7710 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# VDD 0.10fF
C7711 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/S 0.06fF
C7712 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# Ad_b 0.00fF
C7713 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# Bd_b 0.01fF
C7714 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X Bd_b 0.00fF
C7715 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.13fF
C7716 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C7717 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C7718 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C7719 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C7720 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.05fF
C7721 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C7722 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.01fF
C7723 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.08fF
C7724 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.04fF
C7725 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.04fF
C7726 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.00fF
C7727 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C7728 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C7729 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C7730 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C7731 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.01fF
C7732 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.01fF
C7733 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C7734 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.12fF
C7735 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C7736 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C7737 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.02fF
C7738 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.04fF
C7739 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkinv_4_7/A 0.45fF
C7740 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.06fF
C7741 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C7742 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C7743 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# VDD 0.09fF
C7744 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C7745 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C7746 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.06fF
C7747 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.01fF
C7748 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C7749 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C7750 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C7751 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# 0.01fF
C7752 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.01fF
C7753 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.01fF
C7754 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__nand2_1_1/B 0.07fF
C7755 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.01fF
C7756 sky130_fd_sc_hd__clkinv_1_3/A clk 0.00fF
C7757 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.86fF
C7758 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.02fF
C7759 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.02fF
C7760 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.02fF
C7761 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C7762 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.00fF
C7763 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C7764 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C7765 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.02fF
C7766 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.00fF
C7767 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.01fF
C7768 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.02fF
C7769 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C7770 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C7771 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C7772 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C7773 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C7774 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C7775 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.03fF
C7776 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C7777 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.02fF
C7778 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C7779 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# 0.09fF
C7780 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_4_5/Y 0.85fF
C7781 sky130_fd_sc_hd__nand2_1_1/A Ad_b 0.55fF
C7782 sky130_fd_sc_hd__clkinv_1_2/Y sky130_fd_sc_hd__nand2_4_2/A 0.69fF
C7783 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C7784 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.02fF
C7785 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C7786 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.01fF
C7787 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.00fF
C7788 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.00fF
C7789 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C7790 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C7791 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C7792 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C7793 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.01fF
C7794 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.02fF
C7795 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# 0.00fF
C7796 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.95fF
C7797 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VDD 0.15fF
C7798 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C7799 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C7800 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C7801 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C7802 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.02fF
C7803 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C7804 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C7805 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C7806 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C7807 VDD sky130_fd_sc_hd__nand2_1_4/Y 0.45fF
C7808 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C7809 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.00fF
C7810 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.11fF
C7811 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.00fF
C7812 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C7813 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.00fF
C7814 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.02fF
C7815 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C7816 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C7817 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C7818 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C7819 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C7820 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.02fF
C7821 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C7822 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.03fF
C7823 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C7824 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C7825 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.55fF
C7826 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.04fF
C7827 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.00fF
C7828 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.00fF
C7829 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C7830 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C7831 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C7832 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C7833 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.02fF
C7834 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.00fF
C7835 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.02fF
C7836 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.00fF
C7837 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.01fF
C7838 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C7839 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.02fF
C7840 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C7841 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C7842 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C7843 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.02fF
C7844 sky130_fd_sc_hd__nand2_1_2/A clk 0.05fF
C7845 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.01fF
C7846 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C7847 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C7848 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# 0.00fF
C7849 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.01fF
C7850 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.00fF
C7851 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.02fF
C7852 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.04fF
C7853 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.04fF
C7854 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C7855 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C7856 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C7857 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C7858 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.00fF
C7859 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.03fF
C7860 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C7861 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.02fF
C7862 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.02fF
C7863 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.00fF
C7864 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C7865 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C7866 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C7867 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.00fF
C7868 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C7869 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.01fF
C7870 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C7871 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.00fF
C7872 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C7873 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.00fF
C7874 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.01fF
C7875 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.18fF
C7876 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.03fF
C7877 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.00fF
C7878 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.00fF
C7879 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y -0.34fF
C7880 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C7881 p2d p2_b 0.53fF
C7882 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C7883 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C7884 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.02fF
C7885 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_561_413# 0.01fF
C7886 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# 0.84fF
C7887 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.00fF
C7888 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C7889 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C7890 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C7891 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.02fF
C7892 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C7893 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C7894 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.03fF
C7895 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C7896 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C7897 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.00fF
C7898 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C7899 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C7900 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C7901 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C7902 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.03fF
C7903 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C7904 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C7905 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.03fF
C7906 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.01fF
C7907 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C7908 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.02fF
C7909 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.02fF
C7910 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C7911 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.65fF
C7912 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C7913 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C7914 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C7915 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.00fF
C7916 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.14fF
C7917 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__nand2_1_4/Y -0.01fF
C7918 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C7919 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C7920 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.03fF
C7921 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.01fF
C7922 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C7923 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.02fF
C7924 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.01fF
C7925 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.07fF
C7926 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.04fF
C7927 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.04fF
C7928 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.57fF
C7929 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C7930 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkinv_1_1/Y 0.02fF
C7931 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C7932 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.66fF
C7933 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C7934 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C7935 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C7936 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.01fF
C7937 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C7938 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C7939 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C7940 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.00fF
C7941 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# VDD 0.12fF
C7942 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.04fF
C7943 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.02fF
C7944 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.01fF
C7945 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__dfxbp_1_1/D 0.07fF
C7946 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A VDD 0.22fF
C7947 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C7948 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C7949 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C7950 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Bd_b 0.03fF
C7951 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.00fF
C7952 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# 0.00fF
C7953 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# 0.00fF
C7954 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.00fF
C7955 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__mux2_1_0/X 0.00fF
C7956 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C7957 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C7958 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C7959 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C7960 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C7961 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# 0.01fF
C7962 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.03fF
C7963 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C7964 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.00fF
C7965 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C7966 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C7967 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.02fF
C7968 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# Bd 0.02fF
C7969 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C7970 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C7971 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.06fF
C7972 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C7973 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.08fF
C7974 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_1/B 0.95fF
C7975 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C7976 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C7977 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C7978 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C7979 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C7980 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C7981 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C7982 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C7983 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.00fF
C7984 p2 sky130_fd_sc_hd__nand2_4_3/B 0.06fF
C7985 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C7986 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C7987 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.02fF
C7988 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.03fF
C7989 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A VDD 0.51fF
C7990 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C7991 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.12fF
C7992 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C7993 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.02fF
C7994 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C7995 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VDD 0.53fF
C7996 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.05fF
C7997 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C7998 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.04fF
C7999 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.03fF
C8000 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.10fF
C8001 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C8002 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.01fF
C8003 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.08fF
C8004 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C8005 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C8006 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C8007 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C8008 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.01fF
C8009 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C8010 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.16fF
C8011 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.14fF
C8012 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.04fF
C8013 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A -0.37fF
C8014 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VDD 0.60fF
C8015 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.11fF
C8016 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C8017 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C8018 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C8019 p2_b sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.12fF
C8020 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# p2 0.12fF
C8021 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C8022 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.04fF
C8023 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.06fF
C8024 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C8025 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.04fF
C8026 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# VDD 0.31fF
C8027 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.74fF
C8028 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C8029 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C8030 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C8031 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C8032 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C8033 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.00fF
C8034 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# VDD 0.39fF
C8035 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C8036 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.00fF
C8037 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.00fF
C8038 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.00fF
C8039 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.08fF
C8040 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C8041 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C8042 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.04fF
C8043 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.04fF
C8044 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VDD 0.54fF
C8045 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.02fF
C8046 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.02fF
C8047 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C8048 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C8049 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.06fF
C8050 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C8051 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.00fF
C8052 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.00fF
C8053 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.01fF
C8054 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.00fF
C8055 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.02fF
C8056 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C8057 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C8058 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C8059 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C8060 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C8061 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C8062 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C8063 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# VDD 0.13fF
C8064 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C8065 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C8066 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.01fF
C8067 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.03fF
C8068 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C8069 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C8070 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C8071 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C8072 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C8073 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.02fF
C8074 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C8075 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C8076 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.01fF
C8077 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C8078 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# VDD 0.15fF
C8079 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# VDD 0.14fF
C8080 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.02fF
C8081 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_2/A 0.26fF
C8082 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.00fF
C8083 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C8084 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C8085 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.02fF
C8086 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VDD 0.06fF
C8087 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C8088 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C8089 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.00fF
C8090 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.00fF
C8091 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.00fF
C8092 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# VDD 0.45fF
C8093 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C8094 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C8095 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.04fF
C8096 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.04fF
C8097 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.05fF
C8098 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.01fF
C8099 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.01fF
C8100 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C8101 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.02fF
C8102 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.14fF
C8103 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# VDD 0.14fF
C8104 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.04fF
C8105 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.04fF
C8106 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C8107 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C8108 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C8109 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.05fF
C8110 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C8111 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C8112 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C8113 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.03fF
C8114 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# VDD 0.18fF
C8115 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C8116 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C8117 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C8118 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C8119 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.02fF
C8120 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.01fF
C8121 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C8122 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C8123 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C8124 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C8125 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.00fF
C8126 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C8127 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C8128 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C8129 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.01fF
C8130 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C8131 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# VDD 0.30fF
C8132 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C8133 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C8134 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C8135 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.02fF
C8136 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.00fF
C8137 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C8138 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C8139 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.02fF
C8140 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.73fF
C8141 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# 0.01fF
C8142 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C8143 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.04fF
C8144 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.00fF
C8145 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C8146 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C8147 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C8148 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.02fF
C8149 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C8150 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Ad 0.05fF
C8151 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# VDD 0.33fF
C8152 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.01fF
C8153 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.04fF
C8154 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.04fF
C8155 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.01fF
C8156 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/X 0.00fF
C8157 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_592_47# -0.00fF
C8158 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.02fF
C8159 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C8160 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C8161 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.01fF
C8162 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.01fF
C8163 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.03fF
C8164 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.01fF
C8165 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C8166 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1d 0.12fF
C8167 p1d_b sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.12fF
C8168 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.11fF
C8169 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C8170 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.05fF
C8171 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C8172 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.00fF
C8173 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.08fF
C8174 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C8175 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C8176 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C8177 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C8178 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C8179 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.01fF
C8180 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C8181 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.02fF
C8182 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.02fF
C8183 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C8184 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C8185 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C8186 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C8187 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C8188 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X Ad_b 0.02fF
C8189 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.02fF
C8190 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.02fF
C8191 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.02fF
C8192 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VDD 0.54fF
C8193 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C8194 VDD A 1.54fF
C8195 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# 0.09fF
C8196 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C8197 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.07fF
C8198 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C8199 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C8200 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C8201 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C8202 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.03fF
C8203 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C8204 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C8205 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.11fF
C8206 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C8207 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C8208 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VDD 0.51fF
C8209 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C8210 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C8211 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C8212 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.02fF
C8213 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C8214 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C8215 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C8216 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.11fF
C8217 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X -0.00fF
C8218 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C8219 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.01fF
C8220 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.01fF
C8221 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.02fF
C8222 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C8223 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C8224 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C8225 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.05fF
C8226 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.01fF
C8227 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C8228 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.09fF
C8229 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.02fF
C8230 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.01fF
C8231 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# VDD 0.14fF
C8232 VDD sky130_fd_sc_hd__nand2_4_1/A 11.01fF
C8233 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C8234 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.03fF
C8235 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C8236 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C8237 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C8238 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C8239 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C8240 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# VDD 0.12fF
C8241 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C8242 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C8243 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C8244 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C8245 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C8246 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C8247 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C8248 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C8249 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C8250 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C8251 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C8252 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C8253 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_1_2/B 0.03fF
C8254 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C8255 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C8256 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.01fF
C8257 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.01fF
C8258 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.02fF
C8259 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C8260 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# VDD 0.30fF
C8261 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__nand2_1_1/B 0.03fF
C8262 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C8263 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C8264 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C8265 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.03fF
C8266 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C8267 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C8268 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.02fF
C8269 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C8270 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C8271 sky130_fd_sc_hd__nand2_4_3/B Ad_b 0.04fF
C8272 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C8273 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.04fF
C8274 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.03fF
C8275 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.01fF
C8276 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.00fF
C8277 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_4_9/Y 0.02fF
C8278 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clk 0.01fF
C8279 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C8280 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.01fF
C8281 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.01fF
C8282 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C8283 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C8284 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.01fF
C8285 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.01fF
C8286 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.02fF
C8287 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C8288 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C8289 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.02fF
C8290 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C8291 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C8292 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.01fF
C8293 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C8294 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# VDD 0.31fF
C8295 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# VDD 0.14fF
C8296 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# VDD 0.16fF
C8297 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.04fF
C8298 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.00fF
C8299 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C8300 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C8301 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C8302 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.01fF
C8303 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C8304 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C8305 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.00fF
C8306 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.05fF
C8307 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C8308 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.02fF
C8309 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.02fF
C8310 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# VDD 0.14fF
C8311 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.02fF
C8312 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.02fF
C8313 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# VDD 0.33fF
C8314 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.04fF
C8315 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.03fF
C8316 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C8317 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.02fF
C8318 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C8319 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C8320 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C8321 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.00fF
C8322 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C8323 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# 0.01fF
C8324 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C8325 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.00fF
C8326 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkinv_4_1/A 0.01fF
C8327 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C8328 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C8329 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C8330 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C8331 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C8332 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.14fF
C8333 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.07fF
C8334 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.03fF
C8335 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C8336 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C8337 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.00fF
C8338 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.02fF
C8339 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C8340 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.02fF
C8341 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.00fF
C8342 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C8343 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C8344 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C8345 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.01fF
C8346 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_7/A 0.72fF
C8347 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C8348 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.05fF
C8349 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C8350 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C8351 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.02fF
C8352 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C8353 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.00fF
C8354 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C8355 sky130_fd_sc_hd__nand2_1_4/B Bd_b 0.02fF
C8356 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.02fF
C8357 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C8358 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.02fF
C8359 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.01fF
C8360 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.01fF
C8361 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.00fF
C8362 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.03fF
C8363 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C8364 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C8365 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C8366 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C8367 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.02fF
C8368 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.01fF
C8369 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C8370 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_0/B 0.14fF
C8371 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VDD 0.35fF
C8372 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.01fF
C8373 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C8374 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.01fF
C8375 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C8376 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.04fF
C8377 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C8378 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C8379 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C8380 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.00fF
C8381 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.00fF
C8382 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.00fF
C8383 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.00fF
C8384 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.00fF
C8385 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.01fF
C8386 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C8387 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C8388 p1d_b p1_b 0.19fF
C8389 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_175/A 0.69fF
C8390 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C8391 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C8392 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.00fF
C8393 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C8394 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.01fF
C8395 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C8396 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C8397 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C8398 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# VDD 0.19fF
C8399 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.05fF
C8400 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.00fF
C8401 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C8402 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.02fF
C8403 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C8404 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C8405 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.01fF
C8406 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.02fF
C8407 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C8408 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkinv_4_5/Y 0.85fF
C8409 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VDD 0.30fF
C8410 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C8411 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.01fF
C8412 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.01fF
C8413 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# 0.03fF
C8414 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.01fF
C8415 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.30fF
C8416 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C8417 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.01fF
C8418 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# B_b 0.12fF
C8419 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C8420 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD 0.78fF
C8421 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.05fF
C8422 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C8423 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C8424 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C8425 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C8426 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.00fF
C8427 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C8428 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X Bd_b 0.02fF
C8429 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C8430 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C8431 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.05fF
C8432 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C8433 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.01fF
C8434 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C8435 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# VDD 0.13fF
C8436 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# VDD 0.17fF
C8437 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C8438 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C8439 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.00fF
C8440 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C8441 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C8442 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C8443 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C8444 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.01fF
C8445 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C8446 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.07fF
C8447 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# VDD 0.30fF
C8448 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.02fF
C8449 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C8450 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.00fF
C8451 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.00fF
C8452 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.00fF
C8453 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.00fF
C8454 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C8455 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.02fF
C8456 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C8457 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C8458 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.00fF
C8459 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.00fF
C8460 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C8461 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.00fF
C8462 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.00fF
C8463 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.08fF
C8464 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.14fF
C8465 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C8466 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.00fF
C8467 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# 0.08fF
C8468 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C8469 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C8470 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.18fF
C8471 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.06fF
C8472 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.11fF
C8473 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C8474 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# 0.02fF
C8475 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# 0.00fF
C8476 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# 0.01fF
C8477 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C8478 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.34fF
C8479 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C8480 p2 VDD 4.24fF
C8481 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# VDD 0.14fF
C8482 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C8483 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C8484 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.03fF
C8485 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.03fF
C8486 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C8487 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C8488 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkinv_1_2/Y 0.00fF
C8489 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.02fF
C8490 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.01fF
C8491 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.68fF
C8492 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C8493 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C8494 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C8495 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.05fF
C8496 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C8497 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.04fF
C8498 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C8499 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# -0.00fF
C8500 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C8501 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.01fF
C8502 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C8503 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C8504 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.01fF
C8505 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.03fF
C8506 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.00fF
C8507 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C8508 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C8509 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.03fF
C8510 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.02fF
C8511 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C8512 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C8513 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C8514 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VDD 0.60fF
C8515 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_1_3/A 0.04fF
C8516 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C8517 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.03fF
C8518 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.01fF
C8519 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.01fF
C8520 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.01fF
C8521 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.01fF
C8522 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkinv_4_7/A 0.04fF
C8523 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.76fF
C8524 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.08fF
C8525 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C8526 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.03fF
C8527 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.04fF
C8528 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.04fF
C8529 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# 0.07fF
C8530 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C8531 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C8532 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C8533 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.02fF
C8534 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# VDD 0.17fF
C8535 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.00fF
C8536 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.00fF
C8537 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.00fF
C8538 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.19fF
C8539 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.04fF
C8540 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.00fF
C8541 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C8542 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C8543 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C8544 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C8545 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.55fF
C8546 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C8547 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C8548 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.00fF
C8549 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C8550 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C8551 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.01fF
C8552 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A -0.00fF
C8553 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.29fF
C8554 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C8555 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C8556 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C8557 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C8558 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C8559 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C8560 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.03fF
C8561 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C8562 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C8563 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.01fF
C8564 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C8565 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.00fF
C8566 p1 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.06fF
C8567 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1d 0.06fF
C8568 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# 0.02fF
C8569 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# 0.02fF
C8570 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C8571 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C8572 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C8573 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C8574 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.02fF
C8575 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C8576 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.04fF
C8577 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0.04fF
C8578 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C8579 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# 0.00fF
C8580 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# 0.01fF
C8581 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# 0.02fF
C8582 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C8583 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.02fF
C8584 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C8585 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.06fF
C8586 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C8587 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# VDD 0.34fF
C8588 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# VDD 0.14fF
C8589 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# VDD 0.14fF
C8590 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# VDD 0.12fF
C8591 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.01fF
C8592 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C8593 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.01fF
C8594 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C8595 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C8596 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.01fF
C8597 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkinv_4_5/Y 0.03fF
C8598 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C8599 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C8600 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C8601 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C8602 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C8603 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.13fF
C8604 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# VDD 0.16fF
C8605 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C8606 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C8607 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C8608 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C8609 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C8610 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C8611 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.07fF
C8612 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# 0.01fF
C8613 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C8614 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.01fF
C8615 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C8616 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C8617 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C8618 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.19fF
C8619 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.04fF
C8620 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# VDD 0.30fF
C8621 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.00fF
C8622 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C8623 VDD sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.34fF
C8624 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.04fF
C8625 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.04fF
C8626 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C8627 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C8628 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C8629 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.03fF
C8630 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C8631 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C8632 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.32fF
C8633 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# 0.05fF
C8634 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C8635 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C8636 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.03fF
C8637 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C8638 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C8639 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C8640 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C8641 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.01fF
C8642 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C8643 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C8644 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.02fF
C8645 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.02fF
C8646 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C8647 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C8648 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C8649 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C8650 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C8651 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.02fF
C8652 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.02fF
C8653 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C8654 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# 0.01fF
C8655 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C8656 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C8657 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C8658 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.01fF
C8659 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C8660 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C8661 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Bd_b 0.02fF
C8662 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.02fF
C8663 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.02fF
C8664 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.02fF
C8665 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# VDD 0.17fF
C8666 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C8667 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.00fF
C8668 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C8669 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.08fF
C8670 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C8671 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.00fF
C8672 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# p2 0.06fF
C8673 p2d sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.06fF
C8674 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.44fF
C8675 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.01fF
C8676 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.03fF
C8677 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.01fF
C8678 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.04fF
C8679 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.02fF
C8680 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C8681 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.09fF
C8682 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.01fF
C8683 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.01fF
C8684 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.00fF
C8685 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C8686 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.02fF
C8687 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C8688 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.00fF
C8689 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.02fF
C8690 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.02fF
C8691 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.01fF
C8692 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.17fF
C8693 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.05fF
C8694 VDD Ad_b 5.95fF
C8695 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# Bd_b 0.46fF
C8696 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C8697 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C8698 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C8699 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C8700 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C8701 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.30fF
C8702 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.45fF
C8703 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/X 0.00fF
C8704 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C8705 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C8706 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C8707 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.02fF
C8708 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.01fF
C8709 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VDD 0.73fF
C8710 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C8711 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C8712 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.01fF
C8713 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.02fF
C8714 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.06fF
C8715 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# VDD 0.31fF
C8716 Bd B_b 0.53fF
C8717 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C8718 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.00fF
C8719 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.00fF
C8720 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C8721 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.09fF
C8722 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.01fF
C8723 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C8724 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.02fF
C8725 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C8726 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C8727 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/X 0.01fF
C8728 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.55fF
C8729 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C8730 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C8731 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C8732 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C8733 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.02fF
C8734 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.02fF
C8735 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C8736 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.10fF
C8737 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# Bd_b 0.01fF
C8738 sky130_fd_sc_hd__nand2_4_3/a_27_47# VDD 0.05fF
C8739 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C8740 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C8741 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C8742 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C8743 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# VDD 0.14fF
C8744 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# Ad_b 0.01fF
C8745 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# Bd_b 0.01fF
C8746 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.00fF
C8747 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.00fF
C8748 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.00fF
C8749 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C8750 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C8751 p1d_b p2d_b 0.11fF
C8752 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.01fF
C8753 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# A 0.12fF
C8754 A_b sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.12fF
C8755 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.01fF
C8756 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.05fF
C8757 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.01fF
C8758 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.01fF
C8759 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.01fF
C8760 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C8761 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.03fF
C8762 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.01fF
C8763 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/X 0.01fF
C8764 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.00fF
C8765 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C8766 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C8767 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.02fF
C8768 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C8769 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.01fF
C8770 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C8771 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.00fF
C8772 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.16fF
C8773 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.01fF
C8774 p1 p1_b 0.47fF
C8775 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.03fF
C8776 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 1.68fF
C8777 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.03fF
C8778 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C8779 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C8780 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C8781 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.06fF
C8782 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C8783 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.09fF
C8784 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.01fF
C8785 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C8786 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C8787 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# 0.05fF
C8788 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.02fF
C8789 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.02fF
C8790 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.02fF
C8791 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C8792 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/X 0.01fF
C8793 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C8794 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.08fF
C8795 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.03fF
C8796 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C8797 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.06fF
C8798 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.05fF
C8799 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C8800 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.07fF
C8801 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C8802 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.00fF
C8803 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.00fF
C8804 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.02fF
C8805 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.01fF
C8806 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.00fF
C8807 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.69fF
C8808 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C8809 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.01fF
C8810 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.01fF
C8811 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C8812 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C8813 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.02fF
C8814 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C8815 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.04fF
C8816 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C8817 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C8818 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C8819 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C8820 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.02fF
C8821 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.02fF
C8822 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C8823 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C8824 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C8825 sky130_fd_sc_hd__nand2_1_1/A Bd_b 1.60fF
C8826 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.02fF
C8827 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# 0.00fF
C8828 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C8829 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.02fF
C8830 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.84fF
C8831 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.01fF
C8832 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.01fF
C8833 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C8834 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C8835 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C8836 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.02fF
C8837 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C8838 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C8839 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.64fF
C8840 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/A 0.41fF
C8841 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C8842 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C8843 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C8844 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C8845 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.04fF
C8846 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.53fF
C8847 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C8848 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.04fF
C8849 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.05fF
C8850 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C8851 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.31fF
C8852 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C8853 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C8854 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.02fF
C8855 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.02fF
C8856 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.02fF
C8857 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C8858 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.54fF
C8859 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.01fF
C8860 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VDD 0.55fF
C8861 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C8862 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C8863 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.06fF
C8864 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.02fF
C8865 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C8866 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.02fF
C8867 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.01fF
C8868 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.01fF
C8869 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C8870 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C8871 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.11fF
C8872 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# 0.01fF
C8873 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C8874 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.01fF
C8875 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C8876 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.00fF
C8877 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C8878 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C8879 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.00fF
C8880 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.00fF
C8881 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C8882 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C8883 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__mux2_1_0/S 0.05fF
C8884 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.03fF
C8885 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C8886 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C8887 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.00fF
C8888 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.04fF
C8889 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.03fF
C8890 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C8891 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.01fF
C8892 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.01fF
C8893 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.01fF
C8894 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.01fF
C8895 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# 0.01fF
C8896 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.04fF
C8897 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.01fF
C8898 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.02fF
C8899 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.01fF
C8900 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C8901 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_3/A 0.16fF
C8902 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.00fF
C8903 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C8904 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C8905 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.01fF
C8906 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.06fF
C8907 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.01fF
C8908 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkinv_4_7/A 0.11fF
C8909 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C8910 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.03fF
C8911 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C8912 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.14fF
C8913 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C8914 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.00fF
C8915 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C8916 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.01fF
C8917 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.09fF
C8918 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# 0.05fF
C8919 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.02fF
C8920 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C8921 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.03fF
C8922 sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C8923 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/B 0.08fF
C8924 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C8925 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C8926 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C8927 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C8928 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.12fF
C8929 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# 0.15fF
C8930 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.02fF
C8931 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.10fF
C8932 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C8933 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# 0.00fF
C8934 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C8935 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.02fF
C8936 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C8937 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C8938 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C8939 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.01fF
C8940 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C8941 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C8942 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.33fF
C8943 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.04fF
C8944 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.04fF
C8945 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C8946 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.05fF
C8947 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.04fF
C8948 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.05fF
C8949 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C8950 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.32fF
C8951 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# VDD 0.33fF
C8952 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.01fF
C8953 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.00fF
C8954 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C8955 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.08fF
C8956 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.03fF
C8957 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.00fF
C8958 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C8959 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# 0.02fF
C8960 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.00fF
C8961 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C8962 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Ad_b 0.03fF
C8963 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C8964 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C8965 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.00fF
C8966 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C8967 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C8968 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C8969 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.08fF
C8970 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C8971 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_0/A 0.21fF
C8972 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C8973 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.00fF
C8974 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.00fF
C8975 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.04fF
C8976 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C8977 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.01fF
C8978 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# 0.00fF
C8979 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.02fF
C8980 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C8981 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.01fF
C8982 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.01fF
C8983 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C8984 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C8985 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.11fF
C8986 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C8987 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C8988 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.01fF
C8989 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.02fF
C8990 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.01fF
C8991 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.57fF
C8992 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.01fF
C8993 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C8994 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.03fF
C8995 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# 0.00fF
C8996 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.09fF
C8997 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C8998 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C8999 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C9000 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C9001 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C9002 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# VDD 0.06fF
C9003 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/A 0.03fF
C9004 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.00fF
C9005 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.02fF
C9006 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.01fF
C9007 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.02fF
C9008 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.02fF
C9009 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.03fF
C9010 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C9011 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.01fF
C9012 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.09fF
C9013 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.02fF
C9014 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.00fF
C9015 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# 0.00fF
C9016 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# 0.02fF
C9017 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.00fF
C9018 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.53fF
C9019 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C9020 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.82fF
C9021 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C9022 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.66fF
C9023 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.08fF
C9024 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C9025 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C9026 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C9027 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.31fF
C9028 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.01fF
C9029 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C9030 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C9031 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.01fF
C9032 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.03fF
C9033 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# 0.01fF
C9034 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C9035 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C9036 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.02fF
C9037 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C9038 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.01fF
C9039 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C9040 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VDD 0.74fF
C9041 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C9042 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C9043 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C9044 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.00fF
C9045 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C9046 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C9047 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C9048 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C9049 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C9050 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.00fF
C9051 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.02fF
C9052 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# 0.01fF
C9053 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_4/Y 0.04fF
C9054 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C9055 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C9056 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.02fF
C9057 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.03fF
C9058 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C9059 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C9060 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C9061 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.01fF
C9062 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.02fF
C9063 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.15fF
C9064 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C9065 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# Ad_b 0.00fF
C9066 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.03fF
C9067 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C9068 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C9069 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.00fF
C9070 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C9071 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.01fF
C9072 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VDD 0.77fF
C9073 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C9074 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C9075 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.02fF
C9076 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.01fF
C9077 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.00fF
C9078 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C9079 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A VDD 0.57fF
C9080 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C9081 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C9082 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.02fF
C9083 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.03fF
C9084 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.15fF
C9085 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.02fF
C9086 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.06fF
C9087 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C9088 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.03fF
C9089 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C9090 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C9091 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C9092 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# VDD 0.18fF
C9093 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C9094 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.09fF
C9095 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C9096 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C9097 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# VDD 0.22fF
C9098 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.23fF
C9099 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C9100 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.00fF
C9101 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.01fF
C9102 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.00fF
C9103 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.00fF
C9104 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C9105 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.34fF
C9106 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# VDD 0.31fF
C9107 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.05fF
C9108 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.00fF
C9109 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.29fF
C9110 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.01fF
C9111 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.03fF
C9112 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C9113 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.02fF
C9114 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C9115 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/X 0.03fF
C9116 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C9117 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.00fF
C9118 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.01fF
C9119 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.01fF
C9120 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C9121 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C9122 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C9123 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C9124 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.04fF
C9125 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C9126 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.01fF
C9127 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.04fF
C9128 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C9129 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C9130 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.01fF
C9131 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.01fF
C9132 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.03fF
C9133 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.03fF
C9134 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C9135 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# VDD 0.12fF
C9136 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.06fF
C9137 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.01fF
C9138 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C9139 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C9140 sky130_fd_sc_hd__dfxbp_1_0/a_561_413# VDD 0.00fF
C9141 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C9142 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C9143 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.00fF
C9144 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.00fF
C9145 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.00fF
C9146 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# VDD 0.19fF
C9147 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkinv_4_5/Y 0.04fF
C9148 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C9149 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C9150 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C9151 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C9152 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C9153 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C9154 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.06fF
C9155 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.01fF
C9156 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C9157 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C9158 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C9159 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C9160 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C9161 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.01fF
C9162 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.02fF
C9163 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C9164 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.07fF
C9165 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C9166 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C9167 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.02fF
C9168 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C9169 p2 sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C9170 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# VDD 0.14fF
C9171 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.04fF
C9172 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C9173 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C9174 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.00fF
C9175 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C9176 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C9177 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C9178 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C9179 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.01fF
C9180 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.02fF
C9181 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C9182 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.01fF
C9183 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C9184 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C9185 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# VDD 0.11fF
C9186 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C9187 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C9188 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C9189 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C9190 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C9191 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.02fF
C9192 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.02fF
C9193 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C9194 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C9195 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C9196 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.04fF
C9197 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.03fF
C9198 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.01fF
C9199 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.30fF
C9200 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.00fF
C9201 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.00fF
C9202 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.03fF
C9203 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# VDD 0.15fF
C9204 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_3/Y 0.03fF
C9205 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C9206 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C9207 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C9208 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__dfxbp_1_0/a_975_413# 0.01fF
C9209 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.01fF
C9210 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C9211 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C9212 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C9213 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C9214 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C9215 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# VDD 0.30fF
C9216 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_1_2/B 0.05fF
C9217 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C9218 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C9219 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C9220 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.02fF
C9221 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.02fF
C9222 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VDD 0.52fF
C9223 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C9224 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.00fF
C9225 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# 0.02fF
C9226 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# 0.02fF
C9227 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.05fF
C9228 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.02fF
C9229 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C9230 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A sky130_fd_sc_hd__clkinv_1_1/Y 0.02fF
C9231 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.03fF
C9232 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.05fF
C9233 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C9234 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.05fF
C9235 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X Bd_b 0.02fF
C9236 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C9237 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C9238 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A VDD 0.58fF
C9239 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C9240 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.03fF
C9241 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C9242 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C9243 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.01fF
C9244 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.01fF
C9245 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.04fF
C9246 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.00fF
C9247 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VDD 0.73fF
C9248 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.05fF
C9249 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C9250 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.11fF
C9251 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C9252 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C9253 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C9254 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C9255 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C9256 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.00fF
C9257 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C9258 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C9259 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkinv_4_1/A 0.45fF
C9260 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VDD 0.57fF
C9261 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.02fF
C9262 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.02fF
C9263 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C9264 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C9265 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C9266 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.03fF
C9267 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C9268 VDD sky130_fd_sc_hd__nand2_4_2/A 5.81fF
C9269 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C9270 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/A 0.46fF
C9271 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.01fF
C9272 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C9273 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C9274 VDD sky130_fd_sc_hd__nand2_1_0/B 1.07fF
C9275 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.01fF
C9276 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C9277 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C9278 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C9279 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C9280 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C9281 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C9282 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C9283 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C9284 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# VDD 0.11fF
C9285 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C9286 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.01fF
C9287 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C9288 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C9289 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C9290 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# 0.00fF
C9291 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.03fF
C9292 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C9293 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.04fF
C9294 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.04fF
C9295 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C9296 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.01fF
C9297 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.02fF
C9298 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.00fF
C9299 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.02fF
C9300 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.01fF
C9301 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C9302 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.00fF
C9303 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C9304 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C9305 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# VDD 0.16fF
C9306 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C9307 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C9308 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.02fF
C9309 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C9310 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C9311 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C9312 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C9313 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C9314 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.02fF
C9315 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C9316 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.06fF
C9317 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C9318 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Ad_b 0.02fF
C9319 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C9320 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.02fF
C9321 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# VDD 0.34fF
C9322 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.02fF
C9323 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.02fF
C9324 sky130_fd_sc_hd__nand2_4_3/B Bd_b 0.03fF
C9325 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.02fF
C9326 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C9327 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.01fF
C9328 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C9329 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# VDD 0.14fF
C9330 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C9331 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C9332 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C9333 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C9334 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C9335 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.00fF
C9336 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.02fF
C9337 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# VDD 0.15fF
C9338 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C9339 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C9340 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.02fF
C9341 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# VDD 0.12fF
C9342 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C9343 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C9344 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# VDD 0.17fF
C9345 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C9346 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.02fF
C9347 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C9348 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C9349 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.01fF
C9350 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# Ad_b 0.16fF
C9351 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.01fF
C9352 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C9353 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# 0.00fF
C9354 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# 0.00fF
C9355 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C9356 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C9357 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# VDD 0.22fF
C9358 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.00fF
C9359 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# VDD 0.33fF
C9360 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.04fF
C9361 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.04fF
C9362 sky130_fd_sc_hd__mux2_1_0/a_76_199# Ad_b 0.02fF
C9363 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/S 0.11fF
C9364 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VDD 0.33fF
C9365 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.06fF
C9366 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C9367 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.02fF
C9368 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.01fF
C9369 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# 0.09fF
C9370 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C9371 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C9372 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.05fF
C9373 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C9374 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C9375 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.11fF
C9376 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.03fF
C9377 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.02fF
C9378 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C9379 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C9380 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C9381 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.00fF
C9382 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C9383 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C9384 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C9385 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C9386 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C9387 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C9388 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.01fF
C9389 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.01fF
C9390 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.01fF
C9391 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C9392 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C9393 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.09fF
C9394 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C9395 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.00fF
C9396 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.02fF
C9397 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C9398 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.02fF
C9399 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.02fF
C9400 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C9401 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C9402 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C9403 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.05fF
C9404 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C9405 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.00fF
C9406 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.00fF
C9407 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VDD 0.19fF
C9408 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_3/Y 0.05fF
C9409 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.34fF
C9410 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C9411 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.01fF
C9412 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.00fF
C9413 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.00fF
C9414 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C9415 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C9416 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.02fF
C9417 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VDD 0.61fF
C9418 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.09fF
C9419 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C9420 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.00fF
C9421 sky130_fd_sc_hd__mux2_1_0/S Ad_b 0.17fF
C9422 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C9423 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C9424 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C9425 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__clkinv_4_5/Y 0.00fF
C9426 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.01fF
C9427 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.38fF
C9428 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C9429 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.02fF
C9430 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C9431 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C9432 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.82fF
C9433 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# VDD 0.15fF
C9434 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C9435 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.01fF
C9436 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C9437 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C9438 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.56fF
C9439 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C9440 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C9441 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.08fF
C9442 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.02fF
C9443 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C9444 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.00fF
C9445 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.03fF
C9446 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VDD 0.18fF
C9447 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C9448 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C9449 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.02fF
C9450 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.05fF
C9451 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.04fF
C9452 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.04fF
C9453 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C9454 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.01fF
C9455 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C9456 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.01fF
C9457 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.00fF
C9458 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.03fF
C9459 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.01fF
C9460 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C9461 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C9462 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.00fF
C9463 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.00fF
C9464 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C9465 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.02fF
C9466 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.01fF
C9467 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.02fF
C9468 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C9469 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.00fF
C9470 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__nand2_4_0/Y 0.09fF
C9471 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C9472 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# VDD 0.14fF
C9473 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C9474 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A sky130_fd_sc_hd__nand2_1_1/A 0.02fF
C9475 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C9476 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C9477 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C9478 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C9479 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.01fF
C9480 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C9481 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.06fF
C9482 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.08fF
C9483 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.23fF
C9484 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C9485 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# VDD 0.16fF
C9486 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.03fF
C9487 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.01fF
C9488 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.15fF
C9489 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.01fF
C9490 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C9491 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C9492 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.01fF
C9493 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# VDD 0.29fF
C9494 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.00fF
C9495 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.00fF
C9496 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.00fF
C9497 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.00fF
C9498 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C9499 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# 0.05fF
C9500 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.04fF
C9501 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C9502 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.15fF
C9503 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.02fF
C9504 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C9505 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.02fF
C9506 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.07fF
C9507 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.03fF
C9508 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.03fF
C9509 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C9510 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C9511 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C9512 VDD sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.25fF
C9513 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.15fF
C9514 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C9515 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# 0.01fF
C9516 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# 0.01fF
C9517 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.11fF
C9518 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.08fF
C9519 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.56fF
C9520 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C9521 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.04fF
C9522 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_110/A 0.09fF
C9523 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C9524 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C9525 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.08fF
C9526 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.70fF
C9527 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.11fF
C9528 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C9529 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.03fF
C9530 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# 0.30fF
C9531 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.07fF
C9532 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.01fF
C9533 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.02fF
C9534 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C9535 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C9536 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.01fF
C9537 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.02fF
C9538 sky130_fd_sc_hd__nand2_4_0/Y Bd_b 0.00fF
C9539 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C9540 Ad_b sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C9541 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.00fF
C9542 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.00fF
C9543 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C9544 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C9545 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C9546 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.01fF
C9547 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/A 0.03fF
C9548 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C9549 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C9550 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C9551 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.11fF
C9552 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.04fF
C9553 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C9554 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.01fF
C9555 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VDD 0.55fF
C9556 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.02fF
C9557 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C9558 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# VDD 0.30fF
C9559 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.02fF
C9560 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.00fF
C9561 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C9562 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.03fF
C9563 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.01fF
C9564 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VDD 0.57fF
C9565 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C9566 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C9567 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.14fF
C9568 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# 0.00fF
C9569 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C9570 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# -0.08fF
C9571 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C9572 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C9573 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C9574 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C9575 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C9576 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# p1_b 0.10fF
C9577 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.08fF
C9578 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# VDD 0.45fF
C9579 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.56fF
C9580 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C9581 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C9582 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C9583 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.03fF
C9584 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C9585 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.15fF
C9586 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C9587 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C9588 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.02fF
C9589 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.00fF
C9590 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C9591 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# VDD 0.14fF
C9592 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.02fF
C9593 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.00fF
C9594 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.02fF
C9595 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.02fF
C9596 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C9597 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# 0.10fF
C9598 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C9599 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C9600 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C9601 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C9602 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.00fF
C9603 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.00fF
C9604 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.00fF
C9605 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.01fF
C9606 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.15fF
C9607 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C9608 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C9609 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C9610 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.00fF
C9611 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C9612 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.02fF
C9613 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.03fF
C9614 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.29fF
C9615 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C9616 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__mux2_1_0/X 0.07fF
C9617 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.01fF
C9618 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C9619 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.01fF
C9620 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C9621 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C9622 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C9623 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.02fF
C9624 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.04fF
C9625 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.04fF
C9626 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.01fF
C9627 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/B 0.16fF
C9628 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C9629 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.01fF
C9630 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.01fF
C9631 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0.01fF
C9632 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.00fF
C9633 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.01fF
C9634 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C9635 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.04fF
C9636 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# 0.01fF
C9637 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# 0.01fF
C9638 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.01fF
C9639 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C9640 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.00fF
C9641 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C9642 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.02fF
C9643 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# VDD 0.34fF
C9644 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C9645 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C9646 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# VDD 0.17fF
C9647 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.70fF
C9648 p2 A 0.02fF
C9649 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C9650 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C9651 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.01fF
C9652 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.01fF
C9653 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.00fF
C9654 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# 0.00fF
C9655 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.04fF
C9656 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.04fF
C9657 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# VDD 0.30fF
C9658 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VDD 0.50fF
C9659 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.02fF
C9660 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.84fF
C9661 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# VDD 0.15fF
C9662 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C9663 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C9664 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C9665 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# 0.02fF
C9666 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# 0.02fF
C9667 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C9668 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C9669 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C9670 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# 0.00fF
C9671 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C9672 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C9673 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.04fF
C9674 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.15fF
C9675 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# VDD 0.15fF
C9676 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C9677 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.02fF
C9678 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.01fF
C9679 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.01fF
C9680 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.02fF
C9681 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C9682 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C9683 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C9684 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.05fF
C9685 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.05fF
C9686 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.01fF
C9687 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.34fF
C9688 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C9689 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C9690 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C9691 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.06fF
C9692 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.14fF
C9693 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C9694 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C9695 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C9696 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.02fF
C9697 p2 sky130_fd_sc_hd__nand2_4_1/A 0.17fF
C9698 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C9699 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.02fF
C9700 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.29fF
C9701 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C9702 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C9703 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.04fF
C9704 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C9705 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C9706 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C9707 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C9708 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C9709 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.00fF
C9710 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.02fF
C9711 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0.09fF
C9712 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C9713 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.01fF
C9714 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.02fF
C9715 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C9716 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.05fF
C9717 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.02fF
C9718 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# 0.00fF
C9719 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.03fF
C9720 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.00fF
C9721 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# VDD 0.15fF
C9722 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C9723 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# -0.07fF
C9724 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C9725 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.01fF
C9726 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.00fF
C9727 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.00fF
C9728 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.00fF
C9729 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# 0.00fF
C9730 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.00fF
C9731 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/A 0.01fF
C9732 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C9733 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.00fF
C9734 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.00fF
C9735 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C9736 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.10fF
C9737 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C9738 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.03fF
C9739 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Ad_b 0.04fF
C9740 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C9741 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.04fF
C9742 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.04fF
C9743 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.01fF
C9744 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C9745 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C9746 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C9747 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VDD 0.33fF
C9748 VDD Bd_b 8.00fF
C9749 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C9750 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.14fF
C9751 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.02fF
C9752 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C9753 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C9754 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C9755 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C9756 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.02fF
C9757 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C9758 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C9759 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.01fF
C9760 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.16fF
C9761 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C9762 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C9763 B_b sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.06fF
C9764 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C9765 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.02fF
C9766 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.02fF
C9767 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C9768 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.23fF
C9769 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.00fF
C9770 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.02fF
C9771 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.01fF
C9772 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# VDD 0.19fF
C9773 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VDD 0.52fF
C9774 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# VDD 0.29fF
C9775 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X Ad_b 0.02fF
C9776 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.00fF
C9777 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.00fF
C9778 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C9779 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C9780 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C9781 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.00fF
C9782 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.04fF
C9783 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C9784 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.00fF
C9785 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.00fF
C9786 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C9787 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C9788 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C9789 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A -0.00fF
C9790 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.00fF
C9791 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C9792 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C9793 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C9794 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C9795 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__nand2_4_3/A 0.05fF
C9796 sky130_fd_sc_hd__nand2_4_3/A clk 0.03fF
C9797 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C9798 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C9799 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C9800 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.00fF
C9801 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.00fF
C9802 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.07fF
C9803 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# Bd_b 0.01fF
C9804 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.11fF
C9805 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C9806 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C9807 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.01fF
C9808 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.02fF
C9809 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.04fF
C9810 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.00fF
C9811 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C9812 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X sky130_fd_sc_hd__clkinv_4_9/Y 0.03fF
C9813 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.02fF
C9814 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.02fF
C9815 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C9816 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.07fF
C9817 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.00fF
C9818 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C9819 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.01fF
C9820 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C9821 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.00fF
C9822 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.02fF
C9823 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C9824 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.01fF
C9825 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.02fF
C9826 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C9827 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.03fF
C9828 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C9829 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C9830 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# 0.03fF
C9831 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C9832 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# 0.09fF
C9833 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C9834 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.02fF
C9835 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.01fF
C9836 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C9837 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.01fF
C9838 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C9839 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C9840 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/A 0.01fF
C9841 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.02fF
C9842 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C9843 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C9844 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.04fF
C9845 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.04fF
C9846 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C9847 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C9848 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C9849 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.02fF
C9850 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C9851 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VDD 0.35fF
C9852 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.03fF
C9853 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_4_5/Y 0.14fF
C9854 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C9855 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C9856 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C9857 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# 0.00fF
C9858 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.00fF
C9859 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.00fF
C9860 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.00fF
C9861 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C9862 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.02fF
C9863 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# 0.01fF
C9864 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.02fF
C9865 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# 0.04fF
C9866 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_70/X 0.01fF
C9867 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkinv_4_1/A 0.08fF
C9868 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.03fF
C9869 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C9870 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.00fF
C9871 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C9872 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.01fF
C9873 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.04fF
C9874 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.04fF
C9875 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C9876 VDD sky130_fd_sc_hd__nand2_1_0/A 1.27fF
C9877 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.01fF
C9878 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C9879 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C9880 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C9881 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C9882 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_1_3/Y 0.04fF
C9883 A Ad_b 0.26fF
C9884 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.01fF
C9885 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C9886 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C9887 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C9888 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.01fF
C9889 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.02fF
C9890 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.01fF
C9891 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.03fF
C9892 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C9893 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C9894 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# 0.01fF
C9895 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C9896 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.63fF
C9897 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C9898 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C9899 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.02fF
C9900 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C9901 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__clkinv_4_7/A 0.01fF
C9902 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C9903 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.02fF
C9904 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.01fF
C9905 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C9906 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C9907 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C9908 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C9909 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C9910 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C9911 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.01fF
C9912 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.02fF
C9913 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.02fF
C9914 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C9915 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_12/X 0.02fF
C9916 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_119/X 0.56fF
C9917 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.55fF
C9918 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C9919 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.05fF
C9920 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.03fF
C9921 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.09fF
C9922 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0.01fF
C9923 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C9924 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C9925 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C9926 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.02fF
C9927 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C9928 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C9929 sky130_fd_sc_hd__nand2_4_1/A Ad_b 0.48fF
C9930 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.01fF
C9931 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C9932 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C9933 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.03fF
C9934 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.01fF
C9935 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.02fF
C9936 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.02fF
C9937 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C9938 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_98/X 0.01fF
C9939 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C9940 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C9941 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.01fF
C9942 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.01fF
C9943 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.01fF
C9944 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C9945 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.00fF
C9946 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.00fF
C9947 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.02fF
C9948 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_51/X 0.01fF
C9949 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.01fF
C9950 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C9951 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.03fF
C9952 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.00fF
C9953 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_592_47# 0.00fF
C9954 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.07fF
C9955 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.12fF
C9956 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.02fF
C9957 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C9958 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C9959 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.01fF
C9960 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C9961 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C9962 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C9963 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C9964 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.17fF
C9965 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.02fF
C9966 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C9967 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C9968 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C9969 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.04fF
C9970 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# 0.02fF
C9971 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C9972 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.02fF
C9973 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.28fF
C9974 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# VDD 0.15fF
C9975 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/X 0.02fF
C9976 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.14fF
C9977 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# 0.01fF
C9978 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.01fF
C9979 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C9980 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C9981 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Bd_b 0.02fF
C9982 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C9983 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.01fF
C9984 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C9985 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.04fF
C9986 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.04fF
C9987 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C9988 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# VDD 0.30fF
C9989 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.30fF
C9990 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.43fF
C9991 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.00fF
C9992 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.00fF
C9993 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.00fF
C9994 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.00fF
C9995 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_1_3/A 0.03fF
C9996 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.00fF
C9997 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.00fF
C9998 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C9999 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.02fF
C10000 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.01fF
C10001 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# 0.01fF
C10002 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C10003 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C10004 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C10005 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C10006 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.06fF
C10007 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.05fF
C10008 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.04fF
C10009 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/Y 0.02fF
C10010 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C10011 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C10012 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C10013 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C10014 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C10015 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.02fF
C10016 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.00fF
C10017 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C10018 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.02fF
C10019 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.04fF
C10020 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.02fF
C10021 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C10022 sky130_fd_sc_hd__dfxbp_1_1/a_561_413# VDD 0.01fF
C10023 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VDD -0.70fF
C10024 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.00fF
C10025 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C10026 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.01fF
C10027 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.01fF
C10028 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.00fF
C10029 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C10030 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# 0.00fF
C10031 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# 0.00fF
C10032 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.00fF
C10033 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.00fF
C10034 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.03fF
C10035 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# VDD 0.37fF
C10036 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.03fF
C10037 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.04fF
C10038 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.02fF
C10039 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C10040 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C10041 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.03fF
C10042 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C10043 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C10044 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C10045 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VDD 0.59fF
C10046 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C10047 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.84fF
C10048 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.02fF
C10049 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# 0.01fF
C10050 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.01fF
C10051 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.01fF
C10052 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.01fF
C10053 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C10054 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# 0.01fF
C10055 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C10056 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C10057 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.01fF
C10058 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_9/X 0.84fF
C10059 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C10060 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.04fF
C10061 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# 0.01fF
C10062 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.01fF
C10063 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C10064 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.02fF
C10065 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.03fF
C10066 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.01fF
C10067 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# Bd_b 0.00fF
C10068 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.02fF
C10069 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.01fF
C10070 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C10071 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.01fF
C10072 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C10073 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C10074 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C10075 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C10076 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.04fF
C10077 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.01fF
C10078 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.03fF
C10079 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# 0.02fF
C10080 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.00fF
C10081 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C10082 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.01fF
C10083 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.02fF
C10084 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.01fF
C10085 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C10086 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C10087 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C10088 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C10089 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C10090 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C10091 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C10092 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.01fF
C10093 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C10094 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.01fF
C10095 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.03fF
C10096 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# sky130_fd_sc_hd__clkinv_4_7/A 0.06fF
C10097 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.08fF
C10098 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/Y 0.05fF
C10099 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C10100 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C10101 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.11fF
C10102 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# 0.01fF
C10103 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C10104 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C10105 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.04fF
C10106 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.04fF
C10107 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# VDD 0.13fF
C10108 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.14fF
C10109 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.01fF
C10110 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# VDD 0.14fF
C10111 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.02fF
C10112 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C10113 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.01fF
C10114 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.00fF
C10115 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.00fF
C10116 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.17fF
C10117 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# VDD 0.18fF
C10118 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.15fF
C10119 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.01fF
C10120 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/A 0.01fF
C10121 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C10122 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.04fF
C10123 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.04fF
C10124 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.02fF
C10125 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.02fF
C10126 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkinv_1_2/Y 0.00fF
C10127 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C10128 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.01fF
C10129 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.01fF
C10130 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.09fF
C10131 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__nand2_4_0/A 0.05fF
C10132 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.02fF
C10133 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# VDD 0.29fF
C10134 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.03fF
C10135 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# -0.33fF
C10136 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C10137 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.31fF
C10138 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# 0.09fF
C10139 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.01fF
C10140 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.00fF
C10141 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C10142 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C10143 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C10144 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C10145 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.00fF
C10146 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.06fF
C10147 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.03fF
C10148 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VDD 0.59fF
C10149 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C10150 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.12fF
C10151 sky130_fd_sc_hd__dfxbp_1_0/a_975_413# VDD 0.00fF
C10152 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C10153 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C10154 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C10155 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.01fF
C10156 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C10157 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.00fF
C10158 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.00fF
C10159 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# VDD 0.14fF
C10160 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C10161 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C10162 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C10163 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.02fF
C10164 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C10165 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__nand2_1_1/A 0.02fF
C10166 p2_b sky130_fd_sc_hd__clkinv_4_10/Y 0.03fF
C10167 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.01fF
C10168 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C10169 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C10170 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.00fF
C10171 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.02fF
C10172 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.02fF
C10173 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.04fF
C10174 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C10175 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.06fF
C10176 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C10177 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.00fF
C10178 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.04fF
C10179 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.04fF
C10180 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C10181 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C10182 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C10183 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C10184 p2 Ad_b 1.13fF
C10185 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.02fF
C10186 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.01fF
C10187 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.04fF
C10188 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.04fF
C10189 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/A 0.01fF
C10190 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/A 0.00fF
C10191 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C10192 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C10193 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.02fF
C10194 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.01fF
C10195 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.01fF
C10196 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/A 0.00fF
C10197 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C10198 B Bd_b 0.08fF
C10199 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C10200 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# VDD 0.14fF
C10201 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# 0.01fF
C10202 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.01fF
C10203 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# VDD 0.29fF
C10204 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/A 0.01fF
C10205 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C10206 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.00fF
C10207 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# 0.11fF
C10208 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C10209 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C10210 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C10211 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.02fF
C10212 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.02fF
C10213 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C10214 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.01fF
C10215 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.15fF
C10216 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C10217 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/X 0.03fF
C10218 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.01fF
C10219 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.00fF
C10220 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C10221 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.07fF
C10222 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# VDD 0.15fF
C10223 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A VDD 0.57fF
C10224 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.04fF
C10225 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.04fF
C10226 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C10227 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C10228 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C10229 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C10230 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C10231 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.08fF
C10232 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C10233 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.03fF
C10234 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.29fF
C10235 sky130_fd_sc_hd__dfxbp_1_0/Q_N VDD 0.20fF
C10236 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# VDD 0.19fF
C10237 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# 0.09fF
C10238 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C10239 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C10240 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.00fF
C10241 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C10242 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.02fF
C10243 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# VDD 0.40fF
C10244 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C10245 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C10246 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VDD 0.41fF
C10247 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.04fF
C10248 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.04fF
C10249 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.01fF
C10250 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.00fF
C10251 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/Y 0.73fF
C10252 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# 0.05fF
C10253 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.02fF
C10254 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.01fF
C10255 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/X 0.01fF
C10256 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C10257 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.68fF
C10258 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C10259 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C10260 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.00fF
C10261 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C10262 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C10263 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C10264 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.00fF
C10265 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.00fF
C10266 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C10267 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C10268 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C10269 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C10270 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.01fF
C10271 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.04fF
C10272 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.02fF
C10273 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C10274 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C10275 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.19fF
C10276 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_1_1/A 0.02fF
C10277 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C10278 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C10279 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C10280 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.03fF
C10281 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C10282 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.01fF
C10283 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C10284 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C10285 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C10286 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C10287 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# p1d 0.05fF
C10288 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.11fF
C10289 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C10290 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C10291 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.00fF
C10292 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C10293 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.04fF
C10294 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.03fF
C10295 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C10296 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374# 0.01fF
C10297 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C10298 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.01fF
C10299 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/A 0.01fF
C10300 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C10301 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C10302 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.00fF
C10303 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.00fF
C10304 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.00fF
C10305 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.00fF
C10306 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C10307 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_7/A 0.68fF
C10308 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/X 0.01fF
C10309 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C10310 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.09fF
C10311 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C10312 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C10313 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C10314 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.01fF
C10315 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.01fF
C10316 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.01fF
C10317 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.01fF
C10318 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C10319 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C10320 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.00fF
C10321 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# 0.02fF
C10322 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.01fF
C10323 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# VDD 0.15fF
C10324 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.03fF
C10325 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.01fF
C10326 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.06fF
C10327 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C10328 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C10329 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C10330 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Bd_b 0.02fF
C10331 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C10332 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C10333 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C10334 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C10335 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C10336 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# VDD 0.20fF
C10337 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.00fF
C10338 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C10339 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C10340 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# VDD 0.14fF
C10341 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VDD 0.47fF
C10342 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C10343 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C10344 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C10345 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C10346 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.09fF
C10347 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.12fF
C10348 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.03fF
C10349 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.01fF
C10350 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A -0.00fF
C10351 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.01fF
C10352 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C10353 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C10354 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C10355 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# VDD 0.14fF
C10356 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C10357 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.01fF
C10358 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C10359 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C10360 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.01fF
C10361 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# Bd_b 0.10fF
C10362 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# 0.00fF
C10363 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# 0.00fF
C10364 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.03fF
C10365 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.05fF
C10366 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# 0.02fF
C10367 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.00fF
C10368 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C10369 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# VDD 0.09fF
C10370 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C10371 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C10372 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C10373 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# VDD 0.17fF
C10374 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VDD 0.18fF
C10375 sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C10376 sky130_fd_sc_hd__mux2_1_0/a_76_199# Bd_b 0.02fF
C10377 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C10378 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C10379 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C10380 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.04fF
C10381 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.04fF
C10382 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A VDD 0.58fF
C10383 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.11fF
C10384 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/X 0.06fF
C10385 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# VDD 0.28fF
C10386 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# VDD 0.28fF
C10387 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X sky130_fd_sc_hd__clkinv_4_2/Y 0.04fF
C10388 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.04fF
C10389 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.05fF
C10390 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.05fF
C10391 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.01fF
C10392 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_4_5/Y 0.37fF
C10393 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C10394 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.02fF
C10395 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C10396 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.00fF
C10397 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C10398 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.02fF
C10399 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.08fF
C10400 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C10401 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C10402 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.02fF
C10403 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C10404 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C10405 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C10406 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.09fF
C10407 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.04fF
C10408 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.02fF
C10409 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__nand2_1_0/A 0.02fF
C10410 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.01fF
C10411 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.00fF
C10412 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.00fF
C10413 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__nand2_4_0/Y 0.09fF
C10414 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C10415 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C10416 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_110/X 0.03fF
C10417 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C10418 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.00fF
C10419 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.00fF
C10420 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.00fF
C10421 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C10422 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.44fF
C10423 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VDD 0.56fF
C10424 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VDD 0.14fF
C10425 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.02fF
C10426 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C10427 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C10428 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.00fF
C10429 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C10430 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2d_b 0.12fF
C10431 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.04fF
C10432 sky130_fd_sc_hd__mux2_1_0/S Bd_b 0.12fF
C10433 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C10434 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C10435 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C10436 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.00fF
C10437 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.00fF
C10438 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.00fF
C10439 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# 0.00fF
C10440 Bd_b sky130_fd_sc_hd__clkinv_4_2/Y 0.10fF
C10441 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C10442 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.02fF
C10443 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C10444 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.00fF
C10445 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C10446 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C10447 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.02fF
C10448 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C10449 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C10450 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C10451 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C10452 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C10453 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.01fF
C10454 sky130_fd_sc_hd__clkinv_4_7/Y VDD 0.55fF
C10455 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C10456 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C10457 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.00fF
C10458 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.00fF
C10459 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.01fF
C10460 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# 0.01fF
C10461 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VDD 0.14fF
C10462 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_166/A 0.06fF
C10463 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C10464 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C10465 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C10466 sky130_fd_sc_hd__clkinv_4_1/A VDD 4.36fF
C10467 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C10468 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.01fF
C10469 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_160/A 0.01fF
C10470 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# 0.01fF
C10471 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C10472 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C10473 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C10474 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.02fF
C10475 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# 0.01fF
C10476 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C10477 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C10478 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C10479 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.03fF
C10480 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_124/X 0.01fF
C10481 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C10482 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.01fF
C10483 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.05fF
C10484 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.00fF
C10485 p2d sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C10486 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# 0.01fF
C10487 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C10488 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C10489 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.00fF
C10490 p1_b p1d 0.52fF
C10491 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.11fF
C10492 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.06fF
C10493 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C10494 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C10495 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.06fF
C10496 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VDD 0.53fF
C10497 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.00fF
C10498 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C10499 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C10500 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.03fF
C10501 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/X 0.00fF
C10502 B sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.06fF
C10503 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# Bd 0.06fF
C10504 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.05fF
C10505 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.04fF
C10506 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.05fF
C10507 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# VDD 0.15fF
C10508 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C10509 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.00fF
C10510 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.00fF
C10511 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.01fF
C10512 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C10513 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VDD 0.53fF
C10514 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C10515 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.01fF
C10516 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# 0.03fF
C10517 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.01fF
C10518 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.00fF
C10519 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.00fF
C10520 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.00fF
C10521 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# 0.00fF
C10522 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# VDD 0.15fF
C10523 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.00fF
C10524 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.01fF
C10525 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_155/X 0.01fF
C10526 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.03fF
C10527 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C10528 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.08fF
C10529 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VDD 0.53fF
C10530 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.15fF
C10531 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__nand2_4_0/A 2.21fF
C10532 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C10533 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C10534 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.82fF
C10535 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.04fF
C10536 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# 0.01fF
C10537 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C10538 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.03fF
C10539 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# 0.14fF
C10540 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.01fF
C10541 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.08fF
C10542 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.07fF
C10543 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.04fF
C10544 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VDD 0.59fF
C10545 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# 0.18fF
C10546 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.00fF
C10547 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C10548 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.01fF
C10549 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.01fF
C10550 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_111/X 0.03fF
C10551 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C10552 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.02fF
C10553 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.01fF
C10554 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C10555 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.09fF
C10556 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.00fF
C10557 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.08fF
C10558 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.02fF
C10559 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.01fF
C10560 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C10561 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/X 0.00fF
C10562 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.11fF
C10563 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.04fF
C10564 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# 0.04fF
C10565 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.29fF
C10566 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.01fF
C10567 sky130_fd_sc_hd__nand2_1_1/B clk 0.00fF
C10568 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.06fF
C10569 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C10570 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.03fF
C10571 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.03fF
C10572 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.59fF
C10573 Bd_b sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C10574 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# 0.01fF
C10575 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# VDD 0.43fF
C10576 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# 0.00fF
C10577 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# 0.00fF
C10578 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# 0.00fF
C10579 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# 0.00fF
C10580 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.11fF
C10581 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X sky130_fd_sc_hd__clkinv_4_7/A 0.84fF
C10582 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C10583 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C10584 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C10585 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C10586 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C10587 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.02fF
C10588 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Ad_b 0.02fF
C10589 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.09fF
C10590 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# VDD 0.33fF
C10591 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.11fF
C10592 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.05fF
C10593 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.01fF
C10594 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# 0.04fF
C10595 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# 0.04fF
C10596 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.01fF
C10597 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# VDD 0.18fF
C10598 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C10599 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.02fF
C10600 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.00fF
C10601 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C10602 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C10603 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C10604 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C10605 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.03fF
C10606 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# VDD 0.43fF
C10607 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VDD 0.62fF
C10608 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VDD 0.60fF
C10609 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.10fF
C10610 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C10611 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.05fF
C10612 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C10613 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C10614 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# 0.05fF
C10615 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# VDD 0.18fF
C10616 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C10617 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C10618 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C10619 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.01fF
C10620 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A VDD 0.56fF
C10621 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C10622 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C10623 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.02fF
C10624 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C10625 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C10626 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C10627 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.03fF
C10628 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C10629 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.03fF
C10630 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# 0.04fF
C10631 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# VDD 0.27fF
C10632 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C10633 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C10634 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# 0.01fF
C10635 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# 0.00fF
C10636 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# 0.00fF
C10637 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.01fF
C10638 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/A 0.01fF
C10639 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.12fF
C10640 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.01fF
C10641 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C10642 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C10643 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C10644 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C10645 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.16fF
C10646 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.03fF
C10647 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.03fF
C10648 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.01fF
C10649 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/X 0.01fF
C10650 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C10651 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C10652 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.02fF
C10653 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C10654 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C10655 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.02fF
C10656 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C10657 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C10658 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C10659 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C10660 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.02fF
C10661 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.32fF
C10662 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C10663 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.01fF
C10664 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.09fF
C10665 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.02fF
C10666 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.02fF
C10667 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# 0.01fF
C10668 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.02fF
C10669 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.01fF
C10670 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.15fF
C10671 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C10672 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C10673 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# 0.01fF
C10674 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C10675 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.02fF
C10676 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/A 0.01fF
C10677 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.01fF
C10678 VDD Ad 1.64fF
C10679 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# VDD 0.17fF
C10680 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.01fF
C10681 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# VDD 0.14fF
C10682 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.00fF
C10683 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# 0.00fF
C10684 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# 0.00fF
C10685 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# 0.00fF
C10686 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C10687 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C10688 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C10689 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C10690 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C10691 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/Y 0.73fF
C10692 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C10693 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# VDD 0.28fF
C10694 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/B 0.07fF
C10695 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.01fF
C10696 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.01fF
C10697 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.02fF
C10698 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# VDD 0.16fF
C10699 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# VDD 0.29fF
C10700 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_1_0/A 0.06fF
C10701 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.00fF
C10702 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C10703 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C10704 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.01fF
C10705 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C10706 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# VDD 0.22fF
C10707 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.57fF
C10708 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# 0.00fF
C10709 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C10710 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/A 0.04fF
C10711 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.02fF
C10712 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.06fF
C10713 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.02fF
C10714 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# VDD 0.14fF
C10715 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C10716 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.02fF
C10717 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.02fF
C10718 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C10719 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C10720 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.06fF
C10721 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.08fF
C10722 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# 0.02fF
C10723 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.01fF
C10724 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# 0.01fF
C10725 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C10726 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.06fF
C10727 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A VDD 0.56fF
C10728 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C10729 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C10730 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.01fF
C10731 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C10732 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.14fF
C10733 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C10734 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C10735 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.17fF
C10736 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C10737 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C10738 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C10739 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C10740 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C10741 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VDD 0.34fF
C10742 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C10743 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.01fF
C10744 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C10745 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_3/A 2.16fF
C10746 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.15fF
C10747 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.29fF
C10748 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# 0.11fF
C10749 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.06fF
C10750 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A sky130_fd_sc_hd__clkdlybuf4s50_1_120/A 0.04fF
C10751 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.00fF
C10752 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.01fF
C10753 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.02fF
C10754 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C10755 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C10756 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C10757 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.07fF
C10758 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A sky130_fd_sc_hd__clkinv_1_3/Y 0.02fF
C10759 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/X 0.01fF
C10760 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.00fF
C10761 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# 0.04fF
C10762 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# 0.04fF
C10763 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C10764 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.10fF
C10765 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C10766 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.09fF
C10767 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C10768 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.03fF
C10769 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.00fF
C10770 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# 0.01fF
C10771 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.02fF
C10772 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.02fF
C10773 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# 0.00fF
C10774 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# 0.00fF
C10775 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# 0.00fF
C10776 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.07fF
C10777 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Bd_b 0.05fF
C10778 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.01fF
C10779 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# 0.05fF
C10780 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C10781 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C10782 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# 0.02fF
C10783 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# 0.01fF
C10784 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# 0.01fF
C10785 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.03fF
C10786 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C10787 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C10788 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.02fF
C10789 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VDD 0.17fF
C10790 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X sky130_fd_sc_hd__nand2_4_1/A 0.05fF
C10791 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.00fF
C10792 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C10793 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C10794 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.15fF
C10795 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.02fF
C10796 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C10797 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C10798 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C10799 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C10800 VDD sky130_fd_sc_hd__clkinv_1_3/Y 0.29fF
C10801 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.01fF
C10802 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C10803 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C10804 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C10805 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.00fF
C10806 B_b VDD 0.77fF
C10807 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C10808 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.00fF
C10809 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# 0.01fF
C10810 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# 0.02fF
C10811 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.07fF
C10812 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C10813 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.11fF
C10814 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C10815 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# VDD 0.15fF
C10816 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C10817 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# 0.02fF
C10818 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# 0.01fF
C10819 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X Bd_b 0.03fF
C10820 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# VDD 0.15fF
C10821 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.05fF
C10822 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.05fF
C10823 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C10824 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# 0.05fF
C10825 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# VDD 0.35fF
C10826 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.02fF
C10827 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# 0.00fF
C10828 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.00fF
C10829 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# 0.01fF
C10830 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C10831 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0.01fF
C10832 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.11fF
C10833 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C10834 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C10835 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C10836 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/A 0.03fF
C10837 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.00fF
C10838 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C10839 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.00fF
C10840 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.01fF
C10841 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.03fF
C10842 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C10843 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_130/X 0.03fF
C10844 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C10845 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C10846 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.09fF
C10847 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C10848 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.01fF
C10849 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C10850 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C10851 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C10852 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_35/X 0.01fF
C10853 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C10854 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.01fF
C10855 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# 0.00fF
C10856 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.02fF
C10857 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# 0.00fF
C10858 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# 0.00fF
C10859 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.03fF
C10860 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C10861 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.01fF
C10862 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C10863 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.02fF
C10864 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.01fF
C10865 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C10866 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C10867 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C10868 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C10869 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# 0.00fF
C10870 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# 0.01fF
C10871 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# 0.02fF
C10872 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.06fF
C10873 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/A 0.00fF
C10874 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C10875 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.03fF
C10876 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.03fF
C10877 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.03fF
C10878 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.01fF
C10879 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.02fF
C10880 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# 0.03fF
C10881 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C10882 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.05fF
C10883 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.05fF
C10884 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.05fF
C10885 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.02fF
C10886 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.00fF
C10887 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# 0.00fF
C10888 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# 0.00fF
C10889 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C10890 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# 0.01fF
C10891 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# 0.01fF
C10892 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# 0.01fF
C10893 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.00fF
C10894 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.01fF
C10895 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C10896 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C10897 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C10898 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.00fF
C10899 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.02fF
C10900 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C10901 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_139/A 0.06fF
C10902 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/X 0.03fF
C10903 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C10904 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C10905 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VDD 0.19fF
C10906 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.04fF
C10907 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C10908 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.01fF
C10909 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C10910 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C10911 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C10912 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.00fF
C10913 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# 0.00fF
C10914 VDD sky130_fd_sc_hd__clkinv_4_9/Y 1.49fF
C10915 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.01fF
C10916 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.01fF
C10917 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.04fF
C10918 sky130_fd_sc_hd__clkinv_4_1/A B 0.00fF
C10919 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C10920 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.01fF
C10921 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/S 0.05fF
C10922 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.04fF
C10923 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.04fF
C10924 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C10925 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C10926 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C10927 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C10928 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.00fF
C10929 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C10930 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkinv_4_7/A 0.00fF
C10931 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.04fF
C10932 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.04fF
C10933 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C10934 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# 0.05fF
C10935 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_4_3/A 0.69fF
C10936 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C10937 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.00fF
C10938 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# 0.00fF
C10939 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C10940 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# 0.00fF
C10941 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# 0.00fF
C10942 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.09fF
C10943 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.02fF
C10944 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.01fF
C10945 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C10946 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.01fF
C10947 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.00fF
C10948 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.00fF
C10949 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C10950 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C10951 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# 0.02fF
C10952 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.00fF
C10953 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.01fF
C10954 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C10955 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C10956 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C10957 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.01fF
C10958 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C10959 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# 0.01fF
C10960 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# 0.02fF
C10961 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# 0.00fF
C10962 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.59fF
C10963 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.04fF
C10964 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.04fF
C10965 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C10966 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C10967 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C10968 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.00fF
C10969 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# 0.01fF
C10970 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# 0.02fF
C10971 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.06fF
C10972 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# 0.04fF
C10973 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.04fF
C10974 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.08fF
C10975 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C10976 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.00fF
C10977 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C10978 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.02fF
C10979 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C10980 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.11fF
C10981 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# 0.04fF
C10982 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# 0.04fF
C10983 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C10984 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C10985 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.00fF
C10986 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# 0.01fF
C10987 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/A 0.51fF
C10988 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VDD 0.34fF
C10989 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.04fF
C10990 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.04fF
C10991 sky130_fd_sc_hd__nand2_4_1/A Bd_b 0.66fF
C10992 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.01fF
C10993 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.02fF
C10994 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# 0.00fF
C10995 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# 0.00fF
C10996 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# 0.00fF
C10997 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.03fF
C10998 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.00fF
C10999 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/X 0.00fF
C11000 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.09fF
C11001 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A 1.25fF
C11002 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# 0.12fF
C11003 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.06fF
C11004 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C11005 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C11006 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.01fF
C11007 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# 0.02fF
C11008 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_19/A 0.03fF
C11009 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.05fF
C11010 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.02fF
C11011 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C11012 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.04fF
C11013 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.04fF
C11014 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.08fF
C11015 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C11016 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/a_975_413# 0.00fF
C11017 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.06fF
C11018 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.07fF
C11019 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.03fF
C11020 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# VDD 0.44fF
C11021 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C11022 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# 0.14fF
C11023 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.09fF
C11024 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# 0.02fF
C11025 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# 0.02fF
C11026 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# 0.01fF
C11027 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.12fF
C11028 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C11029 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C11030 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.04fF
C11031 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.14fF
C11032 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C11033 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# VDD 0.14fF
C11034 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C11035 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.03fF
C11036 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C11037 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.01fF
C11038 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# 0.01fF
C11039 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.04fF
C11040 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.04fF
C11041 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_10/Y 0.32fF
C11042 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C11043 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C11044 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C11045 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.44fF
C11046 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.03fF
C11047 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C11048 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C11049 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C11050 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C11051 sky130_fd_sc_hd__nand2_1_4/B clk 0.07fF
C11052 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.17fF
C11053 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# 0.14fF
C11054 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.02fF
C11055 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# VDD 0.18fF
C11056 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# 0.01fF
C11057 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# 0.00fF
C11058 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.00fF
C11059 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# 0.01fF
C11060 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.02fF
C11061 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.03fF
C11062 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# 0.02fF
C11063 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.04fF
C11064 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.04fF
C11065 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.11fF
C11066 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.06fF
C11067 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.32fF
C11068 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# VDD 0.31fF
C11069 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C11070 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C11071 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# 0.01fF
C11072 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C11073 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.03fF
C11074 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_74/X 0.03fF
C11075 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.00fF
C11076 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.02fF
C11077 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C11078 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C11079 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.01fF
C11080 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.02fF
C11081 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.05fF
C11082 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_28/A 0.01fF
C11083 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C11084 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.03fF
C11085 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.01fF
C11086 sky130_fd_sc_hd__dfxbp_1_1/a_975_413# VDD 0.01fF
C11087 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# 0.03fF
C11088 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_60/A 0.01fF
C11089 p1d_b sky130_fd_sc_hd__clkinv_4_8/Y 0.03fF
C11090 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.01fF
C11091 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.01fF
C11092 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C11093 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C11094 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# 0.00fF
C11095 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.02fF
C11096 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.05fF
C11097 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_26/A 0.00fF
C11098 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# 0.00fF
C11099 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# 0.00fF
C11100 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.09fF
C11101 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.01fF
C11102 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A VDD 0.58fF
C11103 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.06fF
C11104 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C11105 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/X 0.03fF
C11106 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.02fF
C11107 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# 0.03fF
C11108 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C11109 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.00fF
C11110 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.00fF
C11111 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# 0.01fF
C11112 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.08fF
C11113 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C11114 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_148/X 0.00fF
C11115 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C11116 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_9/A 0.01fF
C11117 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.02fF
C11118 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.04fF
C11119 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.01fF
C11120 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# 0.01fF
C11121 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# 0.02fF
C11122 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# 0.00fF
C11123 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/Y 0.16fF
C11124 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.02fF
C11125 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# 0.01fF
C11126 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C11127 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.02fF
C11128 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C11129 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C11130 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C11131 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# 0.01fF
C11132 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.01fF
C11133 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C11134 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.02fF
C11135 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Ad_b 0.02fF
C11136 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_151/X 0.03fF
C11137 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.06fF
C11138 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_64/A 0.02fF
C11139 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.04fF
C11140 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C11141 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C11142 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C11143 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.00fF
C11144 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.02fF
C11145 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# 0.00fF
C11146 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.01fF
C11147 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# 0.02fF
C11148 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C11149 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.02fF
C11150 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# 0.00fF
C11151 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# 0.02fF
C11152 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# 0.01fF
C11153 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C11154 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/Y 0.05fF
C11155 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/A 0.00fF
C11156 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.00fF
C11157 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.02fF
C11158 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C11159 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# 0.04fF
C11160 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# 0.04fF
C11161 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C11162 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.00fF
C11163 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C11164 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C11165 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.03fF
C11166 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkinv_4_8/Y 0.03fF
C11167 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.01fF
C11168 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# 0.01fF
C11169 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# 0.01fF
C11170 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# 0.01fF
C11171 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# 0.00fF
C11172 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# 0.02fF
C11173 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C11174 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_2/Y 0.68fF
C11175 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C11176 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C11177 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X sky130_fd_sc_hd__clkdlybuf4s50_1_128/X 0.04fF
C11178 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_45/X 0.03fF
C11179 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C11180 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_170/X 0.00fF
C11181 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# 0.00fF
C11182 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# 0.02fF
C11183 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# 0.01fF
C11184 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# 0.01fF
C11185 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C11186 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C11187 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_76/X 0.03fF
C11188 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/A 0.08fF
C11189 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# 0.05fF
C11190 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C11191 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# 0.01fF
C11192 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# 0.01fF
C11193 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# 0.01fF
C11194 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# 0.01fF
C11195 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.11fF
C11196 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C11197 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# 0.02fF
C11198 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# 0.01fF
C11199 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.02fF
C11200 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C11201 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VDD 0.28fF
C11202 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C11203 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A sky130_fd_sc_hd__clkdlybuf4s50_1_43/X 0.02fF
C11204 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C11205 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.14fF
C11206 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.56fF
C11207 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/X 0.01fF
C11208 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C11209 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# VDD 0.14fF
C11210 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.12fF
C11211 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# 0.03fF
C11212 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C11213 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# 0.01fF
C11214 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# 0.02fF
C11215 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# 0.01fF
C11216 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.00fF
C11217 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C11218 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_40/X 0.04fF
C11219 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/A 0.49fF
C11220 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C11221 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C11222 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C11223 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C11224 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# VDD 0.11fF
C11225 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VDD 0.36fF
C11226 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# 0.09fF
C11227 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_46/A 0.01fF
C11228 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_175/X 0.01fF
C11229 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.00fF
C11230 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# 0.07fF
C11231 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X sky130_fd_sc_hd__clkdlybuf4s50_1_62/A 0.00fF
C11232 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/Y 0.02fF
C11233 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_41/A 0.01fF
C11234 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# 0.00fF
C11235 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C11236 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C11237 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.06fF
C11238 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C11239 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_14/X 0.00fF
C11240 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.00fF
C11241 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# VDD 0.30fF
C11242 VDD sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.11fF
C11243 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C11244 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_185/A 0.03fF
C11245 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.07fF
C11246 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C11247 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C11248 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C11249 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_592_47# 0.01fF
C11250 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.02fF
C11251 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_57/X 0.00fF
C11252 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C11253 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C11254 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.01fF
C11255 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C11256 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# 0.00fF
C11257 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C11258 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# 0.01fF
C11259 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.00fF
C11260 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# 0.00fF
C11261 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C11262 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C11263 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C11264 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# 0.00fF
C11265 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# 0.00fF
C11266 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C11267 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.01fF
C11268 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C11269 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.04fF
C11270 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C11271 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# 0.01fF
C11272 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_30/A 0.06fF
C11273 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# 0.01fF
C11274 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# 0.01fF
C11275 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C11276 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C11277 sky130_fd_sc_hd__nand2_4_2/Y p1d 0.00fF
C11278 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C11279 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# 0.00fF
C11280 sky130_fd_sc_hd__nand2_4_2/A VSS 17.09fF
C11281 sky130_fd_sc_hd__clkinv_4_7/A VSS 79.29fF
C11282 sky130_fd_sc_hd__clkinv_4_9/Y VSS 75.42fF
C11283 sky130_fd_sc_hd__clkinv_4_5/Y VSS 117.98fF
C11284 sky130_fd_sc_hd__clkinv_4_2/Y VSS 38.91fF
C11285 clk VSS 17.23fF
C11286 p1d VSS 14.97fF
C11287 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# VSS 1.46fF
C11288 sky130_fd_sc_hd__nand2_1_0/B VSS 20.35fF
C11289 sky130_fd_sc_hd__nand2_1_4/Y VSS 34.19fF
C11290 Bd_b VSS 36.75fF
C11291 Ad_b VSS 11.70fF
C11292 sky130_fd_sc_hd__mux2_1_0/S VSS 10.43fF
C11293 sky130_fd_sc_hd__mux2_1_0/a_439_47# VSS 0.01fF
C11294 sky130_fd_sc_hd__mux2_1_0/a_218_47# VSS 0.01fF
C11295 sky130_fd_sc_hd__mux2_1_0/a_505_21# VSS 0.30fF
C11296 sky130_fd_sc_hd__mux2_1_0/a_76_199# VSS 0.28fF
C11297 sky130_fd_sc_hd__clkinv_1_3/Y VSS 32.97fF
C11298 sky130_fd_sc_hd__mux2_1_0/X VSS 43.22fF
C11299 sky130_fd_sc_hd__nand2_1_4/a_113_47# VSS 0.01fF
C11300 sky130_fd_sc_hd__clkinv_1_2/Y VSS 25.04fF
C11301 sky130_fd_sc_hd__nand2_4_3/A VSS 25.82fF
C11302 sky130_fd_sc_hd__nand2_1_3/A VSS 19.61fF
C11303 sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS -0.00fF
C11304 sky130_fd_sc_hd__clkdlybuf4s50_1_111/X VSS 8.53fF
C11305 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# VSS 0.20fF
C11306 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# VSS 0.27fF
C11307 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# VSS 0.36fF
C11308 sky130_fd_sc_hd__clkinv_1_1/Y VSS 32.89fF
C11309 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS 12.26fF
C11310 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_390_47# VSS 0.19fF
C11311 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_283_47# VSS 0.26fF
C11312 sky130_fd_sc_hd__clkdlybuf4s50_1_19/a_27_47# VSS 0.40fF
C11313 sky130_fd_sc_hd__nand2_1_2/A VSS 10.59fF
C11314 sky130_fd_sc_hd__nand2_1_2/B VSS 11.61fF
C11315 sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_390_47# VSS 0.21fF
C11316 sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_283_47# VSS 0.28fF
C11317 sky130_fd_sc_hd__clkdlybuf4s50_1_119/a_27_47# VSS 0.42fF
C11318 sky130_fd_sc_hd__clkdlybuf4s50_1_110/X VSS 6.20fF
C11319 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# VSS 0.19fF
C11320 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# VSS 0.27fF
C11321 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# VSS 0.37fF
C11322 sky130_fd_sc_hd__clkdlybuf4s50_1_30/A VSS 24.18fF
C11323 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# VSS 0.19fF
C11324 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# VSS 0.26fF
C11325 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# VSS 0.41fF
C11326 sky130_fd_sc_hd__clkdlybuf4s50_1_19/A VSS 35.56fF
C11327 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# VSS 0.19fF
C11328 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# VSS 0.26fF
C11329 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# VSS 0.40fF
C11330 sky130_fd_sc_hd__clkinv_1_0/Y VSS 32.90fF
C11331 p1_b VSS 15.64fF
C11332 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# VSS 1.58fF
C11333 sky130_fd_sc_hd__nand2_4_1/A VSS 25.68fF
C11334 sky130_fd_sc_hd__nand2_1_1/B VSS 13.67fF
C11335 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.01fF
C11336 sky130_fd_sc_hd__clkdlybuf4s50_1_130/X VSS 20.16fF
C11337 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# VSS 0.21fF
C11338 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# VSS 0.27fF
C11339 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# VSS 0.37fF
C11340 sky130_fd_sc_hd__clkdlybuf4s50_1_120/A VSS 22.45fF
C11341 sky130_fd_sc_hd__clkdlybuf4s50_1_119/X VSS 20.78fF
C11342 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# VSS 0.21fF
C11343 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# VSS 0.28fF
C11344 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# VSS 0.42fF
C11345 sky130_fd_sc_hd__clkdlybuf4s50_1_107/A VSS 10.35fF
C11346 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# VSS 0.19fF
C11347 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# VSS 0.27fF
C11348 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# VSS 0.35fF
C11349 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS 28.21fF
C11350 sky130_fd_sc_hd__clkdlybuf4s50_1_40/X VSS 47.97fF
C11351 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# VSS 0.22fF
C11352 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# VSS 0.30fF
C11353 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# VSS 0.40fF
C11354 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS 19.06fF
C11355 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_390_47# VSS 0.20fF
C11356 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_283_47# VSS 0.26fF
C11357 sky130_fd_sc_hd__clkdlybuf4s50_1_28/a_27_47# VSS 0.41fF
C11358 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS 14.40fF
C11359 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# VSS 0.21fF
C11360 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# VSS 0.27fF
C11361 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# VSS 0.35fF
C11362 p1 VSS 7.25fF
C11363 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# VSS 1.41fF
C11364 sky130_fd_sc_hd__nand2_4_0/A VSS 22.52fF
C11365 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS -0.00fF
C11366 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS 24.55fF
C11367 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_390_47# VSS 0.19fF
C11368 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_283_47# VSS 0.27fF
C11369 sky130_fd_sc_hd__clkdlybuf4s50_1_139/a_27_47# VSS 0.40fF
C11370 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS 20.48fF
C11371 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_390_47# VSS 0.20fF
C11372 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_283_47# VSS 0.28fF
C11373 sky130_fd_sc_hd__clkdlybuf4s50_1_128/a_27_47# VSS 0.38fF
C11374 sky130_fd_sc_hd__clkdlybuf4s50_1_119/A VSS 14.76fF
C11375 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# VSS 0.21fF
C11376 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# VSS 0.28fF
C11377 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# VSS 0.41fF
C11378 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS 6.50fF
C11379 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_390_47# VSS 0.19fF
C11380 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_283_47# VSS 0.27fF
C11381 sky130_fd_sc_hd__clkdlybuf4s50_1_106/a_27_47# VSS 0.37fF
C11382 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS 23.36fF
C11383 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# VSS 0.21fF
C11384 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# VSS 0.27fF
C11385 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# VSS 0.35fF
C11386 sky130_fd_sc_hd__clkdlybuf4s50_1_28/A VSS 14.77fF
C11387 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# VSS 0.20fF
C11388 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# VSS 0.26fF
C11389 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# VSS 0.40fF
C11390 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# VSS 0.23fF
C11391 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# VSS 0.35fF
C11392 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# VSS 0.81fF
C11393 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS 20.17fF
C11394 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_390_47# VSS 0.20fF
C11395 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_283_47# VSS 0.28fF
C11396 sky130_fd_sc_hd__clkdlybuf4s50_1_16/a_27_47# VSS 0.36fF
C11397 A VSS 28.24fF
C11398 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# VSS 1.45fF
C11399 sky130_fd_sc_hd__clkdlybuf4s50_1_151/X VSS 7.60fF
C11400 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# VSS 0.21fF
C11401 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# VSS 0.30fF
C11402 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# VSS 0.39fF
C11403 sky130_fd_sc_hd__clkdlybuf4s50_1_139/A VSS 24.18fF
C11404 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# VSS 0.21fF
C11405 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# VSS 0.28fF
C11406 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# VSS 0.42fF
C11407 sky130_fd_sc_hd__clkdlybuf4s50_1_128/X VSS 14.52fF
C11408 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# VSS 0.20fF
C11409 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# VSS 0.28fF
C11410 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# VSS 0.38fF
C11411 sky130_fd_sc_hd__clkdlybuf4s50_1_116/X VSS 20.88fF
C11412 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# VSS 0.20fF
C11413 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# VSS 0.28fF
C11414 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# VSS 0.40fF
C11415 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS 10.08fF
C11416 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_390_47# VSS 0.19fF
C11417 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_283_47# VSS 0.27fF
C11418 sky130_fd_sc_hd__clkdlybuf4s50_1_105/a_27_47# VSS 0.42fF
C11419 sky130_fd_sc_hd__clkdlybuf4s50_1_60/A VSS 20.32fF
C11420 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# VSS 0.21fF
C11421 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# VSS 0.28fF
C11422 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# VSS 0.41fF
C11423 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS 40.22fF
C11424 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_390_47# VSS 0.20fF
C11425 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_283_47# VSS 0.28fF
C11426 sky130_fd_sc_hd__clkdlybuf4s50_1_37/a_27_47# VSS 0.36fF
C11427 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS 15.15fF
C11428 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_390_47# VSS 0.19fF
C11429 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_283_47# VSS 0.26fF
C11430 sky130_fd_sc_hd__clkdlybuf4s50_1_26/a_27_47# VSS 0.40fF
C11431 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS 23.92fF
C11432 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# VSS 0.21fF
C11433 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# VSS 0.29fF
C11434 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# VSS 0.39fF
C11435 sky130_fd_sc_hd__clkdlybuf4s50_1_16/X VSS 20.10fF
C11436 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# VSS 0.22fF
C11437 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# VSS 0.30fF
C11438 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# VSS 0.39fF
C11439 A_b VSS 15.73fF
C11440 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# VSS 1.58fF
C11441 sky130_fd_sc_hd__clkdlybuf4s50_1_160/A VSS 41.64fF
C11442 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS 23.71fF
C11443 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# VSS 0.20fF
C11444 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# VSS 0.27fF
C11445 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# VSS 0.40fF
C11446 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS 25.00fF
C11447 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_390_47# VSS 0.20fF
C11448 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_283_47# VSS 0.27fF
C11449 sky130_fd_sc_hd__clkdlybuf4s50_1_148/a_27_47# VSS 0.38fF
C11450 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS 19.05fF
C11451 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_390_47# VSS 0.21fF
C11452 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_283_47# VSS 0.28fF
C11453 sky130_fd_sc_hd__clkdlybuf4s50_1_137/a_27_47# VSS 0.41fF
C11454 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS 14.79fF
C11455 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_390_47# VSS 0.20fF
C11456 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_283_47# VSS 0.28fF
C11457 sky130_fd_sc_hd__clkdlybuf4s50_1_126/a_27_47# VSS 0.38fF
C11458 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS 8.14fF
C11459 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_390_47# VSS 0.20fF
C11460 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_283_47# VSS 0.28fF
C11461 sky130_fd_sc_hd__clkdlybuf4s50_1_115/a_27_47# VSS 0.41fF
C11462 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS 11.05fF
C11463 sky130_fd_sc_hd__clkdlybuf4s50_1_105/X VSS 4.33fF
C11464 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# VSS 0.20fF
C11465 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# VSS 0.29fF
C11466 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# VSS 0.37fF
C11467 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS 14.27fF
C11468 sky130_fd_sc_hd__clkdlybuf4s50_1_70/X VSS 23.97fF
C11469 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# VSS 0.20fF
C11470 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# VSS 0.27fF
C11471 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# VSS 0.38fF
C11472 sky130_fd_sc_hd__clkdlybuf4s50_1_37/X VSS 40.31fF
C11473 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# VSS 0.22fF
C11474 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# VSS 0.30fF
C11475 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# VSS 0.39fF
C11476 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# VSS 0.20fF
C11477 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# VSS 0.26fF
C11478 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# VSS 0.35fF
C11479 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS 20.33fF
C11480 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS 14.28fF
C11481 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# VSS 0.20fF
C11482 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# VSS 0.27fF
C11483 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# VSS 0.40fF
C11484 sky130_fd_sc_hd__clkdlybuf4s50_1_26/A VSS 13.93fF
C11485 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# VSS 0.19fF
C11486 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# VSS 0.26fF
C11487 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# VSS 0.39fF
C11488 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS 20.43fF
C11489 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_390_47# VSS 0.22fF
C11490 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_283_47# VSS 0.30fF
C11491 sky130_fd_sc_hd__clkdlybuf4s50_1_14/a_27_47# VSS 0.39fF
C11492 Ad VSS 12.34fF
C11493 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# VSS 1.46fF
C11494 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# VSS 0.20fF
C11495 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# VSS 0.26fF
C11496 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# VSS 0.35fF
C11497 sky130_fd_sc_hd__clkdlybuf4s50_1_148/X VSS 41.58fF
C11498 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# VSS 0.20fF
C11499 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# VSS 0.27fF
C11500 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# VSS 0.37fF
C11501 sky130_fd_sc_hd__clkdlybuf4s50_1_137/A VSS 14.76fF
C11502 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# VSS 0.21fF
C11503 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# VSS 0.28fF
C11504 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# VSS 0.41fF
C11505 sky130_fd_sc_hd__clkdlybuf4s50_1_126/X VSS 9.74fF
C11506 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# VSS 0.20fF
C11507 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# VSS 0.27fF
C11508 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# VSS 0.37fF
C11509 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS 20.67fF
C11510 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_390_47# VSS 0.20fF
C11511 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_283_47# VSS 0.28fF
C11512 sky130_fd_sc_hd__clkdlybuf4s50_1_114/a_27_47# VSS 0.41fF
C11513 sky130_fd_sc_hd__nand2_4_2/B VSS 55.13fF
C11514 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# VSS 0.18fF
C11515 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# VSS 0.25fF
C11516 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# VSS 0.37fF
C11517 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# VSS 0.23fF
C11518 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# VSS 0.35fF
C11519 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# VSS 0.81fF
C11520 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS 20.68fF
C11521 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_390_47# VSS 0.20fF
C11522 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_283_47# VSS 0.28fF
C11523 sky130_fd_sc_hd__clkdlybuf4s50_1_79/a_27_47# VSS 0.41fF
C11524 sky130_fd_sc_hd__nand2_1_0/A VSS 15.19fF
C11525 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS 23.06fF
C11526 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# VSS 0.22fF
C11527 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# VSS 0.35fF
C11528 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# VSS 0.82fF
C11529 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS 41.09fF
C11530 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_390_47# VSS 0.22fF
C11531 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_283_47# VSS 0.30fF
C11532 sky130_fd_sc_hd__clkdlybuf4s50_1_35/a_27_47# VSS 0.39fF
C11533 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS 20.19fF
C11534 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_390_47# VSS 0.19fF
C11535 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_283_47# VSS 0.26fF
C11536 sky130_fd_sc_hd__clkdlybuf4s50_1_57/a_27_47# VSS 0.35fF
C11537 sky130_fd_sc_hd__clkdlybuf4s50_1_46/A VSS 23.84fF
C11538 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_390_47# VSS 0.21fF
C11539 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_283_47# VSS 0.29fF
C11540 sky130_fd_sc_hd__clkdlybuf4s50_1_46/a_27_47# VSS 0.45fF
C11541 sky130_fd_sc_hd__clkdlybuf4s50_1_14/X VSS 14.47fF
C11542 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# VSS 0.21fF
C11543 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# VSS 0.30fF
C11544 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# VSS 0.39fF
C11545 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# VSS 0.18fF
C11546 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# VSS 0.25fF
C11547 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# VSS 0.39fF
C11548 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# VSS 1.64fF
C11549 sky130_fd_sc_hd__clkdlybuf4s50_1_170/X VSS 23.92fF
C11550 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# VSS 0.21fF
C11551 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# VSS 0.29fF
C11552 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# VSS 0.39fF
C11553 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS 20.67fF
C11554 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_390_47# VSS 0.19fF
C11555 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_283_47# VSS 0.26fF
C11556 sky130_fd_sc_hd__clkdlybuf4s50_1_179/a_27_47# VSS 0.40fF
C11557 sky130_fd_sc_hd__clkdlybuf4s50_1_146/A VSS 24.60fF
C11558 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# VSS 0.21fF
C11559 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# VSS 0.29fF
C11560 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# VSS 0.38fF
C11561 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS 15.14fF
C11562 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_390_47# VSS 0.20fF
C11563 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_283_47# VSS 0.28fF
C11564 sky130_fd_sc_hd__clkdlybuf4s50_1_135/a_27_47# VSS 0.41fF
C11565 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS 23.89fF
C11566 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_390_47# VSS 0.20fF
C11567 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_283_47# VSS 0.27fF
C11568 sky130_fd_sc_hd__clkdlybuf4s50_1_124/a_27_47# VSS 0.44fF
C11569 sky130_fd_sc_hd__clkdlybuf4s50_1_114/A VSS 20.32fF
C11570 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# VSS 0.21fF
C11571 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# VSS 0.28fF
C11572 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# VSS 0.41fF
C11573 VDD VSS -38123.39fF
C11574 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS 18.11fF
C11575 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# VSS 0.19fF
C11576 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# VSS 0.25fF
C11577 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# VSS 0.37fF
C11578 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# VSS 0.21fF
C11579 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# VSS 0.27fF
C11580 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# VSS 0.35fF
C11581 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS 12.29fF
C11582 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# VSS 0.22fF
C11583 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# VSS 0.35fF
C11584 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# VSS 0.56fF
C11585 sky130_fd_sc_hd__clkdlybuf4s50_1_79/A VSS 20.32fF
C11586 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# VSS 0.21fF
C11587 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# VSS 0.29fF
C11588 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# VSS 0.41fF
C11589 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS 14.36fF
C11590 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# VSS 0.19fF
C11591 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# VSS 0.26fF
C11592 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# VSS 0.40fF
C11593 sky130_fd_sc_hd__clkdlybuf4s50_1_35/X VSS 14.73fF
C11594 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# VSS 0.21fF
C11595 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# VSS 0.30fF
C11596 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# VSS 0.39fF
C11597 sky130_fd_sc_hd__clkdlybuf4s50_1_57/X VSS 20.18fF
C11598 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# VSS 0.21fF
C11599 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# VSS 0.28fF
C11600 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# VSS 0.38fF
C11601 sky130_fd_sc_hd__clkdlybuf4s50_1_45/X VSS 20.68fF
C11602 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_390_47# VSS 0.19fF
C11603 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_283_47# VSS 0.26fF
C11604 sky130_fd_sc_hd__clkdlybuf4s50_1_45/a_27_47# VSS 0.39fF
C11605 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS 14.74fF
C11606 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_390_47# VSS 0.21fF
C11607 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_283_47# VSS 0.29fF
C11608 sky130_fd_sc_hd__clkdlybuf4s50_1_12/a_27_47# VSS 0.39fF
C11609 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS 41.04fF
C11610 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_390_47# VSS 0.18fF
C11611 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_283_47# VSS 0.25fF
C11612 sky130_fd_sc_hd__clkdlybuf4s50_1_23/a_27_47# VSS 0.39fF
C11613 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VSS 1.56fF
C11614 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS 14.82fF
C11615 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_390_47# VSS 0.21fF
C11616 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_283_47# VSS 0.29fF
C11617 sky130_fd_sc_hd__clkdlybuf4s50_1_145/a_27_47# VSS 0.39fF
C11618 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS 34.63fF
C11619 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_390_47# VSS 0.19fF
C11620 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_283_47# VSS 0.26fF
C11621 sky130_fd_sc_hd__clkdlybuf4s50_1_156/a_27_47# VSS 0.35fF
C11622 sky130_fd_sc_hd__clkdlybuf4s50_1_135/A VSS 13.93fF
C11623 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# VSS 0.20fF
C11624 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# VSS 0.27fF
C11625 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# VSS 0.40fF
C11626 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS 14.27fF
C11627 sky130_fd_sc_hd__clkdlybuf4s50_1_124/X VSS 23.97fF
C11628 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# VSS 0.20fF
C11629 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# VSS 0.27fF
C11630 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# VSS 0.38fF
C11631 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS 19.57fF
C11632 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# VSS 0.19fF
C11633 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# VSS 0.25fF
C11634 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# VSS 0.36fF
C11635 sky130_fd_sc_hd__clkinv_4_8/Y VSS 11.48fF
C11636 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# VSS 0.19fF
C11637 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# VSS 0.24fF
C11638 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# VSS 0.32fF
C11639 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS 19.93fF
C11640 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# VSS 0.18fF
C11641 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# VSS 0.25fF
C11642 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# VSS 0.40fF
C11643 sky130_fd_sc_hd__clkdlybuf4s50_1_179/A VSS 20.32fF
C11644 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS 20.13fF
C11645 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# VSS 0.20fF
C11646 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# VSS 0.27fF
C11647 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# VSS 0.41fF
C11648 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS 24.88fF
C11649 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_390_47# VSS 0.21fF
C11650 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_283_47# VSS 0.30fF
C11651 sky130_fd_sc_hd__clkdlybuf4s50_1_189/a_27_47# VSS 0.40fF
C11652 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS 47.99fF
C11653 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_390_47# VSS 0.20fF
C11654 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_283_47# VSS 0.28fF
C11655 sky130_fd_sc_hd__clkdlybuf4s50_1_88/a_27_47# VSS 0.44fF
C11656 sky130_fd_sc_hd__clkinv_4_3/Y VSS 43.40fF
C11657 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# VSS 0.19fF
C11658 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# VSS 0.24fF
C11659 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# VSS 0.33fF
C11660 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# VSS 0.19fF
C11661 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# VSS 0.24fF
C11662 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# VSS 0.34fF
C11663 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS 24.55fF
C11664 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_390_47# VSS 0.19fF
C11665 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_283_47# VSS 0.27fF
C11666 sky130_fd_sc_hd__clkdlybuf4s50_1_66/a_27_47# VSS 0.40fF
C11667 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS 29.20fF
C11668 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_390_47# VSS 0.21fF
C11669 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_283_47# VSS 0.29fF
C11670 sky130_fd_sc_hd__clkdlybuf4s50_1_33/a_27_47# VSS 0.39fF
C11671 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS 20.51fF
C11672 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_390_47# VSS 0.21fF
C11673 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_283_47# VSS 0.28fF
C11674 sky130_fd_sc_hd__clkdlybuf4s50_1_55/a_27_47# VSS 0.38fF
C11675 sky130_fd_sc_hd__clkdlybuf4s50_1_12/X VSS 9.69fF
C11676 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# VSS 0.21fF
C11677 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# VSS 0.29fF
C11678 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# VSS 0.38fF
C11679 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS 34.89fF
C11680 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS 20.30fF
C11681 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# VSS 0.20fF
C11682 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# VSS 0.27fF
C11683 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# VSS 0.41fF
C11684 sky130_fd_sc_hd__clkdlybuf4s50_1_23/A VSS 36.99fF
C11685 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# VSS 0.19fF
C11686 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# VSS 0.26fF
C11687 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# VSS 0.41fF
C11688 B_b VSS 21.34fF
C11689 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# VSS 1.52fF
C11690 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS 36.62fF
C11691 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_390_47# VSS 0.20fF
C11692 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_283_47# VSS 0.27fF
C11693 sky130_fd_sc_hd__clkdlybuf4s50_1_144/a_27_47# VSS 0.44fF
C11694 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS 20.68fF
C11695 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_390_47# VSS 0.20fF
C11696 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_283_47# VSS 0.28fF
C11697 sky130_fd_sc_hd__clkdlybuf4s50_1_133/a_27_47# VSS 0.40fF
C11698 sky130_fd_sc_hd__nand2_1_4/B VSS 40.86fF
C11699 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS 23.05fF
C11700 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# VSS 0.22fF
C11701 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# VSS 0.33fF
C11702 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# VSS 0.80fF
C11703 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS 8.39fF
C11704 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# VSS 0.20fF
C11705 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# VSS 0.27fF
C11706 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# VSS 0.49fF
C11707 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS 8.58fF
C11708 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_390_47# VSS 0.18fF
C11709 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_283_47# VSS 0.25fF
C11710 sky130_fd_sc_hd__clkdlybuf4s50_1_111/a_27_47# VSS 0.33fF
C11711 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS 49.56fF
C11712 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_390_47# VSS 0.18fF
C11713 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_283_47# VSS 0.25fF
C11714 sky130_fd_sc_hd__clkdlybuf4s50_1_166/a_27_47# VSS 0.39fF
C11715 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS 20.17fF
C11716 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_390_47# VSS 0.20fF
C11717 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_283_47# VSS 0.28fF
C11718 sky130_fd_sc_hd__clkdlybuf4s50_1_155/a_27_47# VSS 0.36fF
C11719 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS 14.39fF
C11720 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# VSS 0.21fF
C11721 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# VSS 0.27fF
C11722 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# VSS 0.35fF
C11723 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS 40.25fF
C11724 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_390_47# VSS 0.22fF
C11725 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_283_47# VSS 0.31fF
C11726 sky130_fd_sc_hd__clkdlybuf4s50_1_188/a_27_47# VSS 0.45fF
C11727 sky130_fd_sc_hd__nand2_4_3/B VSS 73.00fF
C11728 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VSS 0.19fF
C11729 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VSS 0.26fF
C11730 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# VSS 0.39fF
C11731 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS 19.82fF
C11732 sky130_fd_sc_hd__clkdlybuf4s50_1_88/X VSS 18.82fF
C11733 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# VSS 0.21fF
C11734 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# VSS 0.29fF
C11735 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# VSS 0.40fF
C11736 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS 40.46fF
C11737 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_390_47# VSS 0.19fF
C11738 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_283_47# VSS 0.26fF
C11739 sky130_fd_sc_hd__clkdlybuf4s50_1_98/a_27_47# VSS 0.34fF
C11740 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS 20.22fF
C11741 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_390_47# VSS 0.19fF
C11742 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_283_47# VSS 0.26fF
C11743 sky130_fd_sc_hd__clkdlybuf4s50_1_76/a_27_47# VSS 0.35fF
C11744 sky130_fd_sc_hd__clkdlybuf4s50_1_66/A VSS 24.18fF
C11745 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# VSS 0.21fF
C11746 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# VSS 0.28fF
C11747 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# VSS 0.42fF
C11748 sky130_fd_sc_hd__clkdlybuf4s50_1_33/X VSS 49.24fF
C11749 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# VSS 0.21fF
C11750 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# VSS 0.29fF
C11751 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# VSS 0.38fF
C11752 sky130_fd_sc_hd__clkdlybuf4s50_1_55/X VSS 7.58fF
C11753 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# VSS 0.20fF
C11754 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# VSS 0.28fF
C11755 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# VSS 0.38fF
C11756 sky130_fd_sc_hd__clkdlybuf4s50_1_43/X VSS 35.04fF
C11757 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_390_47# VSS 0.19fF
C11758 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_283_47# VSS 0.26fF
C11759 sky130_fd_sc_hd__clkdlybuf4s50_1_43/a_27_47# VSS 0.40fF
C11760 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS 35.49fF
C11761 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_390_47# VSS 0.20fF
C11762 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_283_47# VSS 0.26fF
C11763 sky130_fd_sc_hd__clkdlybuf4s50_1_21/a_27_47# VSS 0.41fF
C11764 sky130_fd_sc_hd__clkdlybuf4s50_1_9/X VSS 24.59fF
C11765 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# VSS 0.20fF
C11766 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# VSS 0.29fF
C11767 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# VSS 0.38fF
C11768 Bd VSS 15.05fF
C11769 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# VSS 1.51fF
C11770 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS 22.18fF
C11771 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_390_47# VSS 0.21fF
C11772 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_283_47# VSS 0.29fF
C11773 sky130_fd_sc_hd__clkdlybuf4s50_1_143/a_27_47# VSS 0.45fF
C11774 sky130_fd_sc_hd__clkdlybuf4s50_1_156/X VSS 34.73fF
C11775 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# VSS 0.21fF
C11776 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# VSS 0.28fF
C11777 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# VSS 0.38fF
C11778 sky130_fd_sc_hd__clkdlybuf4s50_1_133/A VSS 20.32fF
C11779 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# VSS 0.21fF
C11780 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# VSS 0.28fF
C11781 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# VSS 0.41fF
C11782 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS 14.43fF
C11783 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# VSS 0.19fF
C11784 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# VSS 0.26fF
C11785 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# VSS 0.40fF
C11786 sky130_fd_sc_hd__clkdlybuf4s50_1_110/A VSS 8.60fF
C11787 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_390_47# VSS 0.19fF
C11788 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_283_47# VSS 0.27fF
C11789 sky130_fd_sc_hd__clkdlybuf4s50_1_110/a_27_47# VSS 0.36fF
C11790 sky130_fd_sc_hd__clkdlybuf4s50_1_165/X VSS 38.85fF
C11791 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_390_47# VSS 0.20fF
C11792 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_283_47# VSS 0.26fF
C11793 sky130_fd_sc_hd__clkdlybuf4s50_1_165/a_27_47# VSS 0.41fF
C11794 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS 20.17fF
C11795 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_390_47# VSS 0.20fF
C11796 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_283_47# VSS 0.28fF
C11797 sky130_fd_sc_hd__clkdlybuf4s50_1_176/a_27_47# VSS 0.36fF
C11798 sky130_fd_sc_hd__clkdlybuf4s50_1_188/X VSS 13.67fF
C11799 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# VSS 0.22fF
C11800 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# VSS 0.31fF
C11801 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# VSS 0.41fF
C11802 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS 24.15fF
C11803 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VSS 0.22fF
C11804 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VSS 0.31fF
C11805 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VSS 0.45fF
C11806 sky130_fd_sc_hd__nand2_4_1/B VSS 72.93fF
C11807 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# VSS 0.21fF
C11808 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# VSS 0.27fF
C11809 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# VSS 0.40fF
C11810 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS 14.40fF
C11811 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# VSS 0.19fF
C11812 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# VSS 0.26fF
C11813 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# VSS 0.40fF
C11814 sky130_fd_sc_hd__clkdlybuf4s50_1_76/X VSS 20.16fF
C11815 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# VSS 0.21fF
C11816 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# VSS 0.27fF
C11817 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# VSS 0.37fF
C11818 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS 19.05fF
C11819 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_390_47# VSS 0.21fF
C11820 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_283_47# VSS 0.28fF
C11821 sky130_fd_sc_hd__clkdlybuf4s50_1_64/a_27_47# VSS 0.41fF
C11822 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS 14.80fF
C11823 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_390_47# VSS 0.20fF
C11824 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_283_47# VSS 0.27fF
C11825 sky130_fd_sc_hd__clkdlybuf4s50_1_53/a_27_47# VSS 0.38fF
C11826 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# VSS 0.18fF
C11827 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# VSS 0.25fF
C11828 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# VSS 0.40fF
C11829 sky130_fd_sc_hd__clkdlybuf4s50_1_21/A VSS 24.91fF
C11830 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# VSS 0.20fF
C11831 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# VSS 0.26fF
C11832 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# VSS 0.40fF
C11833 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS 9.64fF
C11834 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# VSS 0.21fF
C11835 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# VSS 0.30fF
C11836 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# VSS 0.39fF
C11837 B VSS 14.98fF
C11838 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# VSS 1.49fF
C11839 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS 35.38fF
C11840 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_390_47# VSS 0.21fF
C11841 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_283_47# VSS 0.28fF
C11842 sky130_fd_sc_hd__clkdlybuf4s50_1_153/a_27_47# VSS 0.38fF
C11843 sky130_fd_sc_hd__clkdlybuf4s50_1_144/X VSS 40.66fF
C11844 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# VSS 0.21fF
C11845 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# VSS 0.28fF
C11846 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# VSS 0.39fF
C11847 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# VSS 0.19fF
C11848 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# VSS 0.24fF
C11849 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# VSS 0.34fF
C11850 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS 24.55fF
C11851 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_390_47# VSS 0.19fF
C11852 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_283_47# VSS 0.27fF
C11853 sky130_fd_sc_hd__clkdlybuf4s50_1_120/a_27_47# VSS 0.40fF
C11854 sky130_fd_sc_hd__clkdlybuf4s50_1_166/A VSS 49.58fF
C11855 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# VSS 0.19fF
C11856 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# VSS 0.26fF
C11857 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# VSS 0.41fF
C11858 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_390_47# VSS 0.22fF
C11859 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_283_47# VSS 0.30fF
C11860 sky130_fd_sc_hd__clkdlybuf4s50_1_175/a_27_47# VSS 0.39fF
C11861 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# VSS 0.18fF
C11862 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# VSS 0.25fF
C11863 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# VSS 0.40fF
C11864 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS 25.83fF
C11865 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# VSS 0.20fF
C11866 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# VSS 0.26fF
C11867 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# VSS 0.39fF
C11868 sky130_fd_sc_hd__clkdlybuf4s50_1_98/X VSS 40.42fF
C11869 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# VSS 0.21fF
C11870 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# VSS 0.28fF
C11871 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# VSS 0.38fF
C11872 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS 24.55fF
C11873 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_390_47# VSS 0.19fF
C11874 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_283_47# VSS 0.27fF
C11875 sky130_fd_sc_hd__clkdlybuf4s50_1_85/a_27_47# VSS 0.40fF
C11876 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS 20.48fF
C11877 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_390_47# VSS 0.20fF
C11878 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_283_47# VSS 0.28fF
C11879 sky130_fd_sc_hd__clkdlybuf4s50_1_74/a_27_47# VSS 0.38fF
C11880 sky130_fd_sc_hd__clkdlybuf4s50_1_64/A VSS 14.76fF
C11881 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# VSS 0.21fF
C11882 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# VSS 0.28fF
C11883 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# VSS 0.41fF
C11884 sky130_fd_sc_hd__clkdlybuf4s50_1_53/X VSS 24.59fF
C11885 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# VSS 0.20fF
C11886 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# VSS 0.27fF
C11887 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# VSS 0.37fF
C11888 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS 24.55fF
C11889 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_390_47# VSS 0.18fF
C11890 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_283_47# VSS 0.25fF
C11891 sky130_fd_sc_hd__clkdlybuf4s50_1_30/a_27_47# VSS 0.39fF
C11892 sky130_fd_sc_hd__clkdlybuf4s50_1_41/A VSS 23.90fF
C11893 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_390_47# VSS 0.20fF
C11894 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_283_47# VSS 0.29fF
C11895 sky130_fd_sc_hd__clkdlybuf4s50_1_41/a_27_47# VSS 0.44fF
C11896 sky130_fd_sc_hd__clkdlybuf4s50_1_165/A VSS 29.90fF
C11897 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# VSS 0.20fF
C11898 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# VSS 0.26fF
C11899 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# VSS 0.40fF
C11900 sky130_fd_sc_hd__clkdlybuf4s50_1_155/X VSS 20.20fF
C11901 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# VSS 0.22fF
C11902 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# VSS 0.30fF
C11903 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# VSS 0.39fF
C11904 sky130_fd_sc_hd__clkdlybuf4s50_1_175/A VSS 20.43fF
C11905 sky130_fd_sc_hd__clkdlybuf4s50_1_176/X VSS 20.10fF
C11906 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# VSS 0.22fF
C11907 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# VSS 0.30fF
C11908 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# VSS 0.39fF
C11909 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS 24.53fF
C11910 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_390_47# VSS 0.18fF
C11911 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_283_47# VSS 0.25fF
C11912 sky130_fd_sc_hd__clkdlybuf4s50_1_185/a_27_47# VSS 0.39fF
C11913 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS 12.67fF
C11914 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# VSS 0.20fF
C11915 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# VSS 0.28fF
C11916 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VSS 0.53fF
C11917 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS 22.84fF
C11918 sky130_fd_sc_hd__clkdlybuf4s50_1_143/X VSS 23.95fF
C11919 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# VSS 0.22fF
C11920 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# VSS 0.30fF
C11921 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# VSS 0.40fF
C11922 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS 20.22fF
C11923 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_390_47# VSS 0.19fF
C11924 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_283_47# VSS 0.26fF
C11925 sky130_fd_sc_hd__clkdlybuf4s50_1_130/a_27_47# VSS 0.35fF
C11926 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS 24.09fF
C11927 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# VSS 0.23fF
C11928 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# VSS 0.32fF
C11929 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# VSS 0.45fF
C11930 sky130_fd_sc_hd__clkdlybuf4s50_1_85/A VSS 22.46fF
C11931 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# VSS 0.21fF
C11932 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# VSS 0.28fF
C11933 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# VSS 0.43fF
C11934 sky130_fd_sc_hd__clkdlybuf4s50_1_74/X VSS 14.52fF
C11935 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# VSS 0.20fF
C11936 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# VSS 0.28fF
C11937 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# VSS 0.38fF
C11938 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS 15.14fF
C11939 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_390_47# VSS 0.20fF
C11940 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_283_47# VSS 0.28fF
C11941 sky130_fd_sc_hd__clkdlybuf4s50_1_62/a_27_47# VSS 0.41fF
C11942 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS 22.17fF
C11943 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_390_47# VSS 0.20fF
C11944 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_283_47# VSS 0.27fF
C11945 sky130_fd_sc_hd__clkdlybuf4s50_1_51/a_27_47# VSS 0.44fF
C11946 sky130_fd_sc_hd__clkdlybuf4s50_1_40/A VSS 44.24fF
C11947 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_390_47# VSS 0.21fF
C11948 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_283_47# VSS 0.29fF
C11949 sky130_fd_sc_hd__clkdlybuf4s50_1_40/a_27_47# VSS 0.45fF
C11950 sky130_fd_sc_hd__clkdlybuf4s50_1_162/X VSS 27.79fF
C11951 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# VSS 0.19fF
C11952 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# VSS 0.26fF
C11953 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# VSS 0.39fF
C11954 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS 20.42fF
C11955 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# VSS 0.19fF
C11956 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# VSS 0.26fF
C11957 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# VSS 0.40fF
C11958 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS 20.53fF
C11959 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_390_47# VSS 0.22fF
C11960 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_283_47# VSS 0.30fF
C11961 sky130_fd_sc_hd__clkdlybuf4s50_1_151/a_27_47# VSS 0.39fF
C11962 sky130_fd_sc_hd__clkdlybuf4s50_1_175/X VSS 14.47fF
C11963 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# VSS 0.21fF
C11964 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# VSS 0.30fF
C11965 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# VSS 0.39fF
C11966 sky130_fd_sc_hd__clkdlybuf4s50_1_185/A VSS 22.44fF
C11967 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# VSS 0.20fF
C11968 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# VSS 0.27fF
C11969 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# VSS 0.41fF
C11970 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# VSS 0.21fF
C11971 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# VSS 0.27fF
C11972 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# VSS 0.35fF
C11973 sky130_fd_sc_hd__dfxbp_1_1/D VSS 8.30fF
C11974 sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# VSS -0.00fF
C11975 sky130_fd_sc_hd__dfxbp_1_1/a_592_47# VSS -0.00fF
C11976 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# VSS 0.05fF
C11977 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# VSS 0.16fF
C11978 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# VSS 0.19fF
C11979 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# VSS 0.36fF
C11980 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# VSS 0.16fF
C11981 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# VSS 0.04fF
C11982 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VSS 0.33fF
C11983 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VSS 0.53fF
C11984 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS 41.20fF
C11985 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_390_47# VSS 0.20fF
C11986 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_283_47# VSS 0.28fF
C11987 sky130_fd_sc_hd__clkdlybuf4s50_1_94/a_27_47# VSS 0.38fF
C11988 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS 20.78fF
C11989 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_390_47# VSS 0.21fF
C11990 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_283_47# VSS 0.29fF
C11991 sky130_fd_sc_hd__clkdlybuf4s50_1_83/a_27_47# VSS 0.42fF
C11992 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS 14.79fF
C11993 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_390_47# VSS 0.20fF
C11994 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_283_47# VSS 0.28fF
C11995 sky130_fd_sc_hd__clkdlybuf4s50_1_72/a_27_47# VSS 0.38fF
C11996 sky130_fd_sc_hd__clkdlybuf4s50_1_62/A VSS 13.93fF
C11997 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# VSS 0.20fF
C11998 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# VSS 0.27fF
C11999 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# VSS 0.40fF
C12000 sky130_fd_sc_hd__clkdlybuf4s50_1_51/X VSS 24.00fF
C12001 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# VSS 0.21fF
C12002 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# VSS 0.28fF
C12003 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# VSS 0.39fF
C12004 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS 30.28fF
C12005 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_390_47# VSS 0.19fF
C12006 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_283_47# VSS 0.26fF
C12007 sky130_fd_sc_hd__clkdlybuf4s50_1_161/a_27_47# VSS 0.40fF
C12008 sky130_fd_sc_hd__clkdlybuf4s50_1_153/X VSS 11.72fF
C12009 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# VSS 0.20fF
C12010 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# VSS 0.28fF
C12011 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# VSS 0.38fF
C12012 sky130_fd_sc_hd__clkdlybuf4s50_1_172/A VSS 9.69fF
C12013 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# VSS 0.21fF
C12014 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# VSS 0.29fF
C12015 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# VSS 0.38fF
C12016 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS 20.77fF
C12017 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_390_47# VSS 0.20fF
C12018 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_283_47# VSS 0.26fF
C12019 sky130_fd_sc_hd__clkdlybuf4s50_1_183/a_27_47# VSS 0.41fF
C12020 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS 34.52fF
C12021 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_390_47# VSS 0.20fF
C12022 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_283_47# VSS 0.28fF
C12023 sky130_fd_sc_hd__clkdlybuf4s50_1_194/a_27_47# VSS 0.36fF
C12024 sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS 0.22fF
C12025 sky130_fd_sc_hd__nand2_1_1/A VSS 49.47fF
C12026 sky130_fd_sc_hd__dfxbp_1_0/a_1017_47# VSS 0.22fF
C12027 sky130_fd_sc_hd__dfxbp_1_0/a_592_47# VSS 0.01fF
C12028 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VSS 0.07fF
C12029 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VSS 0.16fF
C12030 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VSS 0.21fF
C12031 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VSS 0.36fF
C12032 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VSS 0.18fF
C12033 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VSS 0.19fF
C12034 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VSS 0.38fF
C12035 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VSS 0.56fF
C12036 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS 25.77fF
C12037 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# VSS 0.23fF
C12038 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# VSS 0.32fF
C12039 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# VSS 0.44fF
C12040 sky130_fd_sc_hd__clkdlybuf4s50_1_83/A VSS 14.76fF
C12041 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# VSS 0.21fF
C12042 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# VSS 0.29fF
C12043 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# VSS 0.41fF
C12044 sky130_fd_sc_hd__clkdlybuf4s50_1_72/X VSS 9.74fF
C12045 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# VSS 0.20fF
C12046 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# VSS 0.27fF
C12047 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# VSS 0.37fF
C12048 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS 20.68fF
C12049 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_390_47# VSS 0.20fF
C12050 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_283_47# VSS 0.28fF
C12051 sky130_fd_sc_hd__clkdlybuf4s50_1_60/a_27_47# VSS 0.40fF
C12052 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS 41.71fF
C12053 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_390_47# VSS 0.19fF
C12054 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_283_47# VSS 0.26fF
C12055 sky130_fd_sc_hd__clkdlybuf4s50_1_160/a_27_47# VSS 0.39fF
C12056 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS 14.74fF
C12057 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_390_47# VSS 0.21fF
C12058 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_283_47# VSS 0.29fF
C12059 sky130_fd_sc_hd__clkdlybuf4s50_1_171/a_27_47# VSS 0.39fF
C12060 sky130_fd_sc_hd__clkdlybuf4s50_1_183/A VSS 14.76fF
C12061 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# VSS 0.20fF
C12062 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# VSS 0.27fF
C12063 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# VSS 0.41fF
C12064 sky130_fd_sc_hd__clkdlybuf4s50_1_194/X VSS 34.45fF
C12065 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# VSS 0.23fF
C12066 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# VSS 0.30fF
C12067 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# VSS 0.39fF
C12068 sky130_fd_sc_hd__nand2_4_3/Y VSS 112.17fF
C12069 sky130_fd_sc_hd__clkdlybuf4s50_1_94/X VSS 29.01fF
C12070 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# VSS 0.20fF
C12071 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# VSS 0.28fF
C12072 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# VSS 0.38fF
C12073 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS 8.15fF
C12074 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_390_47# VSS 0.21fF
C12075 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_283_47# VSS 0.28fF
C12076 sky130_fd_sc_hd__clkdlybuf4s50_1_81/a_27_47# VSS 0.41fF
C12077 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS 23.89fF
C12078 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_390_47# VSS 0.20fF
C12079 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_283_47# VSS 0.27fF
C12080 sky130_fd_sc_hd__clkdlybuf4s50_1_70/a_27_47# VSS 0.44fF
C12081 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS 23.84fF
C12082 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_390_47# VSS 0.21fF
C12083 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_283_47# VSS 0.29fF
C12084 sky130_fd_sc_hd__clkdlybuf4s50_1_170/a_27_47# VSS 0.45fF
C12085 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS 8.14fF
C12086 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_390_47# VSS 0.19fF
C12087 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_283_47# VSS 0.26fF
C12088 sky130_fd_sc_hd__clkdlybuf4s50_1_181/a_27_47# VSS 0.40fF
C12089 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS 35.11fF
C12090 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_390_47# VSS 0.22fF
C12091 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_283_47# VSS 0.30fF
C12092 sky130_fd_sc_hd__clkdlybuf4s50_1_192/a_27_47# VSS 0.39fF
C12093 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS 29.33fF
C12094 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_390_47# VSS 0.20fF
C12095 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_283_47# VSS 0.28fF
C12096 sky130_fd_sc_hd__clkdlybuf4s50_1_91/a_27_47# VSS 0.39fF
C12097 sky130_fd_sc_hd__clkdlybuf4s50_1_81/A VSS 20.88fF
C12098 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VSS 0.20fF
C12099 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VSS 0.28fF
C12100 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VSS 0.41fF
C12101 sky130_fd_sc_hd__clkdlybuf4s50_1_181/A VSS 20.88fF
C12102 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VSS 0.19fF
C12103 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VSS 0.26fF
C12104 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VSS 0.40fF
C12105 sky130_fd_sc_hd__clkdlybuf4s50_1_192/X VSS 24.58fF
C12106 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VSS 0.22fF
C12107 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VSS 0.31fF
C12108 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VSS 0.40fF
C12109 sky130_fd_sc_hd__clkinv_4_7/Y VSS 28.94fF
C12110 sky130_fd_sc_hd__clkdlybuf4s50_1_91/X VSS 49.41fF
C12111 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VSS 0.19fF
C12112 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VSS 0.28fF
C12113 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VSS 0.38fF
C12114 sky130_fd_sc_hd__clkdlybuf4s50_1_190/A VSS 41.43fF
C12115 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VSS 0.21fF
C12116 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VSS 0.30fF
C12117 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VSS 0.39fF
C12118 sky130_fd_sc_hd__clkdlybuf4s50_1_9/A VSS 14.82fF
C12119 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_390_47# VSS 0.21fF
C12120 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_283_47# VSS 0.30fF
C12121 sky130_fd_sc_hd__clkdlybuf4s50_1_9/a_27_47# VSS 0.39fF
C12122 sky130_fd_sc_hd__clkinv_4_4/Y VSS 28.94fF
C12123 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS 14.52fF
C12124 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VSS 0.21fF
C12125 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VSS 0.30fF
C12126 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VSS 0.39fF
C12127 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_390_47# VSS 0.21fF
C12128 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_283_47# VSS 0.29fF
C12129 sky130_fd_sc_hd__clkdlybuf4s50_1_7/a_27_47# VSS 0.38fF
C12130 sky130_fd_sc_hd__nand2_4_0/Y VSS 64.76fF
C12131 sky130_fd_sc_hd__clkdlybuf4s50_1_7/A VSS 20.48fF
C12132 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS 20.15fF
C12133 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VSS 0.21fF
C12134 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VSS 0.29fF
C12135 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VSS 0.38fF
C12136 sky130_fd_sc_hd__nand2_4_3/a_27_47# VSS 0.38fF
C12137 sky130_fd_sc_hd__clkinv_4_1/Y VSS 58.23fF
C12138 sky130_fd_sc_hd__clkinv_4_1/A VSS 127.09fF
C12139 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VSS 0.20fF
C12140 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VSS 0.26fF
C12141 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VSS 0.34fF
C12142 sky130_fd_sc_hd__nand2_4_2/Y VSS 64.29fF
C12143 sky130_fd_sc_hd__nand2_4_2/a_27_47# VSS 0.35fF
C12144 sky130_fd_sc_hd__clkdlybuf4s50_1_5/X VSS 20.20fF
C12145 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_390_47# VSS 0.20fF
C12146 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_283_47# VSS 0.28fF
C12147 sky130_fd_sc_hd__clkdlybuf4s50_1_4/a_27_47# VSS 0.36fF
C12148 sky130_fd_sc_hd__nand2_4_1/Y VSS 66.78fF
C12149 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.40fF
C12150 sky130_fd_sc_hd__nand2_4_0/B VSS 72.94fF
C12151 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VSS 0.18fF
C12152 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VSS 0.25fF
C12153 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VSS 0.37fF
C12154 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.35fF
C12155 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS 24.11fF
C12156 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VSS 0.19fF
C12157 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VSS 0.25fF
C12158 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VSS 0.38fF
C12159 p2 VSS 59.01fF
C12160 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VSS 1.52fF
C12161 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS 25.77fF
C12162 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VSS 0.19fF
C12163 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VSS 0.25fF
C12164 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VSS 0.37fF
C12165 sky130_fd_sc_hd__clkinv_4_10/Y VSS 29.07fF
C12166 sky130_fd_sc_hd__clkinv_1_3/A VSS 100.50fF
C12167 p2_b VSS 15.65fF
C12168 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VSS 1.52fF
C12169 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS 12.52fF
C12170 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VSS 0.19fF
C12171 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VSS 0.27fF
C12172 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VSS 0.49fF
C12173 p2d VSS 15.07fF
C12174 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VSS 1.51fF
C12175 p2d_b VSS 23.55fF
C12176 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VSS 1.57fF
C12177 p1d_b VSS 12.85fF
C12178 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VSS 1.63fF
.ends

