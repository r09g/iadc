* NGSPICE file created from _flat.ext - technology: sky130A


* Top level circuit _flat

.end

