magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< error_p >>
rect -1469 172 -1411 178
rect -1277 172 -1219 178
rect -1085 172 -1027 178
rect -893 172 -835 178
rect -701 172 -643 178
rect -509 172 -451 178
rect -317 172 -259 178
rect -125 172 -67 178
rect 67 172 125 178
rect 259 172 317 178
rect 451 172 509 178
rect 643 172 701 178
rect 835 172 893 178
rect 1027 172 1085 178
rect 1219 172 1277 178
rect 1411 172 1469 178
rect -1469 138 -1457 172
rect -1277 138 -1265 172
rect -1085 138 -1073 172
rect -893 138 -881 172
rect -701 138 -689 172
rect -509 138 -497 172
rect -317 138 -305 172
rect -125 138 -113 172
rect 67 138 79 172
rect 259 138 271 172
rect 451 138 463 172
rect 643 138 655 172
rect 835 138 847 172
rect 1027 138 1039 172
rect 1219 138 1231 172
rect 1411 138 1423 172
rect -1469 132 -1411 138
rect -1277 132 -1219 138
rect -1085 132 -1027 138
rect -893 132 -835 138
rect -701 132 -643 138
rect -509 132 -451 138
rect -317 132 -259 138
rect -125 132 -67 138
rect 67 132 125 138
rect 259 132 317 138
rect 451 132 509 138
rect 643 132 701 138
rect 835 132 893 138
rect 1027 132 1085 138
rect 1219 132 1277 138
rect 1411 132 1469 138
<< pwell >>
rect -1799 -310 1799 310
<< nmos >>
rect -1599 -100 -1569 100
rect -1503 -100 -1473 100
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
rect 1473 -100 1503 100
rect 1569 -100 1599 100
<< ndiff >>
rect -1661 88 -1599 100
rect -1661 -88 -1649 88
rect -1615 -88 -1599 88
rect -1661 -100 -1599 -88
rect -1569 88 -1503 100
rect -1569 -88 -1553 88
rect -1519 -88 -1503 88
rect -1569 -100 -1503 -88
rect -1473 88 -1407 100
rect -1473 -88 -1457 88
rect -1423 -88 -1407 88
rect -1473 -100 -1407 -88
rect -1377 88 -1311 100
rect -1377 -88 -1361 88
rect -1327 -88 -1311 88
rect -1377 -100 -1311 -88
rect -1281 88 -1215 100
rect -1281 -88 -1265 88
rect -1231 -88 -1215 88
rect -1281 -100 -1215 -88
rect -1185 88 -1119 100
rect -1185 -88 -1169 88
rect -1135 -88 -1119 88
rect -1185 -100 -1119 -88
rect -1089 88 -1023 100
rect -1089 -88 -1073 88
rect -1039 -88 -1023 88
rect -1089 -100 -1023 -88
rect -993 88 -927 100
rect -993 -88 -977 88
rect -943 -88 -927 88
rect -993 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 993 100
rect 927 -88 943 88
rect 977 -88 993 88
rect 927 -100 993 -88
rect 1023 88 1089 100
rect 1023 -88 1039 88
rect 1073 -88 1089 88
rect 1023 -100 1089 -88
rect 1119 88 1185 100
rect 1119 -88 1135 88
rect 1169 -88 1185 88
rect 1119 -100 1185 -88
rect 1215 88 1281 100
rect 1215 -88 1231 88
rect 1265 -88 1281 88
rect 1215 -100 1281 -88
rect 1311 88 1377 100
rect 1311 -88 1327 88
rect 1361 -88 1377 88
rect 1311 -100 1377 -88
rect 1407 88 1473 100
rect 1407 -88 1423 88
rect 1457 -88 1473 88
rect 1407 -100 1473 -88
rect 1503 88 1569 100
rect 1503 -88 1519 88
rect 1553 -88 1569 88
rect 1503 -100 1569 -88
rect 1599 88 1661 100
rect 1599 -88 1615 88
rect 1649 -88 1661 88
rect 1599 -100 1661 -88
<< ndiffc >>
rect -1649 -88 -1615 88
rect -1553 -88 -1519 88
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect 1519 -88 1553 88
rect 1615 -88 1649 88
<< psubdiff >>
rect -1763 240 -1667 274
rect 1667 240 1763 274
rect -1763 178 -1729 240
rect 1729 178 1763 240
rect -1763 -240 -1729 -178
rect 1729 -240 1763 -178
rect -1763 -274 -1667 -240
rect 1667 -274 1763 -240
<< psubdiffcont >>
rect -1667 240 1667 274
rect -1763 -178 -1729 178
rect 1729 -178 1763 178
rect -1667 -274 1667 -240
<< poly >>
rect -1521 172 1521 188
rect -1521 138 -1457 172
rect -1423 138 -1265 172
rect -1231 138 -1073 172
rect -1039 138 -881 172
rect -847 138 -689 172
rect -655 138 -497 172
rect -463 138 -305 172
rect -271 138 -113 172
rect -79 138 79 172
rect 113 138 271 172
rect 305 138 463 172
rect 497 138 655 172
rect 689 138 847 172
rect 881 138 1039 172
rect 1073 138 1231 172
rect 1265 138 1423 172
rect 1457 138 1521 172
rect -1599 100 -1569 126
rect -1521 122 1521 138
rect -1503 100 -1473 122
rect -1407 100 -1377 122
rect -1311 100 -1281 122
rect -1215 100 -1185 122
rect -1119 100 -1089 122
rect -1023 100 -993 122
rect -927 100 -897 122
rect -831 100 -801 122
rect -735 100 -705 122
rect -639 100 -609 122
rect -543 100 -513 122
rect -447 100 -417 122
rect -351 100 -321 122
rect -255 100 -225 122
rect -159 100 -129 122
rect -63 100 -33 122
rect 33 100 63 122
rect 129 100 159 122
rect 225 100 255 122
rect 321 100 351 122
rect 417 100 447 122
rect 513 100 543 122
rect 609 100 639 122
rect 705 100 735 122
rect 801 100 831 122
rect 897 100 927 122
rect 993 100 1023 122
rect 1089 100 1119 122
rect 1185 100 1215 122
rect 1281 100 1311 122
rect 1377 100 1407 122
rect 1473 100 1503 122
rect 1569 100 1599 126
rect -1599 -122 -1569 -100
rect -1617 -138 -1551 -122
rect -1503 -126 -1473 -100
rect -1407 -126 -1377 -100
rect -1311 -126 -1281 -100
rect -1215 -126 -1185 -100
rect -1119 -126 -1089 -100
rect -1023 -126 -993 -100
rect -927 -126 -897 -100
rect -831 -126 -801 -100
rect -735 -126 -705 -100
rect -639 -126 -609 -100
rect -543 -126 -513 -100
rect -447 -126 -417 -100
rect -351 -126 -321 -100
rect -255 -126 -225 -100
rect -159 -126 -129 -100
rect -63 -126 -33 -100
rect 33 -126 63 -100
rect 129 -126 159 -100
rect 225 -126 255 -100
rect 321 -126 351 -100
rect 417 -126 447 -100
rect 513 -126 543 -100
rect 609 -126 639 -100
rect 705 -126 735 -100
rect 801 -126 831 -100
rect 897 -126 927 -100
rect 993 -126 1023 -100
rect 1089 -126 1119 -100
rect 1185 -126 1215 -100
rect 1281 -126 1311 -100
rect 1377 -126 1407 -100
rect 1473 -126 1503 -100
rect 1569 -126 1599 -100
rect -1617 -172 -1601 -138
rect -1567 -172 -1551 -138
rect -1617 -188 -1551 -172
rect 1551 -142 1617 -126
rect 1551 -176 1567 -142
rect 1601 -176 1617 -142
rect 1551 -192 1617 -176
<< polycont >>
rect -1457 138 -1423 172
rect -1265 138 -1231 172
rect -1073 138 -1039 172
rect -881 138 -847 172
rect -689 138 -655 172
rect -497 138 -463 172
rect -305 138 -271 172
rect -113 138 -79 172
rect 79 138 113 172
rect 271 138 305 172
rect 463 138 497 172
rect 655 138 689 172
rect 847 138 881 172
rect 1039 138 1073 172
rect 1231 138 1265 172
rect 1423 138 1457 172
rect -1601 -172 -1567 -138
rect 1567 -176 1601 -142
<< locali >>
rect -1763 240 -1667 274
rect 1667 240 1763 274
rect -1763 178 -1729 240
rect 1729 178 1763 240
rect -1473 138 -1457 172
rect -1423 138 -1407 172
rect -1281 138 -1265 172
rect -1231 138 -1215 172
rect -1089 138 -1073 172
rect -1039 138 -1023 172
rect -897 138 -881 172
rect -847 138 -831 172
rect -705 138 -689 172
rect -655 138 -639 172
rect -513 138 -497 172
rect -463 138 -447 172
rect -321 138 -305 172
rect -271 138 -255 172
rect -129 138 -113 172
rect -79 138 -63 172
rect 63 138 79 172
rect 113 138 129 172
rect 255 138 271 172
rect 305 138 321 172
rect 447 138 463 172
rect 497 138 513 172
rect 639 138 655 172
rect 689 138 705 172
rect 831 138 847 172
rect 881 138 897 172
rect 1023 138 1039 172
rect 1073 138 1089 172
rect 1215 138 1231 172
rect 1265 138 1281 172
rect 1407 138 1423 172
rect 1457 138 1473 172
rect -1763 -240 -1729 -178
rect -1649 88 -1615 104
rect -1649 -138 -1615 -88
rect -1553 88 -1519 104
rect -1553 -104 -1519 -88
rect -1457 88 -1423 104
rect -1457 -104 -1423 -88
rect -1361 88 -1327 104
rect -1361 -104 -1327 -88
rect -1265 88 -1231 104
rect -1265 -104 -1231 -88
rect -1169 88 -1135 104
rect -1169 -104 -1135 -88
rect -1073 88 -1039 104
rect -1073 -104 -1039 -88
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect 1039 88 1073 104
rect 1039 -104 1073 -88
rect 1135 88 1169 104
rect 1135 -104 1169 -88
rect 1231 88 1265 104
rect 1231 -104 1265 -88
rect 1327 88 1361 104
rect 1327 -104 1361 -88
rect 1423 88 1457 104
rect 1423 -104 1457 -88
rect 1519 88 1553 104
rect 1519 -104 1553 -88
rect 1615 88 1649 104
rect -1649 -172 -1601 -138
rect -1567 -172 -1551 -138
rect 1615 -142 1649 -88
rect -1649 -240 -1615 -172
rect 1551 -176 1567 -142
rect 1601 -176 1649 -142
rect 1615 -240 1649 -176
rect 1729 -240 1763 -178
rect -1763 -274 -1667 -240
rect 1667 -274 1763 -240
<< viali >>
rect -1457 138 -1423 172
rect -1265 138 -1231 172
rect -1073 138 -1039 172
rect -881 138 -847 172
rect -689 138 -655 172
rect -497 138 -463 172
rect -305 138 -271 172
rect -113 138 -79 172
rect 79 138 113 172
rect 271 138 305 172
rect 463 138 497 172
rect 655 138 689 172
rect 847 138 881 172
rect 1039 138 1073 172
rect 1231 138 1265 172
rect 1423 138 1457 172
<< metal1 >>
rect -1469 172 -1411 178
rect -1469 138 -1457 172
rect -1423 138 -1411 172
rect -1469 132 -1411 138
rect -1277 172 -1219 178
rect -1277 138 -1265 172
rect -1231 138 -1219 172
rect -1277 132 -1219 138
rect -1085 172 -1027 178
rect -1085 138 -1073 172
rect -1039 138 -1027 172
rect -1085 132 -1027 138
rect -893 172 -835 178
rect -893 138 -881 172
rect -847 138 -835 172
rect -893 132 -835 138
rect -701 172 -643 178
rect -701 138 -689 172
rect -655 138 -643 172
rect -701 132 -643 138
rect -509 172 -451 178
rect -509 138 -497 172
rect -463 138 -451 172
rect -509 132 -451 138
rect -317 172 -259 178
rect -317 138 -305 172
rect -271 138 -259 172
rect -317 132 -259 138
rect -125 172 -67 178
rect -125 138 -113 172
rect -79 138 -67 172
rect -125 132 -67 138
rect 67 172 125 178
rect 67 138 79 172
rect 113 138 125 172
rect 67 132 125 138
rect 259 172 317 178
rect 259 138 271 172
rect 305 138 317 172
rect 259 132 317 138
rect 451 172 509 178
rect 451 138 463 172
rect 497 138 509 172
rect 451 132 509 138
rect 643 172 701 178
rect 643 138 655 172
rect 689 138 701 172
rect 643 132 701 138
rect 835 172 893 178
rect 835 138 847 172
rect 881 138 893 172
rect 835 132 893 138
rect 1027 172 1085 178
rect 1027 138 1039 172
rect 1073 138 1085 172
rect 1027 132 1085 138
rect 1219 172 1277 178
rect 1219 138 1231 172
rect 1265 138 1277 172
rect 1219 132 1277 138
rect 1411 172 1469 178
rect 1411 138 1423 172
rect 1457 138 1469 172
rect 1411 132 1469 138
<< properties >>
string FIXED_BBOX -1746 -256 1746 256
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 34 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
