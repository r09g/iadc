* user analog project wrapper gold spice netlist

.include "sky130_fd_sc_hd.spice"

.subckt user_analog_project_wrapper_gold vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0] user_clock2
+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0] io_clamp_high[2],io_clamp_high[1],io_clamp_high[0] io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
+ user_irq[2],user_irq[1],user_irq[0]
+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
*.iopin vdda1
*.iopin vdda2
*.iopin vssa1
*.iopin vssa2
*.iopin vccd1
*.iopin vccd2
*.iopin vssd1
*.iopin vssd2
*.ipin wb_clk_i
*.ipin wb_rst_i
*.ipin wbs_stb_i
*.ipin wbs_cyc_i
*.ipin wbs_we_i
*.ipin wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
*.ipin
*+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
*.ipin
*+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0]
*.opin wbs_ack_o
*.opin
*+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
*.ipin
*+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
*.opin
*+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
*.ipin
*+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
*.ipin
*+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0]
*.ipin user_clock2
*.opin
*+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
*.opin
*+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
*.iopin
*+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
*.iopin
*+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
*.iopin
*+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0]
*.iopin io_clamp_high[2],io_clamp_high[1],io_clamp_high[0]
*.iopin io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
*.opin user_irq[2],user_irq[1],user_irq[0]
*.ipin
*+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
x1 mod_clk io_analog[10] io_analog[9] mod_rst io_analog[8] io_analog[1] la_data_in[101]
+ la_data_in[100] la_data_in[99] la_data_in[63] la_data_in[62] la_data_in[65] la_data_in[64] io_out_7_buf[23]
+ io_analog[2] io_analog[0] io_analog[7] io_analog[3] io_out_26_buf[38] la_data_in[61] la_data_in[60] vccd1 vssd1
+ VDD VSS analog_top
x2 vccd1 vssd1 vssd1 io_out_7_buf[23] df_clk df_rst io_in_12_buf[0] io_in_11_buf[0] io_out[8]
+ io_out_13_buf[20] io_out[25] io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17]
+ io_out[16] io_out[15] io_out[14] digital_filter
x3[38] io_out_26_buf[38] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[37] sky130_fd_sc_hd__clkbuf_4
x3[37] io_out_26_buf[37] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[36] sky130_fd_sc_hd__clkbuf_4
x3[36] io_out_26_buf[36] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[35] sky130_fd_sc_hd__clkbuf_4
x3[35] io_out_26_buf[35] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[34] sky130_fd_sc_hd__clkbuf_4
x3[34] io_out_26_buf[34] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[33] sky130_fd_sc_hd__clkbuf_4
x3[33] io_out_26_buf[33] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[32] sky130_fd_sc_hd__clkbuf_4
x3[32] io_out_26_buf[32] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[31] sky130_fd_sc_hd__clkbuf_4
x3[31] io_out_26_buf[31] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[30] sky130_fd_sc_hd__clkbuf_4
x3[30] io_out_26_buf[30] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[29] sky130_fd_sc_hd__clkbuf_4
x3[29] io_out_26_buf[29] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[28] sky130_fd_sc_hd__clkbuf_4
x3[28] io_out_26_buf[28] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[27] sky130_fd_sc_hd__clkbuf_4
x3[27] io_out_26_buf[27] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[26] sky130_fd_sc_hd__clkbuf_4
x3[26] io_out_26_buf[26] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[25] sky130_fd_sc_hd__clkbuf_4
x3[25] io_out_26_buf[25] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[24] sky130_fd_sc_hd__clkbuf_4
x3[24] io_out_26_buf[24] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[23] sky130_fd_sc_hd__clkbuf_4
x3[23] io_out_26_buf[23] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[22] sky130_fd_sc_hd__clkbuf_4
x3[22] io_out_26_buf[22] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[21] sky130_fd_sc_hd__clkbuf_4
x3[21] io_out_26_buf[21] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[20] sky130_fd_sc_hd__clkbuf_4
x3[20] io_out_26_buf[20] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[19] sky130_fd_sc_hd__clkbuf_4
x3[19] io_out_26_buf[19] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[18] sky130_fd_sc_hd__clkbuf_4
x3[18] io_out_26_buf[18] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[17] sky130_fd_sc_hd__clkbuf_4
x3[17] io_out_26_buf[17] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[16] sky130_fd_sc_hd__clkbuf_4
x3[16] io_out_26_buf[16] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[15] sky130_fd_sc_hd__clkbuf_4
x3[15] io_out_26_buf[15] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[14] sky130_fd_sc_hd__clkbuf_4
x3[14] io_out_26_buf[14] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[13] sky130_fd_sc_hd__clkbuf_4
x3[13] io_out_26_buf[13] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[12] sky130_fd_sc_hd__clkbuf_4
x3[12] io_out_26_buf[12] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[11] sky130_fd_sc_hd__clkbuf_4
x3[11] io_out_26_buf[11] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[10] sky130_fd_sc_hd__clkbuf_4
x3[10] io_out_26_buf[10] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[9] sky130_fd_sc_hd__clkbuf_4
x3[9] io_out_26_buf[9] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[8] sky130_fd_sc_hd__clkbuf_4
x3[8] io_out_26_buf[8] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[7] sky130_fd_sc_hd__clkbuf_4
x3[7] io_out_26_buf[7] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[6] sky130_fd_sc_hd__clkbuf_4
x3[6] io_out_26_buf[6] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[5] sky130_fd_sc_hd__clkbuf_4
x3[5] io_out_26_buf[5] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[4] sky130_fd_sc_hd__clkbuf_4
x3[4] io_out_26_buf[4] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[3] sky130_fd_sc_hd__clkbuf_4
x3[3] io_out_26_buf[3] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[2] sky130_fd_sc_hd__clkbuf_4
x3[2] io_out_26_buf[2] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[1] sky130_fd_sc_hd__clkbuf_4
x3[1] io_out_26_buf[1] vssd1 vssd1 vccd1 vccd1 io_out_26_buf[0] sky130_fd_sc_hd__clkbuf_4
x3[0] io_out_26_buf[0] vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__clkbuf_4
x1[23] io_out_7_buf[23] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[22] sky130_fd_sc_hd__clkbuf_4
x1[22] io_out_7_buf[22] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[21] sky130_fd_sc_hd__clkbuf_4
x1[21] io_out_7_buf[21] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[20] sky130_fd_sc_hd__clkbuf_4
x1[20] io_out_7_buf[20] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[19] sky130_fd_sc_hd__clkbuf_4
x1[19] io_out_7_buf[19] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[18] sky130_fd_sc_hd__clkbuf_4
x1[18] io_out_7_buf[18] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[17] sky130_fd_sc_hd__clkbuf_4
x1[17] io_out_7_buf[17] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[16] sky130_fd_sc_hd__clkbuf_4
x1[16] io_out_7_buf[16] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[15] sky130_fd_sc_hd__clkbuf_4
x1[15] io_out_7_buf[15] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[14] sky130_fd_sc_hd__clkbuf_4
x1[14] io_out_7_buf[14] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[13] sky130_fd_sc_hd__clkbuf_4
x1[13] io_out_7_buf[13] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[12] sky130_fd_sc_hd__clkbuf_4
x1[12] io_out_7_buf[12] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[11] sky130_fd_sc_hd__clkbuf_4
x1[11] io_out_7_buf[11] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[10] sky130_fd_sc_hd__clkbuf_4
x1[10] io_out_7_buf[10] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[9] sky130_fd_sc_hd__clkbuf_4
x1[9] io_out_7_buf[9] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[8] sky130_fd_sc_hd__clkbuf_4
x1[8] io_out_7_buf[8] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[7] sky130_fd_sc_hd__clkbuf_4
x1[7] io_out_7_buf[7] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[6] sky130_fd_sc_hd__clkbuf_4
x1[6] io_out_7_buf[6] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[5] sky130_fd_sc_hd__clkbuf_4
x1[5] io_out_7_buf[5] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[4] sky130_fd_sc_hd__clkbuf_4
x1[4] io_out_7_buf[4] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[3] sky130_fd_sc_hd__clkbuf_4
x1[3] io_out_7_buf[3] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[2] sky130_fd_sc_hd__clkbuf_4
x1[2] io_out_7_buf[2] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[1] sky130_fd_sc_hd__clkbuf_4
x1[1] io_out_7_buf[1] vssd1 vssd1 vccd1 vccd1 io_out_7_buf[0] sky130_fd_sc_hd__clkbuf_4
x1[0] io_out_7_buf[0] vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__clkbuf_4
x1[14] io_in[10] vssd1 vssd1 vccd1 vccd1 clk_net[14] sky130_fd_sc_hd__clkbuf_4
x1[13] clk_net[14] vssd1 vssd1 vccd1 vccd1 clk_net[13] sky130_fd_sc_hd__clkbuf_4
x1[12] clk_net[13] vssd1 vssd1 vccd1 vccd1 clk_net[12] sky130_fd_sc_hd__clkbuf_4
x1[11] clk_net[12] vssd1 vssd1 vccd1 vccd1 clk_net[11] sky130_fd_sc_hd__clkbuf_4
x1[10] clk_net[11] vssd1 vssd1 vccd1 vccd1 clk_net[10] sky130_fd_sc_hd__clkbuf_4
x1[9] clk_net[10] vssd1 vssd1 vccd1 vccd1 clk_net[9] sky130_fd_sc_hd__clkbuf_4
x1[8] clk_net[9] vssd1 vssd1 vccd1 vccd1 clk_net[8] sky130_fd_sc_hd__clkbuf_4
x1[7] clk_net[8] vssd1 vssd1 vccd1 vccd1 clk_net[7] sky130_fd_sc_hd__clkbuf_4
x1[6] clk_net[7] vssd1 vssd1 vccd1 vccd1 clk_net[6] sky130_fd_sc_hd__clkbuf_4
x1[5] clk_net[6] vssd1 vssd1 vccd1 vccd1 clk_net[5] sky130_fd_sc_hd__clkbuf_4
x1[4] clk_net[5] vssd1 vssd1 vccd1 vccd1 clk_net[4] sky130_fd_sc_hd__clkbuf_4
x1[3] clk_net[4] vssd1 vssd1 vccd1 vccd1 clk_net[3] sky130_fd_sc_hd__clkbuf_4
x1[2] clk_net[3] vssd1 vssd1 vccd1 vccd1 clk_net[2] sky130_fd_sc_hd__clkbuf_4
x1[1] clk_net[2] vssd1 vssd1 vccd1 vccd1 clk_net[1] sky130_fd_sc_hd__clkbuf_4
x1[0] clk_net[1] vssd1 vssd1 vccd1 vccd1 clk_net[0] sky130_fd_sc_hd__clkbuf_4
x4 clk_net[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
x3 clk_net[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
x5 net1 vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
x6 net3 vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_4
x7 net4 vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_4
x8 net5 vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
x9 net6 vssd1 vssd1 vccd1 vccd1 df_clk sky130_fd_sc_hd__clkbuf_4
x10 net2 vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_4
x11 net7 vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
x12 net8 vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_4
x13 net9 vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_4
x14 net10 vssd1 vssd1 vccd1 vccd1 mod_clk sky130_fd_sc_hd__clkbuf_4
x2[14] io_in[9] vssd1 vssd1 vccd1 vccd1 rst_net[14] sky130_fd_sc_hd__clkbuf_4
x2[13] rst_net[14] vssd1 vssd1 vccd1 vccd1 rst_net[13] sky130_fd_sc_hd__clkbuf_4
x2[12] rst_net[13] vssd1 vssd1 vccd1 vccd1 rst_net[12] sky130_fd_sc_hd__clkbuf_4
x2[11] rst_net[12] vssd1 vssd1 vccd1 vccd1 rst_net[11] sky130_fd_sc_hd__clkbuf_4
x2[10] rst_net[11] vssd1 vssd1 vccd1 vccd1 rst_net[10] sky130_fd_sc_hd__clkbuf_4
x2[9] rst_net[10] vssd1 vssd1 vccd1 vccd1 rst_net[9] sky130_fd_sc_hd__clkbuf_4
x2[8] rst_net[9] vssd1 vssd1 vccd1 vccd1 rst_net[8] sky130_fd_sc_hd__clkbuf_4
x2[7] rst_net[8] vssd1 vssd1 vccd1 vccd1 rst_net[7] sky130_fd_sc_hd__clkbuf_4
x2[6] rst_net[7] vssd1 vssd1 vccd1 vccd1 rst_net[6] sky130_fd_sc_hd__clkbuf_4
x2[5] rst_net[6] vssd1 vssd1 vccd1 vccd1 rst_net[5] sky130_fd_sc_hd__clkbuf_4
x2[4] rst_net[5] vssd1 vssd1 vccd1 vccd1 rst_net[4] sky130_fd_sc_hd__clkbuf_4
x2[3] rst_net[4] vssd1 vssd1 vccd1 vccd1 rst_net[3] sky130_fd_sc_hd__clkbuf_4
x2[2] rst_net[3] vssd1 vssd1 vccd1 vccd1 rst_net[2] sky130_fd_sc_hd__clkbuf_4
x2[1] rst_net[2] vssd1 vssd1 vccd1 vccd1 rst_net[1] sky130_fd_sc_hd__clkbuf_4
x2[0] rst_net[1] vssd1 vssd1 vccd1 vccd1 rst_net[0] sky130_fd_sc_hd__clkbuf_4
x15 rst_net[0] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_4
x16 rst_net[0] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
x17 net11 vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_4
x18 net13 vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_4
x19 net14 vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_4
x20 net15 vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
x21 net16 vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_4
x22 net12 vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
x23 net18 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_4
x24 net19 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_4
x25 net20 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_4
x26 net21 vssd1 vssd1 vccd1 vccd1 mod_rst sky130_fd_sc_hd__clkbuf_4
x27 net17 vssd1 vssd1 vccd1 vccd1 df_rst sky130_fd_sc_hd__clkbuf_4
XC1 vccd1 vssd1 sky130_fd_pr__cap_mim_m3_1 W=29.99 L=29.99 MF=96 m=96
x2[20] io_out_13_buf[20] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[19] sky130_fd_sc_hd__clkbuf_4
x2[19] io_out_13_buf[19] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[18] sky130_fd_sc_hd__clkbuf_4
x2[18] io_out_13_buf[18] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[17] sky130_fd_sc_hd__clkbuf_4
x2[17] io_out_13_buf[17] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[16] sky130_fd_sc_hd__clkbuf_4
x2[16] io_out_13_buf[16] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[15] sky130_fd_sc_hd__clkbuf_4
x2[15] io_out_13_buf[15] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[14] sky130_fd_sc_hd__clkbuf_4
x2[14] io_out_13_buf[14] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[13] sky130_fd_sc_hd__clkbuf_4
x2[13] io_out_13_buf[13] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[12] sky130_fd_sc_hd__clkbuf_4
x2[12] io_out_13_buf[12] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[11] sky130_fd_sc_hd__clkbuf_4
x2[11] io_out_13_buf[11] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[10] sky130_fd_sc_hd__clkbuf_4
x2[10] io_out_13_buf[10] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[9] sky130_fd_sc_hd__clkbuf_4
x2[9] io_out_13_buf[9] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[8] sky130_fd_sc_hd__clkbuf_4
x2[8] io_out_13_buf[8] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[7] sky130_fd_sc_hd__clkbuf_4
x2[7] io_out_13_buf[7] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[6] sky130_fd_sc_hd__clkbuf_4
x2[6] io_out_13_buf[6] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[5] sky130_fd_sc_hd__clkbuf_4
x2[5] io_out_13_buf[5] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[4] sky130_fd_sc_hd__clkbuf_4
x2[4] io_out_13_buf[4] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[3] sky130_fd_sc_hd__clkbuf_4
x2[3] io_out_13_buf[3] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[2] sky130_fd_sc_hd__clkbuf_4
x2[2] io_out_13_buf[2] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[1] sky130_fd_sc_hd__clkbuf_4
x2[1] io_out_13_buf[1] vssd1 vssd1 vccd1 vccd1 io_out_13_buf[0] sky130_fd_sc_hd__clkbuf_4
x2[0] io_out_13_buf[0] vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__clkbuf_4
x1[20] io_in[12] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[20] sky130_fd_sc_hd__clkbuf_4
x1[19] io_in_12_buf[20] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[19] sky130_fd_sc_hd__clkbuf_4
x1[18] io_in_12_buf[19] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[18] sky130_fd_sc_hd__clkbuf_4
x1[17] io_in_12_buf[18] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[17] sky130_fd_sc_hd__clkbuf_4
x1[16] io_in_12_buf[17] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[16] sky130_fd_sc_hd__clkbuf_4
x1[15] io_in_12_buf[16] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[15] sky130_fd_sc_hd__clkbuf_4
x1[14] io_in_12_buf[15] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[14] sky130_fd_sc_hd__clkbuf_4
x1[13] io_in_12_buf[14] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[13] sky130_fd_sc_hd__clkbuf_4
x1[12] io_in_12_buf[13] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[12] sky130_fd_sc_hd__clkbuf_4
x1[11] io_in_12_buf[12] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[11] sky130_fd_sc_hd__clkbuf_4
x1[10] io_in_12_buf[11] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[10] sky130_fd_sc_hd__clkbuf_4
x1[9] io_in_12_buf[10] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[9] sky130_fd_sc_hd__clkbuf_4
x1[8] io_in_12_buf[9] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[8] sky130_fd_sc_hd__clkbuf_4
x1[7] io_in_12_buf[8] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[7] sky130_fd_sc_hd__clkbuf_4
x1[6] io_in_12_buf[7] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[6] sky130_fd_sc_hd__clkbuf_4
x1[5] io_in_12_buf[6] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[5] sky130_fd_sc_hd__clkbuf_4
x1[4] io_in_12_buf[5] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[4] sky130_fd_sc_hd__clkbuf_4
x1[3] io_in_12_buf[4] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[3] sky130_fd_sc_hd__clkbuf_4
x1[2] io_in_12_buf[3] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[2] sky130_fd_sc_hd__clkbuf_4
x1[1] io_in_12_buf[2] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[1] sky130_fd_sc_hd__clkbuf_4
x1[0] io_in_12_buf[1] vssd1 vssd1 vccd1 vccd1 io_in_12_buf[0] sky130_fd_sc_hd__clkbuf_4
x3[20] io_in[11] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[20] sky130_fd_sc_hd__clkbuf_4
x3[19] io_in_11_buf[20] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[19] sky130_fd_sc_hd__clkbuf_4
x3[18] io_in_11_buf[19] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[18] sky130_fd_sc_hd__clkbuf_4
x3[17] io_in_11_buf[18] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[17] sky130_fd_sc_hd__clkbuf_4
x3[16] io_in_11_buf[17] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[16] sky130_fd_sc_hd__clkbuf_4
x3[15] io_in_11_buf[16] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[15] sky130_fd_sc_hd__clkbuf_4
x3[14] io_in_11_buf[15] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[14] sky130_fd_sc_hd__clkbuf_4
x3[13] io_in_11_buf[14] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[13] sky130_fd_sc_hd__clkbuf_4
x3[12] io_in_11_buf[13] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[12] sky130_fd_sc_hd__clkbuf_4
x3[11] io_in_11_buf[12] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[11] sky130_fd_sc_hd__clkbuf_4
x3[10] io_in_11_buf[11] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[10] sky130_fd_sc_hd__clkbuf_4
x3[9] io_in_11_buf[10] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[9] sky130_fd_sc_hd__clkbuf_4
x3[8] io_in_11_buf[9] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[8] sky130_fd_sc_hd__clkbuf_4
x3[7] io_in_11_buf[8] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[7] sky130_fd_sc_hd__clkbuf_4
x3[6] io_in_11_buf[7] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[6] sky130_fd_sc_hd__clkbuf_4
x3[5] io_in_11_buf[6] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[5] sky130_fd_sc_hd__clkbuf_4
x3[4] io_in_11_buf[5] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[4] sky130_fd_sc_hd__clkbuf_4
x3[3] io_in_11_buf[4] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[3] sky130_fd_sc_hd__clkbuf_4
x3[2] io_in_11_buf[3] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[2] sky130_fd_sc_hd__clkbuf_4
x3[1] io_in_11_buf[2] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[1] sky130_fd_sc_hd__clkbuf_4
x3[0] io_in_11_buf[1] vssd1 vssd1 vccd1 vccd1 io_in_11_buf[0] sky130_fd_sc_hd__clkbuf_4
.ends

* expanding   symbol:  analog_top.sym # of pins=23
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/analog_top.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/analog_top.sch
.subckt analog_top  clk ip in rst_n i_bias_1 i_bias_2 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1 debug
+ d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 op a_probe_0 a_probe_1 a_probe_2 a_probe_3
+ d_probe d_probe_ctrl_0 d_probe_ctrl_1 VDD VSS
*.ipin ip
*.ipin in
*.ipin rst_n
*.ipin i_bias_1
*.ipin i_bias_2
*.ipin a_mod_grp_ctrl_0
*.ipin a_mod_grp_ctrl_1
*.ipin debug
*.opin op
*.opin a_probe_0
*.opin a_probe_1
*.opin a_probe_2
*.opin a_probe_3
*.ipin clk
*.opin d_probe
*.ipin d_clk_grp_1_ctrl_0
*.ipin d_clk_grp_1_ctrl_1
*.ipin d_clk_grp_2_ctrl_0
*.ipin d_clk_grp_2_ctrl_1
*.ipin d_probe_ctrl_0
*.ipin d_probe_ctrl_1
*.iopin VDD
*.iopin VSS
x1 ip in A A_b Ad Ad_b B B_b Bd Bd_b p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b rst_n rst_n_b i_bias_1
+ i_bias_2 op bias_a bias_b bias_c bias_d cm1 cmc op2 op1 on1 on2 VDD VSS modulator_w_test
x2 a_mod_grp_ctrl_1 a_mod_grp_ctrl_0 debug cm1 bias_b cmc net1 a_probe_2 VDD VSS a_mux4_en
x3 a_mod_grp_ctrl_1 a_mod_grp_ctrl_0 debug bias_a bias_c bias_d net2 a_probe_3 VDD VSS a_mux4_en
x4 a_mod_grp_ctrl_0 debug op1 on1 a_probe_0 VDD VSS a_mux2_en
x5 a_mod_grp_ctrl_0 debug op2 on2 a_probe_1 VDD VSS a_mux2_en
x8 a_probe_0 VDD VSS esd_cell
x9 a_probe_1 VDD VSS esd_cell
x10 a_probe_2 VDD VSS esd_cell
x11 a_probe_3 VDD VSS esd_cell
x12 i_bias_1 VDD VSS esd_cell
x13 i_bias_2 VDD VSS esd_cell
x14 ip VDD VSS esd_cell
x15 in VDD VSS esd_cell
x6 A A_b Ad Ad_b Bd_b Bd B_b B p2 p2_b p2d clk p2d_b p1d_b p1d p1_b p1 VDD VSS clock_v2
x16 p1 A p1_b A_b d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 VSS VSS VDD VDD net3 sky130_fd_sc_hd__mux4_1
x17 p2 B p2_b B_b d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 VSS VSS VDD VDD net4 sky130_fd_sc_hd__mux4_1
x18 p1d Ad p1d_b Ad_b d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VSS VDD VDD net5
+ sky130_fd_sc_hd__mux4_1
x19 p2d Bd p2d_b Bd_b d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VSS VDD VDD net6
+ sky130_fd_sc_hd__mux4_1
x20 net3 VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkinv_4
x21 net7 VSS VSS VDD VDD d_probe_0 sky130_fd_sc_hd__clkinv_16
x22 net4 VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkinv_4
x23 net8 VSS VSS VDD VDD d_probe_1 sky130_fd_sc_hd__clkinv_16
x24 net5 VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkinv_4
x25 net9 VSS VSS VDD VDD d_probe_2 sky130_fd_sc_hd__clkinv_16
x26 net6 VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkinv_4
x27 net10 VSS VSS VDD VDD d_probe_3 sky130_fd_sc_hd__clkinv_16
x7 rst_n VSS VSS VDD VDD rst_n_b sky130_fd_sc_hd__clkinv_16
x28 d_probe_3 d_probe_2 d_probe_1 d_probe_0 d_probe_ctrl_0 d_probe_ctrl_1 VSS VSS VDD VDD net11
+ sky130_fd_sc_hd__mux4_1
x29 net11 VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkinv_4
x30 net12 VSS VSS VDD VDD d_probe sky130_fd_sc_hd__clkinv_16
.ends


.subckt digital_filter  VDD VSS VSUBS data_in clk rst_n sclk cs_n new_data serial_data_out
+ data_out[11] data_out[10] data_out[9] data_out[8] data_out[7] data_out[6] data_out[5] data_out[4] data_out[3]
+ data_out[2] data_out[1] data_out[0]
Xsky130_fd_sc_hd__decap_6_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__ha_2_11 sky130_fd_sc_hd__ha_2_11/A sky130_fd_sc_hd__ha_2_11/B VSS
+ VDD sky130_fd_sc_hd__ha_2_10/B sky130_fd_sc_hd__ha_2_11/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkinv_1_7 sky130_fd_sc_hd__o21a_1_9/B1 VSS VDD sky130_fd_sc_hd__o21a_1_8/A1
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_97 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_54/X
+ VSS VDD sky130_fd_sc_hd__fa_2_0/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_64 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_5/X
+ VSS VDD sky130_fd_sc_hd__ha_2_3/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_86 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_27/X
+ VSS VDD sky130_fd_sc_hd__fa_2_0/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_42 sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__fa_2_7/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_42/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_20 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_17/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_20/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_53 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__ha_2_11/A
+ VSS VDD data_out[6] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_31 sky130_fd_sc_hd__clkinv_8_3/Y sclk VSS VDD sky130_fd_sc_hd__o21ai_1_0/A1
+ VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_75 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_16/X
+ VSS VDD sky130_fd_sc_hd__fa_2_11/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_36 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_47 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_58 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_4 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_1/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_4/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_9 sky130_fd_sc_hd__nor2_1_6/Y sky130_fd_sc_hd__fa_2_20/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_5/B VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__fa_2_20 sky130_fd_sc_hd__fa_2_20/A sky130_fd_sc_hd__fa_2_20/B sky130_fd_sc_hd__fa_2_20/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_19/CIN sky130_fd_sc_hd__fa_2_20/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_12_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__dfxtp_1_120 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_58/X
+ VSS VDD sky130_fd_sc_hd__fa_2_23/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_8_1 sky130_fd_sc_hd__clkinv_8_1/A VSS VDD sky130_fd_sc_hd__clkinv_8_4/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_6_36 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__ha_2_12 sky130_fd_sc_hd__ha_2_12/A sky130_fd_sc_hd__ha_2_12/B VSS
+ VDD sky130_fd_sc_hd__ha_2_11/B sky130_fd_sc_hd__ha_2_12/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__clkinv_1_8 sky130_fd_sc_hd__fa_2_23/B VSS VDD sky130_fd_sc_hd__nor2_1_7/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_98 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_53/X
+ VSS VDD sky130_fd_sc_hd__fa_2_2/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_65 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_6/X
+ VSS VDD sky130_fd_sc_hd__ha_2_2/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_87 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_28/X
+ VSS VDD sky130_fd_sc_hd__ha_2_14/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_43 sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__fa_2_6/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_43/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_10 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_7/X
+ VSS VDD sky130_fd_sc_hd__a22o_1_6/B1 VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_21 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_18/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_21/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_32 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__ha_2_15/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_32/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_76 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_17/X
+ VSS VDD sky130_fd_sc_hd__fa_2_10/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_54 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__ha_2_10/A
+ VSS VDD data_out[7] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_48 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_37 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_59 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_5 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_2/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_5/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22o_1_0 data_out[11] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_4/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_0/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__fa_2_21 sky130_fd_sc_hd__fa_2_21/A sky130_fd_sc_hd__fa_2_21/B sky130_fd_sc_hd__fa_2_21/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_20/CIN sky130_fd_sc_hd__fa_2_21/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_10 sky130_fd_sc_hd__fa_2_18/A sky130_fd_sc_hd__fa_2_10/B sky130_fd_sc_hd__fa_2_10/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_9/CIN sky130_fd_sc_hd__fa_2_10/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_121 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_57/X
+ VSS VDD sky130_fd_sc_hd__fa_2_24/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_110 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_41/X
+ VSS VDD sky130_fd_sc_hd__fa_2_22/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_8_2 sky130_fd_sc_hd__clkinv_8_4/A VSS VDD sky130_fd_sc_hd__clkinv_8_2/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_6_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__ha_2_13 sky130_fd_sc_hd__ha_2_13/A sky130_fd_sc_hd__ha_2_13/B VSS
+ VDD sky130_fd_sc_hd__ha_2_12/B sky130_fd_sc_hd__ha_2_13/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_6_37 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_9 sky130_fd_sc_hd__fa_2_21/B VSS VDD sky130_fd_sc_hd__nor2_1_6/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_11 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_8/X
+ VSS VDD sky130_fd_sc_hd__a22o_1_7/B1 VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_22 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_19/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_22/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_33 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__fa_2_16/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_33/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_99 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_52/X
+ VSS VDD sky130_fd_sc_hd__fa_2_3/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_44 sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__fa_2_5/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_44/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_66 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_7/X
+ VSS VDD sky130_fd_sc_hd__ha_2_1/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_88 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_29/X
+ VSS VDD sky130_fd_sc_hd__ha_2_13/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_77 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_18/X
+ VSS VDD sky130_fd_sc_hd__fa_2_9/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_55 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__ha_2_9/A
+ VSS VDD data_out[8] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_49 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_38 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_6 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_3/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_6/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_1_10 sky130_fd_sc_hd__fa_2_19/B VSS VDD sky130_fd_sc_hd__nor2_1_5/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__a22o_1_1 data_out[10] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_5/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_1/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__fa_2_11 sky130_fd_sc_hd__fa_2_19/A sky130_fd_sc_hd__fa_2_11/B sky130_fd_sc_hd__fa_2_11/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_10/CIN sky130_fd_sc_hd__fa_2_11/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_22 sky130_fd_sc_hd__fa_2_22/A sky130_fd_sc_hd__fa_2_22/B sky130_fd_sc_hd__fa_2_22/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_21/CIN sky130_fd_sc_hd__fa_2_22/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_100 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_51/X
+ VSS VDD sky130_fd_sc_hd__fa_2_4/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_111 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_40/X
+ VSS VDD sky130_fd_sc_hd__fa_2_23/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_122 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_56/X
+ VSS VDD sky130_fd_sc_hd__nor2_1_1/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_8_3 sky130_fd_sc_hd__clkinv_8_4/A VSS VDD sky130_fd_sc_hd__clkinv_8_3/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__ha_2_14 sky130_fd_sc_hd__ha_2_14/A sky130_fd_sc_hd__ha_2_14/B VSS
+ VDD sky130_fd_sc_hd__ha_2_13/B sky130_fd_sc_hd__ha_2_14/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_6_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__dfxtp_1_45 sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__fa_2_4/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_45/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_12 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_9/X
+ VSS VDD sky130_fd_sc_hd__a22o_1_8/B1 VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_67 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_8/X
+ VSS VDD sky130_fd_sc_hd__ha_2_0/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_34 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__fa_2_15/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_34/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_56 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__ha_2_8/A
+ VSS VDD data_out[9] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_23 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_20/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_23/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_89 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_30/X
+ VSS VDD sky130_fd_sc_hd__ha_2_12/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_78 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_19/X
+ VSS VDD sky130_fd_sc_hd__fa_2_8/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_39 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_7 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_4/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_7/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22o_1_2 data_out[9] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_6/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_2/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_60 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_23 sky130_fd_sc_hd__fa_2_23/A sky130_fd_sc_hd__fa_2_23/B sky130_fd_sc_hd__fa_2_23/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_22/CIN sky130_fd_sc_hd__fa_2_23/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_12 sky130_fd_sc_hd__fa_2_20/A sky130_fd_sc_hd__fa_2_12/B sky130_fd_sc_hd__fa_2_12/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_11/CIN sky130_fd_sc_hd__fa_2_12/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__dfxtp_1_101 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_50/X
+ VSS VDD sky130_fd_sc_hd__fa_2_5/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_112 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_39/X
+ VSS VDD sky130_fd_sc_hd__fa_2_24/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_8_4 sky130_fd_sc_hd__clkinv_8_4/A VSS VDD sky130_fd_sc_hd__clkinv_8_4/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_8
Xsky130_fd_sc_hd__decap_6_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__ha_2_15 sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__ha_2_15/B VSS
+ VDD sky130_fd_sc_hd__fa_2_16/CIN sky130_fd_sc_hd__ha_2_15/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__dfxtp_1_46 sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__fa_2_3/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_46/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_13 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_10/X
+ VSS VDD sky130_fd_sc_hd__a22o_1_9/B1 VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_68 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_9/X
+ VSS VDD sky130_fd_sc_hd__xor2_1_0/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_79 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_20/X
+ VSS VDD sky130_fd_sc_hd__fa_2_7/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_35 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__fa_2_14/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_35/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_24 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_21/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_24/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_57 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__ha_2_7/A
+ VSS VDD data_out[10] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_8 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_5/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_8/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__a22o_1_3 data_out[8] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_7/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_3/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_50 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_24 sky130_fd_sc_hd__fa_2_24/A sky130_fd_sc_hd__fa_2_24/B sky130_fd_sc_hd__nor2_1_0/A
+ VSS VDD sky130_fd_sc_hd__fa_2_23/CIN sky130_fd_sc_hd__fa_2_24/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__fa_2_13 sky130_fd_sc_hd__fa_2_21/A sky130_fd_sc_hd__fa_2_13/B sky130_fd_sc_hd__fa_2_13/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_12/CIN sky130_fd_sc_hd__fa_2_13/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_61 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_102 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_48/X
+ VSS VDD sky130_fd_sc_hd__fa_2_6/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_113 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_38/X
+ VSS VDD sky130_fd_sc_hd__ha_2_15/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_6_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__o21a_1_0 sky130_fd_sc_hd__nor2_1_2/Y sky130_fd_sc_hd__fa_2_1/A sky130_fd_sc_hd__xnor2_1_0/B
+ VSS VDD sky130_fd_sc_hd__o21a_1_0/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_47 sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__fa_2_2/B
+ VSS VDD data_out[0] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_14 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_11/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_14/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_69 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_10/X
+ VSS VDD sky130_fd_sc_hd__ha_2_15/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_36 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__fa_2_13/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_36/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_58 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__xor2_1_1/B
+ VSS VDD data_out[11] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_25 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_22/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_25/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_9 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_6/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_9/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_0 sky130_fd_sc_hd__fa_2_0/A sky130_fd_sc_hd__fa_2_0/B sky130_fd_sc_hd__fa_2_0/CIN
+ VSS VDD sky130_fd_sc_hd__ha_2_14/B sky130_fd_sc_hd__fa_2_0/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_4 data_out[7] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_8/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_4/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand4_1_0 sky130_fd_sc_hd__ha_2_6/B sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__ha_2_2/A
+ sky130_fd_sc_hd__ha_2_6/A VSS VDD sky130_fd_sc_hd__nor3_1_0/C VSUBS VDD sky130_fd_sc_hd__nand4_1
Xsky130_fd_sc_hd__decap_4_51 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_14 sky130_fd_sc_hd__fa_2_22/A sky130_fd_sc_hd__fa_2_14/B sky130_fd_sc_hd__fa_2_14/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_13/CIN sky130_fd_sc_hd__fa_2_14/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_62 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_40 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/A sky130_fd_sc_hd__nor2_1_1/Y
+ VSS VDD sky130_fd_sc_hd__nor2_1_0/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_103 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_49/X
+ VSS VDD sky130_fd_sc_hd__fa_2_7/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_114 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_63/X
+ VSS VDD sky130_fd_sc_hd__fa_2_18/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_6_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__o21a_1_1 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__fa_2_3/A sky130_fd_sc_hd__nor2_1_2/B
+ VSS VDD sky130_fd_sc_hd__o21a_1_1/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__xnor2_1_0 sky130_fd_sc_hd__fa_2_0/A sky130_fd_sc_hd__xnor2_1_0/B
+ VSS VDD sky130_fd_sc_hd__xnor2_1_0/Y VSUBS VDD sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_15 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_12/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_15/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_48 sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__fa_2_1/B
+ VSS VDD data_out[1] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_59 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_1/X
+ VSS VDD new_data VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_37 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__fa_2_12/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_37/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_26 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_23/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_26/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__clkinv_4_0/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__fa_2_1 sky130_fd_sc_hd__fa_2_1/A sky130_fd_sc_hd__fa_2_1/B sky130_fd_sc_hd__fa_2_1/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_0/CIN sky130_fd_sc_hd__fa_2_1/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_5 data_out[6] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_9/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_5/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_52 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_63 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_15 sky130_fd_sc_hd__fa_2_23/A sky130_fd_sc_hd__fa_2_15/B sky130_fd_sc_hd__fa_2_15/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_14/CIN sky130_fd_sc_hd__fa_2_15/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_41 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__nor2_1_1/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_1/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_104 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_47/X
+ VSS VDD sky130_fd_sc_hd__fa_2_8/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_115 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_64/X
+ VSS VDD sky130_fd_sc_hd__fa_2_17/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21a_1_2 sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__nor2_1_3/B
+ VSS VDD sky130_fd_sc_hd__o21a_1_2/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__xnor2_1_1 sky130_fd_sc_hd__fa_2_17/B sky130_fd_sc_hd__xnor2_1_1/B
+ VSS VDD sky130_fd_sc_hd__xnor2_1_1/Y VSUBS VDD sky130_fd_sc_hd__xnor2_1
Xsky130_fd_sc_hd__dfxtp_1_49 sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__fa_2_0/B
+ VSS VDD data_out[2] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_16 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_13/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_16/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_27 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_24/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_27/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_38 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__fa_2_11/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_38/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__fa_2_2 sky130_fd_sc_hd__fa_2_2/A sky130_fd_sc_hd__fa_2_2/B sky130_fd_sc_hd__fa_2_2/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_1/CIN sky130_fd_sc_hd__fa_2_2/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_6 data_out[5] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_6/B1
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_6/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_16 sky130_fd_sc_hd__fa_2_24/A sky130_fd_sc_hd__fa_2_16/B sky130_fd_sc_hd__fa_2_16/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_15/CIN sky130_fd_sc_hd__fa_2_16/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_53 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__nor2_1_2/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_2/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_105 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_46/X
+ VSS VDD sky130_fd_sc_hd__fa_2_9/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_116 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_62/X
+ VSS VDD sky130_fd_sc_hd__fa_2_19/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__o21a_1_3 sky130_fd_sc_hd__o21a_1_3/A1 sky130_fd_sc_hd__fa_2_7/A
+ sky130_fd_sc_hd__nor2_1_4/B VSS VDD sky130_fd_sc_hd__o21a_1_3/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_17 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_14/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_17/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_28 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_25/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_28/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_39 sky130_fd_sc_hd__dfxtp_1_55/CLK sky130_fd_sc_hd__fa_2_10/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_39/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_3 sky130_fd_sc_hd__fa_2_3/A sky130_fd_sc_hd__fa_2_3/B sky130_fd_sc_hd__fa_2_3/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_2/CIN sky130_fd_sc_hd__fa_2_3/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_7 data_out[4] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_7/B1
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_7/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_20 sky130_fd_sc_hd__dfxtp_1_38/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_24/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_20/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__nand2_1_10 sky130_fd_sc_hd__nor2_1_7/Y sky130_fd_sc_hd__fa_2_22/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_6/B VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_17 sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__fa_2_17/B sky130_fd_sc_hd__fa_2_17/CIN
+ VSS VDD sky130_fd_sc_hd__o21a_1_4/A1 sky130_fd_sc_hd__fa_2_17/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__nor2_1_3/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_3/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__sdlclkp_4_0 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__o21ai_1_0/Y
+ sky130_fd_sc_hd__conb_1_0/LO VSS VDD sky130_fd_sc_hd__dfxtp_1_9/CLK VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__dfxtp_1_117 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_61/X
+ VSS VDD sky130_fd_sc_hd__fa_2_20/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_106 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_45/X
+ VSS VDD sky130_fd_sc_hd__fa_2_18/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_4 sky130_fd_sc_hd__o21a_1_4/A1 sky130_fd_sc_hd__fa_2_8/A
+ sky130_fd_sc_hd__o21a_1_4/B1 VSS VDD sky130_fd_sc_hd__o21a_1_4/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_18 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__a22o_1_15/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_18/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_29 sky130_fd_sc_hd__dfxtp_1_7/CLK sky130_fd_sc_hd__a22o_1_26/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_29/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_4 sky130_fd_sc_hd__fa_2_4/A sky130_fd_sc_hd__fa_2_4/B sky130_fd_sc_hd__fa_2_4/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_3/CIN sky130_fd_sc_hd__fa_2_4/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_10 data_out[1] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_14/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_10/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_8 data_out[3] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_8/B1
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_8/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_21 sky130_fd_sc_hd__dfxtp_1_37/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_25/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_21/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__clkinv_2_0 clk VSS VDD sky130_fd_sc_hd__clkinv_8_0/A VSUBS VDD sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_18 sky130_fd_sc_hd__fa_2_18/A sky130_fd_sc_hd__fa_2_18/B sky130_fd_sc_hd__fa_2_18/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_17/CIN sky130_fd_sc_hd__fa_2_18/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__sdlclkp_4_1 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__o21ai_1_0/Y
+ sky130_fd_sc_hd__conb_1_0/LO VSS VDD sky130_fd_sc_hd__clkinv_4_0/A VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__nor2_1_4/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_4/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_118 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_60/X
+ VSS VDD sky130_fd_sc_hd__fa_2_21/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_107 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_44/X
+ VSS VDD sky130_fd_sc_hd__fa_2_19/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_5 sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__fa_2_18/B
+ sky130_fd_sc_hd__xnor2_1_1/B VSS VDD sky130_fd_sc_hd__o21a_1_5/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__dfxtp_1_19 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_16/X
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_19/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__fa_2_5 sky130_fd_sc_hd__fa_2_5/A sky130_fd_sc_hd__fa_2_5/B sky130_fd_sc_hd__fa_2_5/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_4/CIN sky130_fd_sc_hd__fa_2_5/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_11 data_out[0] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__dfxtp_1_15/Q
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_11/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_9 data_out[2] sky130_fd_sc_hd__a22o_1_9/A2 sky130_fd_sc_hd__a22o_1_9/B1
+ sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_9/X VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_22 sky130_fd_sc_hd__dfxtp_1_36/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_26/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_22/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_45 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__fa_2_19 sky130_fd_sc_hd__fa_2_19/A sky130_fd_sc_hd__fa_2_19/B sky130_fd_sc_hd__fa_2_19/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_18/CIN sky130_fd_sc_hd__fa_2_19/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__sdlclkp_4_2 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__o21ai_1_0/Y
+ sky130_fd_sc_hd__conb_1_0/LO VSS VDD sky130_fd_sc_hd__dfxtp_1_7/CLK VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__nor2_1_5/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_5/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_119 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_59/X
+ VSS VDD sky130_fd_sc_hd__fa_2_22/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_108 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_43/X
+ VSS VDD sky130_fd_sc_hd__fa_2_20/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_6 sky130_fd_sc_hd__nor2_1_6/Y sky130_fd_sc_hd__fa_2_20/B
+ sky130_fd_sc_hd__nor2_1_5/B VSS VDD sky130_fd_sc_hd__o21a_1_6/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__fa_2_6 sky130_fd_sc_hd__fa_2_6/A sky130_fd_sc_hd__fa_2_6/B sky130_fd_sc_hd__fa_2_6/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_5/CIN sky130_fd_sc_hd__fa_2_6/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_12 sky130_fd_sc_hd__dfxtp_1_46/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_16/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_12/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_23 sky130_fd_sc_hd__dfxtp_1_35/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_27/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_23/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_46 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__sdlclkp_4_3 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__and2_0_1/X
+ sky130_fd_sc_hd__conb_1_1/LO VSS VDD sky130_fd_sc_hd__dfxtp_1_55/CLK VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_6 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__nor2_1_6/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_6/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__dfxtp_1_109 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_42/X
+ VSS VDD sky130_fd_sc_hd__fa_2_21/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_7 sky130_fd_sc_hd__nor2_1_7/Y sky130_fd_sc_hd__fa_2_22/B
+ sky130_fd_sc_hd__nor2_1_6/B VSS VDD sky130_fd_sc_hd__o21a_1_7/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__fa_2_7 sky130_fd_sc_hd__fa_2_7/A sky130_fd_sc_hd__fa_2_7/B sky130_fd_sc_hd__fa_2_7/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_6/CIN sky130_fd_sc_hd__fa_2_7/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_13 sky130_fd_sc_hd__dfxtp_1_45/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_17/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_13/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__o21ai_1_0 sky130_fd_sc_hd__o21ai_1_0/A1 sky130_fd_sc_hd__nand2_1_0/Y
+ sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__o21ai_1_0/Y VSUBS VDD sky130_fd_sc_hd__o21ai_1
Xsky130_fd_sc_hd__a22o_1_24 sky130_fd_sc_hd__dfxtp_1_34/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_28/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_24/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__sdlclkp_4_4 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__and2_0_1/X
+ sky130_fd_sc_hd__conb_1_1/LO VSS VDD sky130_fd_sc_hd__dfxtp_1_45/CLK VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__nor2_1_7 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1_7/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_7/Y VSUBS VDD sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__decap_3_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_8 sky130_fd_sc_hd__o21a_1_8/A1 sky130_fd_sc_hd__fa_2_24/B
+ sky130_fd_sc_hd__nor2_1_7/B VSS VDD sky130_fd_sc_hd__o21a_1_8/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__fa_2_8 sky130_fd_sc_hd__fa_2_8/A sky130_fd_sc_hd__fa_2_8/B sky130_fd_sc_hd__fa_2_8/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_7/CIN sky130_fd_sc_hd__fa_2_8/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_14 sky130_fd_sc_hd__dfxtp_1_44/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_18/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_14/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_25 sky130_fd_sc_hd__dfxtp_1_33/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_29/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_25/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__sdlclkp_4_5 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__and2_0_1/X
+ sky130_fd_sc_hd__conb_1_1/LO VSS VDD sky130_fd_sc_hd__dfxtp_1_58/CLK VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__decap_3_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__o21a_1_9 data_in sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__o21a_1_9/B1
+ VSS VDD sky130_fd_sc_hd__o21a_1_9/X VSUBS VDD sky130_fd_sc_hd__o21a_1
Xsky130_fd_sc_hd__fa_2_9 sky130_fd_sc_hd__fa_2_9/A sky130_fd_sc_hd__fa_2_9/B sky130_fd_sc_hd__fa_2_9/CIN
+ VSS VDD sky130_fd_sc_hd__fa_2_8/CIN sky130_fd_sc_hd__fa_2_9/SUM VSUBS VDD sky130_fd_sc_hd__fa_2
Xsky130_fd_sc_hd__a22o_1_15 sky130_fd_sc_hd__dfxtp_1_43/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_19/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_15/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__a22o_1_26 sky130_fd_sc_hd__dfxtp_1_32/Q sky130_fd_sc_hd__a22o_1_9/A2
+ serial_data_out sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_26/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_38 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__sdlclkp_4_6 sky130_fd_sc_hd__clkinv_8_1/A sky130_fd_sc_hd__and2_0_1/X
+ sky130_fd_sc_hd__conb_1_1/LO VSS VDD sky130_fd_sc_hd__dfxtp_1_51/CLK VSUBS VDD sky130_fd_sc_hd__sdlclkp_4
Xsky130_fd_sc_hd__decap_3_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__a22o_1_16 sky130_fd_sc_hd__dfxtp_1_42/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_20/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_16/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__a22o_1_17 sky130_fd_sc_hd__dfxtp_1_41/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_21/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_17/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_8_60 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand3_1_0 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__ha_2_1/A
+ sky130_fd_sc_hd__ha_2_5/A VSS VDD sky130_fd_sc_hd__nor3_1_0/B VSUBS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__a22o_1_18 sky130_fd_sc_hd__dfxtp_1_40/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_22/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_18/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_8_50 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_61 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand3_1_1 sky130_fd_sc_hd__o21a_1_4/A1 sky130_fd_sc_hd__fa_2_8/A
+ sky130_fd_sc_hd__fa_2_7/A VSS VDD sky130_fd_sc_hd__nor2_1_4/B VSUBS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__a22o_1_19 sky130_fd_sc_hd__dfxtp_1_39/Q sky130_fd_sc_hd__a22o_1_9/A2
+ sky130_fd_sc_hd__dfxtp_1_23/Q sky130_fd_sc_hd__nand2_1_0/B VSS VDD sky130_fd_sc_hd__a22o_1_19/X
+ VSUBS VDD sky130_fd_sc_hd__a22o_1
Xsky130_fd_sc_hd__decap_8_40 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_51 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand3_1_2 data_in sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__fa_2_24/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_7/B VSUBS VDD sky130_fd_sc_hd__nand3_1
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__and2_0_60 sky130_fd_sc_hd__and2_0_60/A rst_n VSS VDD sky130_fd_sc_hd__and2_0_60/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_0 sky130_fd_sc_hd__ha_2_0/A sky130_fd_sc_hd__ha_2_0/B VSS VDD
+ sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__ha_2_0/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_41 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_52 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__and2_0_50 sky130_fd_sc_hd__o21a_1_2/X sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_50/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_61 sky130_fd_sc_hd__o21a_1_6/X rst_n VSS VDD sky130_fd_sc_hd__and2_0_61/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_1 sky130_fd_sc_hd__ha_2_1/A sky130_fd_sc_hd__ha_2_1/B VSS VDD
+ sky130_fd_sc_hd__ha_2_0/B sky130_fd_sc_hd__ha_2_1/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_53 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_42 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__and2_0_51 sky130_fd_sc_hd__and2_0_51/A sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_51/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_40 sky130_fd_sc_hd__fa_2_23/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_40/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_62 sky130_fd_sc_hd__and2_0_62/A rst_n VSS VDD sky130_fd_sc_hd__and2_0_62/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_2 sky130_fd_sc_hd__ha_2_2/A sky130_fd_sc_hd__ha_2_2/B VSS VDD
+ sky130_fd_sc_hd__ha_2_1/B sky130_fd_sc_hd__ha_2_2/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_54 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_43 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_0 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nor2_1_2/Y VSS VDD sky130_fd_sc_hd__and2_0_53/A VSUBS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_52 sky130_fd_sc_hd__o21a_1_1/X sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_52/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_63 sky130_fd_sc_hd__o21a_1_5/X rst_n VSS VDD sky130_fd_sc_hd__and2_0_63/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_41 sky130_fd_sc_hd__fa_2_22/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_41/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_30 sky130_fd_sc_hd__ha_2_12/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_30/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_3 sky130_fd_sc_hd__ha_2_3/A sky130_fd_sc_hd__ha_2_3/B VSS VDD
+ sky130_fd_sc_hd__ha_2_2/B sky130_fd_sc_hd__ha_2_3/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_44 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_55 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_1 sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nor2_1_3/Y VSS VDD sky130_fd_sc_hd__and2_0_51/A VSUBS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_20 sky130_fd_sc_hd__fa_2_7/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_20/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_31 sky130_fd_sc_hd__ha_2_11/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_31/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_53 sky130_fd_sc_hd__and2_0_53/A sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_53/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_64 sky130_fd_sc_hd__xnor2_1_1/Y rst_n VSS VDD sky130_fd_sc_hd__and2_0_64/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_42 sky130_fd_sc_hd__fa_2_21/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_42/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_4 sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__ha_2_4/B VSS VDD
+ sky130_fd_sc_hd__ha_2_3/B sky130_fd_sc_hd__ha_2_4/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_45 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_56 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_2 sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__nor2_1_4/B
+ sky130_fd_sc_hd__nor2_1_4/Y VSS VDD sky130_fd_sc_hd__and2_0_48/A VSUBS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_54 sky130_fd_sc_hd__xnor2_1_0/Y sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_54/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_21 sky130_fd_sc_hd__fa_2_6/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_21/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_10 sky130_fd_sc_hd__ha_2_15/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_10/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_32 sky130_fd_sc_hd__ha_2_10/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_32/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_43 sky130_fd_sc_hd__fa_2_20/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_43/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__ha_2_5 sky130_fd_sc_hd__ha_2_5/A sky130_fd_sc_hd__ha_2_5/B VSS VDD
+ sky130_fd_sc_hd__ha_2_4/B sky130_fd_sc_hd__ha_2_5/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_8_57 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_46 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_3 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__nor2_1_5/B
+ sky130_fd_sc_hd__nor2_1_5/Y VSS VDD sky130_fd_sc_hd__and2_0_62/A VSUBS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_55 sky130_fd_sc_hd__o21a_1_0/X sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_55/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_22 sky130_fd_sc_hd__fa_2_5/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_22/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_11 sky130_fd_sc_hd__fa_2_16/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_11/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_33 sky130_fd_sc_hd__ha_2_9/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_33/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_44 sky130_fd_sc_hd__fa_2_19/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_44/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__ha_2_6 sky130_fd_sc_hd__ha_2_6/A sky130_fd_sc_hd__ha_2_6/B VSS VDD
+ sky130_fd_sc_hd__ha_2_5/B sky130_fd_sc_hd__ha_2_6/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__conb_1_0 VSS VSUBS VDD VDD sky130_fd_sc_hd__conb_1_0/HI sky130_fd_sc_hd__conb_1_0/LO
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_58 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_47 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_36 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_4 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__nor2_1_6/B
+ sky130_fd_sc_hd__nor2_1_6/Y VSS VDD sky130_fd_sc_hd__and2_0_60/A VSUBS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_23 sky130_fd_sc_hd__fa_2_4/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_23/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_56 sky130_fd_sc_hd__o21a_1_9/X rst_n VSS VDD sky130_fd_sc_hd__and2_0_56/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_34 sky130_fd_sc_hd__ha_2_8/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_34/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_12 sky130_fd_sc_hd__fa_2_15/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_12/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_45 sky130_fd_sc_hd__fa_2_18/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_45/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__ha_2_7 sky130_fd_sc_hd__ha_2_7/A sky130_fd_sc_hd__ha_2_7/B VSS VDD
+ sky130_fd_sc_hd__xor2_1_1/A sky130_fd_sc_hd__ha_2_7/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__conb_1_1 VSS VSUBS VDD VDD sky130_fd_sc_hd__conb_1_1/HI sky130_fd_sc_hd__conb_1_1/LO
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_48 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_59 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_37 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__and2_0_0 sky130_fd_sc_hd__and2_0_0/A sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_0/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_8_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__a21oi_1_5 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1_7/B
+ sky130_fd_sc_hd__nor2_1_7/Y VSS VDD sky130_fd_sc_hd__and2_0_58/A VSUBS VDD sky130_fd_sc_hd__a21oi_1
Xsky130_fd_sc_hd__decap_6_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_13 sky130_fd_sc_hd__fa_2_14/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_13/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_24 sky130_fd_sc_hd__fa_2_3/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_24/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_46 sky130_fd_sc_hd__fa_2_17/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_46/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_35 sky130_fd_sc_hd__ha_2_7/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_35/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_57 sky130_fd_sc_hd__o21a_1_8/X rst_n VSS VDD sky130_fd_sc_hd__and2_0_57/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__ha_2_8 sky130_fd_sc_hd__ha_2_8/A sky130_fd_sc_hd__ha_2_8/B VSS VDD
+ sky130_fd_sc_hd__ha_2_7/B sky130_fd_sc_hd__ha_2_8/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_3_60 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_8_38 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_49 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_1_0/Y VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_1 sky130_fd_sc_hd__nor3_1_0/Y sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_1/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_8_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_6_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_25 sky130_fd_sc_hd__fa_2_2/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_25/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_36 sky130_fd_sc_hd__xor2_1_1/X sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_36/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_14 sky130_fd_sc_hd__fa_2_13/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_14/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_47 sky130_fd_sc_hd__o21a_1_4/X sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_47/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_58 sky130_fd_sc_hd__and2_0_58/A rst_n VSS VDD sky130_fd_sc_hd__and2_0_58/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__ha_2_9 sky130_fd_sc_hd__ha_2_9/A sky130_fd_sc_hd__ha_2_9/B VSS VDD
+ sky130_fd_sc_hd__ha_2_8/B sky130_fd_sc_hd__ha_2_9/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_3_61 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_50 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_8_39 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_1 cs_n new_data VSS VDD sky130_fd_sc_hd__nand2_1_1/Y VSUBS
+ VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_2 sky130_fd_sc_hd__ha_2_6/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_2/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__and2_0_48 sky130_fd_sc_hd__and2_0_48/A sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_48/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_26 sky130_fd_sc_hd__fa_2_1/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_26/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_37 sky130_fd_sc_hd__ha_2_15/A sky130_fd_sc_hd__nor2_1_1/B
+ VSS VDD sky130_fd_sc_hd__nor2_1_0/A VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_59 sky130_fd_sc_hd__o21a_1_7/X rst_n VSS VDD sky130_fd_sc_hd__and2_0_59/X
+ VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__nand2_1_1/Y VSS VDD sky130_fd_sc_hd__a22o_1_9/A2
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_15 sky130_fd_sc_hd__fa_2_12/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_15/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_90 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_31/X
+ VSS VDD sky130_fd_sc_hd__ha_2_11/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_40 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_51 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_62 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_8_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__ha_2_4/A sky130_fd_sc_hd__ha_2_0/A VSS
+ VDD sky130_fd_sc_hd__nor3_1_0/A VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_3 sky130_fd_sc_hd__ha_2_5/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_3/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_1 cs_n VSS VDD sky130_fd_sc_hd__nand2_1_0/B VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_27 sky130_fd_sc_hd__fa_2_0/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_27/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_49 sky130_fd_sc_hd__o21a_1_3/X sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_49/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_38 sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_38/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_16 sky130_fd_sc_hd__fa_2_11/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_16/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_91 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_32/X
+ VSS VDD sky130_fd_sc_hd__ha_2_10/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_80 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_21/X
+ VSS VDD sky130_fd_sc_hd__fa_2_6/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_52 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_63 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_41 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_8_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__o21a_1_4/A1 sky130_fd_sc_hd__fa_2_8/A
+ VSS VDD sky130_fd_sc_hd__o21a_1_4/B1 VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_4 sky130_fd_sc_hd__ha_2_4/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_4/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__nor3_1_0 sky130_fd_sc_hd__nor3_1_0/A sky130_fd_sc_hd__nor3_1_0/B
+ sky130_fd_sc_hd__nor3_1_0/C VSS VDD sky130_fd_sc_hd__nor3_1_0/Y VSUBS VDD sky130_fd_sc_hd__nor3_1
Xsky130_fd_sc_hd__decap_6_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__ha_2_6/B VSS VDD sky130_fd_sc_hd__and2_0_0/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_28 sky130_fd_sc_hd__ha_2_14/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_28/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_17 sky130_fd_sc_hd__fa_2_10/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_17/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_39 sky130_fd_sc_hd__fa_2_24/SUM sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_39/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_81 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_22/X
+ VSS VDD sky130_fd_sc_hd__fa_2_5/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_92 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_33/X
+ VSS VDD sky130_fd_sc_hd__ha_2_9/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_70 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_11/X
+ VSS VDD sky130_fd_sc_hd__fa_2_16/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_64 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_42 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_53 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__nor2_1_2/Y sky130_fd_sc_hd__fa_2_1/A
+ VSS VDD sky130_fd_sc_hd__xnor2_1_0/B VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_5 sky130_fd_sc_hd__ha_2_3/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_5/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__fa_2_6/A VSS VDD sky130_fd_sc_hd__nor2_1_4/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_18 sky130_fd_sc_hd__fa_2_9/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_18/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__and2_0_29 sky130_fd_sc_hd__ha_2_13/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_29/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_82 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_23/X
+ VSS VDD sky130_fd_sc_hd__fa_2_4/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_60 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_0/X
+ VSS VDD sky130_fd_sc_hd__ha_2_6/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_71 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_12/X
+ VSS VDD sky130_fd_sc_hd__fa_2_15/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_93 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_34/X
+ VSS VDD sky130_fd_sc_hd__ha_2_8/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_43 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_65 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_54 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_0 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_9/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_5 sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__fa_2_3/A
+ VSS VDD sky130_fd_sc_hd__nor2_1_2/B VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_6 sky130_fd_sc_hd__ha_2_2/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_6/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_6_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__o21a_1_4/B1 VSS VDD sky130_fd_sc_hd__o21a_1_3/A1
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__and2_0_19 sky130_fd_sc_hd__fa_2_8/SUM sky130_fd_sc_hd__dfxtp_1_1/Q
+ VSS VDD sky130_fd_sc_hd__and2_0_19/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_83 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_24/X
+ VSS VDD sky130_fd_sc_hd__fa_2_3/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_61 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_2/X
+ VSS VDD sky130_fd_sc_hd__ha_2_6/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_50 sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__ha_2_14/A
+ VSS VDD data_out[3] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_72 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_13/X
+ VSS VDD sky130_fd_sc_hd__fa_2_14/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_94 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_35/X
+ VSS VDD sky130_fd_sc_hd__ha_2_7/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_44 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_55 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_1 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_1/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_6 sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__fa_2_5/A
+ VSS VDD sky130_fd_sc_hd__nor2_1_3/B VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_7 sky130_fd_sc_hd__ha_2_1/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_7/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/B
+ VSS VDD sky130_fd_sc_hd__xor2_1_0/X VSUBS VDD sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__fa_2_4/A VSS VDD sky130_fd_sc_hd__nor2_1_3/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfxtp_1_51 sky130_fd_sc_hd__dfxtp_1_51/CLK sky130_fd_sc_hd__ha_2_13/A
+ VSS VDD data_out[4] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_40 sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__fa_2_9/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_40/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_84 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_25/X
+ VSS VDD sky130_fd_sc_hd__fa_2_2/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_62 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_3/X
+ VSS VDD sky130_fd_sc_hd__ha_2_5/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_95 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_36/X
+ VSS VDD sky130_fd_sc_hd__xor2_1_1/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_73 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_14/X
+ VSS VDD sky130_fd_sc_hd__fa_2_13/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_45 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_56 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_2 sky130_fd_sc_hd__clkinv_8_3/Y rst_n VSS VDD sky130_fd_sc_hd__dfxtp_1_2/Q
+ VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_7 data_in sky130_fd_sc_hd__nor2_1_1/B VSS VDD sky130_fd_sc_hd__o21a_1_9/B1
+ VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_8 sky130_fd_sc_hd__ha_2_0/SUM sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_8/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__xor2_1_1 sky130_fd_sc_hd__xor2_1_1/A sky130_fd_sc_hd__xor2_1_1/B
+ VSS VDD sky130_fd_sc_hd__xor2_1_1/X VSUBS VDD sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__ha_2_10 sky130_fd_sc_hd__ha_2_10/A sky130_fd_sc_hd__ha_2_10/B VSS
+ VDD sky130_fd_sc_hd__ha_2_9/B sky130_fd_sc_hd__ha_2_10/SUM VSUBS VDD sky130_fd_sc_hd__ha_2
Xsky130_fd_sc_hd__decap_6_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkinv_1_6 sky130_fd_sc_hd__fa_2_2/A VSS VDD sky130_fd_sc_hd__nor2_1_2/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__dfxtp_1_85 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_26/X
+ VSS VDD sky130_fd_sc_hd__fa_2_1/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_63 sky130_fd_sc_hd__clkinv_8_2/Y sky130_fd_sc_hd__and2_0_4/X
+ VSS VDD sky130_fd_sc_hd__ha_2_4/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_41 sky130_fd_sc_hd__dfxtp_1_45/CLK sky130_fd_sc_hd__fa_2_8/B
+ VSS VDD sky130_fd_sc_hd__dfxtp_1_41/Q VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_52 sky130_fd_sc_hd__dfxtp_1_58/CLK sky130_fd_sc_hd__ha_2_12/A
+ VSS VDD data_out[5] VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_30 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__o21ai_1_0/A1
+ VSS VDD sky130_fd_sc_hd__nand2_1_0/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_74 sky130_fd_sc_hd__clkinv_8_3/Y sky130_fd_sc_hd__and2_0_15/X
+ VSS VDD sky130_fd_sc_hd__fa_2_12/B VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__dfxtp_1_96 sky130_fd_sc_hd__clkinv_8_4/Y sky130_fd_sc_hd__and2_0_55/X
+ VSS VDD sky130_fd_sc_hd__fa_2_1/A VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__decap_3_57 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_46 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfxtp_1_3 sky130_fd_sc_hd__dfxtp_1_9/CLK sky130_fd_sc_hd__a22o_1_0/X
+ VSS VDD serial_data_out VSUBS VDD sky130_fd_sc_hd__dfxtp_1
Xsky130_fd_sc_hd__nand2_1_8 sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__fa_2_18/B
+ VSS VDD sky130_fd_sc_hd__xnor2_1_1/B VSUBS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__and2_0_9 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_0_9/B
+ VSS VDD sky130_fd_sc_hd__and2_0_9/X VSUBS VDD sky130_fd_sc_hd__and2_0
Xsky130_fd_sc_hd__clkinv_8_0 sky130_fd_sc_hd__clkinv_8_0/A VSS VDD sky130_fd_sc_hd__clkinv_8_1/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_8
.ends


* expanding   symbol:  modulator_w_test.sym # of pins=33
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/modulator_w_test.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/modulator_w_test.sch
.subckt modulator_w_test  ip in A A_b Ad Ad_b B B_b Bd Bd_b p1 p1_b p1d p1d_b p2 p2_b p2d p2d_b
+ rst_n rst_n_b i_bias_1 i_bias_2 op bias_a bias_b bias_c bias_d cm1 cmc op2 op1 on1 on2  VDD  VSS
*.ipin ip
*.ipin in
*.ipin A
*.ipin A_b
*.ipin Ad
*.ipin Ad_b
*.ipin B
*.ipin B_b
*.ipin Bd
*.ipin Bd_b
*.ipin p1
*.ipin p1_b
*.ipin p1d
*.ipin p1d_b
*.ipin p2
*.ipin p2_b
*.ipin p2d
*.ipin p2d_b
*.ipin rst_n
*.ipin rst_n_b
*.ipin i_bias_1
*.ipin i_bias_2
*.opin op
*.opin bias_a
*.opin bias_b
*.opin bias_c
*.opin bias_d
*.opin cm1
*.opin cmc
*.opin op1
*.opin on1
*.opin op2
*.opin on2
x4 c1r in1 p2 p2_b VDD VSS transmission_gate
x5 net1 ip1 p2 p2_b VDD VSS transmission_gate
x2 c1r cm1 p1 p1_b VDD VSS transmission_gate
x3 net1 cm1 p1 p1_b VDD VSS transmission_gate
x10 ip c1l p1d p1d_b VDD VSS transmission_gate
x11 dac_n net2 p2d p2d_b VDD VSS transmission_gate
x12 VDD VSS op dac_p on VDD VSS 1b_dac
x13 dac_p c1l p2d p2d_b VDD VSS transmission_gate
x14 in net2 p1d p1d_b VDD VSS transmission_gate
x19 on1 op1 rst_n_b rst_n VDD VSS transmission_gate
x20 cm1 in1 rst_n_b rst_n VDD VSS transmission_gate
x21 cm1 ip1 rst_n_b rst_n VDD VSS transmission_gate
x22 op1 c3l p1d p1d_b VDD VSS transmission_gate
x23 on1 net3 p1d p1d_b VDD VSS transmission_gate
x24 net3 c3l p2d p2d_b VDD VSS transmission_gate
x25 c3r cm2 p1 p1_b VDD VSS transmission_gate
x26 net4 cm2 p1 p1_b VDD VSS transmission_gate
x27 ip c4l p1d p1d_b VDD VSS transmission_gate
x28 dac_p c4l p2d p2d_b VDD VSS transmission_gate
x29 c3r in2 p2 p2_b VDD VSS transmission_gate
x30 net4 ip2 p2 p2_b VDD VSS transmission_gate
x32 cm2 in2 rst_n_b rst_n VDD VSS transmission_gate
x33 cm2 ip2 rst_n_b rst_n VDD VSS transmission_gate
x34 on2 op2 rst_n_b rst_n VDD VSS transmission_gate
x36 VSS VDD op dac_n on VDD VSS 1b_dac
x37 in net5 p1d p1d_b VDD VSS transmission_gate
x38 dac_n net5 p2d p2d_b VDD VSS transmission_gate
XC11 c1l c1r sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=2 m=2
XC1 net2 net1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=2 m=2
XC2 op1 in1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=10 m=10
XC3 on1 ip1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=10 m=10
XC4 c3r c4l sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=1 m=1
XC5 c3r c3l sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=2 m=2
XC6 net4 net3 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=2 m=2
XC7 net4 net5 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=1 m=1
XC8 op2 in2 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=14 m=14
XC9 on2 ip2 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=14 m=14
XC10 op2 VSS sky130_fd_pr__cap_mim_m3_1 W=11.6 L=11.6 MF=1 m=1
XC12 on2 VSS sky130_fd_pr__cap_mim_m3_1 W=11.6 L=11.6 MF=1 m=1
x6 in1 in1_c A A_b VDD VSS transmission_gate
x8 ip1 in1_c B B_b VDD VSS transmission_gate
x15 op1_c op1 Ad Ad_b VDD VSS transmission_gate
x16 on1_c on1 Ad Ad_b VDD VSS transmission_gate
x17 op1_c on1 Bd Bd_b VDD VSS transmission_gate
x18 on1_c op1 Bd Bd_b VDD VSS transmission_gate
x7 ip1 ip1_c A A_b VDD VSS transmission_gate
x9 in1 ip1_c B B_b VDD VSS transmission_gate
XC13 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 sky130_fd_pr__cap_mim_m3_1 W=8.8 L=8.8 MF=24 m=24
XC14 __UNCONNECTED_PIN__2 __UNCONNECTED_PIN__3 sky130_fd_pr__cap_mim_m3_1 W=2.1 L=2.1 MF=38 m=38
x35 op2 on2 op p1_b on VDD VSS comparator
XM2 VSS on VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
XM3 VDD on VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=3 m=3 
x1 i_bias_1 ip1_c in1_c p1 p1_b p2 p2_b op1_c on1_c cm1 bias_a bias_b bias_c bias_d cmc VDD VSS
+ ota_w_test
x31 i_bias_2 ip2 in2 p1 p1_b p2 p2_b op2 on2 cm2 VDD VSS ota
.ends


* expanding   symbol:  a_mux4_en.sym # of pins=8
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux4_en.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux4_en.sch
.subckt a_mux4_en  s0 s1 en in0 in1 in2 in3 out  VDD  VSS
*.ipin en
*.ipin s1
*.ipin s0
*.ipin in0
*.ipin in1
*.ipin in2
*.ipin in3
*.opin out
x1 net4 out net5 en3_b VDD VSS switch_5t
x2 net3 out net6 en2_b VDD VSS switch_5t
x3 net2 out net7 en1_b VDD VSS switch_5t
x4 net1 out net8 en0_b VDD VSS switch_5t
x5 en3_b VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x6 en2_b VSS VSS VDD VDD net6 sky130_fd_sc_hd__inv_1
x7 en1_b VSS VSS VDD VDD net7 sky130_fd_sc_hd__inv_1
x8 en0_b VSS VSS VDD VDD net8 sky130_fd_sc_hd__inv_1
x13 s0 VSS VSS VDD VDD s0_b sky130_fd_sc_hd__inv_1
x14 s1 VSS VSS VDD VDD s1_b sky130_fd_sc_hd__inv_1
x9 s1_b s0_b VSS VSS VDD VDD en0_b sky130_fd_sc_hd__nand2_1
x10 s1 s0_b VSS VSS VDD VDD en1_b sky130_fd_sc_hd__nand2_1
x11 s0 s1_b VSS VSS VDD VDD en2_b sky130_fd_sc_hd__nand2_1
x12 s0 s1 VSS VSS VDD VDD en3_b sky130_fd_sc_hd__nand2_1
x15 in0 net1 en en_b VDD VSS transmission_gate
x16 in1 net2 en en_b VDD VSS transmission_gate
x17 in2 net3 en en_b VDD VSS transmission_gate
x18 in3 net4 en en_b VDD VSS transmission_gate
x19 en VSS VSS VDD VDD en_b sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  a_mux2_en.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux2_en.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/a_mux2_en.sch
.subckt a_mux2_en  s0 en in0 in1 out  VDD  VSS
*.ipin en
*.ipin s0
*.ipin in0
*.ipin in1
*.opin out
x3 net2 out s0 s0_b VDD VSS switch_5t
x4 net1 out s0_b s0 VDD VSS switch_5t
x15 in0 net1 en en_b VDD VSS transmission_gate
x16 in1 net2 en en_b VDD VSS transmission_gate
x19 en VSS VSS VDD VDD en_b sky130_fd_sc_hd__inv_1
x1 s0 VSS VSS VDD VDD s0_b sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  esd_cell.sym # of pins=1
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/esd_cell.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/esd_cell.sch
.subckt esd_cell  esd  VDD  VSS
*.iopin esd
XM1 esd VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM2 esd VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
.ends


* expanding   symbol:  clock_v2.sym # of pins=17
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/clock_v2.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/clock_v2.sch
.subckt clock_v2  A A_b Ad Ad_b Bd_b Bd B_b B p2 p2_b p2d clk p2d_b p1d_b p1d p1_b p1  VDD  VSS
*.ipin clk
*.opin p2d_b
*.opin p2d
*.opin p2_b
*.opin p2
*.opin p1d_b
*.opin p1d
*.opin p1_b
*.opin p1
*.opin Ad_b
*.opin Ad
*.opin A_b
*.opin A
*.opin Bd_b
*.opin Bd
*.opin B_b
*.opin B
x2 latch_out clk VSS VSS VDD VDD net1 sky130_fd_sc_hd__nand2_1
x3 net3 net6 VSS VSS VDD VDD net4 sky130_fd_sc_hd__nand2_1
x4 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__clkinv_4
x6 net2 VSS VSS VDD VDD net34 sky130_fd_sc_hd__clkinv_1
x9 net4 VSS VSS VDD VDD net5 sky130_fd_sc_hd__clkinv_4
x11 net5 VSS VSS VDD VDD net35 sky130_fd_sc_hd__clkinv_1
x1 clk VSS VSS VDD VDD net3 sky130_fd_sc_hd__clkinv_1
x20 net36 VSS VSS VDD VDD latch_in sky130_fd_sc_hd__clkdlybuf4s50_1
x21 net37 VSS VSS VDD VDD net6 sky130_fd_sc_hd__clkdlybuf4s50_1
x22 net34 VSS VSS VDD VDD net38 sky130_fd_sc_hd__clkdlybuf4s50_1
x25 net35 VSS VSS VDD VDD net39 sky130_fd_sc_hd__clkdlybuf4s50_1
x7 net40 VSS VSS VDD VDD net36 sky130_fd_sc_hd__clkdlybuf4s50_1
x12 net41 VSS VSS VDD VDD net37 sky130_fd_sc_hd__clkdlybuf4s50_1
x14 net38 VSS VSS VDD VDD net42 sky130_fd_sc_hd__clkdlybuf4s50_1
x15 net39 VSS VSS VDD VDD net43 sky130_fd_sc_hd__clkdlybuf4s50_1
x16 net44 VSS VSS VDD VDD net40 sky130_fd_sc_hd__clkdlybuf4s50_1
x17 net45 VSS VSS VDD VDD net41 sky130_fd_sc_hd__clkdlybuf4s50_1
x18 net42 VSS VSS VDD VDD net46 sky130_fd_sc_hd__clkdlybuf4s50_1
x19 net43 VSS VSS VDD VDD net47 sky130_fd_sc_hd__clkdlybuf4s50_1
x23 net48 VSS VSS VDD VDD net44 sky130_fd_sc_hd__clkdlybuf4s50_1
x24 net49 VSS VSS VDD VDD net45 sky130_fd_sc_hd__clkdlybuf4s50_1
x26 net46 VSS VSS VDD VDD net7 sky130_fd_sc_hd__clkdlybuf4s50_1
x27 net47 VSS VSS VDD VDD net8 sky130_fd_sc_hd__clkdlybuf4s50_1
x28 net50 VSS VSS VDD VDD net48 sky130_fd_sc_hd__clkdlybuf4s50_1
x29 net51 VSS VSS VDD VDD net49 sky130_fd_sc_hd__clkdlybuf4s50_1
x32 net52 VSS VSS VDD VDD net50 sky130_fd_sc_hd__clkdlybuf4s50_1
x33 net53 VSS VSS VDD VDD net51 sky130_fd_sc_hd__clkdlybuf4s50_1
x36 net54 VSS VSS VDD VDD net52 sky130_fd_sc_hd__clkdlybuf4s50_1
x37 net55 VSS VSS VDD VDD net53 sky130_fd_sc_hd__clkdlybuf4s50_1
x40 net56 VSS VSS VDD VDD net54 sky130_fd_sc_hd__clkdlybuf4s50_1
x41 net57 VSS VSS VDD VDD net55 sky130_fd_sc_hd__clkdlybuf4s50_1
x44 net58 VSS VSS VDD VDD net56 sky130_fd_sc_hd__clkdlybuf4s50_1
x45 net59 VSS VSS VDD VDD net57 sky130_fd_sc_hd__clkdlybuf4s50_1
x48 net60 VSS VSS VDD VDD net58 sky130_fd_sc_hd__clkdlybuf4s50_1
x49 net61 VSS VSS VDD VDD net59 sky130_fd_sc_hd__clkdlybuf4s50_1
x52 net62 VSS VSS VDD VDD net60 sky130_fd_sc_hd__clkdlybuf4s50_1
x53 net63 VSS VSS VDD VDD net61 sky130_fd_sc_hd__clkdlybuf4s50_1
x56 net64 VSS VSS VDD VDD net62 sky130_fd_sc_hd__clkdlybuf4s50_1
x57 net65 VSS VSS VDD VDD net63 sky130_fd_sc_hd__clkdlybuf4s50_1
x60 net66 VSS VSS VDD VDD net64 sky130_fd_sc_hd__clkdlybuf4s50_1
x61 net67 VSS VSS VDD VDD net65 sky130_fd_sc_hd__clkdlybuf4s50_1
x64 net68 VSS VSS VDD VDD net66 sky130_fd_sc_hd__clkdlybuf4s50_1
x65 net69 VSS VSS VDD VDD net67 sky130_fd_sc_hd__clkdlybuf4s50_1
x68 net70 VSS VSS VDD VDD net68 sky130_fd_sc_hd__clkdlybuf4s50_1
x69 net71 VSS VSS VDD VDD net69 sky130_fd_sc_hd__clkdlybuf4s50_1
x72 net72 VSS VSS VDD VDD net70 sky130_fd_sc_hd__clkdlybuf4s50_1
x73 net73 VSS VSS VDD VDD net71 sky130_fd_sc_hd__clkdlybuf4s50_1
x76 net74 VSS VSS VDD VDD net72 sky130_fd_sc_hd__clkdlybuf4s50_1
x77 net75 VSS VSS VDD VDD net73 sky130_fd_sc_hd__clkdlybuf4s50_1
x80 net76 VSS VSS VDD VDD net74 sky130_fd_sc_hd__clkdlybuf4s50_1
x81 net77 VSS VSS VDD VDD net75 sky130_fd_sc_hd__clkdlybuf4s50_1
x84 net78 VSS VSS VDD VDD net79 sky130_fd_sc_hd__clkdlybuf4s50_1
x85 net80 VSS VSS VDD VDD net81 sky130_fd_sc_hd__clkdlybuf4s50_1
x86 net82 VSS VSS VDD VDD net78 sky130_fd_sc_hd__clkdlybuf4s50_1
x87 net83 VSS VSS VDD VDD net80 sky130_fd_sc_hd__clkdlybuf4s50_1
x88 net29 VSS VSS VDD VDD net82 sky130_fd_sc_hd__clkdlybuf4s50_1
x89 net28 VSS VSS VDD VDD net83 sky130_fd_sc_hd__clkdlybuf4s50_1
x30 clk_div net17 VSS VSS VDD VDD net9 sky130_fd_sc_hd__nand2_1
x31 net16 net12 VSS VSS VDD VDD net13 sky130_fd_sc_hd__nand2_1
x34 net9 VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkinv_4
x35 net10 VSS VSS VDD VDD net84 sky130_fd_sc_hd__clkinv_1
x38 net13 VSS VSS VDD VDD net14 sky130_fd_sc_hd__clkinv_4
x39 net14 VSS VSS VDD VDD net85 sky130_fd_sc_hd__clkinv_1
x42 clk_div VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkinv_1
x43 net86 VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkdlybuf4s50_1
x46 net87 VSS VSS VDD VDD net16 sky130_fd_sc_hd__clkdlybuf4s50_1
x47 net84 VSS VSS VDD VDD net88 sky130_fd_sc_hd__clkdlybuf4s50_1
x50 net85 VSS VSS VDD VDD net89 sky130_fd_sc_hd__clkdlybuf4s50_1
x51 net90 VSS VSS VDD VDD net86 sky130_fd_sc_hd__clkdlybuf4s50_1
x54 net91 VSS VSS VDD VDD net87 sky130_fd_sc_hd__clkdlybuf4s50_1
x55 net88 VSS VSS VDD VDD net92 sky130_fd_sc_hd__clkdlybuf4s50_1
x58 net89 VSS VSS VDD VDD net93 sky130_fd_sc_hd__clkdlybuf4s50_1
x59 net94 VSS VSS VDD VDD net90 sky130_fd_sc_hd__clkdlybuf4s50_1
x62 net95 VSS VSS VDD VDD net91 sky130_fd_sc_hd__clkdlybuf4s50_1
x63 net92 VSS VSS VDD VDD net96 sky130_fd_sc_hd__clkdlybuf4s50_1
x66 net93 VSS VSS VDD VDD net97 sky130_fd_sc_hd__clkdlybuf4s50_1
x67 net98 VSS VSS VDD VDD net94 sky130_fd_sc_hd__clkdlybuf4s50_1
x70 net99 VSS VSS VDD VDD net95 sky130_fd_sc_hd__clkdlybuf4s50_1
x71 net96 VSS VSS VDD VDD net18 sky130_fd_sc_hd__clkdlybuf4s50_1
x74 net97 VSS VSS VDD VDD net20 sky130_fd_sc_hd__clkdlybuf4s50_1
x75 net100 VSS VSS VDD VDD net98 sky130_fd_sc_hd__clkdlybuf4s50_1
x136 net101 VSS VSS VDD VDD net99 sky130_fd_sc_hd__clkdlybuf4s50_1
x137 net102 VSS VSS VDD VDD net100 sky130_fd_sc_hd__clkdlybuf4s50_1
x138 net103 VSS VSS VDD VDD net101 sky130_fd_sc_hd__clkdlybuf4s50_1
x139 net104 VSS VSS VDD VDD net102 sky130_fd_sc_hd__clkdlybuf4s50_1
x140 net105 VSS VSS VDD VDD net103 sky130_fd_sc_hd__clkdlybuf4s50_1
x141 net106 VSS VSS VDD VDD net104 sky130_fd_sc_hd__clkdlybuf4s50_1
x142 net107 VSS VSS VDD VDD net105 sky130_fd_sc_hd__clkdlybuf4s50_1
x143 net108 VSS VSS VDD VDD net106 sky130_fd_sc_hd__clkdlybuf4s50_1
x144 net109 VSS VSS VDD VDD net107 sky130_fd_sc_hd__clkdlybuf4s50_1
x145 net110 VSS VSS VDD VDD net108 sky130_fd_sc_hd__clkdlybuf4s50_1
x146 net111 VSS VSS VDD VDD net109 sky130_fd_sc_hd__clkdlybuf4s50_1
x147 net112 VSS VSS VDD VDD net110 sky130_fd_sc_hd__clkdlybuf4s50_1
x148 net113 VSS VSS VDD VDD net111 sky130_fd_sc_hd__clkdlybuf4s50_1
x149 net114 VSS VSS VDD VDD net112 sky130_fd_sc_hd__clkdlybuf4s50_1
x150 net115 VSS VSS VDD VDD net113 sky130_fd_sc_hd__clkdlybuf4s50_1
x151 net116 VSS VSS VDD VDD net114 sky130_fd_sc_hd__clkdlybuf4s50_1
x152 net117 VSS VSS VDD VDD net115 sky130_fd_sc_hd__clkdlybuf4s50_1
x153 net118 VSS VSS VDD VDD net116 sky130_fd_sc_hd__clkdlybuf4s50_1
x154 net119 VSS VSS VDD VDD net117 sky130_fd_sc_hd__clkdlybuf4s50_1
x155 net120 VSS VSS VDD VDD net118 sky130_fd_sc_hd__clkdlybuf4s50_1
x156 net121 VSS VSS VDD VDD net119 sky130_fd_sc_hd__clkdlybuf4s50_1
x157 net122 VSS VSS VDD VDD net120 sky130_fd_sc_hd__clkdlybuf4s50_1
x158 net123 VSS VSS VDD VDD net121 sky130_fd_sc_hd__clkdlybuf4s50_1
x195 net9 net18 VSS VSS VDD VDD net23 sky130_fd_sc_hd__nand2_4
x196 net10 VSS VSS VDD VDD net22 sky130_fd_sc_hd__clkinv_4
x197 net14 VSS VSS VDD VDD net21 sky130_fd_sc_hd__clkinv_4
x198 net13 net20 VSS VSS VDD VDD net19 sky130_fd_sc_hd__nand2_4
x223 clk net24 VSS VSS VDD VDD clk_div net24 sky130_fd_sc_hd__dfxbp_1
x224 p2 clk_div VSS VSS VDD VDD net25 net124 sky130_fd_sc_hd__dfxbp_1
x225 Ad_b Bd_b net25 VSS VSS VDD VDD net26 sky130_fd_sc_hd__mux2_1
x226 net26 latch_in VSS VSS VDD VDD net27 sky130_fd_sc_hd__nand2_1
x227 net27 VSS VSS VDD VDD latch_out sky130_fd_sc_hd__clkinv_1
x232 net22 VSS VSS VDD VDD A_b sky130_fd_sc_hd__clkbuf_16
x233 net10 VSS VSS VDD VDD A sky130_fd_sc_hd__clkbuf_16
x234 net11 VSS VSS VDD VDD Ad_b sky130_fd_sc_hd__clkbuf_16
x235 net23 VSS VSS VDD VDD Ad sky130_fd_sc_hd__clkbuf_16
x236 net19 VSS VSS VDD VDD Bd sky130_fd_sc_hd__clkbuf_16
x237 net15 VSS VSS VDD VDD Bd_b sky130_fd_sc_hd__clkbuf_16
x238 net14 VSS VSS VDD VDD B sky130_fd_sc_hd__clkbuf_16
x239 net21 VSS VSS VDD VDD B_b sky130_fd_sc_hd__clkbuf_16
x228 net23 VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkinv_4
x229 net19 VSS VSS VDD VDD net15 sky130_fd_sc_hd__clkinv_4
x5 net1 net7 VSS VSS VDD VDD net33 sky130_fd_sc_hd__nand2_4
x10 net2 VSS VSS VDD VDD net32 sky130_fd_sc_hd__clkinv_4
x116 net5 VSS VSS VDD VDD net31 sky130_fd_sc_hd__clkinv_4
x117 net4 net8 VSS VSS VDD VDD net30 sky130_fd_sc_hd__nand2_4
x230 net32 VSS VSS VDD VDD p2_b sky130_fd_sc_hd__clkbuf_16
x231 net2 VSS VSS VDD VDD p2 sky130_fd_sc_hd__clkbuf_16
x240 net28 VSS VSS VDD VDD p2d_b sky130_fd_sc_hd__clkbuf_16
x241 net33 VSS VSS VDD VDD p2d sky130_fd_sc_hd__clkbuf_16
x242 net30 VSS VSS VDD VDD p1d sky130_fd_sc_hd__clkbuf_16
x243 net29 VSS VSS VDD VDD p1d_b sky130_fd_sc_hd__clkbuf_16
x244 net5 VSS VSS VDD VDD p1 sky130_fd_sc_hd__clkbuf_16
x245 net31 VSS VSS VDD VDD p1_b sky130_fd_sc_hd__clkbuf_16
x246 net33 VSS VSS VDD VDD net28 sky130_fd_sc_hd__clkinv_4
x247 net30 VSS VSS VDD VDD net29 sky130_fd_sc_hd__clkinv_4
x8 net125 VSS VSS VDD VDD net123 sky130_fd_sc_hd__clkdlybuf4s50_1
x13 net126 VSS VSS VDD VDD net122 sky130_fd_sc_hd__clkdlybuf4s50_1
x78 net127 VSS VSS VDD VDD net125 sky130_fd_sc_hd__clkdlybuf4s50_1
x79 net128 VSS VSS VDD VDD net126 sky130_fd_sc_hd__clkdlybuf4s50_1
x82 net129 VSS VSS VDD VDD net130 sky130_fd_sc_hd__clkdlybuf4s50_1
x83 net131 VSS VSS VDD VDD net132 sky130_fd_sc_hd__clkdlybuf4s50_1
x90 net133 VSS VSS VDD VDD net129 sky130_fd_sc_hd__clkdlybuf4s50_1
x91 net134 VSS VSS VDD VDD net131 sky130_fd_sc_hd__clkdlybuf4s50_1
x92 net11 VSS VSS VDD VDD net133 sky130_fd_sc_hd__clkdlybuf4s50_1
x93 net15 VSS VSS VDD VDD net134 sky130_fd_sc_hd__clkdlybuf4s50_1
x94 net135 VSS VSS VDD VDD net128 sky130_fd_sc_hd__clkdlybuf4s50_1
x95 net136 VSS VSS VDD VDD net127 sky130_fd_sc_hd__clkdlybuf4s50_1
x96 net137 VSS VSS VDD VDD net135 sky130_fd_sc_hd__clkdlybuf4s50_1
x97 net138 VSS VSS VDD VDD net136 sky130_fd_sc_hd__clkdlybuf4s50_1
x98 net139 VSS VSS VDD VDD net137 sky130_fd_sc_hd__clkdlybuf4s50_1
x99 net140 VSS VSS VDD VDD net138 sky130_fd_sc_hd__clkdlybuf4s50_1
x100 net141 VSS VSS VDD VDD net140 sky130_fd_sc_hd__clkdlybuf4s50_1
x101 net142 VSS VSS VDD VDD net139 sky130_fd_sc_hd__clkdlybuf4s50_1
x102 net130 VSS VSS VDD VDD net141 sky130_fd_sc_hd__clkdlybuf4s50_1
x103 net132 VSS VSS VDD VDD net142 sky130_fd_sc_hd__clkdlybuf4s50_1
x104 net143 VSS VSS VDD VDD net77 sky130_fd_sc_hd__clkdlybuf4s50_1
x105 net144 VSS VSS VDD VDD net76 sky130_fd_sc_hd__clkdlybuf4s50_1
x106 net145 VSS VSS VDD VDD net143 sky130_fd_sc_hd__clkdlybuf4s50_1
x107 net146 VSS VSS VDD VDD net144 sky130_fd_sc_hd__clkdlybuf4s50_1
x108 net147 VSS VSS VDD VDD net145 sky130_fd_sc_hd__clkdlybuf4s50_1
x109 net148 VSS VSS VDD VDD net146 sky130_fd_sc_hd__clkdlybuf4s50_1
x110 net149 VSS VSS VDD VDD net148 sky130_fd_sc_hd__clkdlybuf4s50_1
x111 net150 VSS VSS VDD VDD net147 sky130_fd_sc_hd__clkdlybuf4s50_1
x112 net79 VSS VSS VDD VDD net149 sky130_fd_sc_hd__clkdlybuf4s50_1
x113 net81 VSS VSS VDD VDD net150 sky130_fd_sc_hd__clkdlybuf4s50_1
.ends


* expanding   symbol:  transmission_gate.sym # of pins=4
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/transmission_gate.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/transmission_gate.sch
.subckt transmission_gate  in out en en_b  VDD  VSS     N=1 W_N=5.3 L_N=0.15 W_P=13.7 L_P=0.15
*.iopin in
*.iopin out
*.ipin en
*.ipin en_b
XM1 out en in VSS sky130_fd_pr__nfet_01v8 L='L_N' W='W_N' nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='N' m='N' 
XM2 out en_b in VDD sky130_fd_pr__pfet_01v8 L='L_P' W='W_P' nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult='N' m='N' 
.ends


* expanding   symbol:  1b_dac.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/1b_dac.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/1b_dac.sch
.subckt 1b_dac  v_hi v_lo v out v_b  VDD  VSS
*.ipin v_hi
*.ipin v_lo
*.ipin v
*.ipin v_b
*.opin out
x1 v_hi out v v_b VDD VSS transmission_gate
x2 v_lo out v_b v VDD VSS transmission_gate
.ends


* expanding   symbol:  comparator.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator.sch
.subckt comparator  ip in outp clk outn  VDD  VSS
*.ipin clk
*.ipin ip
*.ipin in
*.opin outp
*.opin outn
x2 s_b VSS VSS VDD VDD s_b_buf sky130_fd_sc_hd__buf_2
x3 r_b VSS VSS VDD VDD r_b_buf sky130_fd_sc_hd__buf_2
x4 s_b_buf r_b_buf outp outn VDD VSS rs_b_latch
x1 ip in s_b clk r_b VDD VSS comparator_core_large
.ends


* expanding   symbol:  ota_w_test.sym # of pins=15
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota_w_test.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota_w_test.sch
.subckt ota_w_test  i_bias ip in phi1 phi1_b phi2 phi2_b op on cm bias_a bias_b bias_c bias_d cmc
+  VDD  VSS
*.ipin ip
*.ipin in
*.ipin phi1
*.ipin phi1_b
*.ipin phi2
*.ipin phi2_b
*.opin op
*.opin on
*.ipin i_bias
*.opin cm
*.opin bias_a
*.opin bias_b
*.opin bias_c
*.opin bias_d
*.opin cmc
x1 bias_a bias_b bias_c bias_d cm i_bias VDD VSS folded_cascode_3_bias
x3 phi1 phi1_b op on cm bias_a cmc phi2 phi2_b VDD VSS sc_cmfb
x2 cmc ip in bias_a bias_b bias_c bias_d op on VDD VSS folded_cascode_3_core
.ends


* expanding   symbol:  ota.sym # of pins=10
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/ota.sch
.subckt ota  i_bias ip in phi1 phi1_b phi2 phi2_b op on cm  VDD  VSS
*.ipin ip
*.ipin in
*.ipin phi1
*.ipin phi1_b
*.ipin phi2
*.ipin phi2_b
*.opin op
*.opin on
*.ipin i_bias
*.opin cm
x1 bias_a bias_b bias_c bias_d cm i_bias VDD VSS folded_cascode_3_bias
x3 phi1 phi1_b op on cm bias_a cmc phi2 phi2_b VDD VSS sc_cmfb
x2 cmc ip in bias_a bias_b bias_c bias_d op on VDD VSS folded_cascode_3_core
.ends


* expanding   symbol:  switch_5t.sym # of pins=4
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/switch_5t.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/switch_5t.sch
.subckt switch_5t  in out en en_b  VDD  VSS
*.iopin in
*.iopin out
*.ipin en
*.ipin en_b
x1 in net1 en en_b VDD VSS transmission_gate
x2 net1 out en en_b VDD VSS transmission_gate
XM1 net1 en_b VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  rs_b_latch.sym # of pins=4
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/rs_b_latch.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/rs_b_latch.sch
.subckt rs_b_latch  s_b r_b q q_b  VDD  VSS
*.ipin s_b
*.ipin r_b
*.opin q
*.opin q_b
x1 s_b q_b VSS VSS VDD VDD q sky130_fd_sc_hd__nand2_4
x2 r_b q VSS VSS VDD VDD q_b sky130_fd_sc_hd__nand2_4
.ends


* expanding   symbol:  comparator_core_large.sym # of pins=5
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator_core_large.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/comparator_core_large.sch
.subckt comparator_core_large  ip in s_b clk r_b  VDD  VSS
*.ipin clk
*.ipin ip
*.ipin in
*.opin s_b
*.opin r_b
XM1 tail_d clk VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=32 m=32 
XM2 p ip tail_d VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=160 m=160 
XM3 q in tail_d VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=160 m=160 
XM4 s_b r_b p VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=80 m=80 
XM5 r_b s_b q VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=80 m=80 
XM6 s_b r_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=40 m=40 
XM7 r_b s_b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=40 m=40 
XM8 s_b clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM9 r_b clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM10 p clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM11 q clk VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM12 tail_d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM13 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=24 m=24 
XM17 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM14 q VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM15 p VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM16 r_b VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM18 s_b VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
.ends


* expanding   symbol:  folded_cascode_3_bias.sym # of pins=6
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_bias.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_bias.sch
.subckt folded_cascode_3_bias  bias_a bias_b bias_c bias_d bias_e i_bias  VDD  VSS
*.opin bias_a
*.opin bias_b
*.opin bias_c
*.opin bias_d
*.opin bias_e
*.ipin i_bias
XM22 bias_b bias_c m21d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM26 m2d bias_c m25d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM32 bias_e bias_c m31d VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM21 m21d bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM25 m25d bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM31 m31d bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6 
XM1 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=56 m=56 
XM2 m2d m2d bias_d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=50 m=50 
XM3 bias_d m2d bias_a VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM4 bias_a bias_d m5d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM5 m5d bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM6 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM7 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=18 m=18 
XM33 bias_e bias_e net1 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM49 net1 bias_e net2 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM50 net2 bias_e net3 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM63 net3 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM68 bias_e bias_e net4 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM69 net4 bias_e net5 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM70 net5 bias_e net6 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM71 net6 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM72 bias_e bias_e net7 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM73 net7 bias_e net8 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM74 net8 bias_e net9 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM75 net9 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM76 bias_e bias_e net10 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM77 net10 bias_e net11 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM78 net11 bias_e net12 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM79 net12 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM64 bias_e bias_e net13 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM65 net13 bias_e net14 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM66 net14 bias_e net15 VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM67 net15 bias_e VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM44 i_bias VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM8 bias_c VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM9 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=14 m=14 
XM11 m21d VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM12 m25d VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM13 m2d VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM14 m2d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM10 bias_b VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM15 bias_b VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM16 bias_d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM17 bias_a VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM18 m31d VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM19 bias_e VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM20 m5d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
.ends


* expanding   symbol:  sc_cmfb.sym # of pins=9
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/sc_cmfb.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/sc_cmfb.sch
.subckt sc_cmfb  phi1 phi1_b op on cm bias_a cmc phi2 phi2_b  VDD  VSS
*.ipin on
*.ipin cm
*.ipin bias_a
*.ipin op
*.opin cmc
*.ipin phi2_b
*.ipin phi2
*.ipin phi1_b
*.ipin phi1
XC3 op cmc sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=4 m=4
XC4 on cmc sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=4 m=4
x1 net1 op phi2 phi2_b VDD VSS transmission_gate
x2 net2 cmc phi2 phi2_b VDD VSS transmission_gate
x3 net3 on phi2 phi2_b VDD VSS transmission_gate
x4 cm net1 phi1 phi1_b VDD VSS transmission_gate
x5 bias_a net2 phi1 phi1_b VDD VSS transmission_gate
x6 cm net3 phi1 phi1_b VDD VSS transmission_gate
XC1 net1 net2 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
XC2 net3 net2 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
x7 cm net4 phi2 phi2_b VDD VSS transmission_gate
x8 bias_a net5 phi2 phi2_b VDD VSS transmission_gate
x9 cm net6 phi2 phi2_b VDD VSS transmission_gate
x10 net4 op phi1 phi1_b VDD VSS transmission_gate
x11 net5 cmc phi1 phi1_b VDD VSS transmission_gate
x12 net6 on phi1 phi1_b VDD VSS transmission_gate
XC5 net4 net5 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
XC6 net6 net5 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=2 m=2
XCdummy __UNCONNECTED_PIN__4 __UNCONNECTED_PIN__5 sky130_fd_pr__cap_mim_m3_1 W=4.8 L=4.8 MF=20 m=20
.ends


* expanding   symbol:  folded_cascode_3_core.sym # of pins=9
* sym_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_core.sym
* sch_path:
*+ /home/users/rhyang/ee372/incremental_delta_sigma_adc/design/analog_modulator/schematic/folded_cascode_3_core.sch
.subckt folded_cascode_3_core  cmc ip in bias_a bias_b bias_c bias_d op on  VDD  VSS
*.ipin cmc
*.ipin ip
*.ipin in
*.ipin bias_a
*.ipin bias_b
*.ipin bias_c
*.ipin bias_d
*.opin op
*.opin on
XM1 foldp ip tail VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM2 foldn in tail VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM6 tail cmc VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=96 m=96 
XM5 tail bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=96 m=96 
XM11 foldp bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24 
XM12 foldn bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24 
XM1A on bias_c foldp VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM8 op bias_c foldn VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20 
XM3A on bias_d m3d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM7 op bias_d m4d VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM3 m3d bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM4 m4d bias_a VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=36 m=36 
XM17 tail VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=24 m=24 
XM10 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.2 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM9 foldp VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM13 foldn VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4 
XM14 on VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM15 on VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM16 op VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM18 op VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM19 m3d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
XM20 m4d VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.6 W=1.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=6 m=6 
.ends


