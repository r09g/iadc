magic
tech sky130A
magscale 1 2
timestamp 1652665259
<< locali >>
rect -216 891 -166 925
rect -87 430 -53 993
rect 81 891 1107 925
rect -216 396 -53 430
rect 1270 396 1304 430
rect -216 84 -166 118
rect -87 19 -53 396
rect 81 84 1107 118
<< viali >>
rect -87 993 -53 1027
rect -166 891 -132 925
rect 1171 545 1205 931
rect 1236 396 1270 430
rect -166 84 -132 118
rect 1171 81 1205 281
rect -87 -15 -53 19
<< metal1 >>
rect -99 1027 -41 1033
rect -99 993 -87 1027
rect -53 993 995 1027
rect -99 987 -41 993
rect -178 925 -120 931
rect 78 925 150 935
rect -178 891 -166 925
rect -132 891 150 925
rect -178 885 -120 891
rect 78 883 150 891
rect 193 832 227 993
rect 271 883 343 935
rect 385 832 419 993
rect 462 883 534 935
rect 577 832 611 993
rect 654 883 726 935
rect 769 832 803 993
rect 846 883 918 935
rect 961 832 995 993
rect 1038 883 1110 935
rect 1165 931 1211 1063
rect 97 430 131 608
rect 289 430 323 608
rect 481 430 515 608
rect 673 430 707 608
rect 865 430 899 608
rect 1057 430 1091 608
rect 1165 545 1171 931
rect 1205 545 1211 931
rect 1165 533 1211 545
rect 1224 430 1282 436
rect 97 396 1236 430
rect 1270 396 1282 430
rect 97 253 131 396
rect 289 253 323 396
rect 481 253 515 396
rect 673 253 707 396
rect 865 253 899 396
rect 1057 253 1091 396
rect 1224 390 1282 396
rect 1165 281 1211 293
rect -178 118 -120 124
rect 78 118 150 128
rect -178 84 -166 118
rect -132 84 150 118
rect -178 78 -120 84
rect 78 76 150 84
rect -99 19 -41 25
rect 193 19 227 180
rect 269 76 341 128
rect 385 19 419 180
rect 461 76 533 128
rect 577 19 611 180
rect 653 76 725 128
rect 769 19 803 180
rect 846 75 918 127
rect 961 19 995 180
rect 1038 75 1110 127
rect 1165 81 1171 281
rect 1205 81 1211 281
rect -99 -15 -87 19
rect -53 -15 995 19
rect -99 -21 -41 -15
rect 1165 -51 1211 81
use sky130_fd_pr__nfet_01v8_6J4AMR  sky130_fd_pr__nfet_01v8_6J4AMR_0
timestamp 1652660033
transform 1 0 594 0 1 212
box -647 -263 647 201
use sky130_fd_pr__pfet_01v8_UNG2NQ  sky130_fd_pr__pfet_01v8_UNG2NQ_0
timestamp 1652659422
transform -1 0 594 0 -1 707
box -647 -356 647 294
<< labels >>
flabel metal1 1188 -48 1188 -48 1 FreeSans 400 0 0 0 VSS
flabel metal1 1188 1058 1188 1058 5 FreeSans 400 0 0 0 VDD
flabel locali 1301 413 1301 413 7 FreeSans 400 0 0 0 out
flabel locali -213 413 -213 413 3 FreeSans 400 0 0 0 in
flabel locali -213 908 -213 908 3 FreeSans 400 0 0 0 en_b
flabel locali -213 101 -213 101 3 FreeSans 400 0 0 0 en
<< end >>
