magic
tech sky130A
magscale 1 2
timestamp 1654583101
<< pwell >>
rect -3170 -166 3170 166
<< nmos >>
rect -3086 -140 -2966 140
rect -2908 -140 -2788 140
rect -2730 -140 -2610 140
rect -2552 -140 -2432 140
rect -2374 -140 -2254 140
rect -2196 -140 -2076 140
rect -2018 -140 -1898 140
rect -1840 -140 -1720 140
rect -1662 -140 -1542 140
rect -1484 -140 -1364 140
rect -1306 -140 -1186 140
rect -1128 -140 -1008 140
rect -950 -140 -830 140
rect -772 -140 -652 140
rect -594 -140 -474 140
rect -416 -140 -296 140
rect -238 -140 -118 140
rect -60 -140 60 140
rect 118 -140 238 140
rect 296 -140 416 140
rect 474 -140 594 140
rect 652 -140 772 140
rect 830 -140 950 140
rect 1008 -140 1128 140
rect 1186 -140 1306 140
rect 1364 -140 1484 140
rect 1542 -140 1662 140
rect 1720 -140 1840 140
rect 1898 -140 2018 140
rect 2076 -140 2196 140
rect 2254 -140 2374 140
rect 2432 -140 2552 140
rect 2610 -140 2730 140
rect 2788 -140 2908 140
rect 2966 -140 3086 140
<< ndiff >>
rect -3144 119 -3086 140
rect -3144 85 -3132 119
rect -3098 85 -3086 119
rect -3144 51 -3086 85
rect -3144 17 -3132 51
rect -3098 17 -3086 51
rect -3144 -17 -3086 17
rect -3144 -51 -3132 -17
rect -3098 -51 -3086 -17
rect -3144 -85 -3086 -51
rect -3144 -119 -3132 -85
rect -3098 -119 -3086 -85
rect -3144 -140 -3086 -119
rect -2966 119 -2908 140
rect -2966 85 -2954 119
rect -2920 85 -2908 119
rect -2966 51 -2908 85
rect -2966 17 -2954 51
rect -2920 17 -2908 51
rect -2966 -17 -2908 17
rect -2966 -51 -2954 -17
rect -2920 -51 -2908 -17
rect -2966 -85 -2908 -51
rect -2966 -119 -2954 -85
rect -2920 -119 -2908 -85
rect -2966 -140 -2908 -119
rect -2788 119 -2730 140
rect -2788 85 -2776 119
rect -2742 85 -2730 119
rect -2788 51 -2730 85
rect -2788 17 -2776 51
rect -2742 17 -2730 51
rect -2788 -17 -2730 17
rect -2788 -51 -2776 -17
rect -2742 -51 -2730 -17
rect -2788 -85 -2730 -51
rect -2788 -119 -2776 -85
rect -2742 -119 -2730 -85
rect -2788 -140 -2730 -119
rect -2610 119 -2552 140
rect -2610 85 -2598 119
rect -2564 85 -2552 119
rect -2610 51 -2552 85
rect -2610 17 -2598 51
rect -2564 17 -2552 51
rect -2610 -17 -2552 17
rect -2610 -51 -2598 -17
rect -2564 -51 -2552 -17
rect -2610 -85 -2552 -51
rect -2610 -119 -2598 -85
rect -2564 -119 -2552 -85
rect -2610 -140 -2552 -119
rect -2432 119 -2374 140
rect -2432 85 -2420 119
rect -2386 85 -2374 119
rect -2432 51 -2374 85
rect -2432 17 -2420 51
rect -2386 17 -2374 51
rect -2432 -17 -2374 17
rect -2432 -51 -2420 -17
rect -2386 -51 -2374 -17
rect -2432 -85 -2374 -51
rect -2432 -119 -2420 -85
rect -2386 -119 -2374 -85
rect -2432 -140 -2374 -119
rect -2254 119 -2196 140
rect -2254 85 -2242 119
rect -2208 85 -2196 119
rect -2254 51 -2196 85
rect -2254 17 -2242 51
rect -2208 17 -2196 51
rect -2254 -17 -2196 17
rect -2254 -51 -2242 -17
rect -2208 -51 -2196 -17
rect -2254 -85 -2196 -51
rect -2254 -119 -2242 -85
rect -2208 -119 -2196 -85
rect -2254 -140 -2196 -119
rect -2076 119 -2018 140
rect -2076 85 -2064 119
rect -2030 85 -2018 119
rect -2076 51 -2018 85
rect -2076 17 -2064 51
rect -2030 17 -2018 51
rect -2076 -17 -2018 17
rect -2076 -51 -2064 -17
rect -2030 -51 -2018 -17
rect -2076 -85 -2018 -51
rect -2076 -119 -2064 -85
rect -2030 -119 -2018 -85
rect -2076 -140 -2018 -119
rect -1898 119 -1840 140
rect -1898 85 -1886 119
rect -1852 85 -1840 119
rect -1898 51 -1840 85
rect -1898 17 -1886 51
rect -1852 17 -1840 51
rect -1898 -17 -1840 17
rect -1898 -51 -1886 -17
rect -1852 -51 -1840 -17
rect -1898 -85 -1840 -51
rect -1898 -119 -1886 -85
rect -1852 -119 -1840 -85
rect -1898 -140 -1840 -119
rect -1720 119 -1662 140
rect -1720 85 -1708 119
rect -1674 85 -1662 119
rect -1720 51 -1662 85
rect -1720 17 -1708 51
rect -1674 17 -1662 51
rect -1720 -17 -1662 17
rect -1720 -51 -1708 -17
rect -1674 -51 -1662 -17
rect -1720 -85 -1662 -51
rect -1720 -119 -1708 -85
rect -1674 -119 -1662 -85
rect -1720 -140 -1662 -119
rect -1542 119 -1484 140
rect -1542 85 -1530 119
rect -1496 85 -1484 119
rect -1542 51 -1484 85
rect -1542 17 -1530 51
rect -1496 17 -1484 51
rect -1542 -17 -1484 17
rect -1542 -51 -1530 -17
rect -1496 -51 -1484 -17
rect -1542 -85 -1484 -51
rect -1542 -119 -1530 -85
rect -1496 -119 -1484 -85
rect -1542 -140 -1484 -119
rect -1364 119 -1306 140
rect -1364 85 -1352 119
rect -1318 85 -1306 119
rect -1364 51 -1306 85
rect -1364 17 -1352 51
rect -1318 17 -1306 51
rect -1364 -17 -1306 17
rect -1364 -51 -1352 -17
rect -1318 -51 -1306 -17
rect -1364 -85 -1306 -51
rect -1364 -119 -1352 -85
rect -1318 -119 -1306 -85
rect -1364 -140 -1306 -119
rect -1186 119 -1128 140
rect -1186 85 -1174 119
rect -1140 85 -1128 119
rect -1186 51 -1128 85
rect -1186 17 -1174 51
rect -1140 17 -1128 51
rect -1186 -17 -1128 17
rect -1186 -51 -1174 -17
rect -1140 -51 -1128 -17
rect -1186 -85 -1128 -51
rect -1186 -119 -1174 -85
rect -1140 -119 -1128 -85
rect -1186 -140 -1128 -119
rect -1008 119 -950 140
rect -1008 85 -996 119
rect -962 85 -950 119
rect -1008 51 -950 85
rect -1008 17 -996 51
rect -962 17 -950 51
rect -1008 -17 -950 17
rect -1008 -51 -996 -17
rect -962 -51 -950 -17
rect -1008 -85 -950 -51
rect -1008 -119 -996 -85
rect -962 -119 -950 -85
rect -1008 -140 -950 -119
rect -830 119 -772 140
rect -830 85 -818 119
rect -784 85 -772 119
rect -830 51 -772 85
rect -830 17 -818 51
rect -784 17 -772 51
rect -830 -17 -772 17
rect -830 -51 -818 -17
rect -784 -51 -772 -17
rect -830 -85 -772 -51
rect -830 -119 -818 -85
rect -784 -119 -772 -85
rect -830 -140 -772 -119
rect -652 119 -594 140
rect -652 85 -640 119
rect -606 85 -594 119
rect -652 51 -594 85
rect -652 17 -640 51
rect -606 17 -594 51
rect -652 -17 -594 17
rect -652 -51 -640 -17
rect -606 -51 -594 -17
rect -652 -85 -594 -51
rect -652 -119 -640 -85
rect -606 -119 -594 -85
rect -652 -140 -594 -119
rect -474 119 -416 140
rect -474 85 -462 119
rect -428 85 -416 119
rect -474 51 -416 85
rect -474 17 -462 51
rect -428 17 -416 51
rect -474 -17 -416 17
rect -474 -51 -462 -17
rect -428 -51 -416 -17
rect -474 -85 -416 -51
rect -474 -119 -462 -85
rect -428 -119 -416 -85
rect -474 -140 -416 -119
rect -296 119 -238 140
rect -296 85 -284 119
rect -250 85 -238 119
rect -296 51 -238 85
rect -296 17 -284 51
rect -250 17 -238 51
rect -296 -17 -238 17
rect -296 -51 -284 -17
rect -250 -51 -238 -17
rect -296 -85 -238 -51
rect -296 -119 -284 -85
rect -250 -119 -238 -85
rect -296 -140 -238 -119
rect -118 119 -60 140
rect -118 85 -106 119
rect -72 85 -60 119
rect -118 51 -60 85
rect -118 17 -106 51
rect -72 17 -60 51
rect -118 -17 -60 17
rect -118 -51 -106 -17
rect -72 -51 -60 -17
rect -118 -85 -60 -51
rect -118 -119 -106 -85
rect -72 -119 -60 -85
rect -118 -140 -60 -119
rect 60 119 118 140
rect 60 85 72 119
rect 106 85 118 119
rect 60 51 118 85
rect 60 17 72 51
rect 106 17 118 51
rect 60 -17 118 17
rect 60 -51 72 -17
rect 106 -51 118 -17
rect 60 -85 118 -51
rect 60 -119 72 -85
rect 106 -119 118 -85
rect 60 -140 118 -119
rect 238 119 296 140
rect 238 85 250 119
rect 284 85 296 119
rect 238 51 296 85
rect 238 17 250 51
rect 284 17 296 51
rect 238 -17 296 17
rect 238 -51 250 -17
rect 284 -51 296 -17
rect 238 -85 296 -51
rect 238 -119 250 -85
rect 284 -119 296 -85
rect 238 -140 296 -119
rect 416 119 474 140
rect 416 85 428 119
rect 462 85 474 119
rect 416 51 474 85
rect 416 17 428 51
rect 462 17 474 51
rect 416 -17 474 17
rect 416 -51 428 -17
rect 462 -51 474 -17
rect 416 -85 474 -51
rect 416 -119 428 -85
rect 462 -119 474 -85
rect 416 -140 474 -119
rect 594 119 652 140
rect 594 85 606 119
rect 640 85 652 119
rect 594 51 652 85
rect 594 17 606 51
rect 640 17 652 51
rect 594 -17 652 17
rect 594 -51 606 -17
rect 640 -51 652 -17
rect 594 -85 652 -51
rect 594 -119 606 -85
rect 640 -119 652 -85
rect 594 -140 652 -119
rect 772 119 830 140
rect 772 85 784 119
rect 818 85 830 119
rect 772 51 830 85
rect 772 17 784 51
rect 818 17 830 51
rect 772 -17 830 17
rect 772 -51 784 -17
rect 818 -51 830 -17
rect 772 -85 830 -51
rect 772 -119 784 -85
rect 818 -119 830 -85
rect 772 -140 830 -119
rect 950 119 1008 140
rect 950 85 962 119
rect 996 85 1008 119
rect 950 51 1008 85
rect 950 17 962 51
rect 996 17 1008 51
rect 950 -17 1008 17
rect 950 -51 962 -17
rect 996 -51 1008 -17
rect 950 -85 1008 -51
rect 950 -119 962 -85
rect 996 -119 1008 -85
rect 950 -140 1008 -119
rect 1128 119 1186 140
rect 1128 85 1140 119
rect 1174 85 1186 119
rect 1128 51 1186 85
rect 1128 17 1140 51
rect 1174 17 1186 51
rect 1128 -17 1186 17
rect 1128 -51 1140 -17
rect 1174 -51 1186 -17
rect 1128 -85 1186 -51
rect 1128 -119 1140 -85
rect 1174 -119 1186 -85
rect 1128 -140 1186 -119
rect 1306 119 1364 140
rect 1306 85 1318 119
rect 1352 85 1364 119
rect 1306 51 1364 85
rect 1306 17 1318 51
rect 1352 17 1364 51
rect 1306 -17 1364 17
rect 1306 -51 1318 -17
rect 1352 -51 1364 -17
rect 1306 -85 1364 -51
rect 1306 -119 1318 -85
rect 1352 -119 1364 -85
rect 1306 -140 1364 -119
rect 1484 119 1542 140
rect 1484 85 1496 119
rect 1530 85 1542 119
rect 1484 51 1542 85
rect 1484 17 1496 51
rect 1530 17 1542 51
rect 1484 -17 1542 17
rect 1484 -51 1496 -17
rect 1530 -51 1542 -17
rect 1484 -85 1542 -51
rect 1484 -119 1496 -85
rect 1530 -119 1542 -85
rect 1484 -140 1542 -119
rect 1662 119 1720 140
rect 1662 85 1674 119
rect 1708 85 1720 119
rect 1662 51 1720 85
rect 1662 17 1674 51
rect 1708 17 1720 51
rect 1662 -17 1720 17
rect 1662 -51 1674 -17
rect 1708 -51 1720 -17
rect 1662 -85 1720 -51
rect 1662 -119 1674 -85
rect 1708 -119 1720 -85
rect 1662 -140 1720 -119
rect 1840 119 1898 140
rect 1840 85 1852 119
rect 1886 85 1898 119
rect 1840 51 1898 85
rect 1840 17 1852 51
rect 1886 17 1898 51
rect 1840 -17 1898 17
rect 1840 -51 1852 -17
rect 1886 -51 1898 -17
rect 1840 -85 1898 -51
rect 1840 -119 1852 -85
rect 1886 -119 1898 -85
rect 1840 -140 1898 -119
rect 2018 119 2076 140
rect 2018 85 2030 119
rect 2064 85 2076 119
rect 2018 51 2076 85
rect 2018 17 2030 51
rect 2064 17 2076 51
rect 2018 -17 2076 17
rect 2018 -51 2030 -17
rect 2064 -51 2076 -17
rect 2018 -85 2076 -51
rect 2018 -119 2030 -85
rect 2064 -119 2076 -85
rect 2018 -140 2076 -119
rect 2196 119 2254 140
rect 2196 85 2208 119
rect 2242 85 2254 119
rect 2196 51 2254 85
rect 2196 17 2208 51
rect 2242 17 2254 51
rect 2196 -17 2254 17
rect 2196 -51 2208 -17
rect 2242 -51 2254 -17
rect 2196 -85 2254 -51
rect 2196 -119 2208 -85
rect 2242 -119 2254 -85
rect 2196 -140 2254 -119
rect 2374 119 2432 140
rect 2374 85 2386 119
rect 2420 85 2432 119
rect 2374 51 2432 85
rect 2374 17 2386 51
rect 2420 17 2432 51
rect 2374 -17 2432 17
rect 2374 -51 2386 -17
rect 2420 -51 2432 -17
rect 2374 -85 2432 -51
rect 2374 -119 2386 -85
rect 2420 -119 2432 -85
rect 2374 -140 2432 -119
rect 2552 119 2610 140
rect 2552 85 2564 119
rect 2598 85 2610 119
rect 2552 51 2610 85
rect 2552 17 2564 51
rect 2598 17 2610 51
rect 2552 -17 2610 17
rect 2552 -51 2564 -17
rect 2598 -51 2610 -17
rect 2552 -85 2610 -51
rect 2552 -119 2564 -85
rect 2598 -119 2610 -85
rect 2552 -140 2610 -119
rect 2730 119 2788 140
rect 2730 85 2742 119
rect 2776 85 2788 119
rect 2730 51 2788 85
rect 2730 17 2742 51
rect 2776 17 2788 51
rect 2730 -17 2788 17
rect 2730 -51 2742 -17
rect 2776 -51 2788 -17
rect 2730 -85 2788 -51
rect 2730 -119 2742 -85
rect 2776 -119 2788 -85
rect 2730 -140 2788 -119
rect 2908 119 2966 140
rect 2908 85 2920 119
rect 2954 85 2966 119
rect 2908 51 2966 85
rect 2908 17 2920 51
rect 2954 17 2966 51
rect 2908 -17 2966 17
rect 2908 -51 2920 -17
rect 2954 -51 2966 -17
rect 2908 -85 2966 -51
rect 2908 -119 2920 -85
rect 2954 -119 2966 -85
rect 2908 -140 2966 -119
rect 3086 119 3144 140
rect 3086 85 3098 119
rect 3132 85 3144 119
rect 3086 51 3144 85
rect 3086 17 3098 51
rect 3132 17 3144 51
rect 3086 -17 3144 17
rect 3086 -51 3098 -17
rect 3132 -51 3144 -17
rect 3086 -85 3144 -51
rect 3086 -119 3098 -85
rect 3132 -119 3144 -85
rect 3086 -140 3144 -119
<< ndiffc >>
rect -3132 85 -3098 119
rect -3132 17 -3098 51
rect -3132 -51 -3098 -17
rect -3132 -119 -3098 -85
rect -2954 85 -2920 119
rect -2954 17 -2920 51
rect -2954 -51 -2920 -17
rect -2954 -119 -2920 -85
rect -2776 85 -2742 119
rect -2776 17 -2742 51
rect -2776 -51 -2742 -17
rect -2776 -119 -2742 -85
rect -2598 85 -2564 119
rect -2598 17 -2564 51
rect -2598 -51 -2564 -17
rect -2598 -119 -2564 -85
rect -2420 85 -2386 119
rect -2420 17 -2386 51
rect -2420 -51 -2386 -17
rect -2420 -119 -2386 -85
rect -2242 85 -2208 119
rect -2242 17 -2208 51
rect -2242 -51 -2208 -17
rect -2242 -119 -2208 -85
rect -2064 85 -2030 119
rect -2064 17 -2030 51
rect -2064 -51 -2030 -17
rect -2064 -119 -2030 -85
rect -1886 85 -1852 119
rect -1886 17 -1852 51
rect -1886 -51 -1852 -17
rect -1886 -119 -1852 -85
rect -1708 85 -1674 119
rect -1708 17 -1674 51
rect -1708 -51 -1674 -17
rect -1708 -119 -1674 -85
rect -1530 85 -1496 119
rect -1530 17 -1496 51
rect -1530 -51 -1496 -17
rect -1530 -119 -1496 -85
rect -1352 85 -1318 119
rect -1352 17 -1318 51
rect -1352 -51 -1318 -17
rect -1352 -119 -1318 -85
rect -1174 85 -1140 119
rect -1174 17 -1140 51
rect -1174 -51 -1140 -17
rect -1174 -119 -1140 -85
rect -996 85 -962 119
rect -996 17 -962 51
rect -996 -51 -962 -17
rect -996 -119 -962 -85
rect -818 85 -784 119
rect -818 17 -784 51
rect -818 -51 -784 -17
rect -818 -119 -784 -85
rect -640 85 -606 119
rect -640 17 -606 51
rect -640 -51 -606 -17
rect -640 -119 -606 -85
rect -462 85 -428 119
rect -462 17 -428 51
rect -462 -51 -428 -17
rect -462 -119 -428 -85
rect -284 85 -250 119
rect -284 17 -250 51
rect -284 -51 -250 -17
rect -284 -119 -250 -85
rect -106 85 -72 119
rect -106 17 -72 51
rect -106 -51 -72 -17
rect -106 -119 -72 -85
rect 72 85 106 119
rect 72 17 106 51
rect 72 -51 106 -17
rect 72 -119 106 -85
rect 250 85 284 119
rect 250 17 284 51
rect 250 -51 284 -17
rect 250 -119 284 -85
rect 428 85 462 119
rect 428 17 462 51
rect 428 -51 462 -17
rect 428 -119 462 -85
rect 606 85 640 119
rect 606 17 640 51
rect 606 -51 640 -17
rect 606 -119 640 -85
rect 784 85 818 119
rect 784 17 818 51
rect 784 -51 818 -17
rect 784 -119 818 -85
rect 962 85 996 119
rect 962 17 996 51
rect 962 -51 996 -17
rect 962 -119 996 -85
rect 1140 85 1174 119
rect 1140 17 1174 51
rect 1140 -51 1174 -17
rect 1140 -119 1174 -85
rect 1318 85 1352 119
rect 1318 17 1352 51
rect 1318 -51 1352 -17
rect 1318 -119 1352 -85
rect 1496 85 1530 119
rect 1496 17 1530 51
rect 1496 -51 1530 -17
rect 1496 -119 1530 -85
rect 1674 85 1708 119
rect 1674 17 1708 51
rect 1674 -51 1708 -17
rect 1674 -119 1708 -85
rect 1852 85 1886 119
rect 1852 17 1886 51
rect 1852 -51 1886 -17
rect 1852 -119 1886 -85
rect 2030 85 2064 119
rect 2030 17 2064 51
rect 2030 -51 2064 -17
rect 2030 -119 2064 -85
rect 2208 85 2242 119
rect 2208 17 2242 51
rect 2208 -51 2242 -17
rect 2208 -119 2242 -85
rect 2386 85 2420 119
rect 2386 17 2420 51
rect 2386 -51 2420 -17
rect 2386 -119 2420 -85
rect 2564 85 2598 119
rect 2564 17 2598 51
rect 2564 -51 2598 -17
rect 2564 -119 2598 -85
rect 2742 85 2776 119
rect 2742 17 2776 51
rect 2742 -51 2776 -17
rect 2742 -119 2776 -85
rect 2920 85 2954 119
rect 2920 17 2954 51
rect 2920 -51 2954 -17
rect 2920 -119 2954 -85
rect 3098 85 3132 119
rect 3098 17 3132 51
rect 3098 -51 3132 -17
rect 3098 -119 3132 -85
<< poly >>
rect -3064 212 -2988 228
rect -3064 194 -3043 212
rect -3086 178 -3043 194
rect -3009 194 -2988 212
rect -2886 212 -2810 228
rect -2886 194 -2865 212
rect -3009 178 -2966 194
rect -3086 140 -2966 178
rect -2908 178 -2865 194
rect -2831 194 -2810 212
rect -2708 212 -2632 228
rect -2708 194 -2687 212
rect -2831 178 -2788 194
rect -2908 140 -2788 178
rect -2730 178 -2687 194
rect -2653 194 -2632 212
rect -2530 212 -2454 228
rect -2530 194 -2509 212
rect -2653 178 -2610 194
rect -2730 140 -2610 178
rect -2552 178 -2509 194
rect -2475 194 -2454 212
rect -2352 212 -2276 228
rect -2352 194 -2331 212
rect -2475 178 -2432 194
rect -2552 140 -2432 178
rect -2374 178 -2331 194
rect -2297 194 -2276 212
rect -2174 212 -2098 228
rect -2174 194 -2153 212
rect -2297 178 -2254 194
rect -2374 140 -2254 178
rect -2196 178 -2153 194
rect -2119 194 -2098 212
rect -1996 212 -1920 228
rect -1996 194 -1975 212
rect -2119 178 -2076 194
rect -2196 140 -2076 178
rect -2018 178 -1975 194
rect -1941 194 -1920 212
rect -1818 212 -1742 228
rect -1818 194 -1797 212
rect -1941 178 -1898 194
rect -2018 140 -1898 178
rect -1840 178 -1797 194
rect -1763 194 -1742 212
rect -1640 212 -1564 228
rect -1640 194 -1619 212
rect -1763 178 -1720 194
rect -1840 140 -1720 178
rect -1662 178 -1619 194
rect -1585 194 -1564 212
rect -1462 212 -1386 228
rect -1462 194 -1441 212
rect -1585 178 -1542 194
rect -1662 140 -1542 178
rect -1484 178 -1441 194
rect -1407 194 -1386 212
rect -1284 212 -1208 228
rect -1284 194 -1263 212
rect -1407 178 -1364 194
rect -1484 140 -1364 178
rect -1306 178 -1263 194
rect -1229 194 -1208 212
rect -1106 212 -1030 228
rect -1106 194 -1085 212
rect -1229 178 -1186 194
rect -1306 140 -1186 178
rect -1128 178 -1085 194
rect -1051 194 -1030 212
rect -928 212 -852 228
rect -928 194 -907 212
rect -1051 178 -1008 194
rect -1128 140 -1008 178
rect -950 178 -907 194
rect -873 194 -852 212
rect -750 212 -674 228
rect -750 194 -729 212
rect -873 178 -830 194
rect -950 140 -830 178
rect -772 178 -729 194
rect -695 194 -674 212
rect -572 212 -496 228
rect -572 194 -551 212
rect -695 178 -652 194
rect -772 140 -652 178
rect -594 178 -551 194
rect -517 194 -496 212
rect -394 212 -318 228
rect -394 194 -373 212
rect -517 178 -474 194
rect -594 140 -474 178
rect -416 178 -373 194
rect -339 194 -318 212
rect -216 212 -140 228
rect -216 194 -195 212
rect -339 178 -296 194
rect -416 140 -296 178
rect -238 178 -195 194
rect -161 194 -140 212
rect -38 212 38 228
rect -38 194 -17 212
rect -161 178 -118 194
rect -238 140 -118 178
rect -60 178 -17 194
rect 17 194 38 212
rect 140 212 216 228
rect 140 194 161 212
rect 17 178 60 194
rect -60 140 60 178
rect 118 178 161 194
rect 195 194 216 212
rect 318 212 394 228
rect 318 194 339 212
rect 195 178 238 194
rect 118 140 238 178
rect 296 178 339 194
rect 373 194 394 212
rect 496 212 572 228
rect 496 194 517 212
rect 373 178 416 194
rect 296 140 416 178
rect 474 178 517 194
rect 551 194 572 212
rect 674 212 750 228
rect 674 194 695 212
rect 551 178 594 194
rect 474 140 594 178
rect 652 178 695 194
rect 729 194 750 212
rect 852 212 928 228
rect 852 194 873 212
rect 729 178 772 194
rect 652 140 772 178
rect 830 178 873 194
rect 907 194 928 212
rect 1030 212 1106 228
rect 1030 194 1051 212
rect 907 178 950 194
rect 830 140 950 178
rect 1008 178 1051 194
rect 1085 194 1106 212
rect 1208 212 1284 228
rect 1208 194 1229 212
rect 1085 178 1128 194
rect 1008 140 1128 178
rect 1186 178 1229 194
rect 1263 194 1284 212
rect 1386 212 1462 228
rect 1386 194 1407 212
rect 1263 178 1306 194
rect 1186 140 1306 178
rect 1364 178 1407 194
rect 1441 194 1462 212
rect 1564 212 1640 228
rect 1564 194 1585 212
rect 1441 178 1484 194
rect 1364 140 1484 178
rect 1542 178 1585 194
rect 1619 194 1640 212
rect 1742 212 1818 228
rect 1742 194 1763 212
rect 1619 178 1662 194
rect 1542 140 1662 178
rect 1720 178 1763 194
rect 1797 194 1818 212
rect 1920 212 1996 228
rect 1920 194 1941 212
rect 1797 178 1840 194
rect 1720 140 1840 178
rect 1898 178 1941 194
rect 1975 194 1996 212
rect 2098 212 2174 228
rect 2098 194 2119 212
rect 1975 178 2018 194
rect 1898 140 2018 178
rect 2076 178 2119 194
rect 2153 194 2174 212
rect 2276 212 2352 228
rect 2276 194 2297 212
rect 2153 178 2196 194
rect 2076 140 2196 178
rect 2254 178 2297 194
rect 2331 194 2352 212
rect 2454 212 2530 228
rect 2454 194 2475 212
rect 2331 178 2374 194
rect 2254 140 2374 178
rect 2432 178 2475 194
rect 2509 194 2530 212
rect 2632 212 2708 228
rect 2632 194 2653 212
rect 2509 178 2552 194
rect 2432 140 2552 178
rect 2610 178 2653 194
rect 2687 194 2708 212
rect 2810 212 2886 228
rect 2810 194 2831 212
rect 2687 178 2730 194
rect 2610 140 2730 178
rect 2788 178 2831 194
rect 2865 194 2886 212
rect 2988 212 3064 228
rect 2988 194 3009 212
rect 2865 178 2908 194
rect 2788 140 2908 178
rect 2966 178 3009 194
rect 3043 194 3064 212
rect 3043 178 3086 194
rect 2966 140 3086 178
rect -3086 -178 -2966 -140
rect -3086 -194 -3043 -178
rect -3064 -212 -3043 -194
rect -3009 -194 -2966 -178
rect -2908 -178 -2788 -140
rect -2908 -194 -2865 -178
rect -3009 -212 -2988 -194
rect -3064 -228 -2988 -212
rect -2886 -212 -2865 -194
rect -2831 -194 -2788 -178
rect -2730 -178 -2610 -140
rect -2730 -194 -2687 -178
rect -2831 -212 -2810 -194
rect -2886 -228 -2810 -212
rect -2708 -212 -2687 -194
rect -2653 -194 -2610 -178
rect -2552 -178 -2432 -140
rect -2552 -194 -2509 -178
rect -2653 -212 -2632 -194
rect -2708 -228 -2632 -212
rect -2530 -212 -2509 -194
rect -2475 -194 -2432 -178
rect -2374 -178 -2254 -140
rect -2374 -194 -2331 -178
rect -2475 -212 -2454 -194
rect -2530 -228 -2454 -212
rect -2352 -212 -2331 -194
rect -2297 -194 -2254 -178
rect -2196 -178 -2076 -140
rect -2196 -194 -2153 -178
rect -2297 -212 -2276 -194
rect -2352 -228 -2276 -212
rect -2174 -212 -2153 -194
rect -2119 -194 -2076 -178
rect -2018 -178 -1898 -140
rect -2018 -194 -1975 -178
rect -2119 -212 -2098 -194
rect -2174 -228 -2098 -212
rect -1996 -212 -1975 -194
rect -1941 -194 -1898 -178
rect -1840 -178 -1720 -140
rect -1840 -194 -1797 -178
rect -1941 -212 -1920 -194
rect -1996 -228 -1920 -212
rect -1818 -212 -1797 -194
rect -1763 -194 -1720 -178
rect -1662 -178 -1542 -140
rect -1662 -194 -1619 -178
rect -1763 -212 -1742 -194
rect -1818 -228 -1742 -212
rect -1640 -212 -1619 -194
rect -1585 -194 -1542 -178
rect -1484 -178 -1364 -140
rect -1484 -194 -1441 -178
rect -1585 -212 -1564 -194
rect -1640 -228 -1564 -212
rect -1462 -212 -1441 -194
rect -1407 -194 -1364 -178
rect -1306 -178 -1186 -140
rect -1306 -194 -1263 -178
rect -1407 -212 -1386 -194
rect -1462 -228 -1386 -212
rect -1284 -212 -1263 -194
rect -1229 -194 -1186 -178
rect -1128 -178 -1008 -140
rect -1128 -194 -1085 -178
rect -1229 -212 -1208 -194
rect -1284 -228 -1208 -212
rect -1106 -212 -1085 -194
rect -1051 -194 -1008 -178
rect -950 -178 -830 -140
rect -950 -194 -907 -178
rect -1051 -212 -1030 -194
rect -1106 -228 -1030 -212
rect -928 -212 -907 -194
rect -873 -194 -830 -178
rect -772 -178 -652 -140
rect -772 -194 -729 -178
rect -873 -212 -852 -194
rect -928 -228 -852 -212
rect -750 -212 -729 -194
rect -695 -194 -652 -178
rect -594 -178 -474 -140
rect -594 -194 -551 -178
rect -695 -212 -674 -194
rect -750 -228 -674 -212
rect -572 -212 -551 -194
rect -517 -194 -474 -178
rect -416 -178 -296 -140
rect -416 -194 -373 -178
rect -517 -212 -496 -194
rect -572 -228 -496 -212
rect -394 -212 -373 -194
rect -339 -194 -296 -178
rect -238 -178 -118 -140
rect -238 -194 -195 -178
rect -339 -212 -318 -194
rect -394 -228 -318 -212
rect -216 -212 -195 -194
rect -161 -194 -118 -178
rect -60 -178 60 -140
rect -60 -194 -17 -178
rect -161 -212 -140 -194
rect -216 -228 -140 -212
rect -38 -212 -17 -194
rect 17 -194 60 -178
rect 118 -178 238 -140
rect 118 -194 161 -178
rect 17 -212 38 -194
rect -38 -228 38 -212
rect 140 -212 161 -194
rect 195 -194 238 -178
rect 296 -178 416 -140
rect 296 -194 339 -178
rect 195 -212 216 -194
rect 140 -228 216 -212
rect 318 -212 339 -194
rect 373 -194 416 -178
rect 474 -178 594 -140
rect 474 -194 517 -178
rect 373 -212 394 -194
rect 318 -228 394 -212
rect 496 -212 517 -194
rect 551 -194 594 -178
rect 652 -178 772 -140
rect 652 -194 695 -178
rect 551 -212 572 -194
rect 496 -228 572 -212
rect 674 -212 695 -194
rect 729 -194 772 -178
rect 830 -178 950 -140
rect 830 -194 873 -178
rect 729 -212 750 -194
rect 674 -228 750 -212
rect 852 -212 873 -194
rect 907 -194 950 -178
rect 1008 -178 1128 -140
rect 1008 -194 1051 -178
rect 907 -212 928 -194
rect 852 -228 928 -212
rect 1030 -212 1051 -194
rect 1085 -194 1128 -178
rect 1186 -178 1306 -140
rect 1186 -194 1229 -178
rect 1085 -212 1106 -194
rect 1030 -228 1106 -212
rect 1208 -212 1229 -194
rect 1263 -194 1306 -178
rect 1364 -178 1484 -140
rect 1364 -194 1407 -178
rect 1263 -212 1284 -194
rect 1208 -228 1284 -212
rect 1386 -212 1407 -194
rect 1441 -194 1484 -178
rect 1542 -178 1662 -140
rect 1542 -194 1585 -178
rect 1441 -212 1462 -194
rect 1386 -228 1462 -212
rect 1564 -212 1585 -194
rect 1619 -194 1662 -178
rect 1720 -178 1840 -140
rect 1720 -194 1763 -178
rect 1619 -212 1640 -194
rect 1564 -228 1640 -212
rect 1742 -212 1763 -194
rect 1797 -194 1840 -178
rect 1898 -178 2018 -140
rect 1898 -194 1941 -178
rect 1797 -212 1818 -194
rect 1742 -228 1818 -212
rect 1920 -212 1941 -194
rect 1975 -194 2018 -178
rect 2076 -178 2196 -140
rect 2076 -194 2119 -178
rect 1975 -212 1996 -194
rect 1920 -228 1996 -212
rect 2098 -212 2119 -194
rect 2153 -194 2196 -178
rect 2254 -178 2374 -140
rect 2254 -194 2297 -178
rect 2153 -212 2174 -194
rect 2098 -228 2174 -212
rect 2276 -212 2297 -194
rect 2331 -194 2374 -178
rect 2432 -178 2552 -140
rect 2432 -194 2475 -178
rect 2331 -212 2352 -194
rect 2276 -228 2352 -212
rect 2454 -212 2475 -194
rect 2509 -194 2552 -178
rect 2610 -178 2730 -140
rect 2610 -194 2653 -178
rect 2509 -212 2530 -194
rect 2454 -228 2530 -212
rect 2632 -212 2653 -194
rect 2687 -194 2730 -178
rect 2788 -178 2908 -140
rect 2788 -194 2831 -178
rect 2687 -212 2708 -194
rect 2632 -228 2708 -212
rect 2810 -212 2831 -194
rect 2865 -194 2908 -178
rect 2966 -178 3086 -140
rect 2966 -194 3009 -178
rect 2865 -212 2886 -194
rect 2810 -228 2886 -212
rect 2988 -212 3009 -194
rect 3043 -194 3086 -178
rect 3043 -212 3064 -194
rect 2988 -228 3064 -212
<< polycont >>
rect -3043 178 -3009 212
rect -2865 178 -2831 212
rect -2687 178 -2653 212
rect -2509 178 -2475 212
rect -2331 178 -2297 212
rect -2153 178 -2119 212
rect -1975 178 -1941 212
rect -1797 178 -1763 212
rect -1619 178 -1585 212
rect -1441 178 -1407 212
rect -1263 178 -1229 212
rect -1085 178 -1051 212
rect -907 178 -873 212
rect -729 178 -695 212
rect -551 178 -517 212
rect -373 178 -339 212
rect -195 178 -161 212
rect -17 178 17 212
rect 161 178 195 212
rect 339 178 373 212
rect 517 178 551 212
rect 695 178 729 212
rect 873 178 907 212
rect 1051 178 1085 212
rect 1229 178 1263 212
rect 1407 178 1441 212
rect 1585 178 1619 212
rect 1763 178 1797 212
rect 1941 178 1975 212
rect 2119 178 2153 212
rect 2297 178 2331 212
rect 2475 178 2509 212
rect 2653 178 2687 212
rect 2831 178 2865 212
rect 3009 178 3043 212
rect -3043 -212 -3009 -178
rect -2865 -212 -2831 -178
rect -2687 -212 -2653 -178
rect -2509 -212 -2475 -178
rect -2331 -212 -2297 -178
rect -2153 -212 -2119 -178
rect -1975 -212 -1941 -178
rect -1797 -212 -1763 -178
rect -1619 -212 -1585 -178
rect -1441 -212 -1407 -178
rect -1263 -212 -1229 -178
rect -1085 -212 -1051 -178
rect -907 -212 -873 -178
rect -729 -212 -695 -178
rect -551 -212 -517 -178
rect -373 -212 -339 -178
rect -195 -212 -161 -178
rect -17 -212 17 -178
rect 161 -212 195 -178
rect 339 -212 373 -178
rect 517 -212 551 -178
rect 695 -212 729 -178
rect 873 -212 907 -178
rect 1051 -212 1085 -178
rect 1229 -212 1263 -178
rect 1407 -212 1441 -178
rect 1585 -212 1619 -178
rect 1763 -212 1797 -178
rect 1941 -212 1975 -178
rect 2119 -212 2153 -178
rect 2297 -212 2331 -178
rect 2475 -212 2509 -178
rect 2653 -212 2687 -178
rect 2831 -212 2865 -178
rect 3009 -212 3043 -178
<< locali >>
rect -3064 178 -3043 212
rect -3009 178 -2988 212
rect -2886 178 -2865 212
rect -2831 178 -2810 212
rect -2708 178 -2687 212
rect -2653 178 -2632 212
rect -2530 178 -2509 212
rect -2475 178 -2454 212
rect -2352 178 -2331 212
rect -2297 178 -2276 212
rect -2174 178 -2153 212
rect -2119 178 -2098 212
rect -1996 178 -1975 212
rect -1941 178 -1920 212
rect -1818 178 -1797 212
rect -1763 178 -1742 212
rect -1640 178 -1619 212
rect -1585 178 -1564 212
rect -1462 178 -1441 212
rect -1407 178 -1386 212
rect -1284 178 -1263 212
rect -1229 178 -1208 212
rect -1106 178 -1085 212
rect -1051 178 -1030 212
rect -928 178 -907 212
rect -873 178 -852 212
rect -750 178 -729 212
rect -695 178 -674 212
rect -572 178 -551 212
rect -517 178 -496 212
rect -394 178 -373 212
rect -339 178 -318 212
rect -216 178 -195 212
rect -161 178 -140 212
rect -38 178 -17 212
rect 17 178 38 212
rect 140 178 161 212
rect 195 178 216 212
rect 318 178 339 212
rect 373 178 394 212
rect 496 178 517 212
rect 551 178 572 212
rect 674 178 695 212
rect 729 178 750 212
rect 852 178 873 212
rect 907 178 928 212
rect 1030 178 1051 212
rect 1085 178 1106 212
rect 1208 178 1229 212
rect 1263 178 1284 212
rect 1386 178 1407 212
rect 1441 178 1462 212
rect 1564 178 1585 212
rect 1619 178 1640 212
rect 1742 178 1763 212
rect 1797 178 1818 212
rect 1920 178 1941 212
rect 1975 178 1996 212
rect 2098 178 2119 212
rect 2153 178 2174 212
rect 2276 178 2297 212
rect 2331 178 2352 212
rect 2454 178 2475 212
rect 2509 178 2530 212
rect 2632 178 2653 212
rect 2687 178 2708 212
rect 2810 178 2831 212
rect 2865 178 2886 212
rect 2988 178 3009 212
rect 3043 178 3064 212
rect -3132 125 -3098 144
rect -3132 53 -3098 85
rect -3132 -17 -3098 17
rect -3132 -85 -3098 -53
rect -3132 -144 -3098 -125
rect -2954 125 -2920 144
rect -2954 53 -2920 85
rect -2954 -17 -2920 17
rect -2954 -85 -2920 -53
rect -2954 -144 -2920 -125
rect -2776 125 -2742 144
rect -2776 53 -2742 85
rect -2776 -17 -2742 17
rect -2776 -85 -2742 -53
rect -2776 -144 -2742 -125
rect -2598 125 -2564 144
rect -2598 53 -2564 85
rect -2598 -17 -2564 17
rect -2598 -85 -2564 -53
rect -2598 -144 -2564 -125
rect -2420 125 -2386 144
rect -2420 53 -2386 85
rect -2420 -17 -2386 17
rect -2420 -85 -2386 -53
rect -2420 -144 -2386 -125
rect -2242 125 -2208 144
rect -2242 53 -2208 85
rect -2242 -17 -2208 17
rect -2242 -85 -2208 -53
rect -2242 -144 -2208 -125
rect -2064 125 -2030 144
rect -2064 53 -2030 85
rect -2064 -17 -2030 17
rect -2064 -85 -2030 -53
rect -2064 -144 -2030 -125
rect -1886 125 -1852 144
rect -1886 53 -1852 85
rect -1886 -17 -1852 17
rect -1886 -85 -1852 -53
rect -1886 -144 -1852 -125
rect -1708 125 -1674 144
rect -1708 53 -1674 85
rect -1708 -17 -1674 17
rect -1708 -85 -1674 -53
rect -1708 -144 -1674 -125
rect -1530 125 -1496 144
rect -1530 53 -1496 85
rect -1530 -17 -1496 17
rect -1530 -85 -1496 -53
rect -1530 -144 -1496 -125
rect -1352 125 -1318 144
rect -1352 53 -1318 85
rect -1352 -17 -1318 17
rect -1352 -85 -1318 -53
rect -1352 -144 -1318 -125
rect -1174 125 -1140 144
rect -1174 53 -1140 85
rect -1174 -17 -1140 17
rect -1174 -85 -1140 -53
rect -1174 -144 -1140 -125
rect -996 125 -962 144
rect -996 53 -962 85
rect -996 -17 -962 17
rect -996 -85 -962 -53
rect -996 -144 -962 -125
rect -818 125 -784 144
rect -818 53 -784 85
rect -818 -17 -784 17
rect -818 -85 -784 -53
rect -818 -144 -784 -125
rect -640 125 -606 144
rect -640 53 -606 85
rect -640 -17 -606 17
rect -640 -85 -606 -53
rect -640 -144 -606 -125
rect -462 125 -428 144
rect -462 53 -428 85
rect -462 -17 -428 17
rect -462 -85 -428 -53
rect -462 -144 -428 -125
rect -284 125 -250 144
rect -284 53 -250 85
rect -284 -17 -250 17
rect -284 -85 -250 -53
rect -284 -144 -250 -125
rect -106 125 -72 144
rect -106 53 -72 85
rect -106 -17 -72 17
rect -106 -85 -72 -53
rect -106 -144 -72 -125
rect 72 125 106 144
rect 72 53 106 85
rect 72 -17 106 17
rect 72 -85 106 -53
rect 72 -144 106 -125
rect 250 125 284 144
rect 250 53 284 85
rect 250 -17 284 17
rect 250 -85 284 -53
rect 250 -144 284 -125
rect 428 125 462 144
rect 428 53 462 85
rect 428 -17 462 17
rect 428 -85 462 -53
rect 428 -144 462 -125
rect 606 125 640 144
rect 606 53 640 85
rect 606 -17 640 17
rect 606 -85 640 -53
rect 606 -144 640 -125
rect 784 125 818 144
rect 784 53 818 85
rect 784 -17 818 17
rect 784 -85 818 -53
rect 784 -144 818 -125
rect 962 125 996 144
rect 962 53 996 85
rect 962 -17 996 17
rect 962 -85 996 -53
rect 962 -144 996 -125
rect 1140 125 1174 144
rect 1140 53 1174 85
rect 1140 -17 1174 17
rect 1140 -85 1174 -53
rect 1140 -144 1174 -125
rect 1318 125 1352 144
rect 1318 53 1352 85
rect 1318 -17 1352 17
rect 1318 -85 1352 -53
rect 1318 -144 1352 -125
rect 1496 125 1530 144
rect 1496 53 1530 85
rect 1496 -17 1530 17
rect 1496 -85 1530 -53
rect 1496 -144 1530 -125
rect 1674 125 1708 144
rect 1674 53 1708 85
rect 1674 -17 1708 17
rect 1674 -85 1708 -53
rect 1674 -144 1708 -125
rect 1852 125 1886 144
rect 1852 53 1886 85
rect 1852 -17 1886 17
rect 1852 -85 1886 -53
rect 1852 -144 1886 -125
rect 2030 125 2064 144
rect 2030 53 2064 85
rect 2030 -17 2064 17
rect 2030 -85 2064 -53
rect 2030 -144 2064 -125
rect 2208 125 2242 144
rect 2208 53 2242 85
rect 2208 -17 2242 17
rect 2208 -85 2242 -53
rect 2208 -144 2242 -125
rect 2386 125 2420 144
rect 2386 53 2420 85
rect 2386 -17 2420 17
rect 2386 -85 2420 -53
rect 2386 -144 2420 -125
rect 2564 125 2598 144
rect 2564 53 2598 85
rect 2564 -17 2598 17
rect 2564 -85 2598 -53
rect 2564 -144 2598 -125
rect 2742 125 2776 144
rect 2742 53 2776 85
rect 2742 -17 2776 17
rect 2742 -85 2776 -53
rect 2742 -144 2776 -125
rect 2920 125 2954 144
rect 2920 53 2954 85
rect 2920 -17 2954 17
rect 2920 -85 2954 -53
rect 2920 -144 2954 -125
rect 3098 125 3132 144
rect 3098 53 3132 85
rect 3098 -17 3132 17
rect 3098 -85 3132 -53
rect 3098 -144 3132 -125
rect -3064 -212 -3043 -178
rect -3009 -212 -2988 -178
rect -2886 -212 -2865 -178
rect -2831 -212 -2810 -178
rect -2708 -212 -2687 -178
rect -2653 -212 -2632 -178
rect -2530 -212 -2509 -178
rect -2475 -212 -2454 -178
rect -2352 -212 -2331 -178
rect -2297 -212 -2276 -178
rect -2174 -212 -2153 -178
rect -2119 -212 -2098 -178
rect -1996 -212 -1975 -178
rect -1941 -212 -1920 -178
rect -1818 -212 -1797 -178
rect -1763 -212 -1742 -178
rect -1640 -212 -1619 -178
rect -1585 -212 -1564 -178
rect -1462 -212 -1441 -178
rect -1407 -212 -1386 -178
rect -1284 -212 -1263 -178
rect -1229 -212 -1208 -178
rect -1106 -212 -1085 -178
rect -1051 -212 -1030 -178
rect -928 -212 -907 -178
rect -873 -212 -852 -178
rect -750 -212 -729 -178
rect -695 -212 -674 -178
rect -572 -212 -551 -178
rect -517 -212 -496 -178
rect -394 -212 -373 -178
rect -339 -212 -318 -178
rect -216 -212 -195 -178
rect -161 -212 -140 -178
rect -38 -212 -17 -178
rect 17 -212 38 -178
rect 140 -212 161 -178
rect 195 -212 216 -178
rect 318 -212 339 -178
rect 373 -212 394 -178
rect 496 -212 517 -178
rect 551 -212 572 -178
rect 674 -212 695 -178
rect 729 -212 750 -178
rect 852 -212 873 -178
rect 907 -212 928 -178
rect 1030 -212 1051 -178
rect 1085 -212 1106 -178
rect 1208 -212 1229 -178
rect 1263 -212 1284 -178
rect 1386 -212 1407 -178
rect 1441 -212 1462 -178
rect 1564 -212 1585 -178
rect 1619 -212 1640 -178
rect 1742 -212 1763 -178
rect 1797 -212 1818 -178
rect 1920 -212 1941 -178
rect 1975 -212 1996 -178
rect 2098 -212 2119 -178
rect 2153 -212 2174 -178
rect 2276 -212 2297 -178
rect 2331 -212 2352 -178
rect 2454 -212 2475 -178
rect 2509 -212 2530 -178
rect 2632 -212 2653 -178
rect 2687 -212 2708 -178
rect 2810 -212 2831 -178
rect 2865 -212 2886 -178
rect 2988 -212 3009 -178
rect 3043 -212 3064 -178
<< viali >>
rect -3043 178 -3009 212
rect -2865 178 -2831 212
rect -2687 178 -2653 212
rect -2509 178 -2475 212
rect -2331 178 -2297 212
rect -2153 178 -2119 212
rect -1975 178 -1941 212
rect -1797 178 -1763 212
rect -1619 178 -1585 212
rect -1441 178 -1407 212
rect -1263 178 -1229 212
rect -1085 178 -1051 212
rect -907 178 -873 212
rect -729 178 -695 212
rect -551 178 -517 212
rect -373 178 -339 212
rect -195 178 -161 212
rect -17 178 17 212
rect 161 178 195 212
rect 339 178 373 212
rect 517 178 551 212
rect 695 178 729 212
rect 873 178 907 212
rect 1051 178 1085 212
rect 1229 178 1263 212
rect 1407 178 1441 212
rect 1585 178 1619 212
rect 1763 178 1797 212
rect 1941 178 1975 212
rect 2119 178 2153 212
rect 2297 178 2331 212
rect 2475 178 2509 212
rect 2653 178 2687 212
rect 2831 178 2865 212
rect 3009 178 3043 212
rect -3132 119 -3098 125
rect -3132 91 -3098 119
rect -3132 51 -3098 53
rect -3132 19 -3098 51
rect -3132 -51 -3098 -19
rect -3132 -53 -3098 -51
rect -3132 -119 -3098 -91
rect -3132 -125 -3098 -119
rect -2954 119 -2920 125
rect -2954 91 -2920 119
rect -2954 51 -2920 53
rect -2954 19 -2920 51
rect -2954 -51 -2920 -19
rect -2954 -53 -2920 -51
rect -2954 -119 -2920 -91
rect -2954 -125 -2920 -119
rect -2776 119 -2742 125
rect -2776 91 -2742 119
rect -2776 51 -2742 53
rect -2776 19 -2742 51
rect -2776 -51 -2742 -19
rect -2776 -53 -2742 -51
rect -2776 -119 -2742 -91
rect -2776 -125 -2742 -119
rect -2598 119 -2564 125
rect -2598 91 -2564 119
rect -2598 51 -2564 53
rect -2598 19 -2564 51
rect -2598 -51 -2564 -19
rect -2598 -53 -2564 -51
rect -2598 -119 -2564 -91
rect -2598 -125 -2564 -119
rect -2420 119 -2386 125
rect -2420 91 -2386 119
rect -2420 51 -2386 53
rect -2420 19 -2386 51
rect -2420 -51 -2386 -19
rect -2420 -53 -2386 -51
rect -2420 -119 -2386 -91
rect -2420 -125 -2386 -119
rect -2242 119 -2208 125
rect -2242 91 -2208 119
rect -2242 51 -2208 53
rect -2242 19 -2208 51
rect -2242 -51 -2208 -19
rect -2242 -53 -2208 -51
rect -2242 -119 -2208 -91
rect -2242 -125 -2208 -119
rect -2064 119 -2030 125
rect -2064 91 -2030 119
rect -2064 51 -2030 53
rect -2064 19 -2030 51
rect -2064 -51 -2030 -19
rect -2064 -53 -2030 -51
rect -2064 -119 -2030 -91
rect -2064 -125 -2030 -119
rect -1886 119 -1852 125
rect -1886 91 -1852 119
rect -1886 51 -1852 53
rect -1886 19 -1852 51
rect -1886 -51 -1852 -19
rect -1886 -53 -1852 -51
rect -1886 -119 -1852 -91
rect -1886 -125 -1852 -119
rect -1708 119 -1674 125
rect -1708 91 -1674 119
rect -1708 51 -1674 53
rect -1708 19 -1674 51
rect -1708 -51 -1674 -19
rect -1708 -53 -1674 -51
rect -1708 -119 -1674 -91
rect -1708 -125 -1674 -119
rect -1530 119 -1496 125
rect -1530 91 -1496 119
rect -1530 51 -1496 53
rect -1530 19 -1496 51
rect -1530 -51 -1496 -19
rect -1530 -53 -1496 -51
rect -1530 -119 -1496 -91
rect -1530 -125 -1496 -119
rect -1352 119 -1318 125
rect -1352 91 -1318 119
rect -1352 51 -1318 53
rect -1352 19 -1318 51
rect -1352 -51 -1318 -19
rect -1352 -53 -1318 -51
rect -1352 -119 -1318 -91
rect -1352 -125 -1318 -119
rect -1174 119 -1140 125
rect -1174 91 -1140 119
rect -1174 51 -1140 53
rect -1174 19 -1140 51
rect -1174 -51 -1140 -19
rect -1174 -53 -1140 -51
rect -1174 -119 -1140 -91
rect -1174 -125 -1140 -119
rect -996 119 -962 125
rect -996 91 -962 119
rect -996 51 -962 53
rect -996 19 -962 51
rect -996 -51 -962 -19
rect -996 -53 -962 -51
rect -996 -119 -962 -91
rect -996 -125 -962 -119
rect -818 119 -784 125
rect -818 91 -784 119
rect -818 51 -784 53
rect -818 19 -784 51
rect -818 -51 -784 -19
rect -818 -53 -784 -51
rect -818 -119 -784 -91
rect -818 -125 -784 -119
rect -640 119 -606 125
rect -640 91 -606 119
rect -640 51 -606 53
rect -640 19 -606 51
rect -640 -51 -606 -19
rect -640 -53 -606 -51
rect -640 -119 -606 -91
rect -640 -125 -606 -119
rect -462 119 -428 125
rect -462 91 -428 119
rect -462 51 -428 53
rect -462 19 -428 51
rect -462 -51 -428 -19
rect -462 -53 -428 -51
rect -462 -119 -428 -91
rect -462 -125 -428 -119
rect -284 119 -250 125
rect -284 91 -250 119
rect -284 51 -250 53
rect -284 19 -250 51
rect -284 -51 -250 -19
rect -284 -53 -250 -51
rect -284 -119 -250 -91
rect -284 -125 -250 -119
rect -106 119 -72 125
rect -106 91 -72 119
rect -106 51 -72 53
rect -106 19 -72 51
rect -106 -51 -72 -19
rect -106 -53 -72 -51
rect -106 -119 -72 -91
rect -106 -125 -72 -119
rect 72 119 106 125
rect 72 91 106 119
rect 72 51 106 53
rect 72 19 106 51
rect 72 -51 106 -19
rect 72 -53 106 -51
rect 72 -119 106 -91
rect 72 -125 106 -119
rect 250 119 284 125
rect 250 91 284 119
rect 250 51 284 53
rect 250 19 284 51
rect 250 -51 284 -19
rect 250 -53 284 -51
rect 250 -119 284 -91
rect 250 -125 284 -119
rect 428 119 462 125
rect 428 91 462 119
rect 428 51 462 53
rect 428 19 462 51
rect 428 -51 462 -19
rect 428 -53 462 -51
rect 428 -119 462 -91
rect 428 -125 462 -119
rect 606 119 640 125
rect 606 91 640 119
rect 606 51 640 53
rect 606 19 640 51
rect 606 -51 640 -19
rect 606 -53 640 -51
rect 606 -119 640 -91
rect 606 -125 640 -119
rect 784 119 818 125
rect 784 91 818 119
rect 784 51 818 53
rect 784 19 818 51
rect 784 -51 818 -19
rect 784 -53 818 -51
rect 784 -119 818 -91
rect 784 -125 818 -119
rect 962 119 996 125
rect 962 91 996 119
rect 962 51 996 53
rect 962 19 996 51
rect 962 -51 996 -19
rect 962 -53 996 -51
rect 962 -119 996 -91
rect 962 -125 996 -119
rect 1140 119 1174 125
rect 1140 91 1174 119
rect 1140 51 1174 53
rect 1140 19 1174 51
rect 1140 -51 1174 -19
rect 1140 -53 1174 -51
rect 1140 -119 1174 -91
rect 1140 -125 1174 -119
rect 1318 119 1352 125
rect 1318 91 1352 119
rect 1318 51 1352 53
rect 1318 19 1352 51
rect 1318 -51 1352 -19
rect 1318 -53 1352 -51
rect 1318 -119 1352 -91
rect 1318 -125 1352 -119
rect 1496 119 1530 125
rect 1496 91 1530 119
rect 1496 51 1530 53
rect 1496 19 1530 51
rect 1496 -51 1530 -19
rect 1496 -53 1530 -51
rect 1496 -119 1530 -91
rect 1496 -125 1530 -119
rect 1674 119 1708 125
rect 1674 91 1708 119
rect 1674 51 1708 53
rect 1674 19 1708 51
rect 1674 -51 1708 -19
rect 1674 -53 1708 -51
rect 1674 -119 1708 -91
rect 1674 -125 1708 -119
rect 1852 119 1886 125
rect 1852 91 1886 119
rect 1852 51 1886 53
rect 1852 19 1886 51
rect 1852 -51 1886 -19
rect 1852 -53 1886 -51
rect 1852 -119 1886 -91
rect 1852 -125 1886 -119
rect 2030 119 2064 125
rect 2030 91 2064 119
rect 2030 51 2064 53
rect 2030 19 2064 51
rect 2030 -51 2064 -19
rect 2030 -53 2064 -51
rect 2030 -119 2064 -91
rect 2030 -125 2064 -119
rect 2208 119 2242 125
rect 2208 91 2242 119
rect 2208 51 2242 53
rect 2208 19 2242 51
rect 2208 -51 2242 -19
rect 2208 -53 2242 -51
rect 2208 -119 2242 -91
rect 2208 -125 2242 -119
rect 2386 119 2420 125
rect 2386 91 2420 119
rect 2386 51 2420 53
rect 2386 19 2420 51
rect 2386 -51 2420 -19
rect 2386 -53 2420 -51
rect 2386 -119 2420 -91
rect 2386 -125 2420 -119
rect 2564 119 2598 125
rect 2564 91 2598 119
rect 2564 51 2598 53
rect 2564 19 2598 51
rect 2564 -51 2598 -19
rect 2564 -53 2598 -51
rect 2564 -119 2598 -91
rect 2564 -125 2598 -119
rect 2742 119 2776 125
rect 2742 91 2776 119
rect 2742 51 2776 53
rect 2742 19 2776 51
rect 2742 -51 2776 -19
rect 2742 -53 2776 -51
rect 2742 -119 2776 -91
rect 2742 -125 2776 -119
rect 2920 119 2954 125
rect 2920 91 2954 119
rect 2920 51 2954 53
rect 2920 19 2954 51
rect 2920 -51 2954 -19
rect 2920 -53 2954 -51
rect 2920 -119 2954 -91
rect 2920 -125 2954 -119
rect 3098 119 3132 125
rect 3098 91 3132 119
rect 3098 51 3132 53
rect 3098 19 3132 51
rect 3098 -51 3132 -19
rect 3098 -53 3132 -51
rect 3098 -119 3132 -91
rect 3098 -125 3132 -119
rect -3043 -212 -3009 -178
rect -2865 -212 -2831 -178
rect -2687 -212 -2653 -178
rect -2509 -212 -2475 -178
rect -2331 -212 -2297 -178
rect -2153 -212 -2119 -178
rect -1975 -212 -1941 -178
rect -1797 -212 -1763 -178
rect -1619 -212 -1585 -178
rect -1441 -212 -1407 -178
rect -1263 -212 -1229 -178
rect -1085 -212 -1051 -178
rect -907 -212 -873 -178
rect -729 -212 -695 -178
rect -551 -212 -517 -178
rect -373 -212 -339 -178
rect -195 -212 -161 -178
rect -17 -212 17 -178
rect 161 -212 195 -178
rect 339 -212 373 -178
rect 517 -212 551 -178
rect 695 -212 729 -178
rect 873 -212 907 -178
rect 1051 -212 1085 -178
rect 1229 -212 1263 -178
rect 1407 -212 1441 -178
rect 1585 -212 1619 -178
rect 1763 -212 1797 -178
rect 1941 -212 1975 -178
rect 2119 -212 2153 -178
rect 2297 -212 2331 -178
rect 2475 -212 2509 -178
rect 2653 -212 2687 -178
rect 2831 -212 2865 -178
rect 3009 -212 3043 -178
<< metal1 >>
rect -3064 212 -2988 228
rect -3064 178 -3043 212
rect -3009 178 -2988 212
rect -3064 172 -2988 178
rect -2886 212 -2810 228
rect -2886 178 -2865 212
rect -2831 178 -2810 212
rect -2886 172 -2810 178
rect -2708 212 -2632 228
rect -2708 178 -2687 212
rect -2653 178 -2632 212
rect -2708 172 -2632 178
rect -2530 212 -2454 228
rect -2530 178 -2509 212
rect -2475 178 -2454 212
rect -2530 172 -2454 178
rect -2352 212 -2276 228
rect -2352 178 -2331 212
rect -2297 178 -2276 212
rect -2352 172 -2276 178
rect -2174 212 -2098 228
rect -2174 178 -2153 212
rect -2119 178 -2098 212
rect -2174 172 -2098 178
rect -1996 212 -1920 228
rect -1996 178 -1975 212
rect -1941 178 -1920 212
rect -1996 172 -1920 178
rect -1818 212 -1742 228
rect -1818 178 -1797 212
rect -1763 178 -1742 212
rect -1818 172 -1742 178
rect -1640 212 -1564 228
rect -1640 178 -1619 212
rect -1585 178 -1564 212
rect -1640 172 -1564 178
rect -1462 212 -1386 228
rect -1462 178 -1441 212
rect -1407 178 -1386 212
rect -1462 172 -1386 178
rect -1284 212 -1208 228
rect -1284 178 -1263 212
rect -1229 178 -1208 212
rect -1284 172 -1208 178
rect -1106 212 -1030 228
rect -1106 178 -1085 212
rect -1051 178 -1030 212
rect -1106 172 -1030 178
rect -928 212 -852 228
rect -928 178 -907 212
rect -873 178 -852 212
rect -928 172 -852 178
rect -750 212 -674 228
rect -750 178 -729 212
rect -695 178 -674 212
rect -750 172 -674 178
rect -572 212 -496 228
rect -572 178 -551 212
rect -517 178 -496 212
rect -572 172 -496 178
rect -394 212 -318 228
rect -394 178 -373 212
rect -339 178 -318 212
rect -394 172 -318 178
rect -216 212 -140 228
rect -216 178 -195 212
rect -161 178 -140 212
rect -216 172 -140 178
rect -38 212 38 228
rect -38 178 -17 212
rect 17 178 38 212
rect -38 172 38 178
rect 140 212 216 228
rect 140 178 161 212
rect 195 178 216 212
rect 140 172 216 178
rect 318 212 394 228
rect 318 178 339 212
rect 373 178 394 212
rect 318 172 394 178
rect 496 212 572 228
rect 496 178 517 212
rect 551 178 572 212
rect 496 172 572 178
rect 674 212 750 228
rect 674 178 695 212
rect 729 178 750 212
rect 674 172 750 178
rect 852 212 928 228
rect 852 178 873 212
rect 907 178 928 212
rect 852 172 928 178
rect 1030 212 1106 228
rect 1030 178 1051 212
rect 1085 178 1106 212
rect 1030 172 1106 178
rect 1208 212 1284 228
rect 1208 178 1229 212
rect 1263 178 1284 212
rect 1208 172 1284 178
rect 1386 212 1462 228
rect 1386 178 1407 212
rect 1441 178 1462 212
rect 1386 172 1462 178
rect 1564 212 1640 228
rect 1564 178 1585 212
rect 1619 178 1640 212
rect 1564 172 1640 178
rect 1742 212 1818 228
rect 1742 178 1763 212
rect 1797 178 1818 212
rect 1742 172 1818 178
rect 1920 212 1996 228
rect 1920 178 1941 212
rect 1975 178 1996 212
rect 1920 172 1996 178
rect 2098 212 2174 228
rect 2098 178 2119 212
rect 2153 178 2174 212
rect 2098 172 2174 178
rect 2276 212 2352 228
rect 2276 178 2297 212
rect 2331 178 2352 212
rect 2276 172 2352 178
rect 2454 212 2530 228
rect 2454 178 2475 212
rect 2509 178 2530 212
rect 2454 172 2530 178
rect 2632 212 2708 228
rect 2632 178 2653 212
rect 2687 178 2708 212
rect 2632 172 2708 178
rect 2810 212 2886 228
rect 2810 178 2831 212
rect 2865 178 2886 212
rect 2810 172 2886 178
rect 2988 212 3064 228
rect 2988 178 3009 212
rect 3043 178 3064 212
rect 2988 172 3064 178
rect -3138 125 -3092 140
rect -3138 91 -3132 125
rect -3098 91 -3092 125
rect -3138 53 -3092 91
rect -3138 19 -3132 53
rect -3098 19 -3092 53
rect -3138 -19 -3092 19
rect -3138 -53 -3132 -19
rect -3098 -53 -3092 -19
rect -3138 -91 -3092 -53
rect -3138 -125 -3132 -91
rect -3098 -125 -3092 -91
rect -3138 -140 -3092 -125
rect -2960 125 -2914 140
rect -2960 91 -2954 125
rect -2920 91 -2914 125
rect -2960 53 -2914 91
rect -2960 19 -2954 53
rect -2920 19 -2914 53
rect -2960 -19 -2914 19
rect -2960 -53 -2954 -19
rect -2920 -53 -2914 -19
rect -2960 -91 -2914 -53
rect -2960 -125 -2954 -91
rect -2920 -125 -2914 -91
rect -2960 -140 -2914 -125
rect -2782 125 -2736 140
rect -2782 91 -2776 125
rect -2742 91 -2736 125
rect -2782 53 -2736 91
rect -2782 19 -2776 53
rect -2742 19 -2736 53
rect -2782 -19 -2736 19
rect -2782 -53 -2776 -19
rect -2742 -53 -2736 -19
rect -2782 -91 -2736 -53
rect -2782 -125 -2776 -91
rect -2742 -125 -2736 -91
rect -2782 -140 -2736 -125
rect -2604 125 -2558 140
rect -2604 91 -2598 125
rect -2564 91 -2558 125
rect -2604 53 -2558 91
rect -2604 19 -2598 53
rect -2564 19 -2558 53
rect -2604 -19 -2558 19
rect -2604 -53 -2598 -19
rect -2564 -53 -2558 -19
rect -2604 -91 -2558 -53
rect -2604 -125 -2598 -91
rect -2564 -125 -2558 -91
rect -2604 -140 -2558 -125
rect -2426 125 -2380 140
rect -2426 91 -2420 125
rect -2386 91 -2380 125
rect -2426 53 -2380 91
rect -2426 19 -2420 53
rect -2386 19 -2380 53
rect -2426 -19 -2380 19
rect -2426 -53 -2420 -19
rect -2386 -53 -2380 -19
rect -2426 -91 -2380 -53
rect -2426 -125 -2420 -91
rect -2386 -125 -2380 -91
rect -2426 -140 -2380 -125
rect -2248 125 -2202 140
rect -2248 91 -2242 125
rect -2208 91 -2202 125
rect -2248 53 -2202 91
rect -2248 19 -2242 53
rect -2208 19 -2202 53
rect -2248 -19 -2202 19
rect -2248 -53 -2242 -19
rect -2208 -53 -2202 -19
rect -2248 -91 -2202 -53
rect -2248 -125 -2242 -91
rect -2208 -125 -2202 -91
rect -2248 -140 -2202 -125
rect -2070 125 -2024 140
rect -2070 91 -2064 125
rect -2030 91 -2024 125
rect -2070 53 -2024 91
rect -2070 19 -2064 53
rect -2030 19 -2024 53
rect -2070 -19 -2024 19
rect -2070 -53 -2064 -19
rect -2030 -53 -2024 -19
rect -2070 -91 -2024 -53
rect -2070 -125 -2064 -91
rect -2030 -125 -2024 -91
rect -2070 -140 -2024 -125
rect -1892 125 -1846 140
rect -1892 91 -1886 125
rect -1852 91 -1846 125
rect -1892 53 -1846 91
rect -1892 19 -1886 53
rect -1852 19 -1846 53
rect -1892 -19 -1846 19
rect -1892 -53 -1886 -19
rect -1852 -53 -1846 -19
rect -1892 -91 -1846 -53
rect -1892 -125 -1886 -91
rect -1852 -125 -1846 -91
rect -1892 -140 -1846 -125
rect -1714 125 -1668 140
rect -1714 91 -1708 125
rect -1674 91 -1668 125
rect -1714 53 -1668 91
rect -1714 19 -1708 53
rect -1674 19 -1668 53
rect -1714 -19 -1668 19
rect -1714 -53 -1708 -19
rect -1674 -53 -1668 -19
rect -1714 -91 -1668 -53
rect -1714 -125 -1708 -91
rect -1674 -125 -1668 -91
rect -1714 -140 -1668 -125
rect -1536 125 -1490 140
rect -1536 91 -1530 125
rect -1496 91 -1490 125
rect -1536 53 -1490 91
rect -1536 19 -1530 53
rect -1496 19 -1490 53
rect -1536 -19 -1490 19
rect -1536 -53 -1530 -19
rect -1496 -53 -1490 -19
rect -1536 -91 -1490 -53
rect -1536 -125 -1530 -91
rect -1496 -125 -1490 -91
rect -1536 -140 -1490 -125
rect -1358 125 -1312 140
rect -1358 91 -1352 125
rect -1318 91 -1312 125
rect -1358 53 -1312 91
rect -1358 19 -1352 53
rect -1318 19 -1312 53
rect -1358 -19 -1312 19
rect -1358 -53 -1352 -19
rect -1318 -53 -1312 -19
rect -1358 -91 -1312 -53
rect -1358 -125 -1352 -91
rect -1318 -125 -1312 -91
rect -1358 -140 -1312 -125
rect -1180 125 -1134 140
rect -1180 91 -1174 125
rect -1140 91 -1134 125
rect -1180 53 -1134 91
rect -1180 19 -1174 53
rect -1140 19 -1134 53
rect -1180 -19 -1134 19
rect -1180 -53 -1174 -19
rect -1140 -53 -1134 -19
rect -1180 -91 -1134 -53
rect -1180 -125 -1174 -91
rect -1140 -125 -1134 -91
rect -1180 -140 -1134 -125
rect -1002 125 -956 140
rect -1002 91 -996 125
rect -962 91 -956 125
rect -1002 53 -956 91
rect -1002 19 -996 53
rect -962 19 -956 53
rect -1002 -19 -956 19
rect -1002 -53 -996 -19
rect -962 -53 -956 -19
rect -1002 -91 -956 -53
rect -1002 -125 -996 -91
rect -962 -125 -956 -91
rect -1002 -140 -956 -125
rect -824 125 -778 140
rect -824 91 -818 125
rect -784 91 -778 125
rect -824 53 -778 91
rect -824 19 -818 53
rect -784 19 -778 53
rect -824 -19 -778 19
rect -824 -53 -818 -19
rect -784 -53 -778 -19
rect -824 -91 -778 -53
rect -824 -125 -818 -91
rect -784 -125 -778 -91
rect -824 -140 -778 -125
rect -646 125 -600 140
rect -646 91 -640 125
rect -606 91 -600 125
rect -646 53 -600 91
rect -646 19 -640 53
rect -606 19 -600 53
rect -646 -19 -600 19
rect -646 -53 -640 -19
rect -606 -53 -600 -19
rect -646 -91 -600 -53
rect -646 -125 -640 -91
rect -606 -125 -600 -91
rect -646 -140 -600 -125
rect -468 125 -422 140
rect -468 91 -462 125
rect -428 91 -422 125
rect -468 53 -422 91
rect -468 19 -462 53
rect -428 19 -422 53
rect -468 -19 -422 19
rect -468 -53 -462 -19
rect -428 -53 -422 -19
rect -468 -91 -422 -53
rect -468 -125 -462 -91
rect -428 -125 -422 -91
rect -468 -140 -422 -125
rect -290 125 -244 140
rect -290 91 -284 125
rect -250 91 -244 125
rect -290 53 -244 91
rect -290 19 -284 53
rect -250 19 -244 53
rect -290 -19 -244 19
rect -290 -53 -284 -19
rect -250 -53 -244 -19
rect -290 -91 -244 -53
rect -290 -125 -284 -91
rect -250 -125 -244 -91
rect -290 -140 -244 -125
rect -112 125 -66 140
rect -112 91 -106 125
rect -72 91 -66 125
rect -112 53 -66 91
rect -112 19 -106 53
rect -72 19 -66 53
rect -112 -19 -66 19
rect -112 -53 -106 -19
rect -72 -53 -66 -19
rect -112 -91 -66 -53
rect -112 -125 -106 -91
rect -72 -125 -66 -91
rect -112 -140 -66 -125
rect 66 125 112 140
rect 66 91 72 125
rect 106 91 112 125
rect 66 53 112 91
rect 66 19 72 53
rect 106 19 112 53
rect 66 -19 112 19
rect 66 -53 72 -19
rect 106 -53 112 -19
rect 66 -91 112 -53
rect 66 -125 72 -91
rect 106 -125 112 -91
rect 66 -140 112 -125
rect 244 125 290 140
rect 244 91 250 125
rect 284 91 290 125
rect 244 53 290 91
rect 244 19 250 53
rect 284 19 290 53
rect 244 -19 290 19
rect 244 -53 250 -19
rect 284 -53 290 -19
rect 244 -91 290 -53
rect 244 -125 250 -91
rect 284 -125 290 -91
rect 244 -140 290 -125
rect 422 125 468 140
rect 422 91 428 125
rect 462 91 468 125
rect 422 53 468 91
rect 422 19 428 53
rect 462 19 468 53
rect 422 -19 468 19
rect 422 -53 428 -19
rect 462 -53 468 -19
rect 422 -91 468 -53
rect 422 -125 428 -91
rect 462 -125 468 -91
rect 422 -140 468 -125
rect 600 125 646 140
rect 600 91 606 125
rect 640 91 646 125
rect 600 53 646 91
rect 600 19 606 53
rect 640 19 646 53
rect 600 -19 646 19
rect 600 -53 606 -19
rect 640 -53 646 -19
rect 600 -91 646 -53
rect 600 -125 606 -91
rect 640 -125 646 -91
rect 600 -140 646 -125
rect 778 125 824 140
rect 778 91 784 125
rect 818 91 824 125
rect 778 53 824 91
rect 778 19 784 53
rect 818 19 824 53
rect 778 -19 824 19
rect 778 -53 784 -19
rect 818 -53 824 -19
rect 778 -91 824 -53
rect 778 -125 784 -91
rect 818 -125 824 -91
rect 778 -140 824 -125
rect 956 125 1002 140
rect 956 91 962 125
rect 996 91 1002 125
rect 956 53 1002 91
rect 956 19 962 53
rect 996 19 1002 53
rect 956 -19 1002 19
rect 956 -53 962 -19
rect 996 -53 1002 -19
rect 956 -91 1002 -53
rect 956 -125 962 -91
rect 996 -125 1002 -91
rect 956 -140 1002 -125
rect 1134 125 1180 140
rect 1134 91 1140 125
rect 1174 91 1180 125
rect 1134 53 1180 91
rect 1134 19 1140 53
rect 1174 19 1180 53
rect 1134 -19 1180 19
rect 1134 -53 1140 -19
rect 1174 -53 1180 -19
rect 1134 -91 1180 -53
rect 1134 -125 1140 -91
rect 1174 -125 1180 -91
rect 1134 -140 1180 -125
rect 1312 125 1358 140
rect 1312 91 1318 125
rect 1352 91 1358 125
rect 1312 53 1358 91
rect 1312 19 1318 53
rect 1352 19 1358 53
rect 1312 -19 1358 19
rect 1312 -53 1318 -19
rect 1352 -53 1358 -19
rect 1312 -91 1358 -53
rect 1312 -125 1318 -91
rect 1352 -125 1358 -91
rect 1312 -140 1358 -125
rect 1490 125 1536 140
rect 1490 91 1496 125
rect 1530 91 1536 125
rect 1490 53 1536 91
rect 1490 19 1496 53
rect 1530 19 1536 53
rect 1490 -19 1536 19
rect 1490 -53 1496 -19
rect 1530 -53 1536 -19
rect 1490 -91 1536 -53
rect 1490 -125 1496 -91
rect 1530 -125 1536 -91
rect 1490 -140 1536 -125
rect 1668 125 1714 140
rect 1668 91 1674 125
rect 1708 91 1714 125
rect 1668 53 1714 91
rect 1668 19 1674 53
rect 1708 19 1714 53
rect 1668 -19 1714 19
rect 1668 -53 1674 -19
rect 1708 -53 1714 -19
rect 1668 -91 1714 -53
rect 1668 -125 1674 -91
rect 1708 -125 1714 -91
rect 1668 -140 1714 -125
rect 1846 125 1892 140
rect 1846 91 1852 125
rect 1886 91 1892 125
rect 1846 53 1892 91
rect 1846 19 1852 53
rect 1886 19 1892 53
rect 1846 -19 1892 19
rect 1846 -53 1852 -19
rect 1886 -53 1892 -19
rect 1846 -91 1892 -53
rect 1846 -125 1852 -91
rect 1886 -125 1892 -91
rect 1846 -140 1892 -125
rect 2024 125 2070 140
rect 2024 91 2030 125
rect 2064 91 2070 125
rect 2024 53 2070 91
rect 2024 19 2030 53
rect 2064 19 2070 53
rect 2024 -19 2070 19
rect 2024 -53 2030 -19
rect 2064 -53 2070 -19
rect 2024 -91 2070 -53
rect 2024 -125 2030 -91
rect 2064 -125 2070 -91
rect 2024 -140 2070 -125
rect 2202 125 2248 140
rect 2202 91 2208 125
rect 2242 91 2248 125
rect 2202 53 2248 91
rect 2202 19 2208 53
rect 2242 19 2248 53
rect 2202 -19 2248 19
rect 2202 -53 2208 -19
rect 2242 -53 2248 -19
rect 2202 -91 2248 -53
rect 2202 -125 2208 -91
rect 2242 -125 2248 -91
rect 2202 -140 2248 -125
rect 2380 125 2426 140
rect 2380 91 2386 125
rect 2420 91 2426 125
rect 2380 53 2426 91
rect 2380 19 2386 53
rect 2420 19 2426 53
rect 2380 -19 2426 19
rect 2380 -53 2386 -19
rect 2420 -53 2426 -19
rect 2380 -91 2426 -53
rect 2380 -125 2386 -91
rect 2420 -125 2426 -91
rect 2380 -140 2426 -125
rect 2558 125 2604 140
rect 2558 91 2564 125
rect 2598 91 2604 125
rect 2558 53 2604 91
rect 2558 19 2564 53
rect 2598 19 2604 53
rect 2558 -19 2604 19
rect 2558 -53 2564 -19
rect 2598 -53 2604 -19
rect 2558 -91 2604 -53
rect 2558 -125 2564 -91
rect 2598 -125 2604 -91
rect 2558 -140 2604 -125
rect 2736 125 2782 140
rect 2736 91 2742 125
rect 2776 91 2782 125
rect 2736 53 2782 91
rect 2736 19 2742 53
rect 2776 19 2782 53
rect 2736 -19 2782 19
rect 2736 -53 2742 -19
rect 2776 -53 2782 -19
rect 2736 -91 2782 -53
rect 2736 -125 2742 -91
rect 2776 -125 2782 -91
rect 2736 -140 2782 -125
rect 2914 125 2960 140
rect 2914 91 2920 125
rect 2954 91 2960 125
rect 2914 53 2960 91
rect 2914 19 2920 53
rect 2954 19 2960 53
rect 2914 -19 2960 19
rect 2914 -53 2920 -19
rect 2954 -53 2960 -19
rect 2914 -91 2960 -53
rect 2914 -125 2920 -91
rect 2954 -125 2960 -91
rect 2914 -140 2960 -125
rect 3092 125 3138 140
rect 3092 91 3098 125
rect 3132 91 3138 125
rect 3092 53 3138 91
rect 3092 19 3098 53
rect 3132 19 3138 53
rect 3092 -19 3138 19
rect 3092 -53 3098 -19
rect 3132 -53 3138 -19
rect 3092 -91 3138 -53
rect 3092 -125 3098 -91
rect 3132 -125 3138 -91
rect 3092 -140 3138 -125
rect -3064 -178 -2988 -172
rect -3064 -212 -3043 -178
rect -3009 -212 -2988 -178
rect -3064 -228 -2988 -212
rect -2886 -178 -2810 -172
rect -2886 -212 -2865 -178
rect -2831 -212 -2810 -178
rect -2886 -228 -2810 -212
rect -2708 -178 -2632 -172
rect -2708 -212 -2687 -178
rect -2653 -212 -2632 -178
rect -2708 -228 -2632 -212
rect -2530 -178 -2454 -172
rect -2530 -212 -2509 -178
rect -2475 -212 -2454 -178
rect -2530 -228 -2454 -212
rect -2352 -178 -2276 -172
rect -2352 -212 -2331 -178
rect -2297 -212 -2276 -178
rect -2352 -228 -2276 -212
rect -2174 -178 -2098 -172
rect -2174 -212 -2153 -178
rect -2119 -212 -2098 -178
rect -2174 -228 -2098 -212
rect -1996 -178 -1920 -172
rect -1996 -212 -1975 -178
rect -1941 -212 -1920 -178
rect -1996 -228 -1920 -212
rect -1818 -178 -1742 -172
rect -1818 -212 -1797 -178
rect -1763 -212 -1742 -178
rect -1818 -228 -1742 -212
rect -1640 -178 -1564 -172
rect -1640 -212 -1619 -178
rect -1585 -212 -1564 -178
rect -1640 -228 -1564 -212
rect -1462 -178 -1386 -172
rect -1462 -212 -1441 -178
rect -1407 -212 -1386 -178
rect -1462 -228 -1386 -212
rect -1284 -178 -1208 -172
rect -1284 -212 -1263 -178
rect -1229 -212 -1208 -178
rect -1284 -228 -1208 -212
rect -1106 -178 -1030 -172
rect -1106 -212 -1085 -178
rect -1051 -212 -1030 -178
rect -1106 -228 -1030 -212
rect -928 -178 -852 -172
rect -928 -212 -907 -178
rect -873 -212 -852 -178
rect -928 -228 -852 -212
rect -750 -178 -674 -172
rect -750 -212 -729 -178
rect -695 -212 -674 -178
rect -750 -228 -674 -212
rect -572 -178 -496 -172
rect -572 -212 -551 -178
rect -517 -212 -496 -178
rect -572 -228 -496 -212
rect -394 -178 -318 -172
rect -394 -212 -373 -178
rect -339 -212 -318 -178
rect -394 -228 -318 -212
rect -216 -178 -140 -172
rect -216 -212 -195 -178
rect -161 -212 -140 -178
rect -216 -228 -140 -212
rect -38 -178 38 -172
rect -38 -212 -17 -178
rect 17 -212 38 -178
rect -38 -228 38 -212
rect 140 -178 216 -172
rect 140 -212 161 -178
rect 195 -212 216 -178
rect 140 -228 216 -212
rect 318 -178 394 -172
rect 318 -212 339 -178
rect 373 -212 394 -178
rect 318 -228 394 -212
rect 496 -178 572 -172
rect 496 -212 517 -178
rect 551 -212 572 -178
rect 496 -228 572 -212
rect 674 -178 750 -172
rect 674 -212 695 -178
rect 729 -212 750 -178
rect 674 -228 750 -212
rect 852 -178 928 -172
rect 852 -212 873 -178
rect 907 -212 928 -178
rect 852 -228 928 -212
rect 1030 -178 1106 -172
rect 1030 -212 1051 -178
rect 1085 -212 1106 -178
rect 1030 -228 1106 -212
rect 1208 -178 1284 -172
rect 1208 -212 1229 -178
rect 1263 -212 1284 -178
rect 1208 -228 1284 -212
rect 1386 -178 1462 -172
rect 1386 -212 1407 -178
rect 1441 -212 1462 -178
rect 1386 -228 1462 -212
rect 1564 -178 1640 -172
rect 1564 -212 1585 -178
rect 1619 -212 1640 -178
rect 1564 -228 1640 -212
rect 1742 -178 1818 -172
rect 1742 -212 1763 -178
rect 1797 -212 1818 -178
rect 1742 -228 1818 -212
rect 1920 -178 1996 -172
rect 1920 -212 1941 -178
rect 1975 -212 1996 -178
rect 1920 -228 1996 -212
rect 2098 -178 2174 -172
rect 2098 -212 2119 -178
rect 2153 -212 2174 -178
rect 2098 -228 2174 -212
rect 2276 -178 2352 -172
rect 2276 -212 2297 -178
rect 2331 -212 2352 -178
rect 2276 -228 2352 -212
rect 2454 -178 2530 -172
rect 2454 -212 2475 -178
rect 2509 -212 2530 -178
rect 2454 -228 2530 -212
rect 2632 -178 2708 -172
rect 2632 -212 2653 -178
rect 2687 -212 2708 -178
rect 2632 -228 2708 -212
rect 2810 -178 2886 -172
rect 2810 -212 2831 -178
rect 2865 -212 2886 -178
rect 2810 -228 2886 -212
rect 2988 -178 3064 -172
rect 2988 -212 3009 -178
rect 3043 -212 3064 -178
rect 2988 -228 3064 -212
<< end >>
