magic
tech sky130A
magscale 1 2
timestamp 1654426382
<< nwell >>
rect -7706 -1114 -7326 -1106
rect 3340 -1114 3860 -1110
rect -7706 -1544 3968 -1114
rect -7706 -7062 -7326 -1544
rect 2580 -5606 2928 -5240
rect 2576 -6508 2968 -6100
rect 3340 -7062 3860 -1544
rect -7738 -7292 3970 -7062
rect -7706 -7368 -7326 -7292
rect 3340 -7316 3860 -7292
<< psubdiff >>
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect 13619 -7731 13719 -7621
rect -7115 -15087 -6889 -15063
rect -7115 -15265 -7091 -15087
rect -6913 -15265 -6889 -15087
rect -7115 -15289 -6889 -15265
rect -7149 -15448 -6923 -15424
rect -7149 -15626 -7125 -15448
rect -6947 -15626 -6923 -15448
rect -7149 -15650 -6923 -15626
rect -7605 -17459 -7505 -17268
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< nsubdiff >>
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect 3610 -1520 3703 -1353
rect 2626 -5346 2852 -5322
rect 2626 -5524 2650 -5346
rect 2828 -5524 2852 -5346
rect 2626 -5548 2852 -5524
rect 2654 -6231 2880 -6207
rect 2654 -6409 2678 -6231
rect 2856 -6409 2880 -6231
rect 2654 -6433 2880 -6409
rect -7605 -7140 -7512 -6976
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
<< psubdiffcont >>
rect -7264 -7621 13443 -7521
rect -7605 -17268 -7505 -7850
rect -7091 -15265 -6913 -15087
rect -7125 -15626 -6947 -15448
rect 13619 -17149 13719 -7731
rect -7323 -17559 13384 -17459
<< nsubdiffcont >>
rect -7379 -1353 3329 -1260
rect -7605 -6976 -7512 -1507
rect 2650 -5524 2828 -5346
rect 2678 -6409 2856 -6231
rect 3610 -6989 3703 -1520
rect -7282 -7233 3426 -7140
<< locali >>
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect 3610 -1520 3703 -1353
rect 2626 -5346 2852 -5322
rect 2626 -5524 2650 -5346
rect 2828 -5524 2852 -5346
rect 2626 -5548 2852 -5524
rect 2654 -6231 2880 -6207
rect 2654 -6409 2678 -6231
rect 2856 -6409 2880 -6231
rect 2654 -6433 2880 -6409
rect -7605 -7140 -7512 -6976
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect 13619 -7731 13719 -7621
rect -7115 -15087 -6889 -15063
rect -7115 -15265 -7091 -15087
rect -6913 -15265 -6889 -15087
rect -7115 -15289 -6889 -15265
rect -7149 -15448 -6923 -15424
rect -7149 -15626 -7125 -15448
rect -6947 -15626 -6923 -15448
rect -7149 -15650 -6923 -15626
rect -7605 -17459 -7505 -17268
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< viali >>
rect -7379 -1353 3329 -1260
rect 2650 -5524 2828 -5346
rect 2678 -6409 2856 -6231
rect -7091 -15265 -6913 -15087
rect -7125 -15626 -6947 -15448
rect -7323 -17559 13384 -17459
<< metal1 >>
rect 7034 2713 7080 2891
rect 16034 2713 16080 2891
rect 7034 1691 7080 1863
rect 16034 1691 16080 1863
rect 7034 913 7080 1091
rect 16034 913 16080 1091
rect 7034 -109 7080 63
rect 16034 -109 16080 63
rect 7034 -887 7080 -709
rect 16034 -887 16080 -709
rect -7605 -1260 3704 -1200
rect -7605 -1353 -7379 -1260
rect 3329 -1353 3704 -1260
rect -7605 -1467 3704 -1353
rect -5132 -1684 -4948 -1467
rect 7034 -1909 7080 -1737
rect 16034 -1909 16080 -1737
rect 5327 -2258 5337 -2205
rect 5390 -2258 5400 -2205
rect 2638 -5346 2840 -5340
rect 2638 -5524 2650 -5346
rect 2828 -5524 2840 -5346
rect 2638 -5530 2840 -5524
rect 5337 -5527 5390 -2258
rect 6670 -2263 6680 -2199
rect 6744 -2263 6754 -2199
rect 7034 -2687 7080 -2509
rect 16034 -2687 16080 -2509
rect 6212 -3515 6222 -3451
rect 6286 -3515 6296 -3451
rect 7034 -3709 7080 -3537
rect 16034 -3709 16080 -3537
rect 7034 -4487 7080 -4309
rect 16034 -4487 16080 -4309
rect 5604 -5271 5614 -5207
rect 5678 -5271 5688 -5207
rect 7034 -5509 7080 -5337
rect 16034 -5509 16080 -5337
rect 5327 -5580 5337 -5527
rect 5390 -5580 5400 -5527
rect 2666 -6231 2868 -6225
rect 2666 -6409 2678 -6231
rect 2856 -6409 2868 -6231
rect 7034 -6287 7080 -6109
rect 16034 -6287 16080 -6109
rect 2666 -6415 2868 -6409
rect 17826 -6521 17901 -4862
rect 17821 -6585 17831 -6521
rect 17895 -6585 17905 -6521
rect 7034 -7309 7080 -7137
rect 16034 -7309 16080 -7137
rect -6976 -12565 -6590 -12512
rect 18337 -13421 18412 -6747
rect 18327 -13496 18337 -13421
rect 18412 -13496 18422 -13421
rect 18337 -13506 18412 -13496
rect -6976 -13905 -6590 -13852
rect -6965 -14260 -6590 -14226
rect -7103 -15087 -6901 -15081
rect -7103 -15265 -7091 -15087
rect -6913 -15265 -6901 -15087
rect -7103 -15271 -6901 -15265
rect -7137 -15448 -6935 -15442
rect -7137 -15626 -7125 -15448
rect -6947 -15626 -6935 -15448
rect -7137 -15632 -6935 -15626
rect -7605 -17251 -7329 -17250
rect -1736 -17251 -1528 -17248
rect -658 -17251 -450 -17248
rect 408 -17251 616 -17248
rect 1488 -17251 1696 -17248
rect 2547 -17251 2755 -17248
rect 3614 -17251 3822 -17248
rect 9672 -17251 9706 -17248
rect -7605 -17252 -5044 -17251
rect -4766 -17252 12798 -17251
rect 13168 -17252 13720 -17251
rect -7605 -17459 13720 -17252
rect -7605 -17559 -7323 -17459
rect 13384 -17527 13720 -17459
rect 13384 -17559 13719 -17527
rect -7605 -17587 13719 -17559
<< via1 >>
rect 5337 -2258 5390 -2205
rect 6680 -2263 6744 -2199
rect 6222 -3515 6286 -3451
rect 5614 -5271 5678 -5207
rect 5337 -5580 5390 -5527
rect 17831 -6585 17895 -6521
rect 18337 -13496 18412 -13421
<< metal2 >>
rect 5337 -2205 5390 -2195
rect 6680 -2199 6744 -2189
rect 5390 -2258 6680 -2205
rect 5337 -2268 5390 -2258
rect 6744 -2258 6748 -2205
rect 6680 -2273 6744 -2263
rect 6222 -3451 6286 -3441
rect 3336 -3509 6222 -3456
rect 6286 -3509 6297 -3456
rect 6222 -3525 6286 -3515
rect 5614 -5207 5678 -5197
rect 3928 -5266 5614 -5213
rect 5678 -5266 5685 -5213
rect 5614 -5281 5678 -5271
rect 5337 -5527 5390 -5517
rect 5337 -7770 5390 -5580
rect 17831 -6521 17895 -6511
rect 17831 -8716 17895 -6585
rect 13184 -8769 17895 -8716
rect 18337 -13421 18412 -13411
rect 13226 -13486 18337 -13433
rect 18412 -13486 18422 -13433
rect 18337 -13506 18412 -13496
<< metal3 >>
rect 6451 929 6515 2665
rect 6704 121 6768 1857
rect 17697 122 17761 1858
rect 17950 929 18014 2665
rect 6451 -6271 6515 -4535
rect 6704 -5279 6768 -3543
rect 17697 -7078 17761 -5342
rect 17950 -6271 18014 -4535
use sc_cmfb  sc_cmfb_0 ~/EE372/incremental_delta_sigma_adc/design/analog_modulator/layout/sc_cmfb
timestamp 1654408082
transform 1 0 9102 0 1 -5469
box -3494 -1840 9310 8360
<< labels >>
flabel metal1 -7420 -1403 -7420 -1403 1 FreeSans 1200 0 0 0 VDD
flabel metal1 -7407 -17402 -7407 -17402 1 FreeSans 1200 0 0 0 VSS
flabel metal1 -6957 -14245 -6957 -14245 1 FreeSans 1200 0 0 0 i_bias
flabel metal1 -6952 -13880 -6952 -13880 1 FreeSans 1200 0 0 0 in
flabel metal1 7057 2874 7057 2874 1 FreeSans 400 0 0 0 VDD
flabel metal1 7057 1707 7057 1707 1 FreeSans 400 0 0 0 VSS
flabel metal1 7058 -83 7058 -83 1 FreeSans 400 0 0 0 VSS
flabel metal1 7058 -739 7058 -739 1 FreeSans 400 0 0 0 VDD
flabel metal1 7058 -1885 7058 -1885 1 FreeSans 400 0 0 0 VSS
flabel metal1 7058 -2537 7058 -2537 1 FreeSans 400 0 0 0 VDD
flabel metal1 7051 -4329 7051 -4329 1 FreeSans 400 0 0 0 VDD
flabel metal1 7054 -5489 7054 -5489 1 FreeSans 400 0 0 0 VSS
flabel metal1 7054 -7288 7054 -7288 1 FreeSans 400 0 0 0 VSS
flabel metal1 16056 -7290 16056 -7290 1 FreeSans 400 0 0 0 VSS
flabel metal1 16057 -6136 16057 -6136 1 FreeSans 400 0 0 0 VDD
flabel metal1 16055 -5482 16055 -5482 1 FreeSans 400 0 0 0 VSS
flabel metal1 16057 -2529 16057 -2529 1 FreeSans 400 0 0 0 VDD
flabel metal1 16055 -1886 16055 -1886 1 FreeSans 400 0 0 0 VSS
flabel metal1 16057 -86 16057 -86 1 FreeSans 400 0 0 0 VSS
flabel metal1 16057 1070 16057 1070 1 FreeSans 400 0 0 0 VDD
flabel metal1 16057 1716 16057 1716 1 FreeSans 400 0 0 0 VSS
flabel metal1 16057 2870 16057 2870 1 FreeSans 400 0 0 0 VDD
flabel metal3 6479 2585 6479 2585 1 FreeSans 400 0 0 0 p2_b
flabel metal3 6738 1807 6738 1807 1 FreeSans 400 0 0 0 p2
flabel metal3 6486 -6211 6486 -6211 1 FreeSans 400 0 0 0 p1_b
flabel metal3 6735 -5207 6735 -5207 1 FreeSans 400 0 0 0 p1
flabel metal3 17730 1821 17730 1821 1 FreeSans 400 0 0 0 p2
flabel metal3 17980 2631 17980 2631 1 FreeSans 400 0 0 0 p2_b
flabel metal3 17727 -7023 17727 -7023 1 FreeSans 400 0 0 0 p1
flabel metal3 17984 -6236 17984 -6236 1 FreeSans 400 0 0 0 p1_b
flabel metal2 17862 -8732 17862 -8732 1 FreeSans 800 0 0 0 cm
flabel metal1 7058 1058 7058 1058 1 FreeSans 400 0 0 0 VDD
flabel metal1 7058 -3672 7058 -3672 1 FreeSans 400 0 0 0 VSS
flabel metal1 7058 -6144 7058 -6144 1 FreeSans 400 0 0 0 VDD
flabel metal1 16056 -4338 16056 -4338 1 FreeSans 400 0 0 0 VDD
flabel metal1 16056 -3678 16056 -3678 1 FreeSans 400 0 0 0 VSS
flabel metal1 16056 -738 16056 -738 1 FreeSans 400 0 0 0 VDD
flabel metal1 -6950 -12541 -6950 -12541 1 FreeSans 1200 0 0 0 ip
flabel metal2 4134 -3484 4134 -3484 1 FreeSans 1600 0 0 0 on
flabel metal2 4024 -5242 4024 -5242 1 FreeSans 1600 0 0 0 op
flabel metal2 5364 -7430 5364 -7430 1 FreeSans 1600 0 0 0 cmc
flabel metal2 13302 -13462 13302 -13462 1 FreeSans 1600 0 0 0 bias_a
flabel viali -7002 -15176 -7002 -15176 1 FreeSans 400 0 0 0 VSS
flabel viali -7036 -15537 -7036 -15537 1 FreeSans 400 0 0 0 VSS
flabel viali 2767 -6320 2767 -6320 1 FreeSans 400 0 0 0 VDD
flabel viali 2739 -5435 2739 -5435 1 FreeSans 400 0 0 0 VDD
<< end >>
