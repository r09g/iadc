* NGSPICE file created from a_mux2_en.ext - technology: sky130A

.subckt pmos_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136#
M0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38 as=4.488e+11p ps=3.38 w=1.36 l=0.15
M1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38 as=4.488e+11p ps=3.38 w=1.36 l=0.15
M2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38 as=0p ps=0u w=1.36 l=0.15
M3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# pmos ad=0p pd=0u as=4.488e+11p ps=3.38 w=1.36 l=0.15
M4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38 as=4.216e+11p ps=3.34 w=1.36 l=0.15
M5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# pmos ad=0p pd=0u as=0p ps=0u w=1.36 l=0.15
M6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38 as=0p ps=0u w=1.36 l=0.15
M7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# pmos ad=4.216e+11p pd=3.34 as=0p ps=0u w=1.36 l=0.15
M8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# pmos ad=4.488e+11p pd=3.38 as=0p ps=0u w=1.36 l=0.15
M9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# pmos ad=0p pd=0u as=0p ps=0u w=1.36 l=0.15
.ends

.subckt nmos_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
M0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7 as=1.716e+11p ps=1.7 w=0.52 l=0.15
M1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7 as=1.612e+11p ps=1.66 w=0.52 l=0.15
M2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7 as=1.716e+11p ps=1.7 w=0.52 l=0.15
M3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
M4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
M5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7 as=1.716e+11p ps=1.7 w=0.52 l=0.15
M6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# nmos ad=1.716e+11p pd=1.7 as=1.716e+11p ps=1.7 w=0.52 l=0.15
M7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
M8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# nmos ad=1.612e+11p pd=1.66 as=0p ps=0u w=0.52 l=0.15
M9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# nmos ad=0p pd=0u as=0p ps=0u w=0.52 l=0.15
.ends

.subckt transmission_gate out en_b en VSS VDD in
Xpmos_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ pmos_UNG2NQ
Xnmos_6J4AMR_0 out in in out in in VSS out en in out out out nmos_6J4AMR
.ends

.subckt nmos_E56BNL a_n33_33# a_n73_n89# a_15_n89# VSUBS
M0 a_15_n89# a_n33_33# a_n73_n89# VSUBS nmos ad=1.45e+11p pd=1.58 as=1.45e+11p ps=1.58 w=0.50 l=0.15
.ends

.subckt switch_5t out en_b en VDD in VSS
Xtransmission_gate_0 transmission_gate_1_in en_b en VSS VDD in transmission_gate
Xtransmission_gate_1 out en_b en VSS VDD transmission_gate_1_in transmission_gate
Xnmos_E56BNL_0 en_b VSS transmission_gate_1_in VSS nmos_E56BNL
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VPWR Y VNB VPB
M0 Y A VGND VNB nmos ad=1.69e+11p pd=1.82 as=1.69e+11p ps=1.82 w=0.65 l=0.15
M1 Y A VPWR VPB pmos_hvt ad=2.6e+11p pd=2.52 as=2.6e+11p ps=2.52 w=1 l=0.15
.ends

.subckt a_mux2_en en s0 in0 in1 out VDD VSS
Xswitch_5t_0 out switch_5t_1_en s0 VDD switch_5t_0_in VSS switch_5t
Xswitch_5t_1 out s0 switch_5t_1_en VDD switch_5t_1_in VSS switch_5t
Xtransmission_gate_0 switch_5t_1_in transmission_gate_1_en_b en VSS VDD in0 transmission_gate
Xtransmission_gate_1 switch_5t_0_in transmission_gate_1_en_b en VSS VDD in1 transmission_gate
Xsky130_fd_sc_hd__inv_1_1 s0 VSS VDD switch_5t_1_en VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 en VSS VDD transmission_gate_1_en_b VSS VDD sky130_fd_sc_hd__inv_1
.ends

