magic
tech sky130A
magscale 1 2
timestamp 1653690071
<< nwell >>
rect -3266 -716 -1972 -66
rect -1018 -1059 -298 -738
rect -742 -1304 -298 -1059
rect 285 -1180 3100 -530
rect -3266 -2050 -1972 -1400
rect -742 -2071 -298 -1826
rect -1294 -2392 -298 -2071
rect 285 -2514 3100 -1864
rect -3266 -3428 -1972 -2778
rect -1294 -3235 -298 -2914
rect -742 -3480 -298 -3235
rect 285 -3892 3100 -3242
rect -3266 -4806 -1972 -4156
rect -742 -4568 -298 -4002
rect 285 -5270 3100 -4620
<< pwell >>
rect -951 -494 -917 -460
rect -583 -494 -549 -460
rect -938 -498 -917 -494
rect -570 -498 -549 -494
rect -938 -515 -635 -498
rect -938 -525 -615 -515
rect -570 -525 -384 -498
rect -938 -680 -384 -525
rect 285 -528 3100 -66
rect 1553 -530 1809 -528
rect -3266 -1180 -1972 -718
rect -701 -1586 -384 -1362
rect -701 -1768 -337 -1586
rect -3266 -2514 -1972 -2052
rect 285 -1862 3100 -1400
rect 1553 -1864 1809 -1862
rect -1253 -2615 -337 -2450
rect -1241 -2632 -337 -2615
rect -1122 -2636 -1101 -2632
rect -1135 -2670 -1101 -2636
rect -857 -2663 -825 -2641
rect -767 -2665 -735 -2643
rect -1122 -2674 -1101 -2670
rect -584 -2674 -550 -2632
rect -1253 -2701 -1167 -2691
rect -1122 -2701 -936 -2674
rect -701 -2701 -615 -2691
rect -607 -2701 -337 -2674
rect -1253 -2856 -337 -2701
rect -3266 -3892 -1972 -3430
rect 285 -3240 3100 -2778
rect 1553 -3242 1809 -3240
rect -701 -3693 -337 -3538
rect -701 -3703 -615 -3693
rect -607 -3720 -337 -3693
rect -584 -3724 -550 -3720
rect -584 -3758 -549 -3724
rect -570 -3762 -549 -3758
rect -701 -3789 -615 -3779
rect -570 -3789 -384 -3762
rect -702 -3944 -338 -3789
rect 285 -4618 3100 -4156
rect 1553 -4620 1809 -4618
rect -701 -4781 -337 -4626
rect -701 -4791 -615 -4781
rect -570 -4808 -384 -4781
rect -3266 -5270 -1972 -4808
rect -570 -4812 -549 -4808
rect -583 -4846 -549 -4812
<< nmos >>
rect 485 -380 515 -276
rect 581 -380 611 -276
rect 677 -380 707 -276
rect 773 -380 803 -276
rect 869 -380 899 -276
rect 965 -380 995 -276
rect 1061 -380 1091 -276
rect 1157 -380 1187 -276
rect 1253 -380 1283 -276
rect 1349 -380 1379 -276
rect 1662 -384 1692 -284
rect 2006 -380 2036 -276
rect 2102 -380 2132 -276
rect 2198 -380 2228 -276
rect 2294 -380 2324 -276
rect 2390 -380 2420 -276
rect 2486 -380 2516 -276
rect 2582 -380 2612 -276
rect 2678 -380 2708 -276
rect 2774 -380 2804 -276
rect 2870 -380 2900 -276
rect -3066 -970 -3036 -866
rect -2970 -970 -2940 -866
rect -2874 -970 -2844 -866
rect -2778 -970 -2748 -866
rect -2682 -970 -2652 -866
rect -2586 -970 -2556 -866
rect -2490 -970 -2460 -866
rect -2394 -970 -2364 -866
rect -2298 -970 -2268 -866
rect -2202 -970 -2172 -866
rect 485 -1714 515 -1610
rect 581 -1714 611 -1610
rect 677 -1714 707 -1610
rect 773 -1714 803 -1610
rect 869 -1714 899 -1610
rect 965 -1714 995 -1610
rect 1061 -1714 1091 -1610
rect 1157 -1714 1187 -1610
rect 1253 -1714 1283 -1610
rect 1349 -1714 1379 -1610
rect 1662 -1718 1692 -1618
rect 2006 -1714 2036 -1610
rect 2102 -1714 2132 -1610
rect 2198 -1714 2228 -1610
rect 2294 -1714 2324 -1610
rect 2390 -1714 2420 -1610
rect 2486 -1714 2516 -1610
rect 2582 -1714 2612 -1610
rect 2678 -1714 2708 -1610
rect 2774 -1714 2804 -1610
rect 2870 -1714 2900 -1610
rect -3066 -2304 -3036 -2200
rect -2970 -2304 -2940 -2200
rect -2874 -2304 -2844 -2200
rect -2778 -2304 -2748 -2200
rect -2682 -2304 -2652 -2200
rect -2586 -2304 -2556 -2200
rect -2490 -2304 -2460 -2200
rect -2394 -2304 -2364 -2200
rect -2298 -2304 -2268 -2200
rect -2202 -2304 -2172 -2200
rect 485 -3092 515 -2988
rect 581 -3092 611 -2988
rect 677 -3092 707 -2988
rect 773 -3092 803 -2988
rect 869 -3092 899 -2988
rect 965 -3092 995 -2988
rect 1061 -3092 1091 -2988
rect 1157 -3092 1187 -2988
rect 1253 -3092 1283 -2988
rect 1349 -3092 1379 -2988
rect 1662 -3096 1692 -2996
rect 2006 -3092 2036 -2988
rect 2102 -3092 2132 -2988
rect 2198 -3092 2228 -2988
rect 2294 -3092 2324 -2988
rect 2390 -3092 2420 -2988
rect 2486 -3092 2516 -2988
rect 2582 -3092 2612 -2988
rect 2678 -3092 2708 -2988
rect 2774 -3092 2804 -2988
rect 2870 -3092 2900 -2988
rect -3066 -3682 -3036 -3578
rect -2970 -3682 -2940 -3578
rect -2874 -3682 -2844 -3578
rect -2778 -3682 -2748 -3578
rect -2682 -3682 -2652 -3578
rect -2586 -3682 -2556 -3578
rect -2490 -3682 -2460 -3578
rect -2394 -3682 -2364 -3578
rect -2298 -3682 -2268 -3578
rect -2202 -3682 -2172 -3578
rect 485 -4470 515 -4366
rect 581 -4470 611 -4366
rect 677 -4470 707 -4366
rect 773 -4470 803 -4366
rect 869 -4470 899 -4366
rect 965 -4470 995 -4366
rect 1061 -4470 1091 -4366
rect 1157 -4470 1187 -4366
rect 1253 -4470 1283 -4366
rect 1349 -4470 1379 -4366
rect 1662 -4474 1692 -4374
rect 2006 -4470 2036 -4366
rect 2102 -4470 2132 -4366
rect 2198 -4470 2228 -4366
rect 2294 -4470 2324 -4366
rect 2390 -4470 2420 -4366
rect 2486 -4470 2516 -4366
rect 2582 -4470 2612 -4366
rect 2678 -4470 2708 -4366
rect 2774 -4470 2804 -4366
rect 2870 -4470 2900 -4366
rect -3066 -5060 -3036 -4956
rect -2970 -5060 -2940 -4956
rect -2874 -5060 -2844 -4956
rect -2778 -5060 -2748 -4956
rect -2682 -5060 -2652 -4956
rect -2586 -5060 -2556 -4956
rect -2490 -5060 -2460 -4956
rect -2394 -5060 -2364 -4956
rect -2298 -5060 -2268 -4956
rect -2202 -5060 -2172 -4956
<< scnmos >>
rect -860 -654 -830 -524
rect -492 -654 -462 -524
rect -492 -1518 -462 -1388
rect -529 -1742 -499 -1612
rect -445 -1742 -415 -1612
rect -1044 -2606 -1014 -2476
rect -529 -2606 -499 -2476
rect -445 -2606 -415 -2476
rect -1044 -2830 -1014 -2700
rect -529 -2830 -499 -2700
rect -445 -2830 -415 -2700
rect -529 -3694 -499 -3564
rect -445 -3694 -415 -3564
rect -492 -3918 -462 -3788
rect -492 -4782 -462 -4652
<< pmos >>
rect -3066 -558 -3036 -286
rect -2970 -558 -2940 -286
rect -2874 -558 -2844 -286
rect -2778 -558 -2748 -286
rect -2682 -558 -2652 -286
rect -2586 -558 -2556 -286
rect -2490 -558 -2460 -286
rect -2394 -558 -2364 -286
rect -2298 -558 -2268 -286
rect -2202 -558 -2172 -286
rect 485 -960 515 -688
rect 581 -960 611 -688
rect 677 -960 707 -688
rect 773 -960 803 -688
rect 869 -960 899 -688
rect 965 -960 995 -688
rect 1061 -960 1091 -688
rect 1157 -960 1187 -688
rect 1253 -960 1283 -688
rect 1349 -960 1379 -688
rect 2006 -960 2036 -688
rect 2102 -960 2132 -688
rect 2198 -960 2228 -688
rect 2294 -960 2324 -688
rect 2390 -960 2420 -688
rect 2486 -960 2516 -688
rect 2582 -960 2612 -688
rect 2678 -960 2708 -688
rect 2774 -960 2804 -688
rect 2870 -960 2900 -688
rect -3066 -1892 -3036 -1620
rect -2970 -1892 -2940 -1620
rect -2874 -1892 -2844 -1620
rect -2778 -1892 -2748 -1620
rect -2682 -1892 -2652 -1620
rect -2586 -1892 -2556 -1620
rect -2490 -1892 -2460 -1620
rect -2394 -1892 -2364 -1620
rect -2298 -1892 -2268 -1620
rect -2202 -1892 -2172 -1620
rect 485 -2294 515 -2022
rect 581 -2294 611 -2022
rect 677 -2294 707 -2022
rect 773 -2294 803 -2022
rect 869 -2294 899 -2022
rect 965 -2294 995 -2022
rect 1061 -2294 1091 -2022
rect 1157 -2294 1187 -2022
rect 1253 -2294 1283 -2022
rect 1349 -2294 1379 -2022
rect 2006 -2294 2036 -2022
rect 2102 -2294 2132 -2022
rect 2198 -2294 2228 -2022
rect 2294 -2294 2324 -2022
rect 2390 -2294 2420 -2022
rect 2486 -2294 2516 -2022
rect 2582 -2294 2612 -2022
rect 2678 -2294 2708 -2022
rect 2774 -2294 2804 -2022
rect 2870 -2294 2900 -2022
rect -3066 -3270 -3036 -2998
rect -2970 -3270 -2940 -2998
rect -2874 -3270 -2844 -2998
rect -2778 -3270 -2748 -2998
rect -2682 -3270 -2652 -2998
rect -2586 -3270 -2556 -2998
rect -2490 -3270 -2460 -2998
rect -2394 -3270 -2364 -2998
rect -2298 -3270 -2268 -2998
rect -2202 -3270 -2172 -2998
rect 485 -3672 515 -3400
rect 581 -3672 611 -3400
rect 677 -3672 707 -3400
rect 773 -3672 803 -3400
rect 869 -3672 899 -3400
rect 965 -3672 995 -3400
rect 1061 -3672 1091 -3400
rect 1157 -3672 1187 -3400
rect 1253 -3672 1283 -3400
rect 1349 -3672 1379 -3400
rect 2006 -3672 2036 -3400
rect 2102 -3672 2132 -3400
rect 2198 -3672 2228 -3400
rect 2294 -3672 2324 -3400
rect 2390 -3672 2420 -3400
rect 2486 -3672 2516 -3400
rect 2582 -3672 2612 -3400
rect 2678 -3672 2708 -3400
rect 2774 -3672 2804 -3400
rect 2870 -3672 2900 -3400
rect -3066 -4648 -3036 -4376
rect -2970 -4648 -2940 -4376
rect -2874 -4648 -2844 -4376
rect -2778 -4648 -2748 -4376
rect -2682 -4648 -2652 -4376
rect -2586 -4648 -2556 -4376
rect -2490 -4648 -2460 -4376
rect -2394 -4648 -2364 -4376
rect -2298 -4648 -2268 -4376
rect -2202 -4648 -2172 -4376
rect 485 -5050 515 -4778
rect 581 -5050 611 -4778
rect 677 -5050 707 -4778
rect 773 -5050 803 -4778
rect 869 -5050 899 -4778
rect 965 -5050 995 -4778
rect 1061 -5050 1091 -4778
rect 1157 -5050 1187 -4778
rect 1253 -5050 1283 -4778
rect 1349 -5050 1379 -4778
rect 2006 -5050 2036 -4778
rect 2102 -5050 2132 -4778
rect 2198 -5050 2228 -4778
rect 2294 -5050 2324 -4778
rect 2390 -5050 2420 -4778
rect 2486 -5050 2516 -4778
rect 2582 -5050 2612 -4778
rect 2678 -5050 2708 -4778
rect 2774 -5050 2804 -4778
rect 2870 -5050 2900 -4778
<< scpmoshvt >>
rect -860 -974 -830 -774
rect -492 -974 -462 -774
rect -492 -1268 -462 -1068
rect -529 -2062 -499 -1862
rect -445 -2062 -415 -1862
rect -1044 -2356 -1014 -2156
rect -529 -2356 -499 -2156
rect -445 -2356 -415 -2156
rect -1044 -3150 -1014 -2950
rect -529 -3150 -499 -2950
rect -445 -3150 -415 -2950
rect -529 -3444 -499 -3244
rect -445 -3444 -415 -3244
rect -492 -4238 -462 -4038
rect -492 -4532 -462 -4332
<< ndiff >>
rect 423 -288 485 -276
rect 423 -368 435 -288
rect 469 -368 485 -288
rect 423 -380 485 -368
rect 515 -288 581 -276
rect 515 -368 531 -288
rect 565 -368 581 -288
rect 515 -380 581 -368
rect 611 -288 677 -276
rect 611 -368 627 -288
rect 661 -368 677 -288
rect 611 -380 677 -368
rect 707 -288 773 -276
rect 707 -368 723 -288
rect 757 -368 773 -288
rect 707 -380 773 -368
rect 803 -288 869 -276
rect 803 -368 819 -288
rect 853 -368 869 -288
rect 803 -380 869 -368
rect 899 -288 965 -276
rect 899 -368 915 -288
rect 949 -368 965 -288
rect 899 -380 965 -368
rect 995 -288 1061 -276
rect 995 -368 1011 -288
rect 1045 -368 1061 -288
rect 995 -380 1061 -368
rect 1091 -288 1157 -276
rect 1091 -368 1107 -288
rect 1141 -368 1157 -288
rect 1091 -380 1157 -368
rect 1187 -288 1253 -276
rect 1187 -368 1203 -288
rect 1237 -368 1253 -288
rect 1187 -380 1253 -368
rect 1283 -288 1349 -276
rect 1283 -368 1299 -288
rect 1333 -368 1349 -288
rect 1283 -380 1349 -368
rect 1379 -288 1441 -276
rect 1379 -368 1395 -288
rect 1429 -368 1441 -288
rect 1379 -380 1441 -368
rect 1604 -296 1662 -284
rect 1604 -372 1616 -296
rect 1650 -372 1662 -296
rect 1604 -384 1662 -372
rect 1692 -296 1750 -284
rect 1692 -372 1704 -296
rect 1738 -372 1750 -296
rect 1692 -384 1750 -372
rect 1944 -288 2006 -276
rect 1944 -368 1956 -288
rect 1990 -368 2006 -288
rect 1944 -380 2006 -368
rect 2036 -288 2102 -276
rect 2036 -368 2052 -288
rect 2086 -368 2102 -288
rect 2036 -380 2102 -368
rect 2132 -288 2198 -276
rect 2132 -368 2148 -288
rect 2182 -368 2198 -288
rect 2132 -380 2198 -368
rect 2228 -288 2294 -276
rect 2228 -368 2244 -288
rect 2278 -368 2294 -288
rect 2228 -380 2294 -368
rect 2324 -288 2390 -276
rect 2324 -368 2340 -288
rect 2374 -368 2390 -288
rect 2324 -380 2390 -368
rect 2420 -288 2486 -276
rect 2420 -368 2436 -288
rect 2470 -368 2486 -288
rect 2420 -380 2486 -368
rect 2516 -288 2582 -276
rect 2516 -368 2532 -288
rect 2566 -368 2582 -288
rect 2516 -380 2582 -368
rect 2612 -288 2678 -276
rect 2612 -368 2628 -288
rect 2662 -368 2678 -288
rect 2612 -380 2678 -368
rect 2708 -288 2774 -276
rect 2708 -368 2724 -288
rect 2758 -368 2774 -288
rect 2708 -380 2774 -368
rect 2804 -288 2870 -276
rect 2804 -368 2820 -288
rect 2854 -368 2870 -288
rect 2804 -380 2870 -368
rect 2900 -288 2962 -276
rect 2900 -368 2916 -288
rect 2950 -368 2962 -288
rect 2900 -380 2962 -368
rect -912 -540 -860 -524
rect -912 -574 -904 -540
rect -870 -574 -860 -540
rect -912 -608 -860 -574
rect -912 -642 -904 -608
rect -870 -642 -860 -608
rect -912 -654 -860 -642
rect -830 -540 -778 -524
rect -830 -574 -820 -540
rect -786 -574 -778 -540
rect -544 -540 -492 -524
rect -830 -608 -778 -574
rect -830 -642 -820 -608
rect -786 -642 -778 -608
rect -830 -654 -778 -642
rect -544 -574 -536 -540
rect -502 -574 -492 -540
rect -544 -608 -492 -574
rect -544 -642 -536 -608
rect -502 -642 -492 -608
rect -544 -654 -492 -642
rect -462 -540 -410 -524
rect -462 -574 -452 -540
rect -418 -574 -410 -540
rect -462 -608 -410 -574
rect -462 -642 -452 -608
rect -418 -642 -410 -608
rect -462 -654 -410 -642
rect -3128 -878 -3066 -866
rect -3128 -958 -3116 -878
rect -3082 -958 -3066 -878
rect -3128 -970 -3066 -958
rect -3036 -878 -2970 -866
rect -3036 -958 -3020 -878
rect -2986 -958 -2970 -878
rect -3036 -970 -2970 -958
rect -2940 -878 -2874 -866
rect -2940 -958 -2924 -878
rect -2890 -958 -2874 -878
rect -2940 -970 -2874 -958
rect -2844 -878 -2778 -866
rect -2844 -958 -2828 -878
rect -2794 -958 -2778 -878
rect -2844 -970 -2778 -958
rect -2748 -878 -2682 -866
rect -2748 -958 -2732 -878
rect -2698 -958 -2682 -878
rect -2748 -970 -2682 -958
rect -2652 -878 -2586 -866
rect -2652 -958 -2636 -878
rect -2602 -958 -2586 -878
rect -2652 -970 -2586 -958
rect -2556 -878 -2490 -866
rect -2556 -958 -2540 -878
rect -2506 -958 -2490 -878
rect -2556 -970 -2490 -958
rect -2460 -878 -2394 -866
rect -2460 -958 -2444 -878
rect -2410 -958 -2394 -878
rect -2460 -970 -2394 -958
rect -2364 -878 -2298 -866
rect -2364 -958 -2348 -878
rect -2314 -958 -2298 -878
rect -2364 -970 -2298 -958
rect -2268 -878 -2202 -866
rect -2268 -958 -2252 -878
rect -2218 -958 -2202 -878
rect -2268 -970 -2202 -958
rect -2172 -878 -2110 -866
rect -2172 -958 -2156 -878
rect -2122 -958 -2110 -878
rect -2172 -970 -2110 -958
rect -544 -1400 -492 -1388
rect -544 -1434 -536 -1400
rect -502 -1434 -492 -1400
rect -544 -1468 -492 -1434
rect -544 -1502 -536 -1468
rect -502 -1502 -492 -1468
rect -544 -1518 -492 -1502
rect -462 -1400 -410 -1388
rect -462 -1434 -452 -1400
rect -418 -1434 -410 -1400
rect -462 -1468 -410 -1434
rect -462 -1502 -452 -1468
rect -418 -1502 -410 -1468
rect -462 -1518 -410 -1502
rect -581 -1624 -529 -1612
rect -581 -1658 -573 -1624
rect -539 -1658 -529 -1624
rect -581 -1692 -529 -1658
rect -581 -1726 -573 -1692
rect -539 -1726 -529 -1692
rect -581 -1742 -529 -1726
rect -499 -1742 -445 -1612
rect -415 -1624 -363 -1612
rect -415 -1658 -405 -1624
rect -371 -1658 -363 -1624
rect -415 -1692 -363 -1658
rect -415 -1726 -405 -1692
rect -371 -1726 -363 -1692
rect -415 -1742 -363 -1726
rect 423 -1622 485 -1610
rect 423 -1702 435 -1622
rect 469 -1702 485 -1622
rect 423 -1714 485 -1702
rect 515 -1622 581 -1610
rect 515 -1702 531 -1622
rect 565 -1702 581 -1622
rect 515 -1714 581 -1702
rect 611 -1622 677 -1610
rect 611 -1702 627 -1622
rect 661 -1702 677 -1622
rect 611 -1714 677 -1702
rect 707 -1622 773 -1610
rect 707 -1702 723 -1622
rect 757 -1702 773 -1622
rect 707 -1714 773 -1702
rect 803 -1622 869 -1610
rect 803 -1702 819 -1622
rect 853 -1702 869 -1622
rect 803 -1714 869 -1702
rect 899 -1622 965 -1610
rect 899 -1702 915 -1622
rect 949 -1702 965 -1622
rect 899 -1714 965 -1702
rect 995 -1622 1061 -1610
rect 995 -1702 1011 -1622
rect 1045 -1702 1061 -1622
rect 995 -1714 1061 -1702
rect 1091 -1622 1157 -1610
rect 1091 -1702 1107 -1622
rect 1141 -1702 1157 -1622
rect 1091 -1714 1157 -1702
rect 1187 -1622 1253 -1610
rect 1187 -1702 1203 -1622
rect 1237 -1702 1253 -1622
rect 1187 -1714 1253 -1702
rect 1283 -1622 1349 -1610
rect 1283 -1702 1299 -1622
rect 1333 -1702 1349 -1622
rect 1283 -1714 1349 -1702
rect 1379 -1622 1441 -1610
rect 1379 -1702 1395 -1622
rect 1429 -1702 1441 -1622
rect 1379 -1714 1441 -1702
rect 1604 -1630 1662 -1618
rect 1604 -1706 1616 -1630
rect 1650 -1706 1662 -1630
rect 1604 -1718 1662 -1706
rect 1692 -1630 1750 -1618
rect 1692 -1706 1704 -1630
rect 1738 -1706 1750 -1630
rect 1692 -1718 1750 -1706
rect 1944 -1622 2006 -1610
rect 1944 -1702 1956 -1622
rect 1990 -1702 2006 -1622
rect 1944 -1714 2006 -1702
rect 2036 -1622 2102 -1610
rect 2036 -1702 2052 -1622
rect 2086 -1702 2102 -1622
rect 2036 -1714 2102 -1702
rect 2132 -1622 2198 -1610
rect 2132 -1702 2148 -1622
rect 2182 -1702 2198 -1622
rect 2132 -1714 2198 -1702
rect 2228 -1622 2294 -1610
rect 2228 -1702 2244 -1622
rect 2278 -1702 2294 -1622
rect 2228 -1714 2294 -1702
rect 2324 -1622 2390 -1610
rect 2324 -1702 2340 -1622
rect 2374 -1702 2390 -1622
rect 2324 -1714 2390 -1702
rect 2420 -1622 2486 -1610
rect 2420 -1702 2436 -1622
rect 2470 -1702 2486 -1622
rect 2420 -1714 2486 -1702
rect 2516 -1622 2582 -1610
rect 2516 -1702 2532 -1622
rect 2566 -1702 2582 -1622
rect 2516 -1714 2582 -1702
rect 2612 -1622 2678 -1610
rect 2612 -1702 2628 -1622
rect 2662 -1702 2678 -1622
rect 2612 -1714 2678 -1702
rect 2708 -1622 2774 -1610
rect 2708 -1702 2724 -1622
rect 2758 -1702 2774 -1622
rect 2708 -1714 2774 -1702
rect 2804 -1622 2870 -1610
rect 2804 -1702 2820 -1622
rect 2854 -1702 2870 -1622
rect 2804 -1714 2870 -1702
rect 2900 -1622 2962 -1610
rect 2900 -1702 2916 -1622
rect 2950 -1702 2962 -1622
rect 2900 -1714 2962 -1702
rect -3128 -2212 -3066 -2200
rect -3128 -2292 -3116 -2212
rect -3082 -2292 -3066 -2212
rect -3128 -2304 -3066 -2292
rect -3036 -2212 -2970 -2200
rect -3036 -2292 -3020 -2212
rect -2986 -2292 -2970 -2212
rect -3036 -2304 -2970 -2292
rect -2940 -2212 -2874 -2200
rect -2940 -2292 -2924 -2212
rect -2890 -2292 -2874 -2212
rect -2940 -2304 -2874 -2292
rect -2844 -2212 -2778 -2200
rect -2844 -2292 -2828 -2212
rect -2794 -2292 -2778 -2212
rect -2844 -2304 -2778 -2292
rect -2748 -2212 -2682 -2200
rect -2748 -2292 -2732 -2212
rect -2698 -2292 -2682 -2212
rect -2748 -2304 -2682 -2292
rect -2652 -2212 -2586 -2200
rect -2652 -2292 -2636 -2212
rect -2602 -2292 -2586 -2212
rect -2652 -2304 -2586 -2292
rect -2556 -2212 -2490 -2200
rect -2556 -2292 -2540 -2212
rect -2506 -2292 -2490 -2212
rect -2556 -2304 -2490 -2292
rect -2460 -2212 -2394 -2200
rect -2460 -2292 -2444 -2212
rect -2410 -2292 -2394 -2212
rect -2460 -2304 -2394 -2292
rect -2364 -2212 -2298 -2200
rect -2364 -2292 -2348 -2212
rect -2314 -2292 -2298 -2212
rect -2364 -2304 -2298 -2292
rect -2268 -2212 -2202 -2200
rect -2268 -2292 -2252 -2212
rect -2218 -2292 -2202 -2212
rect -2268 -2304 -2202 -2292
rect -2172 -2212 -2110 -2200
rect -2172 -2292 -2156 -2212
rect -2122 -2292 -2110 -2212
rect -2172 -2304 -2110 -2292
rect -1096 -2488 -1044 -2476
rect -1096 -2522 -1088 -2488
rect -1054 -2522 -1044 -2488
rect -1096 -2556 -1044 -2522
rect -1096 -2590 -1088 -2556
rect -1054 -2590 -1044 -2556
rect -1096 -2606 -1044 -2590
rect -1014 -2488 -962 -2476
rect -1014 -2522 -1004 -2488
rect -970 -2522 -962 -2488
rect -1014 -2556 -962 -2522
rect -1014 -2590 -1004 -2556
rect -970 -2590 -962 -2556
rect -581 -2492 -529 -2476
rect -581 -2526 -573 -2492
rect -539 -2526 -529 -2492
rect -581 -2560 -529 -2526
rect -1014 -2606 -962 -2590
rect -581 -2594 -573 -2560
rect -539 -2594 -529 -2560
rect -581 -2606 -529 -2594
rect -499 -2606 -445 -2476
rect -415 -2492 -363 -2476
rect -415 -2526 -405 -2492
rect -371 -2526 -363 -2492
rect -415 -2560 -363 -2526
rect -415 -2594 -405 -2560
rect -371 -2594 -363 -2560
rect -415 -2606 -363 -2594
rect -1096 -2716 -1044 -2700
rect -1096 -2750 -1088 -2716
rect -1054 -2750 -1044 -2716
rect -1096 -2784 -1044 -2750
rect -1096 -2818 -1088 -2784
rect -1054 -2818 -1044 -2784
rect -1096 -2830 -1044 -2818
rect -1014 -2716 -962 -2700
rect -1014 -2750 -1004 -2716
rect -970 -2750 -962 -2716
rect -581 -2712 -529 -2700
rect -1014 -2784 -962 -2750
rect -1014 -2818 -1004 -2784
rect -970 -2818 -962 -2784
rect -1014 -2830 -962 -2818
rect -581 -2746 -573 -2712
rect -539 -2746 -529 -2712
rect -581 -2780 -529 -2746
rect -581 -2814 -573 -2780
rect -539 -2814 -529 -2780
rect -581 -2830 -529 -2814
rect -499 -2830 -445 -2700
rect -415 -2712 -363 -2700
rect -415 -2746 -405 -2712
rect -371 -2746 -363 -2712
rect -415 -2780 -363 -2746
rect -415 -2814 -405 -2780
rect -371 -2814 -363 -2780
rect -415 -2830 -363 -2814
rect 423 -3000 485 -2988
rect 423 -3080 435 -3000
rect 469 -3080 485 -3000
rect 423 -3092 485 -3080
rect 515 -3000 581 -2988
rect 515 -3080 531 -3000
rect 565 -3080 581 -3000
rect 515 -3092 581 -3080
rect 611 -3000 677 -2988
rect 611 -3080 627 -3000
rect 661 -3080 677 -3000
rect 611 -3092 677 -3080
rect 707 -3000 773 -2988
rect 707 -3080 723 -3000
rect 757 -3080 773 -3000
rect 707 -3092 773 -3080
rect 803 -3000 869 -2988
rect 803 -3080 819 -3000
rect 853 -3080 869 -3000
rect 803 -3092 869 -3080
rect 899 -3000 965 -2988
rect 899 -3080 915 -3000
rect 949 -3080 965 -3000
rect 899 -3092 965 -3080
rect 995 -3000 1061 -2988
rect 995 -3080 1011 -3000
rect 1045 -3080 1061 -3000
rect 995 -3092 1061 -3080
rect 1091 -3000 1157 -2988
rect 1091 -3080 1107 -3000
rect 1141 -3080 1157 -3000
rect 1091 -3092 1157 -3080
rect 1187 -3000 1253 -2988
rect 1187 -3080 1203 -3000
rect 1237 -3080 1253 -3000
rect 1187 -3092 1253 -3080
rect 1283 -3000 1349 -2988
rect 1283 -3080 1299 -3000
rect 1333 -3080 1349 -3000
rect 1283 -3092 1349 -3080
rect 1379 -3000 1441 -2988
rect 1379 -3080 1395 -3000
rect 1429 -3080 1441 -3000
rect 1379 -3092 1441 -3080
rect 1604 -3008 1662 -2996
rect 1604 -3084 1616 -3008
rect 1650 -3084 1662 -3008
rect 1604 -3096 1662 -3084
rect 1692 -3008 1750 -2996
rect 1692 -3084 1704 -3008
rect 1738 -3084 1750 -3008
rect 1692 -3096 1750 -3084
rect 1944 -3000 2006 -2988
rect 1944 -3080 1956 -3000
rect 1990 -3080 2006 -3000
rect 1944 -3092 2006 -3080
rect 2036 -3000 2102 -2988
rect 2036 -3080 2052 -3000
rect 2086 -3080 2102 -3000
rect 2036 -3092 2102 -3080
rect 2132 -3000 2198 -2988
rect 2132 -3080 2148 -3000
rect 2182 -3080 2198 -3000
rect 2132 -3092 2198 -3080
rect 2228 -3000 2294 -2988
rect 2228 -3080 2244 -3000
rect 2278 -3080 2294 -3000
rect 2228 -3092 2294 -3080
rect 2324 -3000 2390 -2988
rect 2324 -3080 2340 -3000
rect 2374 -3080 2390 -3000
rect 2324 -3092 2390 -3080
rect 2420 -3000 2486 -2988
rect 2420 -3080 2436 -3000
rect 2470 -3080 2486 -3000
rect 2420 -3092 2486 -3080
rect 2516 -3000 2582 -2988
rect 2516 -3080 2532 -3000
rect 2566 -3080 2582 -3000
rect 2516 -3092 2582 -3080
rect 2612 -3000 2678 -2988
rect 2612 -3080 2628 -3000
rect 2662 -3080 2678 -3000
rect 2612 -3092 2678 -3080
rect 2708 -3000 2774 -2988
rect 2708 -3080 2724 -3000
rect 2758 -3080 2774 -3000
rect 2708 -3092 2774 -3080
rect 2804 -3000 2870 -2988
rect 2804 -3080 2820 -3000
rect 2854 -3080 2870 -3000
rect 2804 -3092 2870 -3080
rect 2900 -3000 2962 -2988
rect 2900 -3080 2916 -3000
rect 2950 -3080 2962 -3000
rect 2900 -3092 2962 -3080
rect -3128 -3590 -3066 -3578
rect -3128 -3670 -3116 -3590
rect -3082 -3670 -3066 -3590
rect -3128 -3682 -3066 -3670
rect -3036 -3590 -2970 -3578
rect -3036 -3670 -3020 -3590
rect -2986 -3670 -2970 -3590
rect -3036 -3682 -2970 -3670
rect -2940 -3590 -2874 -3578
rect -2940 -3670 -2924 -3590
rect -2890 -3670 -2874 -3590
rect -2940 -3682 -2874 -3670
rect -2844 -3590 -2778 -3578
rect -2844 -3670 -2828 -3590
rect -2794 -3670 -2778 -3590
rect -2844 -3682 -2778 -3670
rect -2748 -3590 -2682 -3578
rect -2748 -3670 -2732 -3590
rect -2698 -3670 -2682 -3590
rect -2748 -3682 -2682 -3670
rect -2652 -3590 -2586 -3578
rect -2652 -3670 -2636 -3590
rect -2602 -3670 -2586 -3590
rect -2652 -3682 -2586 -3670
rect -2556 -3590 -2490 -3578
rect -2556 -3670 -2540 -3590
rect -2506 -3670 -2490 -3590
rect -2556 -3682 -2490 -3670
rect -2460 -3590 -2394 -3578
rect -2460 -3670 -2444 -3590
rect -2410 -3670 -2394 -3590
rect -2460 -3682 -2394 -3670
rect -2364 -3590 -2298 -3578
rect -2364 -3670 -2348 -3590
rect -2314 -3670 -2298 -3590
rect -2364 -3682 -2298 -3670
rect -2268 -3590 -2202 -3578
rect -2268 -3670 -2252 -3590
rect -2218 -3670 -2202 -3590
rect -2268 -3682 -2202 -3670
rect -2172 -3590 -2110 -3578
rect -2172 -3670 -2156 -3590
rect -2122 -3670 -2110 -3590
rect -2172 -3682 -2110 -3670
rect -581 -3580 -529 -3564
rect -581 -3614 -573 -3580
rect -539 -3614 -529 -3580
rect -581 -3648 -529 -3614
rect -581 -3682 -573 -3648
rect -539 -3682 -529 -3648
rect -581 -3694 -529 -3682
rect -499 -3694 -445 -3564
rect -415 -3580 -363 -3564
rect -415 -3614 -405 -3580
rect -371 -3614 -363 -3580
rect -415 -3648 -363 -3614
rect -415 -3682 -405 -3648
rect -371 -3682 -363 -3648
rect -415 -3694 -363 -3682
rect -544 -3804 -492 -3788
rect -544 -3838 -536 -3804
rect -502 -3838 -492 -3804
rect -544 -3872 -492 -3838
rect -544 -3906 -536 -3872
rect -502 -3906 -492 -3872
rect -544 -3918 -492 -3906
rect -462 -3804 -410 -3788
rect -462 -3838 -452 -3804
rect -418 -3838 -410 -3804
rect -462 -3872 -410 -3838
rect -462 -3906 -452 -3872
rect -418 -3906 -410 -3872
rect -462 -3918 -410 -3906
rect 423 -4378 485 -4366
rect 423 -4458 435 -4378
rect 469 -4458 485 -4378
rect 423 -4470 485 -4458
rect 515 -4378 581 -4366
rect 515 -4458 531 -4378
rect 565 -4458 581 -4378
rect 515 -4470 581 -4458
rect 611 -4378 677 -4366
rect 611 -4458 627 -4378
rect 661 -4458 677 -4378
rect 611 -4470 677 -4458
rect 707 -4378 773 -4366
rect 707 -4458 723 -4378
rect 757 -4458 773 -4378
rect 707 -4470 773 -4458
rect 803 -4378 869 -4366
rect 803 -4458 819 -4378
rect 853 -4458 869 -4378
rect 803 -4470 869 -4458
rect 899 -4378 965 -4366
rect 899 -4458 915 -4378
rect 949 -4458 965 -4378
rect 899 -4470 965 -4458
rect 995 -4378 1061 -4366
rect 995 -4458 1011 -4378
rect 1045 -4458 1061 -4378
rect 995 -4470 1061 -4458
rect 1091 -4378 1157 -4366
rect 1091 -4458 1107 -4378
rect 1141 -4458 1157 -4378
rect 1091 -4470 1157 -4458
rect 1187 -4378 1253 -4366
rect 1187 -4458 1203 -4378
rect 1237 -4458 1253 -4378
rect 1187 -4470 1253 -4458
rect 1283 -4378 1349 -4366
rect 1283 -4458 1299 -4378
rect 1333 -4458 1349 -4378
rect 1283 -4470 1349 -4458
rect 1379 -4378 1441 -4366
rect 1379 -4458 1395 -4378
rect 1429 -4458 1441 -4378
rect 1379 -4470 1441 -4458
rect 1604 -4386 1662 -4374
rect 1604 -4462 1616 -4386
rect 1650 -4462 1662 -4386
rect 1604 -4474 1662 -4462
rect 1692 -4386 1750 -4374
rect 1692 -4462 1704 -4386
rect 1738 -4462 1750 -4386
rect 1692 -4474 1750 -4462
rect 1944 -4378 2006 -4366
rect 1944 -4458 1956 -4378
rect 1990 -4458 2006 -4378
rect 1944 -4470 2006 -4458
rect 2036 -4378 2102 -4366
rect 2036 -4458 2052 -4378
rect 2086 -4458 2102 -4378
rect 2036 -4470 2102 -4458
rect 2132 -4378 2198 -4366
rect 2132 -4458 2148 -4378
rect 2182 -4458 2198 -4378
rect 2132 -4470 2198 -4458
rect 2228 -4378 2294 -4366
rect 2228 -4458 2244 -4378
rect 2278 -4458 2294 -4378
rect 2228 -4470 2294 -4458
rect 2324 -4378 2390 -4366
rect 2324 -4458 2340 -4378
rect 2374 -4458 2390 -4378
rect 2324 -4470 2390 -4458
rect 2420 -4378 2486 -4366
rect 2420 -4458 2436 -4378
rect 2470 -4458 2486 -4378
rect 2420 -4470 2486 -4458
rect 2516 -4378 2582 -4366
rect 2516 -4458 2532 -4378
rect 2566 -4458 2582 -4378
rect 2516 -4470 2582 -4458
rect 2612 -4378 2678 -4366
rect 2612 -4458 2628 -4378
rect 2662 -4458 2678 -4378
rect 2612 -4470 2678 -4458
rect 2708 -4378 2774 -4366
rect 2708 -4458 2724 -4378
rect 2758 -4458 2774 -4378
rect 2708 -4470 2774 -4458
rect 2804 -4378 2870 -4366
rect 2804 -4458 2820 -4378
rect 2854 -4458 2870 -4378
rect 2804 -4470 2870 -4458
rect 2900 -4378 2962 -4366
rect 2900 -4458 2916 -4378
rect 2950 -4458 2962 -4378
rect 2900 -4470 2962 -4458
rect -544 -4664 -492 -4652
rect -544 -4698 -536 -4664
rect -502 -4698 -492 -4664
rect -544 -4732 -492 -4698
rect -544 -4766 -536 -4732
rect -502 -4766 -492 -4732
rect -544 -4782 -492 -4766
rect -462 -4664 -410 -4652
rect -462 -4698 -452 -4664
rect -418 -4698 -410 -4664
rect -462 -4732 -410 -4698
rect -462 -4766 -452 -4732
rect -418 -4766 -410 -4732
rect -462 -4782 -410 -4766
rect -3128 -4968 -3066 -4956
rect -3128 -5048 -3116 -4968
rect -3082 -5048 -3066 -4968
rect -3128 -5060 -3066 -5048
rect -3036 -4968 -2970 -4956
rect -3036 -5048 -3020 -4968
rect -2986 -5048 -2970 -4968
rect -3036 -5060 -2970 -5048
rect -2940 -4968 -2874 -4956
rect -2940 -5048 -2924 -4968
rect -2890 -5048 -2874 -4968
rect -2940 -5060 -2874 -5048
rect -2844 -4968 -2778 -4956
rect -2844 -5048 -2828 -4968
rect -2794 -5048 -2778 -4968
rect -2844 -5060 -2778 -5048
rect -2748 -4968 -2682 -4956
rect -2748 -5048 -2732 -4968
rect -2698 -5048 -2682 -4968
rect -2748 -5060 -2682 -5048
rect -2652 -4968 -2586 -4956
rect -2652 -5048 -2636 -4968
rect -2602 -5048 -2586 -4968
rect -2652 -5060 -2586 -5048
rect -2556 -4968 -2490 -4956
rect -2556 -5048 -2540 -4968
rect -2506 -5048 -2490 -4968
rect -2556 -5060 -2490 -5048
rect -2460 -4968 -2394 -4956
rect -2460 -5048 -2444 -4968
rect -2410 -5048 -2394 -4968
rect -2460 -5060 -2394 -5048
rect -2364 -4968 -2298 -4956
rect -2364 -5048 -2348 -4968
rect -2314 -5048 -2298 -4968
rect -2364 -5060 -2298 -5048
rect -2268 -4968 -2202 -4956
rect -2268 -5048 -2252 -4968
rect -2218 -5048 -2202 -4968
rect -2268 -5060 -2202 -5048
rect -2172 -4968 -2110 -4956
rect -2172 -5048 -2156 -4968
rect -2122 -5048 -2110 -4968
rect -2172 -5060 -2110 -5048
<< pdiff >>
rect -3128 -298 -3066 -286
rect -3128 -546 -3116 -298
rect -3082 -546 -3066 -298
rect -3128 -558 -3066 -546
rect -3036 -298 -2970 -286
rect -3036 -546 -3020 -298
rect -2986 -546 -2970 -298
rect -3036 -558 -2970 -546
rect -2940 -298 -2874 -286
rect -2940 -546 -2924 -298
rect -2890 -546 -2874 -298
rect -2940 -558 -2874 -546
rect -2844 -298 -2778 -286
rect -2844 -546 -2828 -298
rect -2794 -546 -2778 -298
rect -2844 -558 -2778 -546
rect -2748 -298 -2682 -286
rect -2748 -546 -2732 -298
rect -2698 -546 -2682 -298
rect -2748 -558 -2682 -546
rect -2652 -298 -2586 -286
rect -2652 -546 -2636 -298
rect -2602 -546 -2586 -298
rect -2652 -558 -2586 -546
rect -2556 -298 -2490 -286
rect -2556 -546 -2540 -298
rect -2506 -546 -2490 -298
rect -2556 -558 -2490 -546
rect -2460 -298 -2394 -286
rect -2460 -546 -2444 -298
rect -2410 -546 -2394 -298
rect -2460 -558 -2394 -546
rect -2364 -298 -2298 -286
rect -2364 -546 -2348 -298
rect -2314 -546 -2298 -298
rect -2364 -558 -2298 -546
rect -2268 -298 -2202 -286
rect -2268 -546 -2252 -298
rect -2218 -546 -2202 -298
rect -2268 -558 -2202 -546
rect -2172 -298 -2110 -286
rect -2172 -546 -2156 -298
rect -2122 -546 -2110 -298
rect -2172 -558 -2110 -546
rect -912 -792 -860 -774
rect -912 -826 -904 -792
rect -870 -826 -860 -792
rect -912 -860 -860 -826
rect -912 -894 -904 -860
rect -870 -894 -860 -860
rect -912 -928 -860 -894
rect -912 -962 -904 -928
rect -870 -962 -860 -928
rect -912 -974 -860 -962
rect -830 -792 -778 -774
rect -830 -826 -820 -792
rect -786 -826 -778 -792
rect -830 -860 -778 -826
rect -830 -894 -820 -860
rect -786 -894 -778 -860
rect -830 -928 -778 -894
rect -830 -962 -820 -928
rect -786 -962 -778 -928
rect -544 -792 -492 -774
rect -544 -826 -536 -792
rect -502 -826 -492 -792
rect -544 -860 -492 -826
rect -544 -894 -536 -860
rect -502 -894 -492 -860
rect -544 -928 -492 -894
rect -830 -974 -778 -962
rect -544 -962 -536 -928
rect -502 -962 -492 -928
rect -544 -974 -492 -962
rect -462 -792 -410 -774
rect -462 -826 -452 -792
rect -418 -826 -410 -792
rect -462 -860 -410 -826
rect -462 -894 -452 -860
rect -418 -894 -410 -860
rect -462 -928 -410 -894
rect -462 -962 -452 -928
rect -418 -962 -410 -928
rect -462 -974 -410 -962
rect 423 -700 485 -688
rect 423 -948 435 -700
rect 469 -948 485 -700
rect 423 -960 485 -948
rect 515 -700 581 -688
rect 515 -948 531 -700
rect 565 -948 581 -700
rect 515 -960 581 -948
rect 611 -700 677 -688
rect 611 -948 627 -700
rect 661 -948 677 -700
rect 611 -960 677 -948
rect 707 -700 773 -688
rect 707 -948 723 -700
rect 757 -948 773 -700
rect 707 -960 773 -948
rect 803 -700 869 -688
rect 803 -948 819 -700
rect 853 -948 869 -700
rect 803 -960 869 -948
rect 899 -700 965 -688
rect 899 -948 915 -700
rect 949 -948 965 -700
rect 899 -960 965 -948
rect 995 -700 1061 -688
rect 995 -948 1011 -700
rect 1045 -948 1061 -700
rect 995 -960 1061 -948
rect 1091 -700 1157 -688
rect 1091 -948 1107 -700
rect 1141 -948 1157 -700
rect 1091 -960 1157 -948
rect 1187 -700 1253 -688
rect 1187 -948 1203 -700
rect 1237 -948 1253 -700
rect 1187 -960 1253 -948
rect 1283 -700 1349 -688
rect 1283 -948 1299 -700
rect 1333 -948 1349 -700
rect 1283 -960 1349 -948
rect 1379 -700 1441 -688
rect 1379 -948 1395 -700
rect 1429 -948 1441 -700
rect 1379 -960 1441 -948
rect -544 -1080 -492 -1068
rect -544 -1114 -536 -1080
rect -502 -1114 -492 -1080
rect -544 -1148 -492 -1114
rect -544 -1182 -536 -1148
rect -502 -1182 -492 -1148
rect -544 -1216 -492 -1182
rect -544 -1250 -536 -1216
rect -502 -1250 -492 -1216
rect -544 -1268 -492 -1250
rect -462 -1080 -410 -1068
rect -462 -1114 -452 -1080
rect -418 -1114 -410 -1080
rect -462 -1148 -410 -1114
rect 1944 -700 2006 -688
rect 1944 -948 1956 -700
rect 1990 -948 2006 -700
rect 1944 -960 2006 -948
rect 2036 -700 2102 -688
rect 2036 -948 2052 -700
rect 2086 -948 2102 -700
rect 2036 -960 2102 -948
rect 2132 -700 2198 -688
rect 2132 -948 2148 -700
rect 2182 -948 2198 -700
rect 2132 -960 2198 -948
rect 2228 -700 2294 -688
rect 2228 -948 2244 -700
rect 2278 -948 2294 -700
rect 2228 -960 2294 -948
rect 2324 -700 2390 -688
rect 2324 -948 2340 -700
rect 2374 -948 2390 -700
rect 2324 -960 2390 -948
rect 2420 -700 2486 -688
rect 2420 -948 2436 -700
rect 2470 -948 2486 -700
rect 2420 -960 2486 -948
rect 2516 -700 2582 -688
rect 2516 -948 2532 -700
rect 2566 -948 2582 -700
rect 2516 -960 2582 -948
rect 2612 -700 2678 -688
rect 2612 -948 2628 -700
rect 2662 -948 2678 -700
rect 2612 -960 2678 -948
rect 2708 -700 2774 -688
rect 2708 -948 2724 -700
rect 2758 -948 2774 -700
rect 2708 -960 2774 -948
rect 2804 -700 2870 -688
rect 2804 -948 2820 -700
rect 2854 -948 2870 -700
rect 2804 -960 2870 -948
rect 2900 -700 2962 -688
rect 2900 -948 2916 -700
rect 2950 -948 2962 -700
rect 2900 -960 2962 -948
rect -462 -1182 -452 -1148
rect -418 -1182 -410 -1148
rect -462 -1216 -410 -1182
rect -462 -1250 -452 -1216
rect -418 -1250 -410 -1216
rect -462 -1268 -410 -1250
rect -3128 -1632 -3066 -1620
rect -3128 -1880 -3116 -1632
rect -3082 -1880 -3066 -1632
rect -3128 -1892 -3066 -1880
rect -3036 -1632 -2970 -1620
rect -3036 -1880 -3020 -1632
rect -2986 -1880 -2970 -1632
rect -3036 -1892 -2970 -1880
rect -2940 -1632 -2874 -1620
rect -2940 -1880 -2924 -1632
rect -2890 -1880 -2874 -1632
rect -2940 -1892 -2874 -1880
rect -2844 -1632 -2778 -1620
rect -2844 -1880 -2828 -1632
rect -2794 -1880 -2778 -1632
rect -2844 -1892 -2778 -1880
rect -2748 -1632 -2682 -1620
rect -2748 -1880 -2732 -1632
rect -2698 -1880 -2682 -1632
rect -2748 -1892 -2682 -1880
rect -2652 -1632 -2586 -1620
rect -2652 -1880 -2636 -1632
rect -2602 -1880 -2586 -1632
rect -2652 -1892 -2586 -1880
rect -2556 -1632 -2490 -1620
rect -2556 -1880 -2540 -1632
rect -2506 -1880 -2490 -1632
rect -2556 -1892 -2490 -1880
rect -2460 -1632 -2394 -1620
rect -2460 -1880 -2444 -1632
rect -2410 -1880 -2394 -1632
rect -2460 -1892 -2394 -1880
rect -2364 -1632 -2298 -1620
rect -2364 -1880 -2348 -1632
rect -2314 -1880 -2298 -1632
rect -2364 -1892 -2298 -1880
rect -2268 -1632 -2202 -1620
rect -2268 -1880 -2252 -1632
rect -2218 -1880 -2202 -1632
rect -2268 -1892 -2202 -1880
rect -2172 -1632 -2110 -1620
rect -2172 -1880 -2156 -1632
rect -2122 -1880 -2110 -1632
rect -2172 -1892 -2110 -1880
rect -581 -1880 -529 -1862
rect -581 -1914 -573 -1880
rect -539 -1914 -529 -1880
rect -581 -1948 -529 -1914
rect -581 -1982 -573 -1948
rect -539 -1982 -529 -1948
rect -581 -2016 -529 -1982
rect -581 -2050 -573 -2016
rect -539 -2050 -529 -2016
rect -581 -2062 -529 -2050
rect -499 -1880 -445 -1862
rect -499 -1914 -489 -1880
rect -455 -1914 -445 -1880
rect -499 -1948 -445 -1914
rect -499 -1982 -489 -1948
rect -455 -1982 -445 -1948
rect -499 -2016 -445 -1982
rect -499 -2050 -489 -2016
rect -455 -2050 -445 -2016
rect -499 -2062 -445 -2050
rect -415 -1880 -363 -1862
rect -415 -1914 -405 -1880
rect -371 -1914 -363 -1880
rect -415 -1948 -363 -1914
rect -415 -1982 -405 -1948
rect -371 -1982 -363 -1948
rect -415 -2016 -363 -1982
rect -415 -2050 -405 -2016
rect -371 -2050 -363 -2016
rect -415 -2062 -363 -2050
rect -1096 -2168 -1044 -2156
rect -1096 -2202 -1088 -2168
rect -1054 -2202 -1044 -2168
rect -1096 -2236 -1044 -2202
rect -1096 -2270 -1088 -2236
rect -1054 -2270 -1044 -2236
rect -1096 -2304 -1044 -2270
rect -1096 -2338 -1088 -2304
rect -1054 -2338 -1044 -2304
rect -1096 -2356 -1044 -2338
rect -1014 -2168 -962 -2156
rect -1014 -2202 -1004 -2168
rect -970 -2202 -962 -2168
rect -581 -2168 -529 -2156
rect -1014 -2236 -962 -2202
rect -1014 -2270 -1004 -2236
rect -970 -2270 -962 -2236
rect -1014 -2304 -962 -2270
rect -1014 -2338 -1004 -2304
rect -970 -2338 -962 -2304
rect -1014 -2356 -962 -2338
rect -581 -2202 -573 -2168
rect -539 -2202 -529 -2168
rect -581 -2236 -529 -2202
rect -581 -2270 -573 -2236
rect -539 -2270 -529 -2236
rect -581 -2304 -529 -2270
rect -581 -2338 -573 -2304
rect -539 -2338 -529 -2304
rect -581 -2356 -529 -2338
rect -499 -2168 -445 -2156
rect -499 -2202 -489 -2168
rect -455 -2202 -445 -2168
rect -499 -2236 -445 -2202
rect -499 -2270 -489 -2236
rect -455 -2270 -445 -2236
rect -499 -2304 -445 -2270
rect -499 -2338 -489 -2304
rect -455 -2338 -445 -2304
rect -499 -2356 -445 -2338
rect -415 -2168 -363 -2156
rect -415 -2202 -405 -2168
rect -371 -2202 -363 -2168
rect -415 -2236 -363 -2202
rect -415 -2270 -405 -2236
rect -371 -2270 -363 -2236
rect -415 -2304 -363 -2270
rect -415 -2338 -405 -2304
rect -371 -2338 -363 -2304
rect -415 -2356 -363 -2338
rect 423 -2034 485 -2022
rect 423 -2282 435 -2034
rect 469 -2282 485 -2034
rect 423 -2294 485 -2282
rect 515 -2034 581 -2022
rect 515 -2282 531 -2034
rect 565 -2282 581 -2034
rect 515 -2294 581 -2282
rect 611 -2034 677 -2022
rect 611 -2282 627 -2034
rect 661 -2282 677 -2034
rect 611 -2294 677 -2282
rect 707 -2034 773 -2022
rect 707 -2282 723 -2034
rect 757 -2282 773 -2034
rect 707 -2294 773 -2282
rect 803 -2034 869 -2022
rect 803 -2282 819 -2034
rect 853 -2282 869 -2034
rect 803 -2294 869 -2282
rect 899 -2034 965 -2022
rect 899 -2282 915 -2034
rect 949 -2282 965 -2034
rect 899 -2294 965 -2282
rect 995 -2034 1061 -2022
rect 995 -2282 1011 -2034
rect 1045 -2282 1061 -2034
rect 995 -2294 1061 -2282
rect 1091 -2034 1157 -2022
rect 1091 -2282 1107 -2034
rect 1141 -2282 1157 -2034
rect 1091 -2294 1157 -2282
rect 1187 -2034 1253 -2022
rect 1187 -2282 1203 -2034
rect 1237 -2282 1253 -2034
rect 1187 -2294 1253 -2282
rect 1283 -2034 1349 -2022
rect 1283 -2282 1299 -2034
rect 1333 -2282 1349 -2034
rect 1283 -2294 1349 -2282
rect 1379 -2034 1441 -2022
rect 1379 -2282 1395 -2034
rect 1429 -2282 1441 -2034
rect 1379 -2294 1441 -2282
rect 1944 -2034 2006 -2022
rect 1944 -2282 1956 -2034
rect 1990 -2282 2006 -2034
rect 1944 -2294 2006 -2282
rect 2036 -2034 2102 -2022
rect 2036 -2282 2052 -2034
rect 2086 -2282 2102 -2034
rect 2036 -2294 2102 -2282
rect 2132 -2034 2198 -2022
rect 2132 -2282 2148 -2034
rect 2182 -2282 2198 -2034
rect 2132 -2294 2198 -2282
rect 2228 -2034 2294 -2022
rect 2228 -2282 2244 -2034
rect 2278 -2282 2294 -2034
rect 2228 -2294 2294 -2282
rect 2324 -2034 2390 -2022
rect 2324 -2282 2340 -2034
rect 2374 -2282 2390 -2034
rect 2324 -2294 2390 -2282
rect 2420 -2034 2486 -2022
rect 2420 -2282 2436 -2034
rect 2470 -2282 2486 -2034
rect 2420 -2294 2486 -2282
rect 2516 -2034 2582 -2022
rect 2516 -2282 2532 -2034
rect 2566 -2282 2582 -2034
rect 2516 -2294 2582 -2282
rect 2612 -2034 2678 -2022
rect 2612 -2282 2628 -2034
rect 2662 -2282 2678 -2034
rect 2612 -2294 2678 -2282
rect 2708 -2034 2774 -2022
rect 2708 -2282 2724 -2034
rect 2758 -2282 2774 -2034
rect 2708 -2294 2774 -2282
rect 2804 -2034 2870 -2022
rect 2804 -2282 2820 -2034
rect 2854 -2282 2870 -2034
rect 2804 -2294 2870 -2282
rect 2900 -2034 2962 -2022
rect 2900 -2282 2916 -2034
rect 2950 -2282 2962 -2034
rect 2900 -2294 2962 -2282
rect -3128 -3010 -3066 -2998
rect -3128 -3258 -3116 -3010
rect -3082 -3258 -3066 -3010
rect -3128 -3270 -3066 -3258
rect -3036 -3010 -2970 -2998
rect -3036 -3258 -3020 -3010
rect -2986 -3258 -2970 -3010
rect -3036 -3270 -2970 -3258
rect -2940 -3010 -2874 -2998
rect -2940 -3258 -2924 -3010
rect -2890 -3258 -2874 -3010
rect -2940 -3270 -2874 -3258
rect -2844 -3010 -2778 -2998
rect -2844 -3258 -2828 -3010
rect -2794 -3258 -2778 -3010
rect -2844 -3270 -2778 -3258
rect -2748 -3010 -2682 -2998
rect -2748 -3258 -2732 -3010
rect -2698 -3258 -2682 -3010
rect -2748 -3270 -2682 -3258
rect -2652 -3010 -2586 -2998
rect -2652 -3258 -2636 -3010
rect -2602 -3258 -2586 -3010
rect -2652 -3270 -2586 -3258
rect -2556 -3010 -2490 -2998
rect -2556 -3258 -2540 -3010
rect -2506 -3258 -2490 -3010
rect -2556 -3270 -2490 -3258
rect -2460 -3010 -2394 -2998
rect -2460 -3258 -2444 -3010
rect -2410 -3258 -2394 -3010
rect -2460 -3270 -2394 -3258
rect -2364 -3010 -2298 -2998
rect -2364 -3258 -2348 -3010
rect -2314 -3258 -2298 -3010
rect -2364 -3270 -2298 -3258
rect -2268 -3010 -2202 -2998
rect -2268 -3258 -2252 -3010
rect -2218 -3258 -2202 -3010
rect -2268 -3270 -2202 -3258
rect -2172 -3010 -2110 -2998
rect -2172 -3258 -2156 -3010
rect -2122 -3258 -2110 -3010
rect -2172 -3270 -2110 -3258
rect -1096 -2968 -1044 -2950
rect -1096 -3002 -1088 -2968
rect -1054 -3002 -1044 -2968
rect -1096 -3036 -1044 -3002
rect -1096 -3070 -1088 -3036
rect -1054 -3070 -1044 -3036
rect -1096 -3104 -1044 -3070
rect -1096 -3138 -1088 -3104
rect -1054 -3138 -1044 -3104
rect -1096 -3150 -1044 -3138
rect -1014 -2968 -962 -2950
rect -1014 -3002 -1004 -2968
rect -970 -3002 -962 -2968
rect -1014 -3036 -962 -3002
rect -1014 -3070 -1004 -3036
rect -970 -3070 -962 -3036
rect -1014 -3104 -962 -3070
rect -1014 -3138 -1004 -3104
rect -970 -3138 -962 -3104
rect -581 -2968 -529 -2950
rect -581 -3002 -573 -2968
rect -539 -3002 -529 -2968
rect -581 -3036 -529 -3002
rect -581 -3070 -573 -3036
rect -539 -3070 -529 -3036
rect -581 -3104 -529 -3070
rect -1014 -3150 -962 -3138
rect -581 -3138 -573 -3104
rect -539 -3138 -529 -3104
rect -581 -3150 -529 -3138
rect -499 -2968 -445 -2950
rect -499 -3002 -489 -2968
rect -455 -3002 -445 -2968
rect -499 -3036 -445 -3002
rect -499 -3070 -489 -3036
rect -455 -3070 -445 -3036
rect -499 -3104 -445 -3070
rect -499 -3138 -489 -3104
rect -455 -3138 -445 -3104
rect -499 -3150 -445 -3138
rect -415 -2968 -363 -2950
rect -415 -3002 -405 -2968
rect -371 -3002 -363 -2968
rect -415 -3036 -363 -3002
rect -415 -3070 -405 -3036
rect -371 -3070 -363 -3036
rect -415 -3104 -363 -3070
rect -415 -3138 -405 -3104
rect -371 -3138 -363 -3104
rect -415 -3150 -363 -3138
rect -581 -3256 -529 -3244
rect -581 -3290 -573 -3256
rect -539 -3290 -529 -3256
rect -581 -3324 -529 -3290
rect -581 -3358 -573 -3324
rect -539 -3358 -529 -3324
rect -581 -3392 -529 -3358
rect -581 -3426 -573 -3392
rect -539 -3426 -529 -3392
rect -581 -3444 -529 -3426
rect -499 -3256 -445 -3244
rect -499 -3290 -489 -3256
rect -455 -3290 -445 -3256
rect -499 -3324 -445 -3290
rect -499 -3358 -489 -3324
rect -455 -3358 -445 -3324
rect -499 -3392 -445 -3358
rect -499 -3426 -489 -3392
rect -455 -3426 -445 -3392
rect -499 -3444 -445 -3426
rect -415 -3256 -363 -3244
rect -415 -3290 -405 -3256
rect -371 -3290 -363 -3256
rect -415 -3324 -363 -3290
rect -415 -3358 -405 -3324
rect -371 -3358 -363 -3324
rect -415 -3392 -363 -3358
rect -415 -3426 -405 -3392
rect -371 -3426 -363 -3392
rect -415 -3444 -363 -3426
rect 423 -3412 485 -3400
rect 423 -3660 435 -3412
rect 469 -3660 485 -3412
rect 423 -3672 485 -3660
rect 515 -3412 581 -3400
rect 515 -3660 531 -3412
rect 565 -3660 581 -3412
rect 515 -3672 581 -3660
rect 611 -3412 677 -3400
rect 611 -3660 627 -3412
rect 661 -3660 677 -3412
rect 611 -3672 677 -3660
rect 707 -3412 773 -3400
rect 707 -3660 723 -3412
rect 757 -3660 773 -3412
rect 707 -3672 773 -3660
rect 803 -3412 869 -3400
rect 803 -3660 819 -3412
rect 853 -3660 869 -3412
rect 803 -3672 869 -3660
rect 899 -3412 965 -3400
rect 899 -3660 915 -3412
rect 949 -3660 965 -3412
rect 899 -3672 965 -3660
rect 995 -3412 1061 -3400
rect 995 -3660 1011 -3412
rect 1045 -3660 1061 -3412
rect 995 -3672 1061 -3660
rect 1091 -3412 1157 -3400
rect 1091 -3660 1107 -3412
rect 1141 -3660 1157 -3412
rect 1091 -3672 1157 -3660
rect 1187 -3412 1253 -3400
rect 1187 -3660 1203 -3412
rect 1237 -3660 1253 -3412
rect 1187 -3672 1253 -3660
rect 1283 -3412 1349 -3400
rect 1283 -3660 1299 -3412
rect 1333 -3660 1349 -3412
rect 1283 -3672 1349 -3660
rect 1379 -3412 1441 -3400
rect 1379 -3660 1395 -3412
rect 1429 -3660 1441 -3412
rect 1379 -3672 1441 -3660
rect 1944 -3412 2006 -3400
rect 1944 -3660 1956 -3412
rect 1990 -3660 2006 -3412
rect 1944 -3672 2006 -3660
rect 2036 -3412 2102 -3400
rect 2036 -3660 2052 -3412
rect 2086 -3660 2102 -3412
rect 2036 -3672 2102 -3660
rect 2132 -3412 2198 -3400
rect 2132 -3660 2148 -3412
rect 2182 -3660 2198 -3412
rect 2132 -3672 2198 -3660
rect 2228 -3412 2294 -3400
rect 2228 -3660 2244 -3412
rect 2278 -3660 2294 -3412
rect 2228 -3672 2294 -3660
rect 2324 -3412 2390 -3400
rect 2324 -3660 2340 -3412
rect 2374 -3660 2390 -3412
rect 2324 -3672 2390 -3660
rect 2420 -3412 2486 -3400
rect 2420 -3660 2436 -3412
rect 2470 -3660 2486 -3412
rect 2420 -3672 2486 -3660
rect 2516 -3412 2582 -3400
rect 2516 -3660 2532 -3412
rect 2566 -3660 2582 -3412
rect 2516 -3672 2582 -3660
rect 2612 -3412 2678 -3400
rect 2612 -3660 2628 -3412
rect 2662 -3660 2678 -3412
rect 2612 -3672 2678 -3660
rect 2708 -3412 2774 -3400
rect 2708 -3660 2724 -3412
rect 2758 -3660 2774 -3412
rect 2708 -3672 2774 -3660
rect 2804 -3412 2870 -3400
rect 2804 -3660 2820 -3412
rect 2854 -3660 2870 -3412
rect 2804 -3672 2870 -3660
rect 2900 -3412 2962 -3400
rect 2900 -3660 2916 -3412
rect 2950 -3660 2962 -3412
rect 2900 -3672 2962 -3660
rect -544 -4056 -492 -4038
rect -544 -4090 -536 -4056
rect -502 -4090 -492 -4056
rect -544 -4124 -492 -4090
rect -544 -4158 -536 -4124
rect -502 -4158 -492 -4124
rect -544 -4192 -492 -4158
rect -544 -4226 -536 -4192
rect -502 -4226 -492 -4192
rect -544 -4238 -492 -4226
rect -462 -4056 -410 -4038
rect -462 -4090 -452 -4056
rect -418 -4090 -410 -4056
rect -462 -4124 -410 -4090
rect -462 -4158 -452 -4124
rect -418 -4158 -410 -4124
rect -462 -4192 -410 -4158
rect -462 -4226 -452 -4192
rect -418 -4226 -410 -4192
rect -462 -4238 -410 -4226
rect -3128 -4388 -3066 -4376
rect -3128 -4636 -3116 -4388
rect -3082 -4636 -3066 -4388
rect -3128 -4648 -3066 -4636
rect -3036 -4388 -2970 -4376
rect -3036 -4636 -3020 -4388
rect -2986 -4636 -2970 -4388
rect -3036 -4648 -2970 -4636
rect -2940 -4388 -2874 -4376
rect -2940 -4636 -2924 -4388
rect -2890 -4636 -2874 -4388
rect -2940 -4648 -2874 -4636
rect -2844 -4388 -2778 -4376
rect -2844 -4636 -2828 -4388
rect -2794 -4636 -2778 -4388
rect -2844 -4648 -2778 -4636
rect -2748 -4388 -2682 -4376
rect -2748 -4636 -2732 -4388
rect -2698 -4636 -2682 -4388
rect -2748 -4648 -2682 -4636
rect -2652 -4388 -2586 -4376
rect -2652 -4636 -2636 -4388
rect -2602 -4636 -2586 -4388
rect -2652 -4648 -2586 -4636
rect -2556 -4388 -2490 -4376
rect -2556 -4636 -2540 -4388
rect -2506 -4636 -2490 -4388
rect -2556 -4648 -2490 -4636
rect -2460 -4388 -2394 -4376
rect -2460 -4636 -2444 -4388
rect -2410 -4636 -2394 -4388
rect -2460 -4648 -2394 -4636
rect -2364 -4388 -2298 -4376
rect -2364 -4636 -2348 -4388
rect -2314 -4636 -2298 -4388
rect -2364 -4648 -2298 -4636
rect -2268 -4388 -2202 -4376
rect -2268 -4636 -2252 -4388
rect -2218 -4636 -2202 -4388
rect -2268 -4648 -2202 -4636
rect -2172 -4388 -2110 -4376
rect -2172 -4636 -2156 -4388
rect -2122 -4636 -2110 -4388
rect -2172 -4648 -2110 -4636
rect -544 -4344 -492 -4332
rect -544 -4378 -536 -4344
rect -502 -4378 -492 -4344
rect -544 -4412 -492 -4378
rect -544 -4446 -536 -4412
rect -502 -4446 -492 -4412
rect -544 -4480 -492 -4446
rect -544 -4514 -536 -4480
rect -502 -4514 -492 -4480
rect -544 -4532 -492 -4514
rect -462 -4344 -410 -4332
rect -462 -4378 -452 -4344
rect -418 -4378 -410 -4344
rect -462 -4412 -410 -4378
rect -462 -4446 -452 -4412
rect -418 -4446 -410 -4412
rect -462 -4480 -410 -4446
rect -462 -4514 -452 -4480
rect -418 -4514 -410 -4480
rect -462 -4532 -410 -4514
rect 423 -4790 485 -4778
rect 423 -5038 435 -4790
rect 469 -5038 485 -4790
rect 423 -5050 485 -5038
rect 515 -4790 581 -4778
rect 515 -5038 531 -4790
rect 565 -5038 581 -4790
rect 515 -5050 581 -5038
rect 611 -4790 677 -4778
rect 611 -5038 627 -4790
rect 661 -5038 677 -4790
rect 611 -5050 677 -5038
rect 707 -4790 773 -4778
rect 707 -5038 723 -4790
rect 757 -5038 773 -4790
rect 707 -5050 773 -5038
rect 803 -4790 869 -4778
rect 803 -5038 819 -4790
rect 853 -5038 869 -4790
rect 803 -5050 869 -5038
rect 899 -4790 965 -4778
rect 899 -5038 915 -4790
rect 949 -5038 965 -4790
rect 899 -5050 965 -5038
rect 995 -4790 1061 -4778
rect 995 -5038 1011 -4790
rect 1045 -5038 1061 -4790
rect 995 -5050 1061 -5038
rect 1091 -4790 1157 -4778
rect 1091 -5038 1107 -4790
rect 1141 -5038 1157 -4790
rect 1091 -5050 1157 -5038
rect 1187 -4790 1253 -4778
rect 1187 -5038 1203 -4790
rect 1237 -5038 1253 -4790
rect 1187 -5050 1253 -5038
rect 1283 -4790 1349 -4778
rect 1283 -5038 1299 -4790
rect 1333 -5038 1349 -4790
rect 1283 -5050 1349 -5038
rect 1379 -4790 1441 -4778
rect 1379 -5038 1395 -4790
rect 1429 -5038 1441 -4790
rect 1379 -5050 1441 -5038
rect 1944 -4790 2006 -4778
rect 1944 -5038 1956 -4790
rect 1990 -5038 2006 -4790
rect 1944 -5050 2006 -5038
rect 2036 -4790 2102 -4778
rect 2036 -5038 2052 -4790
rect 2086 -5038 2102 -4790
rect 2036 -5050 2102 -5038
rect 2132 -4790 2198 -4778
rect 2132 -5038 2148 -4790
rect 2182 -5038 2198 -4790
rect 2132 -5050 2198 -5038
rect 2228 -4790 2294 -4778
rect 2228 -5038 2244 -4790
rect 2278 -5038 2294 -4790
rect 2228 -5050 2294 -5038
rect 2324 -4790 2390 -4778
rect 2324 -5038 2340 -4790
rect 2374 -5038 2390 -4790
rect 2324 -5050 2390 -5038
rect 2420 -4790 2486 -4778
rect 2420 -5038 2436 -4790
rect 2470 -5038 2486 -4790
rect 2420 -5050 2486 -5038
rect 2516 -4790 2582 -4778
rect 2516 -5038 2532 -4790
rect 2566 -5038 2582 -4790
rect 2516 -5050 2582 -5038
rect 2612 -4790 2678 -4778
rect 2612 -5038 2628 -4790
rect 2662 -5038 2678 -4790
rect 2612 -5050 2678 -5038
rect 2708 -4790 2774 -4778
rect 2708 -5038 2724 -4790
rect 2758 -5038 2774 -4790
rect 2708 -5050 2774 -5038
rect 2804 -4790 2870 -4778
rect 2804 -5038 2820 -4790
rect 2854 -5038 2870 -4790
rect 2804 -5050 2870 -5038
rect 2900 -4790 2962 -4778
rect 2900 -5038 2916 -4790
rect 2950 -5038 2962 -4790
rect 2900 -5050 2962 -5038
<< ndiffc >>
rect 435 -368 469 -288
rect 531 -368 565 -288
rect 627 -368 661 -288
rect 723 -368 757 -288
rect 819 -368 853 -288
rect 915 -368 949 -288
rect 1011 -368 1045 -288
rect 1107 -368 1141 -288
rect 1203 -368 1237 -288
rect 1299 -368 1333 -288
rect 1395 -368 1429 -288
rect 1616 -372 1650 -296
rect 1704 -372 1738 -296
rect 1956 -368 1990 -288
rect 2052 -368 2086 -288
rect 2148 -368 2182 -288
rect 2244 -368 2278 -288
rect 2340 -368 2374 -288
rect 2436 -368 2470 -288
rect 2532 -368 2566 -288
rect 2628 -368 2662 -288
rect 2724 -368 2758 -288
rect 2820 -368 2854 -288
rect 2916 -368 2950 -288
rect -904 -574 -870 -540
rect -904 -642 -870 -608
rect -820 -574 -786 -540
rect -820 -642 -786 -608
rect -536 -574 -502 -540
rect -536 -642 -502 -608
rect -452 -574 -418 -540
rect -452 -642 -418 -608
rect -3116 -958 -3082 -878
rect -3020 -958 -2986 -878
rect -2924 -958 -2890 -878
rect -2828 -958 -2794 -878
rect -2732 -958 -2698 -878
rect -2636 -958 -2602 -878
rect -2540 -958 -2506 -878
rect -2444 -958 -2410 -878
rect -2348 -958 -2314 -878
rect -2252 -958 -2218 -878
rect -2156 -958 -2122 -878
rect -536 -1434 -502 -1400
rect -536 -1502 -502 -1468
rect -452 -1434 -418 -1400
rect -452 -1502 -418 -1468
rect -573 -1658 -539 -1624
rect -573 -1726 -539 -1692
rect -405 -1658 -371 -1624
rect -405 -1726 -371 -1692
rect 435 -1702 469 -1622
rect 531 -1702 565 -1622
rect 627 -1702 661 -1622
rect 723 -1702 757 -1622
rect 819 -1702 853 -1622
rect 915 -1702 949 -1622
rect 1011 -1702 1045 -1622
rect 1107 -1702 1141 -1622
rect 1203 -1702 1237 -1622
rect 1299 -1702 1333 -1622
rect 1395 -1702 1429 -1622
rect 1616 -1706 1650 -1630
rect 1704 -1706 1738 -1630
rect 1956 -1702 1990 -1622
rect 2052 -1702 2086 -1622
rect 2148 -1702 2182 -1622
rect 2244 -1702 2278 -1622
rect 2340 -1702 2374 -1622
rect 2436 -1702 2470 -1622
rect 2532 -1702 2566 -1622
rect 2628 -1702 2662 -1622
rect 2724 -1702 2758 -1622
rect 2820 -1702 2854 -1622
rect 2916 -1702 2950 -1622
rect -3116 -2292 -3082 -2212
rect -3020 -2292 -2986 -2212
rect -2924 -2292 -2890 -2212
rect -2828 -2292 -2794 -2212
rect -2732 -2292 -2698 -2212
rect -2636 -2292 -2602 -2212
rect -2540 -2292 -2506 -2212
rect -2444 -2292 -2410 -2212
rect -2348 -2292 -2314 -2212
rect -2252 -2292 -2218 -2212
rect -2156 -2292 -2122 -2212
rect -1088 -2522 -1054 -2488
rect -1088 -2590 -1054 -2556
rect -1004 -2522 -970 -2488
rect -1004 -2590 -970 -2556
rect -573 -2526 -539 -2492
rect -573 -2594 -539 -2560
rect -405 -2526 -371 -2492
rect -405 -2594 -371 -2560
rect -1088 -2750 -1054 -2716
rect -1088 -2818 -1054 -2784
rect -1004 -2750 -970 -2716
rect -1004 -2818 -970 -2784
rect -573 -2746 -539 -2712
rect -573 -2814 -539 -2780
rect -405 -2746 -371 -2712
rect -405 -2814 -371 -2780
rect 435 -3080 469 -3000
rect 531 -3080 565 -3000
rect 627 -3080 661 -3000
rect 723 -3080 757 -3000
rect 819 -3080 853 -3000
rect 915 -3080 949 -3000
rect 1011 -3080 1045 -3000
rect 1107 -3080 1141 -3000
rect 1203 -3080 1237 -3000
rect 1299 -3080 1333 -3000
rect 1395 -3080 1429 -3000
rect 1616 -3084 1650 -3008
rect 1704 -3084 1738 -3008
rect 1956 -3080 1990 -3000
rect 2052 -3080 2086 -3000
rect 2148 -3080 2182 -3000
rect 2244 -3080 2278 -3000
rect 2340 -3080 2374 -3000
rect 2436 -3080 2470 -3000
rect 2532 -3080 2566 -3000
rect 2628 -3080 2662 -3000
rect 2724 -3080 2758 -3000
rect 2820 -3080 2854 -3000
rect 2916 -3080 2950 -3000
rect -3116 -3670 -3082 -3590
rect -3020 -3670 -2986 -3590
rect -2924 -3670 -2890 -3590
rect -2828 -3670 -2794 -3590
rect -2732 -3670 -2698 -3590
rect -2636 -3670 -2602 -3590
rect -2540 -3670 -2506 -3590
rect -2444 -3670 -2410 -3590
rect -2348 -3670 -2314 -3590
rect -2252 -3670 -2218 -3590
rect -2156 -3670 -2122 -3590
rect -573 -3614 -539 -3580
rect -573 -3682 -539 -3648
rect -405 -3614 -371 -3580
rect -405 -3682 -371 -3648
rect -536 -3838 -502 -3804
rect -536 -3906 -502 -3872
rect -452 -3838 -418 -3804
rect -452 -3906 -418 -3872
rect 435 -4458 469 -4378
rect 531 -4458 565 -4378
rect 627 -4458 661 -4378
rect 723 -4458 757 -4378
rect 819 -4458 853 -4378
rect 915 -4458 949 -4378
rect 1011 -4458 1045 -4378
rect 1107 -4458 1141 -4378
rect 1203 -4458 1237 -4378
rect 1299 -4458 1333 -4378
rect 1395 -4458 1429 -4378
rect 1616 -4462 1650 -4386
rect 1704 -4462 1738 -4386
rect 1956 -4458 1990 -4378
rect 2052 -4458 2086 -4378
rect 2148 -4458 2182 -4378
rect 2244 -4458 2278 -4378
rect 2340 -4458 2374 -4378
rect 2436 -4458 2470 -4378
rect 2532 -4458 2566 -4378
rect 2628 -4458 2662 -4378
rect 2724 -4458 2758 -4378
rect 2820 -4458 2854 -4378
rect 2916 -4458 2950 -4378
rect -536 -4698 -502 -4664
rect -536 -4766 -502 -4732
rect -452 -4698 -418 -4664
rect -452 -4766 -418 -4732
rect -3116 -5048 -3082 -4968
rect -3020 -5048 -2986 -4968
rect -2924 -5048 -2890 -4968
rect -2828 -5048 -2794 -4968
rect -2732 -5048 -2698 -4968
rect -2636 -5048 -2602 -4968
rect -2540 -5048 -2506 -4968
rect -2444 -5048 -2410 -4968
rect -2348 -5048 -2314 -4968
rect -2252 -5048 -2218 -4968
rect -2156 -5048 -2122 -4968
<< pdiffc >>
rect -3116 -546 -3082 -298
rect -3020 -546 -2986 -298
rect -2924 -546 -2890 -298
rect -2828 -546 -2794 -298
rect -2732 -546 -2698 -298
rect -2636 -546 -2602 -298
rect -2540 -546 -2506 -298
rect -2444 -546 -2410 -298
rect -2348 -546 -2314 -298
rect -2252 -546 -2218 -298
rect -2156 -546 -2122 -298
rect -904 -826 -870 -792
rect -904 -894 -870 -860
rect -904 -962 -870 -928
rect -820 -826 -786 -792
rect -820 -894 -786 -860
rect -820 -962 -786 -928
rect -536 -826 -502 -792
rect -536 -894 -502 -860
rect -536 -962 -502 -928
rect -452 -826 -418 -792
rect -452 -894 -418 -860
rect -452 -962 -418 -928
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect -536 -1114 -502 -1080
rect -536 -1182 -502 -1148
rect -536 -1250 -502 -1216
rect -452 -1114 -418 -1080
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect -452 -1182 -418 -1148
rect -452 -1250 -418 -1216
rect -3116 -1880 -3082 -1632
rect -3020 -1880 -2986 -1632
rect -2924 -1880 -2890 -1632
rect -2828 -1880 -2794 -1632
rect -2732 -1880 -2698 -1632
rect -2636 -1880 -2602 -1632
rect -2540 -1880 -2506 -1632
rect -2444 -1880 -2410 -1632
rect -2348 -1880 -2314 -1632
rect -2252 -1880 -2218 -1632
rect -2156 -1880 -2122 -1632
rect -573 -1914 -539 -1880
rect -573 -1982 -539 -1948
rect -573 -2050 -539 -2016
rect -489 -1914 -455 -1880
rect -489 -1982 -455 -1948
rect -489 -2050 -455 -2016
rect -405 -1914 -371 -1880
rect -405 -1982 -371 -1948
rect -405 -2050 -371 -2016
rect -1088 -2202 -1054 -2168
rect -1088 -2270 -1054 -2236
rect -1088 -2338 -1054 -2304
rect -1004 -2202 -970 -2168
rect -1004 -2270 -970 -2236
rect -1004 -2338 -970 -2304
rect -573 -2202 -539 -2168
rect -573 -2270 -539 -2236
rect -573 -2338 -539 -2304
rect -489 -2202 -455 -2168
rect -489 -2270 -455 -2236
rect -489 -2338 -455 -2304
rect -405 -2202 -371 -2168
rect -405 -2270 -371 -2236
rect -405 -2338 -371 -2304
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
rect -3116 -3258 -3082 -3010
rect -3020 -3258 -2986 -3010
rect -2924 -3258 -2890 -3010
rect -2828 -3258 -2794 -3010
rect -2732 -3258 -2698 -3010
rect -2636 -3258 -2602 -3010
rect -2540 -3258 -2506 -3010
rect -2444 -3258 -2410 -3010
rect -2348 -3258 -2314 -3010
rect -2252 -3258 -2218 -3010
rect -2156 -3258 -2122 -3010
rect -1088 -3002 -1054 -2968
rect -1088 -3070 -1054 -3036
rect -1088 -3138 -1054 -3104
rect -1004 -3002 -970 -2968
rect -1004 -3070 -970 -3036
rect -1004 -3138 -970 -3104
rect -573 -3002 -539 -2968
rect -573 -3070 -539 -3036
rect -573 -3138 -539 -3104
rect -489 -3002 -455 -2968
rect -489 -3070 -455 -3036
rect -489 -3138 -455 -3104
rect -405 -3002 -371 -2968
rect -405 -3070 -371 -3036
rect -405 -3138 -371 -3104
rect -573 -3290 -539 -3256
rect -573 -3358 -539 -3324
rect -573 -3426 -539 -3392
rect -489 -3290 -455 -3256
rect -489 -3358 -455 -3324
rect -489 -3426 -455 -3392
rect -405 -3290 -371 -3256
rect -405 -3358 -371 -3324
rect -405 -3426 -371 -3392
rect 435 -3660 469 -3412
rect 531 -3660 565 -3412
rect 627 -3660 661 -3412
rect 723 -3660 757 -3412
rect 819 -3660 853 -3412
rect 915 -3660 949 -3412
rect 1011 -3660 1045 -3412
rect 1107 -3660 1141 -3412
rect 1203 -3660 1237 -3412
rect 1299 -3660 1333 -3412
rect 1395 -3660 1429 -3412
rect 1956 -3660 1990 -3412
rect 2052 -3660 2086 -3412
rect 2148 -3660 2182 -3412
rect 2244 -3660 2278 -3412
rect 2340 -3660 2374 -3412
rect 2436 -3660 2470 -3412
rect 2532 -3660 2566 -3412
rect 2628 -3660 2662 -3412
rect 2724 -3660 2758 -3412
rect 2820 -3660 2854 -3412
rect 2916 -3660 2950 -3412
rect -536 -4090 -502 -4056
rect -536 -4158 -502 -4124
rect -536 -4226 -502 -4192
rect -452 -4090 -418 -4056
rect -452 -4158 -418 -4124
rect -452 -4226 -418 -4192
rect -3116 -4636 -3082 -4388
rect -3020 -4636 -2986 -4388
rect -2924 -4636 -2890 -4388
rect -2828 -4636 -2794 -4388
rect -2732 -4636 -2698 -4388
rect -2636 -4636 -2602 -4388
rect -2540 -4636 -2506 -4388
rect -2444 -4636 -2410 -4388
rect -2348 -4636 -2314 -4388
rect -2252 -4636 -2218 -4388
rect -2156 -4636 -2122 -4388
rect -536 -4378 -502 -4344
rect -536 -4446 -502 -4412
rect -536 -4514 -502 -4480
rect -452 -4378 -418 -4344
rect -452 -4446 -418 -4412
rect -452 -4514 -418 -4480
rect 435 -5038 469 -4790
rect 531 -5038 565 -4790
rect 627 -5038 661 -4790
rect 723 -5038 757 -4790
rect 819 -5038 853 -4790
rect 915 -5038 949 -4790
rect 1011 -5038 1045 -4790
rect 1107 -5038 1141 -4790
rect 1203 -5038 1237 -4790
rect 1299 -5038 1333 -4790
rect 1395 -5038 1429 -4790
rect 1956 -5038 1990 -4790
rect 2052 -5038 2086 -4790
rect 2148 -5038 2182 -4790
rect 2244 -5038 2278 -4790
rect 2340 -5038 2374 -4790
rect 2436 -5038 2470 -4790
rect 2532 -5038 2566 -4790
rect 2628 -5038 2662 -4790
rect 2724 -5038 2758 -4790
rect 2820 -5038 2854 -4790
rect 2916 -5038 2950 -4790
<< psubdiff >>
rect 321 -136 417 -102
rect 1447 -136 1543 -102
rect 321 -198 355 -136
rect 1509 -198 1543 -136
rect 321 -458 355 -396
rect 1842 -136 1938 -102
rect 2968 -136 3064 -102
rect 1842 -198 1876 -136
rect 1509 -458 1543 -396
rect 3030 -198 3064 -136
rect 321 -492 417 -458
rect 1447 -492 1543 -458
rect 1842 -458 1876 -396
rect 3030 -458 3064 -396
rect 1842 -492 1938 -458
rect 2968 -492 3064 -458
rect -675 -588 -641 -541
rect -675 -646 -641 -622
rect -3230 -788 -3134 -754
rect -2104 -788 -2008 -754
rect -3230 -850 -3196 -788
rect -2042 -850 -2008 -788
rect -3230 -1110 -3196 -1048
rect -2042 -1110 -2008 -1048
rect -3230 -1144 -3134 -1110
rect -2104 -1144 -2008 -1110
rect -675 -1420 -641 -1396
rect -675 -1501 -641 -1454
rect 321 -1470 417 -1436
rect 1447 -1470 1543 -1436
rect 321 -1532 355 -1470
rect -675 -1676 -641 -1629
rect -675 -1734 -641 -1710
rect 1509 -1532 1543 -1470
rect 321 -1792 355 -1730
rect 1842 -1470 1938 -1436
rect 2968 -1470 3064 -1436
rect 1842 -1532 1876 -1470
rect 1509 -1792 1543 -1730
rect 3030 -1532 3064 -1470
rect 321 -1826 417 -1792
rect 1447 -1826 1543 -1792
rect 1842 -1792 1876 -1730
rect 3030 -1792 3064 -1730
rect 1842 -1826 1938 -1792
rect 2968 -1826 3064 -1792
rect -3230 -2122 -3134 -2088
rect -2104 -2122 -2008 -2088
rect -3230 -2184 -3196 -2122
rect -2042 -2184 -2008 -2122
rect -3230 -2444 -3196 -2382
rect -2042 -2444 -2008 -2382
rect -3230 -2478 -3134 -2444
rect -2104 -2478 -2008 -2444
rect -1227 -2508 -1193 -2484
rect -1227 -2589 -1193 -2542
rect -675 -2508 -641 -2484
rect -675 -2589 -641 -2542
rect -1227 -2764 -1193 -2717
rect -1227 -2822 -1193 -2798
rect -675 -2764 -641 -2717
rect -675 -2822 -641 -2798
rect 321 -2848 417 -2814
rect 1447 -2848 1543 -2814
rect 321 -2910 355 -2848
rect 1509 -2910 1543 -2848
rect 321 -3170 355 -3108
rect 1842 -2848 1938 -2814
rect 2968 -2848 3064 -2814
rect 1842 -2910 1876 -2848
rect 1509 -3170 1543 -3108
rect 3030 -2910 3064 -2848
rect 321 -3204 417 -3170
rect 1447 -3204 1543 -3170
rect 1842 -3170 1876 -3108
rect 3030 -3170 3064 -3108
rect 1842 -3204 1938 -3170
rect 2968 -3204 3064 -3170
rect -3230 -3500 -3134 -3466
rect -2104 -3500 -2008 -3466
rect -3230 -3562 -3196 -3500
rect -2042 -3562 -2008 -3500
rect -3230 -3822 -3196 -3760
rect -675 -3596 -641 -3572
rect -675 -3677 -641 -3630
rect -2042 -3822 -2008 -3760
rect -3230 -3856 -3134 -3822
rect -2104 -3856 -2008 -3822
rect -675 -3852 -641 -3805
rect -675 -3910 -641 -3886
rect 321 -4226 417 -4192
rect 1447 -4226 1543 -4192
rect 321 -4288 355 -4226
rect 1509 -4288 1543 -4226
rect 321 -4548 355 -4486
rect 1842 -4226 1938 -4192
rect 2968 -4226 3064 -4192
rect 1842 -4288 1876 -4226
rect 1509 -4548 1543 -4486
rect 3030 -4288 3064 -4226
rect 321 -4582 417 -4548
rect 1447 -4582 1543 -4548
rect 1842 -4548 1876 -4486
rect 3030 -4548 3064 -4486
rect 1842 -4582 1938 -4548
rect 2968 -4582 3064 -4548
rect -675 -4684 -641 -4660
rect -675 -4765 -641 -4718
rect -3230 -4878 -3134 -4844
rect -2104 -4878 -2008 -4844
rect -3230 -4940 -3196 -4878
rect -2042 -4940 -2008 -4878
rect -3230 -5200 -3196 -5138
rect -2042 -5200 -2008 -5138
rect -3230 -5234 -3134 -5200
rect -2104 -5234 -2008 -5200
<< nsubdiff >>
rect -3230 -136 -3134 -102
rect -2104 -136 -2008 -102
rect -3230 -198 -3196 -136
rect -2042 -198 -2008 -136
rect -3230 -646 -3196 -584
rect -2042 -646 -2008 -584
rect -3230 -680 -3134 -646
rect -2104 -680 -2008 -646
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect 1509 -662 1543 -600
rect -675 -806 -641 -782
rect -675 -899 -641 -840
rect -675 -957 -641 -933
rect -675 -1109 -641 -1085
rect -675 -1202 -641 -1143
rect -675 -1260 -641 -1236
rect 321 -1110 355 -1048
rect 1509 -1110 1543 -1048
rect 321 -1144 417 -1110
rect 1447 -1144 1543 -1110
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1842 -1110 1876 -1048
rect 3030 -1110 3064 -1048
rect 1842 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect -3230 -1470 -3134 -1436
rect -2104 -1470 -2008 -1436
rect -3230 -1532 -3196 -1470
rect -2042 -1532 -2008 -1470
rect -3230 -1980 -3196 -1918
rect -2042 -1980 -2008 -1918
rect -3230 -2014 -3134 -1980
rect -2104 -2014 -2008 -1980
rect -675 -1894 -641 -1870
rect -675 -1987 -641 -1928
rect -675 -2045 -641 -2021
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect 1509 -1996 1543 -1934
rect -1227 -2197 -1193 -2173
rect -1227 -2290 -1193 -2231
rect -1227 -2348 -1193 -2324
rect -675 -2197 -641 -2173
rect -675 -2290 -641 -2231
rect -675 -2348 -641 -2324
rect 321 -2444 355 -2382
rect 1509 -2444 1543 -2382
rect 321 -2478 417 -2444
rect 1447 -2478 1543 -2444
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1842 -2444 1876 -2382
rect 3030 -2444 3064 -2382
rect 1842 -2478 1938 -2444
rect 2968 -2478 3064 -2444
rect -3230 -2848 -3134 -2814
rect -2104 -2848 -2008 -2814
rect -3230 -2910 -3196 -2848
rect -2042 -2910 -2008 -2848
rect -1227 -2982 -1193 -2958
rect -1227 -3075 -1193 -3016
rect -1227 -3133 -1193 -3109
rect -675 -2982 -641 -2958
rect -675 -3075 -641 -3016
rect -675 -3133 -641 -3109
rect -3230 -3358 -3196 -3296
rect -2042 -3358 -2008 -3296
rect -3230 -3392 -3134 -3358
rect -2104 -3392 -2008 -3358
rect -675 -3285 -641 -3261
rect -675 -3378 -641 -3319
rect -675 -3436 -641 -3412
rect 321 -3312 417 -3278
rect 1447 -3312 1543 -3278
rect 321 -3374 355 -3312
rect 1509 -3374 1543 -3312
rect 321 -3822 355 -3760
rect 1509 -3822 1543 -3760
rect 321 -3856 417 -3822
rect 1447 -3856 1543 -3822
rect 1842 -3312 1938 -3278
rect 2968 -3312 3064 -3278
rect 1842 -3374 1876 -3312
rect 3030 -3374 3064 -3312
rect 1842 -3822 1876 -3760
rect 3030 -3822 3064 -3760
rect 1842 -3856 1938 -3822
rect 2968 -3856 3064 -3822
rect -675 -4070 -641 -4046
rect -675 -4163 -641 -4104
rect -3230 -4226 -3134 -4192
rect -2104 -4226 -2008 -4192
rect -675 -4221 -641 -4197
rect -3230 -4288 -3196 -4226
rect -2042 -4288 -2008 -4226
rect -675 -4373 -641 -4349
rect -675 -4466 -641 -4407
rect -675 -4524 -641 -4500
rect -3230 -4736 -3196 -4674
rect -2042 -4736 -2008 -4674
rect -3230 -4770 -3134 -4736
rect -2104 -4770 -2008 -4736
rect 321 -4690 417 -4656
rect 1447 -4690 1543 -4656
rect 321 -4752 355 -4690
rect 1509 -4752 1543 -4690
rect 321 -5200 355 -5138
rect 1509 -5200 1543 -5138
rect 321 -5234 417 -5200
rect 1447 -5234 1543 -5200
rect 1842 -4690 1938 -4656
rect 2968 -4690 3064 -4656
rect 1842 -4752 1876 -4690
rect 3030 -4752 3064 -4690
rect 1842 -5200 1876 -5138
rect 3030 -5200 3064 -5138
rect 1842 -5234 1938 -5200
rect 2968 -5234 3064 -5200
<< psubdiffcont >>
rect 417 -136 1447 -102
rect 321 -396 355 -198
rect 1509 -396 1543 -198
rect 1938 -136 2968 -102
rect 1842 -396 1876 -198
rect 417 -492 1447 -458
rect 3030 -396 3064 -198
rect 1938 -492 2968 -458
rect -675 -622 -641 -588
rect -3134 -788 -2104 -754
rect -3230 -1048 -3196 -850
rect -2042 -1048 -2008 -850
rect -3134 -1144 -2104 -1110
rect -675 -1454 -641 -1420
rect 417 -1470 1447 -1436
rect -675 -1710 -641 -1676
rect 321 -1730 355 -1532
rect 1509 -1730 1543 -1532
rect 1938 -1470 2968 -1436
rect 1842 -1730 1876 -1532
rect 417 -1826 1447 -1792
rect 3030 -1730 3064 -1532
rect 1938 -1826 2968 -1792
rect -3134 -2122 -2104 -2088
rect -3230 -2382 -3196 -2184
rect -2042 -2382 -2008 -2184
rect -3134 -2478 -2104 -2444
rect -1227 -2542 -1193 -2508
rect -675 -2542 -641 -2508
rect -1227 -2798 -1193 -2764
rect -675 -2798 -641 -2764
rect 417 -2848 1447 -2814
rect 321 -3108 355 -2910
rect 1509 -3108 1543 -2910
rect 1938 -2848 2968 -2814
rect 1842 -3108 1876 -2910
rect 417 -3204 1447 -3170
rect 3030 -3108 3064 -2910
rect 1938 -3204 2968 -3170
rect -3134 -3500 -2104 -3466
rect -3230 -3760 -3196 -3562
rect -2042 -3760 -2008 -3562
rect -675 -3630 -641 -3596
rect -3134 -3856 -2104 -3822
rect -675 -3886 -641 -3852
rect 417 -4226 1447 -4192
rect 321 -4486 355 -4288
rect 1509 -4486 1543 -4288
rect 1938 -4226 2968 -4192
rect 1842 -4486 1876 -4288
rect 417 -4582 1447 -4548
rect 3030 -4486 3064 -4288
rect 1938 -4582 2968 -4548
rect -675 -4718 -641 -4684
rect -3134 -4878 -2104 -4844
rect -3230 -5138 -3196 -4940
rect -2042 -5138 -2008 -4940
rect -3134 -5234 -2104 -5200
<< nsubdiffcont >>
rect -3134 -136 -2104 -102
rect -3230 -584 -3196 -198
rect -2042 -584 -2008 -198
rect -3134 -680 -2104 -646
rect 417 -600 1447 -566
rect -675 -840 -641 -806
rect -675 -933 -641 -899
rect 321 -1048 355 -662
rect -675 -1143 -641 -1109
rect -675 -1236 -641 -1202
rect 1509 -1048 1543 -662
rect 417 -1144 1447 -1110
rect 1938 -600 2968 -566
rect 1842 -1048 1876 -662
rect 3030 -1048 3064 -662
rect 1938 -1144 2968 -1110
rect -3134 -1470 -2104 -1436
rect -3230 -1918 -3196 -1532
rect -2042 -1918 -2008 -1532
rect -3134 -2014 -2104 -1980
rect -675 -1928 -641 -1894
rect -675 -2021 -641 -1987
rect 417 -1934 1447 -1900
rect -1227 -2231 -1193 -2197
rect -1227 -2324 -1193 -2290
rect -675 -2231 -641 -2197
rect -675 -2324 -641 -2290
rect 321 -2382 355 -1996
rect 1509 -2382 1543 -1996
rect 417 -2478 1447 -2444
rect 1938 -1934 2968 -1900
rect 1842 -2382 1876 -1996
rect 3030 -2382 3064 -1996
rect 1938 -2478 2968 -2444
rect -3134 -2848 -2104 -2814
rect -3230 -3296 -3196 -2910
rect -2042 -3296 -2008 -2910
rect -1227 -3016 -1193 -2982
rect -1227 -3109 -1193 -3075
rect -675 -3016 -641 -2982
rect -675 -3109 -641 -3075
rect -3134 -3392 -2104 -3358
rect -675 -3319 -641 -3285
rect -675 -3412 -641 -3378
rect 417 -3312 1447 -3278
rect 321 -3760 355 -3374
rect 1509 -3760 1543 -3374
rect 417 -3856 1447 -3822
rect 1938 -3312 2968 -3278
rect 1842 -3760 1876 -3374
rect 3030 -3760 3064 -3374
rect 1938 -3856 2968 -3822
rect -675 -4104 -641 -4070
rect -3134 -4226 -2104 -4192
rect -675 -4197 -641 -4163
rect -3230 -4674 -3196 -4288
rect -2042 -4674 -2008 -4288
rect -675 -4407 -641 -4373
rect -675 -4500 -641 -4466
rect -3134 -4770 -2104 -4736
rect 417 -4690 1447 -4656
rect 321 -5138 355 -4752
rect 1509 -5138 1543 -4752
rect 417 -5234 1447 -5200
rect 1938 -4690 2968 -4656
rect 1842 -5138 1876 -4752
rect 3030 -5138 3064 -4752
rect 1938 -5234 2968 -5200
<< poly >>
rect -3132 -204 -2106 -188
rect -3132 -238 -3116 -204
rect -3082 -238 -2924 -204
rect -2890 -238 -2732 -204
rect -2698 -238 -2540 -204
rect -2506 -238 -2348 -204
rect -2314 -238 -2156 -204
rect -2122 -238 -2106 -204
rect -3132 -254 -2106 -238
rect -3066 -286 -3036 -254
rect -2970 -286 -2940 -254
rect -2874 -286 -2844 -254
rect -2778 -286 -2748 -254
rect -2682 -286 -2652 -254
rect -2586 -286 -2556 -254
rect -2490 -286 -2460 -254
rect -2394 -286 -2364 -254
rect -2298 -286 -2268 -254
rect -2202 -286 -2172 -254
rect -3066 -584 -3036 -558
rect -2970 -584 -2940 -558
rect -2874 -584 -2844 -558
rect -2778 -584 -2748 -558
rect -2682 -584 -2652 -558
rect -2586 -584 -2556 -558
rect -2490 -584 -2460 -558
rect -2394 -584 -2364 -558
rect -2298 -584 -2268 -558
rect -2202 -584 -2172 -558
rect 419 -200 1445 -188
rect 419 -234 435 -200
rect 469 -234 627 -200
rect 661 -234 819 -200
rect 853 -234 1011 -200
rect 1045 -234 1203 -200
rect 1237 -234 1395 -200
rect 1429 -234 1445 -200
rect 419 -254 1445 -234
rect 485 -276 515 -254
rect 581 -276 611 -254
rect 677 -276 707 -254
rect 773 -276 803 -254
rect 869 -276 899 -254
rect 965 -276 995 -254
rect 1061 -276 1091 -254
rect 1157 -276 1187 -254
rect 1253 -276 1283 -254
rect 1349 -276 1379 -254
rect 485 -406 515 -380
rect 581 -406 611 -380
rect 677 -406 707 -380
rect 773 -406 803 -380
rect 869 -406 899 -380
rect 965 -406 995 -380
rect 1061 -406 1091 -380
rect 1157 -406 1187 -380
rect 1253 -406 1283 -380
rect 1349 -406 1379 -380
rect 1662 -284 1692 -258
rect 1662 -406 1692 -384
rect 1940 -200 2966 -188
rect 1940 -234 1956 -200
rect 1990 -234 2148 -200
rect 2182 -234 2340 -200
rect 2374 -234 2532 -200
rect 2566 -234 2724 -200
rect 2758 -234 2916 -200
rect 2950 -234 2966 -200
rect 1940 -254 2966 -234
rect 2006 -276 2036 -254
rect 2102 -276 2132 -254
rect 2198 -276 2228 -254
rect 2294 -276 2324 -254
rect 2390 -276 2420 -254
rect 2486 -276 2516 -254
rect 2582 -276 2612 -254
rect 2678 -276 2708 -254
rect 2774 -276 2804 -254
rect 2870 -276 2900 -254
rect 1644 -422 1710 -406
rect 1644 -456 1660 -422
rect 1694 -456 1710 -422
rect 1644 -472 1710 -456
rect 2006 -406 2036 -380
rect 2102 -406 2132 -380
rect 2198 -406 2228 -380
rect 2294 -406 2324 -380
rect 2390 -406 2420 -380
rect 2486 -406 2516 -380
rect 2582 -406 2612 -380
rect 2678 -406 2708 -380
rect 2774 -406 2804 -380
rect 2870 -406 2900 -380
rect -860 -524 -830 -498
rect -492 -524 -462 -498
rect -860 -676 -830 -654
rect -492 -676 -462 -654
rect -916 -692 -830 -676
rect -916 -726 -900 -692
rect -866 -726 -830 -692
rect -916 -742 -830 -726
rect -548 -692 -462 -676
rect -548 -726 -532 -692
rect -498 -726 -462 -692
rect -548 -742 -462 -726
rect -860 -774 -830 -742
rect -492 -774 -462 -742
rect -3066 -866 -3036 -840
rect -2970 -866 -2940 -840
rect -2874 -866 -2844 -840
rect -2778 -866 -2748 -840
rect -2682 -866 -2652 -840
rect -2586 -866 -2556 -840
rect -2490 -866 -2460 -840
rect -2394 -866 -2364 -840
rect -2298 -866 -2268 -840
rect -2202 -866 -2172 -840
rect -3066 -992 -3036 -970
rect -2970 -992 -2940 -970
rect -2874 -992 -2844 -970
rect -2778 -992 -2748 -970
rect -2682 -992 -2652 -970
rect -2586 -992 -2556 -970
rect -2490 -992 -2460 -970
rect -2394 -992 -2364 -970
rect -2298 -992 -2268 -970
rect -2202 -992 -2172 -970
rect -3132 -1012 -2106 -992
rect -3132 -1046 -3116 -1012
rect -3082 -1046 -2924 -1012
rect -2890 -1046 -2732 -1012
rect -2698 -1046 -2540 -1012
rect -2506 -1046 -2348 -1012
rect -2314 -1046 -2156 -1012
rect -2122 -1046 -2106 -1012
rect -3132 -1058 -2106 -1046
rect -860 -1000 -830 -974
rect -492 -1000 -462 -974
rect -492 -1068 -462 -1042
rect 485 -688 515 -662
rect 581 -688 611 -662
rect 677 -688 707 -662
rect 773 -688 803 -662
rect 869 -688 899 -662
rect 965 -688 995 -662
rect 1061 -688 1091 -662
rect 1157 -688 1187 -662
rect 1253 -688 1283 -662
rect 1349 -688 1379 -662
rect 485 -992 515 -960
rect 581 -992 611 -960
rect 677 -992 707 -960
rect 773 -992 803 -960
rect 869 -992 899 -960
rect 965 -992 995 -960
rect 1061 -992 1091 -960
rect 1157 -992 1187 -960
rect 1253 -992 1283 -960
rect 1349 -992 1379 -960
rect 419 -1008 1445 -992
rect 419 -1042 435 -1008
rect 469 -1042 627 -1008
rect 661 -1042 819 -1008
rect 853 -1042 1011 -1008
rect 1045 -1042 1203 -1008
rect 1237 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect 419 -1058 1445 -1042
rect 2006 -688 2036 -662
rect 2102 -688 2132 -662
rect 2198 -688 2228 -662
rect 2294 -688 2324 -662
rect 2390 -688 2420 -662
rect 2486 -688 2516 -662
rect 2582 -688 2612 -662
rect 2678 -688 2708 -662
rect 2774 -688 2804 -662
rect 2870 -688 2900 -662
rect 2006 -992 2036 -960
rect 2102 -992 2132 -960
rect 2198 -992 2228 -960
rect 2294 -992 2324 -960
rect 2390 -992 2420 -960
rect 2486 -992 2516 -960
rect 2582 -992 2612 -960
rect 2678 -992 2708 -960
rect 2774 -992 2804 -960
rect 2870 -992 2900 -960
rect 1940 -1008 2966 -992
rect 1940 -1042 1956 -1008
rect 1990 -1042 2148 -1008
rect 2182 -1042 2340 -1008
rect 2374 -1042 2532 -1008
rect 2566 -1042 2724 -1008
rect 2758 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1940 -1058 2966 -1042
rect -492 -1300 -462 -1268
rect -548 -1316 -462 -1300
rect -548 -1350 -532 -1316
rect -498 -1350 -462 -1316
rect -548 -1366 -462 -1350
rect -492 -1388 -462 -1366
rect -3132 -1538 -2106 -1522
rect -3132 -1572 -3116 -1538
rect -3082 -1572 -2924 -1538
rect -2890 -1572 -2732 -1538
rect -2698 -1572 -2540 -1538
rect -2506 -1572 -2348 -1538
rect -2314 -1572 -2156 -1538
rect -2122 -1572 -2106 -1538
rect -3132 -1588 -2106 -1572
rect -3066 -1620 -3036 -1588
rect -2970 -1620 -2940 -1588
rect -2874 -1620 -2844 -1588
rect -2778 -1620 -2748 -1588
rect -2682 -1620 -2652 -1588
rect -2586 -1620 -2556 -1588
rect -2490 -1620 -2460 -1588
rect -2394 -1620 -2364 -1588
rect -2298 -1620 -2268 -1588
rect -2202 -1620 -2172 -1588
rect -3066 -1918 -3036 -1892
rect -2970 -1918 -2940 -1892
rect -2874 -1918 -2844 -1892
rect -2778 -1918 -2748 -1892
rect -2682 -1918 -2652 -1892
rect -2586 -1918 -2556 -1892
rect -2490 -1918 -2460 -1892
rect -2394 -1918 -2364 -1892
rect -2298 -1918 -2268 -1892
rect -2202 -1918 -2172 -1892
rect -492 -1544 -462 -1518
rect -529 -1612 -499 -1586
rect -445 -1612 -415 -1586
rect 419 -1534 1445 -1522
rect 419 -1568 435 -1534
rect 469 -1568 627 -1534
rect 661 -1568 819 -1534
rect 853 -1568 1011 -1534
rect 1045 -1568 1203 -1534
rect 1237 -1568 1395 -1534
rect 1429 -1568 1445 -1534
rect 419 -1588 1445 -1568
rect 485 -1610 515 -1588
rect 581 -1610 611 -1588
rect 677 -1610 707 -1588
rect 773 -1610 803 -1588
rect 869 -1610 899 -1588
rect 965 -1610 995 -1588
rect 1061 -1610 1091 -1588
rect 1157 -1610 1187 -1588
rect 1253 -1610 1283 -1588
rect 1349 -1610 1379 -1588
rect -529 -1764 -499 -1742
rect -591 -1780 -499 -1764
rect -591 -1814 -576 -1780
rect -542 -1814 -499 -1780
rect -591 -1830 -499 -1814
rect -529 -1862 -499 -1830
rect -445 -1764 -415 -1742
rect -445 -1780 -357 -1764
rect -445 -1814 -408 -1780
rect -374 -1814 -357 -1780
rect -445 -1830 -357 -1814
rect 485 -1740 515 -1714
rect 581 -1740 611 -1714
rect 677 -1740 707 -1714
rect 773 -1740 803 -1714
rect 869 -1740 899 -1714
rect 965 -1740 995 -1714
rect 1061 -1740 1091 -1714
rect 1157 -1740 1187 -1714
rect 1253 -1740 1283 -1714
rect 1349 -1740 1379 -1714
rect 1662 -1618 1692 -1592
rect 1662 -1740 1692 -1718
rect 1940 -1534 2966 -1522
rect 1940 -1568 1956 -1534
rect 1990 -1568 2148 -1534
rect 2182 -1568 2340 -1534
rect 2374 -1568 2532 -1534
rect 2566 -1568 2724 -1534
rect 2758 -1568 2916 -1534
rect 2950 -1568 2966 -1534
rect 1940 -1588 2966 -1568
rect 2006 -1610 2036 -1588
rect 2102 -1610 2132 -1588
rect 2198 -1610 2228 -1588
rect 2294 -1610 2324 -1588
rect 2390 -1610 2420 -1588
rect 2486 -1610 2516 -1588
rect 2582 -1610 2612 -1588
rect 2678 -1610 2708 -1588
rect 2774 -1610 2804 -1588
rect 2870 -1610 2900 -1588
rect 1644 -1756 1710 -1740
rect 1644 -1790 1660 -1756
rect 1694 -1790 1710 -1756
rect 1644 -1806 1710 -1790
rect 2006 -1740 2036 -1714
rect 2102 -1740 2132 -1714
rect 2198 -1740 2228 -1714
rect 2294 -1740 2324 -1714
rect 2390 -1740 2420 -1714
rect 2486 -1740 2516 -1714
rect 2582 -1740 2612 -1714
rect 2678 -1740 2708 -1714
rect 2774 -1740 2804 -1714
rect 2870 -1740 2900 -1714
rect -445 -1862 -415 -1830
rect -529 -2088 -499 -2062
rect -445 -2088 -415 -2062
rect -3066 -2200 -3036 -2174
rect -2970 -2200 -2940 -2174
rect -2874 -2200 -2844 -2174
rect -2778 -2200 -2748 -2174
rect -2682 -2200 -2652 -2174
rect -2586 -2200 -2556 -2174
rect -2490 -2200 -2460 -2174
rect -2394 -2200 -2364 -2174
rect -2298 -2200 -2268 -2174
rect -2202 -2200 -2172 -2174
rect -1044 -2156 -1014 -2130
rect -529 -2156 -499 -2130
rect -445 -2156 -415 -2130
rect -3066 -2326 -3036 -2304
rect -2970 -2326 -2940 -2304
rect -2874 -2326 -2844 -2304
rect -2778 -2326 -2748 -2304
rect -2682 -2326 -2652 -2304
rect -2586 -2326 -2556 -2304
rect -2490 -2326 -2460 -2304
rect -2394 -2326 -2364 -2304
rect -2298 -2326 -2268 -2304
rect -2202 -2326 -2172 -2304
rect -3132 -2346 -2106 -2326
rect -3132 -2380 -3116 -2346
rect -3082 -2380 -2924 -2346
rect -2890 -2380 -2732 -2346
rect -2698 -2380 -2540 -2346
rect -2506 -2380 -2348 -2346
rect -2314 -2380 -2156 -2346
rect -2122 -2380 -2106 -2346
rect -3132 -2392 -2106 -2380
rect -1044 -2388 -1014 -2356
rect -529 -2388 -499 -2356
rect -1100 -2404 -1014 -2388
rect -1100 -2438 -1084 -2404
rect -1050 -2438 -1014 -2404
rect -1100 -2454 -1014 -2438
rect -591 -2404 -499 -2388
rect -591 -2438 -576 -2404
rect -542 -2438 -499 -2404
rect -591 -2454 -499 -2438
rect -1044 -2476 -1014 -2454
rect -529 -2476 -499 -2454
rect -445 -2388 -415 -2356
rect 485 -2022 515 -1996
rect 581 -2022 611 -1996
rect 677 -2022 707 -1996
rect 773 -2022 803 -1996
rect 869 -2022 899 -1996
rect 965 -2022 995 -1996
rect 1061 -2022 1091 -1996
rect 1157 -2022 1187 -1996
rect 1253 -2022 1283 -1996
rect 1349 -2022 1379 -1996
rect 485 -2326 515 -2294
rect 581 -2326 611 -2294
rect 677 -2326 707 -2294
rect 773 -2326 803 -2294
rect 869 -2326 899 -2294
rect 965 -2326 995 -2294
rect 1061 -2326 1091 -2294
rect 1157 -2326 1187 -2294
rect 1253 -2326 1283 -2294
rect 1349 -2326 1379 -2294
rect -445 -2404 -357 -2388
rect -445 -2438 -408 -2404
rect -374 -2438 -357 -2404
rect -445 -2454 -357 -2438
rect 419 -2342 1445 -2326
rect 419 -2376 435 -2342
rect 469 -2376 627 -2342
rect 661 -2376 819 -2342
rect 853 -2376 1011 -2342
rect 1045 -2376 1203 -2342
rect 1237 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect 419 -2392 1445 -2376
rect -445 -2476 -415 -2454
rect 2006 -2022 2036 -1996
rect 2102 -2022 2132 -1996
rect 2198 -2022 2228 -1996
rect 2294 -2022 2324 -1996
rect 2390 -2022 2420 -1996
rect 2486 -2022 2516 -1996
rect 2582 -2022 2612 -1996
rect 2678 -2022 2708 -1996
rect 2774 -2022 2804 -1996
rect 2870 -2022 2900 -1996
rect 2006 -2326 2036 -2294
rect 2102 -2326 2132 -2294
rect 2198 -2326 2228 -2294
rect 2294 -2326 2324 -2294
rect 2390 -2326 2420 -2294
rect 2486 -2326 2516 -2294
rect 2582 -2326 2612 -2294
rect 2678 -2326 2708 -2294
rect 2774 -2326 2804 -2294
rect 2870 -2326 2900 -2294
rect 1940 -2342 2966 -2326
rect 1940 -2376 1956 -2342
rect 1990 -2376 2148 -2342
rect 2182 -2376 2340 -2342
rect 2374 -2376 2532 -2342
rect 2566 -2376 2724 -2342
rect 2758 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1940 -2392 2966 -2376
rect -1044 -2632 -1014 -2606
rect -529 -2632 -499 -2606
rect -445 -2632 -415 -2606
rect -1044 -2700 -1014 -2674
rect -529 -2700 -499 -2674
rect -445 -2700 -415 -2674
rect -3132 -2916 -2106 -2900
rect -3132 -2950 -3116 -2916
rect -3082 -2950 -2924 -2916
rect -2890 -2950 -2732 -2916
rect -2698 -2950 -2540 -2916
rect -2506 -2950 -2348 -2916
rect -2314 -2950 -2156 -2916
rect -2122 -2950 -2106 -2916
rect -3132 -2966 -2106 -2950
rect -1044 -2852 -1014 -2830
rect -529 -2852 -499 -2830
rect -3066 -2998 -3036 -2966
rect -2970 -2998 -2940 -2966
rect -2874 -2998 -2844 -2966
rect -2778 -2998 -2748 -2966
rect -2682 -2998 -2652 -2966
rect -2586 -2998 -2556 -2966
rect -2490 -2998 -2460 -2966
rect -2394 -2998 -2364 -2966
rect -2298 -2998 -2268 -2966
rect -2202 -2998 -2172 -2966
rect -3066 -3296 -3036 -3270
rect -2970 -3296 -2940 -3270
rect -2874 -3296 -2844 -3270
rect -2778 -3296 -2748 -3270
rect -2682 -3296 -2652 -3270
rect -2586 -3296 -2556 -3270
rect -2490 -3296 -2460 -3270
rect -2394 -3296 -2364 -3270
rect -2298 -3296 -2268 -3270
rect -2202 -3296 -2172 -3270
rect -1100 -2868 -1014 -2852
rect -1100 -2902 -1084 -2868
rect -1050 -2902 -1014 -2868
rect -1100 -2918 -1014 -2902
rect -591 -2868 -499 -2852
rect -591 -2902 -576 -2868
rect -542 -2902 -499 -2868
rect -591 -2918 -499 -2902
rect -1044 -2950 -1014 -2918
rect -529 -2950 -499 -2918
rect -445 -2852 -415 -2830
rect -445 -2868 -357 -2852
rect -445 -2902 -408 -2868
rect -374 -2902 -357 -2868
rect -445 -2918 -357 -2902
rect -445 -2950 -415 -2918
rect 419 -2912 1445 -2900
rect 419 -2946 435 -2912
rect 469 -2946 627 -2912
rect 661 -2946 819 -2912
rect 853 -2946 1011 -2912
rect 1045 -2946 1203 -2912
rect 1237 -2946 1395 -2912
rect 1429 -2946 1445 -2912
rect 419 -2966 1445 -2946
rect 485 -2988 515 -2966
rect 581 -2988 611 -2966
rect 677 -2988 707 -2966
rect 773 -2988 803 -2966
rect 869 -2988 899 -2966
rect 965 -2988 995 -2966
rect 1061 -2988 1091 -2966
rect 1157 -2988 1187 -2966
rect 1253 -2988 1283 -2966
rect 1349 -2988 1379 -2966
rect -1044 -3176 -1014 -3150
rect -529 -3176 -499 -3150
rect -445 -3176 -415 -3150
rect 485 -3118 515 -3092
rect 581 -3118 611 -3092
rect 677 -3118 707 -3092
rect 773 -3118 803 -3092
rect 869 -3118 899 -3092
rect 965 -3118 995 -3092
rect 1061 -3118 1091 -3092
rect 1157 -3118 1187 -3092
rect 1253 -3118 1283 -3092
rect 1349 -3118 1379 -3092
rect 1662 -2996 1692 -2970
rect 1662 -3118 1692 -3096
rect 1940 -2912 2966 -2900
rect 1940 -2946 1956 -2912
rect 1990 -2946 2148 -2912
rect 2182 -2946 2340 -2912
rect 2374 -2946 2532 -2912
rect 2566 -2946 2724 -2912
rect 2758 -2946 2916 -2912
rect 2950 -2946 2966 -2912
rect 1940 -2966 2966 -2946
rect 2006 -2988 2036 -2966
rect 2102 -2988 2132 -2966
rect 2198 -2988 2228 -2966
rect 2294 -2988 2324 -2966
rect 2390 -2988 2420 -2966
rect 2486 -2988 2516 -2966
rect 2582 -2988 2612 -2966
rect 2678 -2988 2708 -2966
rect 2774 -2988 2804 -2966
rect 2870 -2988 2900 -2966
rect 1644 -3134 1710 -3118
rect 1644 -3168 1660 -3134
rect 1694 -3168 1710 -3134
rect 1644 -3184 1710 -3168
rect 2006 -3118 2036 -3092
rect 2102 -3118 2132 -3092
rect 2198 -3118 2228 -3092
rect 2294 -3118 2324 -3092
rect 2390 -3118 2420 -3092
rect 2486 -3118 2516 -3092
rect 2582 -3118 2612 -3092
rect 2678 -3118 2708 -3092
rect 2774 -3118 2804 -3092
rect 2870 -3118 2900 -3092
rect -529 -3244 -499 -3218
rect -445 -3244 -415 -3218
rect -529 -3476 -499 -3444
rect -3066 -3578 -3036 -3552
rect -2970 -3578 -2940 -3552
rect -2874 -3578 -2844 -3552
rect -2778 -3578 -2748 -3552
rect -2682 -3578 -2652 -3552
rect -2586 -3578 -2556 -3552
rect -2490 -3578 -2460 -3552
rect -2394 -3578 -2364 -3552
rect -2298 -3578 -2268 -3552
rect -2202 -3578 -2172 -3552
rect -591 -3492 -499 -3476
rect -591 -3526 -576 -3492
rect -542 -3526 -499 -3492
rect -591 -3542 -499 -3526
rect -3066 -3704 -3036 -3682
rect -2970 -3704 -2940 -3682
rect -2874 -3704 -2844 -3682
rect -2778 -3704 -2748 -3682
rect -2682 -3704 -2652 -3682
rect -2586 -3704 -2556 -3682
rect -2490 -3704 -2460 -3682
rect -2394 -3704 -2364 -3682
rect -2298 -3704 -2268 -3682
rect -2202 -3704 -2172 -3682
rect -3132 -3724 -2106 -3704
rect -3132 -3758 -3116 -3724
rect -3082 -3758 -2924 -3724
rect -2890 -3758 -2732 -3724
rect -2698 -3758 -2540 -3724
rect -2506 -3758 -2348 -3724
rect -2314 -3758 -2156 -3724
rect -2122 -3758 -2106 -3724
rect -3132 -3770 -2106 -3758
rect -529 -3564 -499 -3542
rect -445 -3476 -415 -3444
rect -445 -3492 -357 -3476
rect -445 -3526 -408 -3492
rect -374 -3526 -357 -3492
rect -445 -3542 -357 -3526
rect -445 -3564 -415 -3542
rect -529 -3720 -499 -3694
rect -445 -3720 -415 -3694
rect 485 -3400 515 -3374
rect 581 -3400 611 -3374
rect 677 -3400 707 -3374
rect 773 -3400 803 -3374
rect 869 -3400 899 -3374
rect 965 -3400 995 -3374
rect 1061 -3400 1091 -3374
rect 1157 -3400 1187 -3374
rect 1253 -3400 1283 -3374
rect 1349 -3400 1379 -3374
rect 485 -3704 515 -3672
rect 581 -3704 611 -3672
rect 677 -3704 707 -3672
rect 773 -3704 803 -3672
rect 869 -3704 899 -3672
rect 965 -3704 995 -3672
rect 1061 -3704 1091 -3672
rect 1157 -3704 1187 -3672
rect 1253 -3704 1283 -3672
rect 1349 -3704 1379 -3672
rect -492 -3788 -462 -3762
rect 419 -3720 1445 -3704
rect 419 -3754 435 -3720
rect 469 -3754 627 -3720
rect 661 -3754 819 -3720
rect 853 -3754 1011 -3720
rect 1045 -3754 1203 -3720
rect 1237 -3754 1395 -3720
rect 1429 -3754 1445 -3720
rect 419 -3770 1445 -3754
rect 2006 -3400 2036 -3374
rect 2102 -3400 2132 -3374
rect 2198 -3400 2228 -3374
rect 2294 -3400 2324 -3374
rect 2390 -3400 2420 -3374
rect 2486 -3400 2516 -3374
rect 2582 -3400 2612 -3374
rect 2678 -3400 2708 -3374
rect 2774 -3400 2804 -3374
rect 2870 -3400 2900 -3374
rect 2006 -3704 2036 -3672
rect 2102 -3704 2132 -3672
rect 2198 -3704 2228 -3672
rect 2294 -3704 2324 -3672
rect 2390 -3704 2420 -3672
rect 2486 -3704 2516 -3672
rect 2582 -3704 2612 -3672
rect 2678 -3704 2708 -3672
rect 2774 -3704 2804 -3672
rect 2870 -3704 2900 -3672
rect 1940 -3720 2966 -3704
rect 1940 -3754 1956 -3720
rect 1990 -3754 2148 -3720
rect 2182 -3754 2340 -3720
rect 2374 -3754 2532 -3720
rect 2566 -3754 2724 -3720
rect 2758 -3754 2916 -3720
rect 2950 -3754 2966 -3720
rect 1940 -3770 2966 -3754
rect -492 -3940 -462 -3918
rect -548 -3956 -462 -3940
rect -548 -3990 -532 -3956
rect -498 -3990 -462 -3956
rect -548 -4006 -462 -3990
rect -492 -4038 -462 -4006
rect -3132 -4294 -2106 -4278
rect -3132 -4328 -3116 -4294
rect -3082 -4328 -2924 -4294
rect -2890 -4328 -2732 -4294
rect -2698 -4328 -2540 -4294
rect -2506 -4328 -2348 -4294
rect -2314 -4328 -2156 -4294
rect -2122 -4328 -2106 -4294
rect -3132 -4344 -2106 -4328
rect -492 -4264 -462 -4238
rect -3066 -4376 -3036 -4344
rect -2970 -4376 -2940 -4344
rect -2874 -4376 -2844 -4344
rect -2778 -4376 -2748 -4344
rect -2682 -4376 -2652 -4344
rect -2586 -4376 -2556 -4344
rect -2490 -4376 -2460 -4344
rect -2394 -4376 -2364 -4344
rect -2298 -4376 -2268 -4344
rect -2202 -4376 -2172 -4344
rect -3066 -4674 -3036 -4648
rect -2970 -4674 -2940 -4648
rect -2874 -4674 -2844 -4648
rect -2778 -4674 -2748 -4648
rect -2682 -4674 -2652 -4648
rect -2586 -4674 -2556 -4648
rect -2490 -4674 -2460 -4648
rect -2394 -4674 -2364 -4648
rect -2298 -4674 -2268 -4648
rect -2202 -4674 -2172 -4648
rect -492 -4332 -462 -4306
rect 419 -4290 1445 -4278
rect 419 -4324 435 -4290
rect 469 -4324 627 -4290
rect 661 -4324 819 -4290
rect 853 -4324 1011 -4290
rect 1045 -4324 1203 -4290
rect 1237 -4324 1395 -4290
rect 1429 -4324 1445 -4290
rect 419 -4344 1445 -4324
rect 485 -4366 515 -4344
rect 581 -4366 611 -4344
rect 677 -4366 707 -4344
rect 773 -4366 803 -4344
rect 869 -4366 899 -4344
rect 965 -4366 995 -4344
rect 1061 -4366 1091 -4344
rect 1157 -4366 1187 -4344
rect 1253 -4366 1283 -4344
rect 1349 -4366 1379 -4344
rect -492 -4564 -462 -4532
rect -548 -4580 -462 -4564
rect -548 -4614 -532 -4580
rect -498 -4614 -462 -4580
rect 485 -4496 515 -4470
rect 581 -4496 611 -4470
rect 677 -4496 707 -4470
rect 773 -4496 803 -4470
rect 869 -4496 899 -4470
rect 965 -4496 995 -4470
rect 1061 -4496 1091 -4470
rect 1157 -4496 1187 -4470
rect 1253 -4496 1283 -4470
rect 1349 -4496 1379 -4470
rect 1662 -4374 1692 -4348
rect 1662 -4496 1692 -4474
rect 1940 -4290 2966 -4278
rect 1940 -4324 1956 -4290
rect 1990 -4324 2148 -4290
rect 2182 -4324 2340 -4290
rect 2374 -4324 2532 -4290
rect 2566 -4324 2724 -4290
rect 2758 -4324 2916 -4290
rect 2950 -4324 2966 -4290
rect 1940 -4344 2966 -4324
rect 2006 -4366 2036 -4344
rect 2102 -4366 2132 -4344
rect 2198 -4366 2228 -4344
rect 2294 -4366 2324 -4344
rect 2390 -4366 2420 -4344
rect 2486 -4366 2516 -4344
rect 2582 -4366 2612 -4344
rect 2678 -4366 2708 -4344
rect 2774 -4366 2804 -4344
rect 2870 -4366 2900 -4344
rect 1644 -4512 1710 -4496
rect 1644 -4546 1660 -4512
rect 1694 -4546 1710 -4512
rect 1644 -4562 1710 -4546
rect 2006 -4496 2036 -4470
rect 2102 -4496 2132 -4470
rect 2198 -4496 2228 -4470
rect 2294 -4496 2324 -4470
rect 2390 -4496 2420 -4470
rect 2486 -4496 2516 -4470
rect 2582 -4496 2612 -4470
rect 2678 -4496 2708 -4470
rect 2774 -4496 2804 -4470
rect 2870 -4496 2900 -4470
rect -548 -4630 -462 -4614
rect -492 -4652 -462 -4630
rect -492 -4808 -462 -4782
rect -3066 -4956 -3036 -4930
rect -2970 -4956 -2940 -4930
rect -2874 -4956 -2844 -4930
rect -2778 -4956 -2748 -4930
rect -2682 -4956 -2652 -4930
rect -2586 -4956 -2556 -4930
rect -2490 -4956 -2460 -4930
rect -2394 -4956 -2364 -4930
rect -2298 -4956 -2268 -4930
rect -2202 -4956 -2172 -4930
rect -3066 -5082 -3036 -5060
rect -2970 -5082 -2940 -5060
rect -2874 -5082 -2844 -5060
rect -2778 -5082 -2748 -5060
rect -2682 -5082 -2652 -5060
rect -2586 -5082 -2556 -5060
rect -2490 -5082 -2460 -5060
rect -2394 -5082 -2364 -5060
rect -2298 -5082 -2268 -5060
rect -2202 -5082 -2172 -5060
rect -3132 -5102 -2106 -5082
rect -3132 -5136 -3116 -5102
rect -3082 -5136 -2924 -5102
rect -2890 -5136 -2732 -5102
rect -2698 -5136 -2540 -5102
rect -2506 -5136 -2348 -5102
rect -2314 -5136 -2156 -5102
rect -2122 -5136 -2106 -5102
rect -3132 -5148 -2106 -5136
rect 485 -4778 515 -4752
rect 581 -4778 611 -4752
rect 677 -4778 707 -4752
rect 773 -4778 803 -4752
rect 869 -4778 899 -4752
rect 965 -4778 995 -4752
rect 1061 -4778 1091 -4752
rect 1157 -4778 1187 -4752
rect 1253 -4778 1283 -4752
rect 1349 -4778 1379 -4752
rect 485 -5082 515 -5050
rect 581 -5082 611 -5050
rect 677 -5082 707 -5050
rect 773 -5082 803 -5050
rect 869 -5082 899 -5050
rect 965 -5082 995 -5050
rect 1061 -5082 1091 -5050
rect 1157 -5082 1187 -5050
rect 1253 -5082 1283 -5050
rect 1349 -5082 1379 -5050
rect 419 -5098 1445 -5082
rect 419 -5132 435 -5098
rect 469 -5132 627 -5098
rect 661 -5132 819 -5098
rect 853 -5132 1011 -5098
rect 1045 -5132 1203 -5098
rect 1237 -5132 1395 -5098
rect 1429 -5132 1445 -5098
rect 419 -5148 1445 -5132
rect 2006 -4778 2036 -4752
rect 2102 -4778 2132 -4752
rect 2198 -4778 2228 -4752
rect 2294 -4778 2324 -4752
rect 2390 -4778 2420 -4752
rect 2486 -4778 2516 -4752
rect 2582 -4778 2612 -4752
rect 2678 -4778 2708 -4752
rect 2774 -4778 2804 -4752
rect 2870 -4778 2900 -4752
rect 2006 -5082 2036 -5050
rect 2102 -5082 2132 -5050
rect 2198 -5082 2228 -5050
rect 2294 -5082 2324 -5050
rect 2390 -5082 2420 -5050
rect 2486 -5082 2516 -5050
rect 2582 -5082 2612 -5050
rect 2678 -5082 2708 -5050
rect 2774 -5082 2804 -5050
rect 2870 -5082 2900 -5050
rect 1940 -5098 2966 -5082
rect 1940 -5132 1956 -5098
rect 1990 -5132 2148 -5098
rect 2182 -5132 2340 -5098
rect 2374 -5132 2532 -5098
rect 2566 -5132 2724 -5098
rect 2758 -5132 2916 -5098
rect 2950 -5132 2966 -5098
rect 1940 -5148 2966 -5132
<< polycont >>
rect -3116 -238 -3082 -204
rect -2924 -238 -2890 -204
rect -2732 -238 -2698 -204
rect -2540 -238 -2506 -204
rect -2348 -238 -2314 -204
rect -2156 -238 -2122 -204
rect 435 -234 469 -200
rect 627 -234 661 -200
rect 819 -234 853 -200
rect 1011 -234 1045 -200
rect 1203 -234 1237 -200
rect 1395 -234 1429 -200
rect 1956 -234 1990 -200
rect 2148 -234 2182 -200
rect 2340 -234 2374 -200
rect 2532 -234 2566 -200
rect 2724 -234 2758 -200
rect 2916 -234 2950 -200
rect 1660 -456 1694 -422
rect -900 -726 -866 -692
rect -532 -726 -498 -692
rect -3116 -1046 -3082 -1012
rect -2924 -1046 -2890 -1012
rect -2732 -1046 -2698 -1012
rect -2540 -1046 -2506 -1012
rect -2348 -1046 -2314 -1012
rect -2156 -1046 -2122 -1012
rect 435 -1042 469 -1008
rect 627 -1042 661 -1008
rect 819 -1042 853 -1008
rect 1011 -1042 1045 -1008
rect 1203 -1042 1237 -1008
rect 1395 -1042 1429 -1008
rect 1956 -1042 1990 -1008
rect 2148 -1042 2182 -1008
rect 2340 -1042 2374 -1008
rect 2532 -1042 2566 -1008
rect 2724 -1042 2758 -1008
rect 2916 -1042 2950 -1008
rect -532 -1350 -498 -1316
rect -3116 -1572 -3082 -1538
rect -2924 -1572 -2890 -1538
rect -2732 -1572 -2698 -1538
rect -2540 -1572 -2506 -1538
rect -2348 -1572 -2314 -1538
rect -2156 -1572 -2122 -1538
rect 435 -1568 469 -1534
rect 627 -1568 661 -1534
rect 819 -1568 853 -1534
rect 1011 -1568 1045 -1534
rect 1203 -1568 1237 -1534
rect 1395 -1568 1429 -1534
rect -576 -1814 -542 -1780
rect -408 -1814 -374 -1780
rect 1956 -1568 1990 -1534
rect 2148 -1568 2182 -1534
rect 2340 -1568 2374 -1534
rect 2532 -1568 2566 -1534
rect 2724 -1568 2758 -1534
rect 2916 -1568 2950 -1534
rect 1660 -1790 1694 -1756
rect -3116 -2380 -3082 -2346
rect -2924 -2380 -2890 -2346
rect -2732 -2380 -2698 -2346
rect -2540 -2380 -2506 -2346
rect -2348 -2380 -2314 -2346
rect -2156 -2380 -2122 -2346
rect -1084 -2438 -1050 -2404
rect -576 -2438 -542 -2404
rect -408 -2438 -374 -2404
rect 435 -2376 469 -2342
rect 627 -2376 661 -2342
rect 819 -2376 853 -2342
rect 1011 -2376 1045 -2342
rect 1203 -2376 1237 -2342
rect 1395 -2376 1429 -2342
rect 1956 -2376 1990 -2342
rect 2148 -2376 2182 -2342
rect 2340 -2376 2374 -2342
rect 2532 -2376 2566 -2342
rect 2724 -2376 2758 -2342
rect 2916 -2376 2950 -2342
rect -3116 -2950 -3082 -2916
rect -2924 -2950 -2890 -2916
rect -2732 -2950 -2698 -2916
rect -2540 -2950 -2506 -2916
rect -2348 -2950 -2314 -2916
rect -2156 -2950 -2122 -2916
rect -1084 -2902 -1050 -2868
rect -576 -2902 -542 -2868
rect -408 -2902 -374 -2868
rect 435 -2946 469 -2912
rect 627 -2946 661 -2912
rect 819 -2946 853 -2912
rect 1011 -2946 1045 -2912
rect 1203 -2946 1237 -2912
rect 1395 -2946 1429 -2912
rect 1956 -2946 1990 -2912
rect 2148 -2946 2182 -2912
rect 2340 -2946 2374 -2912
rect 2532 -2946 2566 -2912
rect 2724 -2946 2758 -2912
rect 2916 -2946 2950 -2912
rect 1660 -3168 1694 -3134
rect -576 -3526 -542 -3492
rect -3116 -3758 -3082 -3724
rect -2924 -3758 -2890 -3724
rect -2732 -3758 -2698 -3724
rect -2540 -3758 -2506 -3724
rect -2348 -3758 -2314 -3724
rect -2156 -3758 -2122 -3724
rect -408 -3526 -374 -3492
rect 435 -3754 469 -3720
rect 627 -3754 661 -3720
rect 819 -3754 853 -3720
rect 1011 -3754 1045 -3720
rect 1203 -3754 1237 -3720
rect 1395 -3754 1429 -3720
rect 1956 -3754 1990 -3720
rect 2148 -3754 2182 -3720
rect 2340 -3754 2374 -3720
rect 2532 -3754 2566 -3720
rect 2724 -3754 2758 -3720
rect 2916 -3754 2950 -3720
rect -532 -3990 -498 -3956
rect -3116 -4328 -3082 -4294
rect -2924 -4328 -2890 -4294
rect -2732 -4328 -2698 -4294
rect -2540 -4328 -2506 -4294
rect -2348 -4328 -2314 -4294
rect -2156 -4328 -2122 -4294
rect 435 -4324 469 -4290
rect 627 -4324 661 -4290
rect 819 -4324 853 -4290
rect 1011 -4324 1045 -4290
rect 1203 -4324 1237 -4290
rect 1395 -4324 1429 -4290
rect -532 -4614 -498 -4580
rect 1956 -4324 1990 -4290
rect 2148 -4324 2182 -4290
rect 2340 -4324 2374 -4290
rect 2532 -4324 2566 -4290
rect 2724 -4324 2758 -4290
rect 2916 -4324 2950 -4290
rect 1660 -4546 1694 -4512
rect -3116 -5136 -3082 -5102
rect -2924 -5136 -2890 -5102
rect -2732 -5136 -2698 -5102
rect -2540 -5136 -2506 -5102
rect -2348 -5136 -2314 -5102
rect -2156 -5136 -2122 -5102
rect 435 -5132 469 -5098
rect 627 -5132 661 -5098
rect 819 -5132 853 -5098
rect 1011 -5132 1045 -5098
rect 1203 -5132 1237 -5098
rect 1395 -5132 1429 -5098
rect 1956 -5132 1990 -5098
rect 2148 -5132 2182 -5098
rect 2340 -5132 2374 -5098
rect 2532 -5132 2566 -5098
rect 2724 -5132 2758 -5098
rect 2916 -5132 2950 -5098
<< locali >>
rect -3230 -136 -3134 -102
rect -2104 -136 -2008 -102
rect -3230 -198 -3196 -136
rect -2042 -198 -2008 -136
rect -3132 -238 -3116 -204
rect -3082 -238 -3066 -204
rect -2940 -238 -2924 -204
rect -2890 -238 -2874 -204
rect -2748 -238 -2732 -204
rect -2698 -238 -2682 -204
rect -2556 -238 -2540 -204
rect -2506 -238 -2490 -204
rect -2364 -238 -2348 -204
rect -2314 -238 -2298 -204
rect -2172 -238 -2156 -204
rect -2122 -238 -2106 -204
rect -3116 -298 -3082 -282
rect -3116 -562 -3082 -546
rect -3020 -298 -2986 -282
rect -3020 -562 -2986 -546
rect -2924 -298 -2890 -282
rect -2924 -562 -2890 -546
rect -2828 -298 -2794 -282
rect -2828 -562 -2794 -546
rect -2732 -298 -2698 -282
rect -2732 -562 -2698 -546
rect -2636 -298 -2602 -282
rect -2636 -562 -2602 -546
rect -2540 -298 -2506 -282
rect -2540 -562 -2506 -546
rect -2444 -298 -2410 -282
rect -2444 -562 -2410 -546
rect -2348 -298 -2314 -282
rect -2348 -562 -2314 -546
rect -2252 -298 -2218 -282
rect -2252 -562 -2218 -546
rect -2156 -298 -2122 -282
rect -2156 -562 -2122 -546
rect -3230 -646 -3196 -584
rect 321 -136 417 -102
rect 1447 -136 1543 -102
rect 321 -198 355 -136
rect 1509 -198 1543 -136
rect 419 -234 435 -200
rect 469 -234 485 -200
rect 611 -234 627 -200
rect 661 -234 677 -200
rect 803 -234 819 -200
rect 853 -234 869 -200
rect 995 -234 1011 -200
rect 1045 -234 1061 -200
rect 1187 -234 1203 -200
rect 1237 -234 1253 -200
rect 1379 -234 1395 -200
rect 1429 -234 1445 -200
rect 435 -288 469 -272
rect 435 -384 469 -368
rect 531 -288 565 -272
rect 531 -384 565 -368
rect 627 -288 661 -272
rect 627 -384 661 -368
rect 723 -288 757 -272
rect 723 -384 757 -368
rect 819 -288 853 -272
rect 819 -384 853 -368
rect 915 -288 949 -272
rect 915 -384 949 -368
rect 1011 -288 1045 -272
rect 1011 -384 1045 -368
rect 1107 -288 1141 -272
rect 1107 -384 1141 -368
rect 1203 -288 1237 -272
rect 1203 -384 1237 -368
rect 1299 -288 1333 -272
rect 1299 -384 1333 -368
rect 1395 -288 1429 -272
rect 1395 -384 1429 -368
rect 321 -458 355 -396
rect 1842 -136 1938 -102
rect 2968 -136 3064 -102
rect 1842 -198 1876 -136
rect 1616 -296 1650 -280
rect 1616 -388 1650 -372
rect 1704 -296 1738 -280
rect 1704 -388 1738 -372
rect 1509 -458 1543 -398
rect 3030 -198 3064 -136
rect 1940 -234 1956 -200
rect 1990 -234 2006 -200
rect 2132 -234 2148 -200
rect 2182 -234 2198 -200
rect 2324 -234 2340 -200
rect 2374 -234 2390 -200
rect 2516 -234 2532 -200
rect 2566 -234 2582 -200
rect 2708 -234 2724 -200
rect 2758 -234 2774 -200
rect 2900 -234 2916 -200
rect 2950 -234 2966 -200
rect 1956 -288 1990 -272
rect 1956 -384 1990 -368
rect 2052 -288 2086 -272
rect 2052 -384 2086 -368
rect 2148 -288 2182 -272
rect 2148 -384 2182 -368
rect 2244 -288 2278 -272
rect 2244 -384 2278 -368
rect 2340 -288 2374 -272
rect 2340 -384 2374 -368
rect 2436 -288 2470 -272
rect 2436 -384 2470 -368
rect 2532 -288 2566 -272
rect 2532 -384 2566 -368
rect 2628 -288 2662 -272
rect 2628 -384 2662 -368
rect 2724 -288 2758 -272
rect 2724 -384 2758 -368
rect 2820 -288 2854 -272
rect 2820 -384 2854 -368
rect 2916 -288 2950 -272
rect 2916 -384 2950 -368
rect 1644 -456 1660 -422
rect 1694 -456 1710 -422
rect -980 -494 -951 -460
rect -917 -494 -859 -460
rect -825 -494 -767 -460
rect -733 -494 -675 -460
rect -641 -494 -583 -460
rect -549 -494 -491 -460
rect -457 -494 -399 -460
rect -365 -494 -336 -460
rect 321 -492 417 -458
rect 1447 -492 1543 -458
rect 1842 -458 1876 -396
rect 3030 -458 3064 -398
rect 1842 -492 1938 -458
rect 2968 -492 3064 -458
rect -2042 -646 -2008 -584
rect -3230 -680 -3134 -646
rect -2104 -680 -2008 -646
rect -916 -540 -870 -494
rect -916 -574 -904 -540
rect -916 -608 -870 -574
rect -916 -642 -904 -608
rect -916 -658 -870 -642
rect -836 -540 -770 -528
rect -836 -574 -820 -540
rect -786 -574 -770 -540
rect -836 -603 -770 -574
rect -836 -637 -822 -603
rect -788 -608 -770 -603
rect -836 -642 -820 -637
rect -786 -642 -770 -608
rect -687 -588 -629 -494
rect -687 -622 -675 -588
rect -641 -622 -629 -588
rect -687 -639 -629 -622
rect -548 -540 -502 -494
rect -548 -574 -536 -540
rect -548 -608 -502 -574
rect -836 -654 -770 -642
rect -916 -698 -900 -692
rect -916 -732 -905 -698
rect -866 -726 -850 -692
rect -871 -732 -850 -726
rect -916 -740 -850 -732
rect -3230 -788 -3134 -754
rect -2104 -788 -2008 -754
rect -816 -774 -770 -654
rect -548 -642 -536 -608
rect -548 -658 -502 -642
rect -468 -540 -402 -528
rect -468 -574 -452 -540
rect -418 -574 -402 -540
rect -468 -594 -402 -574
rect -468 -642 -452 -594
rect -418 -642 -402 -594
rect -468 -654 -402 -642
rect -548 -700 -532 -692
rect -548 -734 -538 -700
rect -498 -726 -482 -692
rect -504 -734 -482 -726
rect -548 -740 -482 -734
rect -3230 -850 -3196 -788
rect -2042 -848 -2008 -788
rect -3116 -878 -3082 -862
rect -3116 -974 -3082 -958
rect -3020 -878 -2986 -862
rect -3020 -974 -2986 -958
rect -2924 -878 -2890 -862
rect -2924 -974 -2890 -958
rect -2828 -878 -2794 -862
rect -2828 -974 -2794 -958
rect -2732 -878 -2698 -862
rect -2732 -974 -2698 -958
rect -2636 -878 -2602 -862
rect -2636 -974 -2602 -958
rect -2540 -878 -2506 -862
rect -2540 -974 -2506 -958
rect -2444 -878 -2410 -862
rect -2444 -974 -2410 -958
rect -2348 -878 -2314 -862
rect -2348 -974 -2314 -958
rect -2252 -878 -2218 -862
rect -2252 -974 -2218 -958
rect -2156 -878 -2122 -862
rect -2156 -974 -2122 -958
rect -3132 -1046 -3116 -1012
rect -3082 -1046 -3066 -1012
rect -2940 -1046 -2924 -1012
rect -2890 -1046 -2874 -1012
rect -2748 -1046 -2732 -1012
rect -2698 -1046 -2682 -1012
rect -2556 -1046 -2540 -1012
rect -2506 -1046 -2490 -1012
rect -2364 -1046 -2348 -1012
rect -2314 -1046 -2298 -1012
rect -2172 -1046 -2156 -1012
rect -2122 -1046 -2106 -1012
rect -3230 -1110 -3196 -1048
rect -912 -792 -870 -776
rect -912 -826 -904 -792
rect -912 -860 -870 -826
rect -912 -894 -904 -860
rect -912 -928 -870 -894
rect -912 -962 -904 -928
rect -912 -1004 -870 -962
rect -836 -792 -770 -774
rect -836 -826 -820 -792
rect -786 -826 -770 -792
rect -836 -860 -770 -826
rect -836 -894 -820 -860
rect -786 -894 -770 -860
rect -836 -928 -770 -894
rect -836 -962 -820 -928
rect -786 -962 -770 -928
rect -836 -970 -770 -962
rect -687 -806 -629 -771
rect -448 -774 -402 -654
rect -687 -840 -675 -806
rect -641 -840 -629 -806
rect -687 -899 -629 -840
rect -687 -933 -675 -899
rect -641 -933 -629 -899
rect -687 -1004 -629 -933
rect -544 -792 -502 -776
rect -544 -826 -536 -792
rect -544 -860 -502 -826
rect -544 -894 -536 -860
rect -544 -928 -502 -894
rect -544 -962 -536 -928
rect -544 -1004 -502 -962
rect -468 -792 -402 -774
rect -468 -826 -452 -792
rect -418 -826 -402 -792
rect -468 -860 -402 -826
rect -468 -894 -452 -860
rect -418 -894 -402 -860
rect -468 -928 -402 -894
rect -468 -962 -452 -928
rect -418 -962 -402 -928
rect -468 -970 -402 -962
rect 321 -600 417 -566
rect 1447 -600 1543 -566
rect 321 -662 355 -600
rect -980 -1038 -951 -1004
rect -917 -1038 -859 -1004
rect -825 -1038 -767 -1004
rect -733 -1038 -675 -1004
rect -641 -1038 -583 -1004
rect -549 -1038 -491 -1004
rect -457 -1038 -399 -1004
rect -365 -1038 -336 -1004
rect -2042 -1110 -2008 -1048
rect -3230 -1144 -3134 -1110
rect -2104 -1144 -2008 -1110
rect -687 -1109 -629 -1038
rect -687 -1143 -675 -1109
rect -641 -1143 -629 -1109
rect -687 -1202 -629 -1143
rect -687 -1236 -675 -1202
rect -641 -1236 -629 -1202
rect -687 -1271 -629 -1236
rect -544 -1080 -502 -1038
rect 1509 -662 1543 -600
rect 435 -700 469 -684
rect 435 -964 469 -948
rect 531 -700 565 -684
rect 531 -964 565 -948
rect 627 -700 661 -684
rect 627 -964 661 -948
rect 723 -700 757 -684
rect 723 -964 757 -948
rect 819 -700 853 -684
rect 819 -964 853 -948
rect 915 -700 949 -684
rect 915 -964 949 -948
rect 1011 -700 1045 -684
rect 1011 -964 1045 -948
rect 1107 -700 1141 -684
rect 1107 -964 1141 -948
rect 1203 -700 1237 -684
rect 1203 -964 1237 -948
rect 1299 -700 1333 -684
rect 1299 -964 1333 -948
rect 1395 -700 1429 -684
rect 1395 -964 1429 -948
rect 419 -1042 435 -1008
rect 469 -1042 485 -1008
rect 611 -1042 627 -1008
rect 661 -1042 677 -1008
rect 803 -1042 819 -1008
rect 853 -1042 869 -1008
rect 995 -1042 1011 -1008
rect 1045 -1042 1061 -1008
rect 1187 -1042 1203 -1008
rect 1237 -1042 1253 -1008
rect 1379 -1042 1395 -1008
rect 1429 -1042 1445 -1008
rect -544 -1114 -536 -1080
rect -544 -1148 -502 -1114
rect -544 -1182 -536 -1148
rect -544 -1216 -502 -1182
rect -544 -1250 -536 -1216
rect -544 -1266 -502 -1250
rect -468 -1080 -402 -1072
rect -468 -1114 -452 -1080
rect -418 -1114 -402 -1080
rect -468 -1148 -402 -1114
rect 321 -1110 355 -1048
rect 1509 -1110 1543 -1048
rect 321 -1144 417 -1110
rect 1447 -1144 1543 -1110
rect 1842 -600 1938 -566
rect 2968 -600 3064 -566
rect 1842 -662 1876 -600
rect 3030 -662 3064 -600
rect 1956 -700 1990 -684
rect 1956 -964 1990 -948
rect 2052 -700 2086 -684
rect 2052 -964 2086 -948
rect 2148 -700 2182 -684
rect 2148 -964 2182 -948
rect 2244 -700 2278 -684
rect 2244 -964 2278 -948
rect 2340 -700 2374 -684
rect 2340 -964 2374 -948
rect 2436 -700 2470 -684
rect 2436 -964 2470 -948
rect 2532 -700 2566 -684
rect 2532 -964 2566 -948
rect 2628 -700 2662 -684
rect 2628 -964 2662 -948
rect 2724 -700 2758 -684
rect 2724 -964 2758 -948
rect 2820 -700 2854 -684
rect 2820 -964 2854 -948
rect 2916 -700 2950 -684
rect 2916 -964 2950 -948
rect 1940 -1042 1956 -1008
rect 1990 -1042 2006 -1008
rect 2132 -1042 2148 -1008
rect 2182 -1042 2198 -1008
rect 2324 -1042 2340 -1008
rect 2374 -1042 2390 -1008
rect 2516 -1042 2532 -1008
rect 2566 -1042 2582 -1008
rect 2708 -1042 2724 -1008
rect 2758 -1042 2774 -1008
rect 2900 -1042 2916 -1008
rect 2950 -1042 2966 -1008
rect 1842 -1110 1876 -1048
rect 3030 -1110 3064 -1048
rect 1842 -1144 1938 -1110
rect 2968 -1144 3064 -1110
rect -468 -1182 -452 -1148
rect -418 -1182 -402 -1148
rect -468 -1197 -402 -1182
rect -468 -1231 -453 -1197
rect -419 -1216 -402 -1197
rect -468 -1250 -452 -1231
rect -418 -1250 -402 -1216
rect -468 -1268 -402 -1250
rect -548 -1312 -482 -1302
rect -548 -1346 -534 -1312
rect -500 -1316 -482 -1312
rect -548 -1350 -532 -1346
rect -498 -1350 -482 -1316
rect -548 -1400 -502 -1384
rect -448 -1388 -402 -1268
rect -687 -1420 -629 -1403
rect -3230 -1470 -3134 -1436
rect -2104 -1470 -2008 -1436
rect -3230 -1532 -3196 -1470
rect -2042 -1532 -2008 -1470
rect -3132 -1572 -3116 -1538
rect -3082 -1572 -3066 -1538
rect -2940 -1572 -2924 -1538
rect -2890 -1572 -2874 -1538
rect -2748 -1572 -2732 -1538
rect -2698 -1572 -2682 -1538
rect -2556 -1572 -2540 -1538
rect -2506 -1572 -2490 -1538
rect -2364 -1572 -2348 -1538
rect -2314 -1572 -2298 -1538
rect -2172 -1572 -2156 -1538
rect -2122 -1572 -2106 -1538
rect -3116 -1632 -3082 -1616
rect -3116 -1896 -3082 -1880
rect -3020 -1632 -2986 -1616
rect -3020 -1896 -2986 -1880
rect -2924 -1632 -2890 -1616
rect -2924 -1896 -2890 -1880
rect -2828 -1632 -2794 -1616
rect -2828 -1896 -2794 -1880
rect -2732 -1632 -2698 -1616
rect -2732 -1896 -2698 -1880
rect -2636 -1632 -2602 -1616
rect -2636 -1896 -2602 -1880
rect -2540 -1632 -2506 -1616
rect -2540 -1896 -2506 -1880
rect -2444 -1632 -2410 -1616
rect -2444 -1896 -2410 -1880
rect -2348 -1632 -2314 -1616
rect -2348 -1896 -2314 -1880
rect -2252 -1632 -2218 -1616
rect -2252 -1896 -2218 -1880
rect -2156 -1632 -2122 -1616
rect -2156 -1896 -2122 -1880
rect -3230 -1980 -3196 -1918
rect -687 -1454 -675 -1420
rect -641 -1454 -629 -1420
rect -687 -1548 -629 -1454
rect -548 -1434 -536 -1400
rect -548 -1468 -502 -1434
rect -548 -1502 -536 -1468
rect -548 -1548 -502 -1502
rect -468 -1400 -402 -1388
rect -468 -1434 -452 -1400
rect -418 -1434 -402 -1400
rect -468 -1468 -402 -1434
rect -468 -1502 -452 -1468
rect -418 -1502 -402 -1468
rect -468 -1514 -402 -1502
rect 321 -1470 417 -1436
rect 1447 -1470 1543 -1436
rect 321 -1532 355 -1470
rect -704 -1582 -675 -1548
rect -641 -1582 -583 -1548
rect -549 -1582 -491 -1548
rect -457 -1582 -399 -1548
rect -365 -1582 -336 -1548
rect -687 -1676 -629 -1582
rect -687 -1710 -675 -1676
rect -641 -1710 -629 -1676
rect -687 -1727 -629 -1710
rect -595 -1624 -533 -1582
rect -595 -1658 -573 -1624
rect -539 -1658 -533 -1624
rect -595 -1692 -533 -1658
rect -595 -1726 -573 -1692
rect -539 -1726 -533 -1692
rect -595 -1742 -533 -1726
rect -492 -1624 -353 -1616
rect -492 -1658 -405 -1624
rect -371 -1658 -353 -1624
rect -492 -1676 -353 -1658
rect -492 -1710 -469 -1676
rect -435 -1692 -353 -1676
rect -435 -1710 -405 -1692
rect -492 -1726 -405 -1710
rect -371 -1726 -353 -1692
rect -492 -1742 -353 -1726
rect 1509 -1532 1543 -1470
rect 419 -1568 435 -1534
rect 469 -1568 485 -1534
rect 611 -1568 627 -1534
rect 661 -1568 677 -1534
rect 803 -1568 819 -1534
rect 853 -1568 869 -1534
rect 995 -1568 1011 -1534
rect 1045 -1568 1061 -1534
rect 1187 -1568 1203 -1534
rect 1237 -1568 1253 -1534
rect 1379 -1568 1395 -1534
rect 1429 -1568 1445 -1534
rect 435 -1622 469 -1606
rect 435 -1718 469 -1702
rect 531 -1622 565 -1606
rect 531 -1718 565 -1702
rect 627 -1622 661 -1606
rect 627 -1718 661 -1702
rect 723 -1622 757 -1606
rect 723 -1718 757 -1702
rect 819 -1622 853 -1606
rect 819 -1718 853 -1702
rect 915 -1622 949 -1606
rect 915 -1718 949 -1702
rect 1011 -1622 1045 -1606
rect 1011 -1718 1045 -1702
rect 1107 -1622 1141 -1606
rect 1107 -1718 1141 -1702
rect 1203 -1622 1237 -1606
rect 1203 -1718 1237 -1702
rect 1299 -1622 1333 -1606
rect 1299 -1718 1333 -1702
rect 1395 -1622 1429 -1606
rect 1395 -1718 1429 -1702
rect -593 -1780 -526 -1776
rect -593 -1784 -576 -1780
rect -593 -1818 -582 -1784
rect -542 -1814 -526 -1780
rect -548 -1818 -526 -1814
rect -593 -1830 -526 -1818
rect -2042 -1980 -2008 -1918
rect -3230 -2014 -3134 -1980
rect -2104 -2014 -2008 -1980
rect -687 -1894 -629 -1859
rect -492 -1862 -458 -1742
rect -424 -1819 -408 -1780
rect -374 -1819 -357 -1780
rect -424 -1830 -357 -1819
rect 321 -1792 355 -1730
rect 1842 -1470 1938 -1436
rect 2968 -1470 3064 -1436
rect 1842 -1532 1876 -1470
rect 1616 -1630 1650 -1614
rect 1616 -1722 1650 -1706
rect 1704 -1630 1738 -1614
rect 1704 -1722 1738 -1706
rect 1509 -1792 1543 -1732
rect 3030 -1532 3064 -1470
rect 1940 -1568 1956 -1534
rect 1990 -1568 2006 -1534
rect 2132 -1568 2148 -1534
rect 2182 -1568 2198 -1534
rect 2324 -1568 2340 -1534
rect 2374 -1568 2390 -1534
rect 2516 -1568 2532 -1534
rect 2566 -1568 2582 -1534
rect 2708 -1568 2724 -1534
rect 2758 -1568 2774 -1534
rect 2900 -1568 2916 -1534
rect 2950 -1568 2966 -1534
rect 1956 -1622 1990 -1606
rect 1956 -1718 1990 -1702
rect 2052 -1622 2086 -1606
rect 2052 -1718 2086 -1702
rect 2148 -1622 2182 -1606
rect 2148 -1718 2182 -1702
rect 2244 -1622 2278 -1606
rect 2244 -1718 2278 -1702
rect 2340 -1622 2374 -1606
rect 2340 -1718 2374 -1702
rect 2436 -1622 2470 -1606
rect 2436 -1718 2470 -1702
rect 2532 -1622 2566 -1606
rect 2532 -1718 2566 -1702
rect 2628 -1622 2662 -1606
rect 2628 -1718 2662 -1702
rect 2724 -1622 2758 -1606
rect 2724 -1718 2758 -1702
rect 2820 -1622 2854 -1606
rect 2820 -1718 2854 -1702
rect 2916 -1622 2950 -1606
rect 2916 -1718 2950 -1702
rect 1644 -1790 1660 -1756
rect 1694 -1790 1710 -1756
rect 321 -1826 417 -1792
rect 1447 -1826 1543 -1792
rect 1842 -1792 1876 -1730
rect 3030 -1792 3064 -1732
rect 1842 -1826 1938 -1792
rect 2968 -1826 3064 -1792
rect -687 -1928 -675 -1894
rect -641 -1928 -629 -1894
rect -687 -1987 -629 -1928
rect -687 -2021 -675 -1987
rect -641 -2021 -629 -1987
rect -3230 -2122 -3134 -2088
rect -2104 -2122 -2008 -2088
rect -687 -2092 -629 -2021
rect -595 -1880 -539 -1864
rect -595 -1914 -573 -1880
rect -595 -1948 -539 -1914
rect -595 -1982 -573 -1948
rect -595 -2016 -539 -1982
rect -595 -2050 -573 -2016
rect -595 -2092 -539 -2050
rect -505 -1880 -439 -1862
rect -505 -1914 -489 -1880
rect -455 -1914 -439 -1880
rect -505 -1948 -439 -1914
rect -505 -1982 -489 -1948
rect -455 -1982 -439 -1948
rect -505 -2016 -439 -1982
rect -505 -2050 -489 -2016
rect -455 -2050 -439 -2016
rect -505 -2058 -439 -2050
rect -405 -1880 -353 -1864
rect -371 -1914 -353 -1880
rect -405 -1948 -353 -1914
rect -371 -1982 -353 -1948
rect -405 -2016 -353 -1982
rect -371 -2050 -353 -2016
rect -405 -2092 -353 -2050
rect 321 -1934 417 -1900
rect 1447 -1934 1543 -1900
rect 321 -1996 355 -1934
rect -3230 -2184 -3196 -2122
rect -2042 -2182 -2008 -2122
rect -1256 -2126 -1227 -2092
rect -1193 -2126 -1135 -2092
rect -1101 -2126 -1043 -2092
rect -1009 -2126 -951 -2092
rect -917 -2126 -859 -2092
rect -825 -2126 -767 -2092
rect -733 -2126 -675 -2092
rect -641 -2126 -583 -2092
rect -549 -2126 -491 -2092
rect -457 -2126 -399 -2092
rect -365 -2126 -336 -2092
rect -3116 -2212 -3082 -2196
rect -3116 -2308 -3082 -2292
rect -3020 -2212 -2986 -2196
rect -3020 -2308 -2986 -2292
rect -2924 -2212 -2890 -2196
rect -2924 -2308 -2890 -2292
rect -2828 -2212 -2794 -2196
rect -2828 -2308 -2794 -2292
rect -2732 -2212 -2698 -2196
rect -2732 -2308 -2698 -2292
rect -2636 -2212 -2602 -2196
rect -2636 -2308 -2602 -2292
rect -2540 -2212 -2506 -2196
rect -2540 -2308 -2506 -2292
rect -2444 -2212 -2410 -2196
rect -2444 -2308 -2410 -2292
rect -2348 -2212 -2314 -2196
rect -2348 -2308 -2314 -2292
rect -2252 -2212 -2218 -2196
rect -2252 -2308 -2218 -2292
rect -2156 -2212 -2122 -2196
rect -2156 -2308 -2122 -2292
rect -3132 -2380 -3116 -2346
rect -3082 -2380 -3066 -2346
rect -2940 -2380 -2924 -2346
rect -2890 -2380 -2874 -2346
rect -2748 -2380 -2732 -2346
rect -2698 -2380 -2682 -2346
rect -2556 -2380 -2540 -2346
rect -2506 -2380 -2490 -2346
rect -2364 -2380 -2348 -2346
rect -2314 -2380 -2298 -2346
rect -2172 -2380 -2156 -2346
rect -2122 -2380 -2106 -2346
rect -3230 -2444 -3196 -2382
rect -1239 -2197 -1181 -2126
rect -1239 -2231 -1227 -2197
rect -1193 -2231 -1181 -2197
rect -1239 -2290 -1181 -2231
rect -1239 -2324 -1227 -2290
rect -1193 -2324 -1181 -2290
rect -1239 -2359 -1181 -2324
rect -1096 -2168 -1054 -2126
rect -1096 -2202 -1088 -2168
rect -1096 -2236 -1054 -2202
rect -1096 -2270 -1088 -2236
rect -1096 -2304 -1054 -2270
rect -1096 -2338 -1088 -2304
rect -1096 -2354 -1054 -2338
rect -1020 -2168 -954 -2160
rect -1020 -2202 -1004 -2168
rect -970 -2202 -954 -2168
rect -1020 -2236 -954 -2202
rect -1020 -2270 -1004 -2236
rect -970 -2270 -954 -2236
rect -1020 -2304 -954 -2270
rect -1020 -2338 -1004 -2304
rect -970 -2338 -954 -2304
rect -1020 -2356 -954 -2338
rect -2042 -2444 -2008 -2382
rect -1100 -2398 -1034 -2390
rect -1100 -2432 -1091 -2398
rect -1057 -2404 -1034 -2398
rect -1100 -2438 -1084 -2432
rect -1050 -2438 -1034 -2404
rect -3230 -2478 -3134 -2444
rect -2104 -2478 -2008 -2444
rect -1100 -2488 -1054 -2472
rect -1000 -2476 -954 -2356
rect -687 -2197 -629 -2126
rect -687 -2231 -675 -2197
rect -641 -2231 -629 -2197
rect -687 -2290 -629 -2231
rect -687 -2324 -675 -2290
rect -641 -2324 -629 -2290
rect -687 -2359 -629 -2324
rect -595 -2168 -539 -2126
rect -595 -2202 -573 -2168
rect -595 -2236 -539 -2202
rect -595 -2270 -573 -2236
rect -595 -2304 -539 -2270
rect -595 -2338 -573 -2304
rect -595 -2354 -539 -2338
rect -505 -2168 -439 -2160
rect -505 -2202 -489 -2168
rect -455 -2202 -439 -2168
rect -505 -2236 -439 -2202
rect -505 -2338 -489 -2236
rect -455 -2338 -439 -2236
rect -505 -2356 -439 -2338
rect -405 -2168 -353 -2126
rect -371 -2202 -353 -2168
rect -405 -2236 -353 -2202
rect -371 -2270 -353 -2236
rect -405 -2304 -353 -2270
rect -371 -2338 -353 -2304
rect -405 -2354 -353 -2338
rect -593 -2398 -526 -2388
rect -593 -2432 -583 -2398
rect -549 -2404 -526 -2398
rect -593 -2438 -576 -2432
rect -542 -2438 -526 -2404
rect -593 -2442 -526 -2438
rect -492 -2476 -458 -2356
rect 1509 -1996 1543 -1934
rect 435 -2034 469 -2018
rect 435 -2298 469 -2282
rect 531 -2034 565 -2018
rect 531 -2298 565 -2282
rect 627 -2034 661 -2018
rect 627 -2298 661 -2282
rect 723 -2034 757 -2018
rect 723 -2298 757 -2282
rect 819 -2034 853 -2018
rect 819 -2298 853 -2282
rect 915 -2034 949 -2018
rect 915 -2298 949 -2282
rect 1011 -2034 1045 -2018
rect 1011 -2298 1045 -2282
rect 1107 -2034 1141 -2018
rect 1107 -2298 1141 -2282
rect 1203 -2034 1237 -2018
rect 1203 -2298 1237 -2282
rect 1299 -2034 1333 -2018
rect 1299 -2298 1333 -2282
rect 1395 -2034 1429 -2018
rect 1395 -2298 1429 -2282
rect 419 -2376 435 -2342
rect 469 -2376 485 -2342
rect 611 -2376 627 -2342
rect 661 -2376 677 -2342
rect 803 -2376 819 -2342
rect 853 -2376 869 -2342
rect 995 -2376 1011 -2342
rect 1045 -2376 1061 -2342
rect 1187 -2376 1203 -2342
rect 1237 -2376 1253 -2342
rect 1379 -2376 1395 -2342
rect 1429 -2376 1445 -2342
rect -424 -2395 -357 -2388
rect -424 -2404 -402 -2395
rect -424 -2438 -408 -2404
rect -368 -2429 -357 -2395
rect -374 -2438 -357 -2429
rect 321 -2444 355 -2382
rect 1509 -2444 1543 -2382
rect -1239 -2508 -1181 -2491
rect -1239 -2542 -1227 -2508
rect -1193 -2542 -1181 -2508
rect -1239 -2636 -1181 -2542
rect -1100 -2522 -1088 -2488
rect -1100 -2556 -1054 -2522
rect -1100 -2590 -1088 -2556
rect -1100 -2636 -1054 -2590
rect -1020 -2488 -954 -2476
rect -1020 -2522 -1004 -2488
rect -970 -2522 -954 -2488
rect -1020 -2556 -954 -2522
rect -1020 -2590 -1004 -2556
rect -970 -2590 -954 -2556
rect -1020 -2602 -954 -2590
rect -687 -2508 -629 -2491
rect -687 -2542 -675 -2508
rect -641 -2542 -629 -2508
rect -687 -2636 -629 -2542
rect -595 -2492 -533 -2476
rect -595 -2526 -573 -2492
rect -539 -2526 -533 -2492
rect -595 -2560 -533 -2526
rect -595 -2594 -573 -2560
rect -539 -2594 -533 -2560
rect -595 -2636 -533 -2594
rect -492 -2492 -353 -2476
rect 321 -2478 417 -2444
rect 1447 -2478 1543 -2444
rect 1842 -1934 1938 -1900
rect 2968 -1934 3064 -1900
rect 1842 -1996 1876 -1934
rect 3030 -1996 3064 -1934
rect 1956 -2034 1990 -2018
rect 1956 -2298 1990 -2282
rect 2052 -2034 2086 -2018
rect 2052 -2298 2086 -2282
rect 2148 -2034 2182 -2018
rect 2148 -2298 2182 -2282
rect 2244 -2034 2278 -2018
rect 2244 -2298 2278 -2282
rect 2340 -2034 2374 -2018
rect 2340 -2298 2374 -2282
rect 2436 -2034 2470 -2018
rect 2436 -2298 2470 -2282
rect 2532 -2034 2566 -2018
rect 2532 -2298 2566 -2282
rect 2628 -2034 2662 -2018
rect 2628 -2298 2662 -2282
rect 2724 -2034 2758 -2018
rect 2724 -2298 2758 -2282
rect 2820 -2034 2854 -2018
rect 2820 -2298 2854 -2282
rect 2916 -2034 2950 -2018
rect 2916 -2298 2950 -2282
rect 1940 -2376 1956 -2342
rect 1990 -2376 2006 -2342
rect 2132 -2376 2148 -2342
rect 2182 -2376 2198 -2342
rect 2324 -2376 2340 -2342
rect 2374 -2376 2390 -2342
rect 2516 -2376 2532 -2342
rect 2566 -2376 2582 -2342
rect 2708 -2376 2724 -2342
rect 2758 -2376 2774 -2342
rect 2900 -2376 2916 -2342
rect 2950 -2376 2966 -2342
rect 1842 -2444 1876 -2382
rect 3030 -2444 3064 -2382
rect 1842 -2478 1938 -2444
rect 2968 -2478 3064 -2444
rect -492 -2526 -405 -2492
rect -371 -2526 -353 -2492
rect -492 -2560 -353 -2526
rect -492 -2594 -405 -2560
rect -371 -2594 -353 -2560
rect -492 -2602 -353 -2594
rect -1256 -2670 -1227 -2636
rect -1193 -2670 -1135 -2636
rect -1101 -2670 -1043 -2636
rect -1009 -2670 -951 -2636
rect -917 -2670 -859 -2636
rect -825 -2670 -767 -2636
rect -733 -2670 -675 -2636
rect -641 -2670 -583 -2636
rect -549 -2670 -491 -2636
rect -457 -2670 -399 -2636
rect -365 -2670 -336 -2636
rect -1239 -2764 -1181 -2670
rect -1239 -2798 -1227 -2764
rect -1193 -2798 -1181 -2764
rect -3230 -2848 -3134 -2814
rect -2104 -2848 -2008 -2814
rect -1239 -2815 -1181 -2798
rect -1100 -2716 -1054 -2670
rect -1100 -2750 -1088 -2716
rect -1100 -2784 -1054 -2750
rect -1100 -2818 -1088 -2784
rect -1100 -2834 -1054 -2818
rect -1020 -2716 -954 -2704
rect -1020 -2750 -1004 -2716
rect -970 -2750 -954 -2716
rect -1020 -2784 -954 -2750
rect -1020 -2818 -1004 -2784
rect -970 -2818 -954 -2784
rect -687 -2764 -629 -2670
rect -687 -2798 -675 -2764
rect -641 -2798 -629 -2764
rect -687 -2815 -629 -2798
rect -595 -2712 -533 -2670
rect -595 -2746 -573 -2712
rect -539 -2746 -533 -2712
rect -595 -2780 -533 -2746
rect -595 -2814 -573 -2780
rect -539 -2814 -533 -2780
rect -1020 -2830 -954 -2818
rect -595 -2830 -533 -2814
rect -492 -2712 -353 -2704
rect -492 -2746 -405 -2712
rect -371 -2746 -353 -2712
rect -492 -2780 -353 -2746
rect -492 -2814 -405 -2780
rect -371 -2814 -353 -2780
rect -492 -2830 -353 -2814
rect -3230 -2910 -3196 -2848
rect -2042 -2910 -2008 -2848
rect -3132 -2950 -3116 -2916
rect -3082 -2950 -3066 -2916
rect -2940 -2950 -2924 -2916
rect -2890 -2950 -2874 -2916
rect -2748 -2950 -2732 -2916
rect -2698 -2950 -2682 -2916
rect -2556 -2950 -2540 -2916
rect -2506 -2950 -2490 -2916
rect -2364 -2950 -2348 -2916
rect -2314 -2950 -2298 -2916
rect -2172 -2950 -2156 -2916
rect -2122 -2950 -2106 -2916
rect -3116 -3010 -3082 -2994
rect -3116 -3274 -3082 -3258
rect -3020 -3010 -2986 -2994
rect -3020 -3274 -2986 -3258
rect -2924 -3010 -2890 -2994
rect -2924 -3274 -2890 -3258
rect -2828 -3010 -2794 -2994
rect -2828 -3274 -2794 -3258
rect -2732 -3010 -2698 -2994
rect -2732 -3274 -2698 -3258
rect -2636 -3010 -2602 -2994
rect -2636 -3274 -2602 -3258
rect -2540 -3010 -2506 -2994
rect -2540 -3274 -2506 -3258
rect -2444 -3010 -2410 -2994
rect -2444 -3274 -2410 -3258
rect -2348 -3010 -2314 -2994
rect -2348 -3274 -2314 -3258
rect -2252 -3010 -2218 -2994
rect -2252 -3274 -2218 -3258
rect -2156 -3010 -2122 -2994
rect -2156 -3274 -2122 -3258
rect -3230 -3358 -3196 -3296
rect -1100 -2874 -1084 -2868
rect -1100 -2908 -1089 -2874
rect -1050 -2902 -1034 -2868
rect -1055 -2908 -1034 -2902
rect -1100 -2916 -1034 -2908
rect -1000 -2874 -954 -2830
rect -1000 -2908 -994 -2874
rect -960 -2908 -954 -2874
rect -1239 -2982 -1181 -2947
rect -1000 -2950 -954 -2908
rect -593 -2868 -526 -2864
rect -593 -2902 -576 -2868
rect -542 -2874 -526 -2868
rect -593 -2908 -574 -2902
rect -540 -2908 -526 -2874
rect -593 -2918 -526 -2908
rect -1239 -3016 -1227 -2982
rect -1193 -3016 -1181 -2982
rect -1239 -3075 -1181 -3016
rect -1239 -3109 -1227 -3075
rect -1193 -3109 -1181 -3075
rect -1239 -3180 -1181 -3109
rect -1096 -2968 -1054 -2952
rect -1096 -3002 -1088 -2968
rect -1096 -3036 -1054 -3002
rect -1096 -3070 -1088 -3036
rect -1096 -3104 -1054 -3070
rect -1096 -3138 -1088 -3104
rect -1096 -3180 -1054 -3138
rect -1020 -2968 -954 -2950
rect -1020 -3002 -1004 -2968
rect -970 -3002 -954 -2968
rect -1020 -3036 -954 -3002
rect -1020 -3070 -1004 -3036
rect -970 -3070 -954 -3036
rect -1020 -3104 -954 -3070
rect -1020 -3138 -1004 -3104
rect -970 -3138 -954 -3104
rect -1020 -3146 -954 -3138
rect -687 -2982 -629 -2947
rect -492 -2950 -458 -2830
rect 321 -2848 417 -2814
rect 1447 -2848 1543 -2814
rect -424 -2902 -408 -2868
rect -374 -2875 -357 -2868
rect -424 -2909 -401 -2902
rect -367 -2909 -357 -2875
rect -424 -2918 -357 -2909
rect 321 -2910 355 -2848
rect -687 -3016 -675 -2982
rect -641 -3016 -629 -2982
rect -687 -3075 -629 -3016
rect -687 -3109 -675 -3075
rect -641 -3109 -629 -3075
rect -687 -3180 -629 -3109
rect -595 -2968 -539 -2952
rect -595 -3002 -573 -2968
rect -595 -3036 -539 -3002
rect -595 -3070 -573 -3036
rect -595 -3104 -539 -3070
rect -595 -3138 -573 -3104
rect -595 -3180 -539 -3138
rect -505 -2968 -439 -2950
rect -505 -3002 -489 -2968
rect -455 -3002 -439 -2968
rect -505 -3036 -439 -3002
rect -505 -3070 -490 -3036
rect -455 -3070 -439 -3036
rect -505 -3104 -439 -3070
rect -505 -3138 -489 -3104
rect -455 -3138 -439 -3104
rect -505 -3146 -439 -3138
rect -405 -2968 -353 -2952
rect -371 -3002 -353 -2968
rect -405 -3036 -353 -3002
rect -371 -3070 -353 -3036
rect -405 -3104 -353 -3070
rect -371 -3138 -353 -3104
rect -405 -3180 -353 -3138
rect 1509 -2910 1543 -2848
rect 419 -2946 435 -2912
rect 469 -2946 485 -2912
rect 611 -2946 627 -2912
rect 661 -2946 677 -2912
rect 803 -2946 819 -2912
rect 853 -2946 869 -2912
rect 995 -2946 1011 -2912
rect 1045 -2946 1061 -2912
rect 1187 -2946 1203 -2912
rect 1237 -2946 1253 -2912
rect 1379 -2946 1395 -2912
rect 1429 -2946 1445 -2912
rect 435 -3000 469 -2984
rect 435 -3096 469 -3080
rect 531 -3000 565 -2984
rect 531 -3096 565 -3080
rect 627 -3000 661 -2984
rect 627 -3096 661 -3080
rect 723 -3000 757 -2984
rect 723 -3096 757 -3080
rect 819 -3000 853 -2984
rect 819 -3096 853 -3080
rect 915 -3000 949 -2984
rect 915 -3096 949 -3080
rect 1011 -3000 1045 -2984
rect 1011 -3096 1045 -3080
rect 1107 -3000 1141 -2984
rect 1107 -3096 1141 -3080
rect 1203 -3000 1237 -2984
rect 1203 -3096 1237 -3080
rect 1299 -3000 1333 -2984
rect 1299 -3096 1333 -3080
rect 1395 -3000 1429 -2984
rect 1395 -3096 1429 -3080
rect 321 -3170 355 -3108
rect 1842 -2848 1938 -2814
rect 2968 -2848 3064 -2814
rect 1842 -2910 1876 -2848
rect 1616 -3008 1650 -2992
rect 1616 -3100 1650 -3084
rect 1704 -3008 1738 -2992
rect 1704 -3100 1738 -3084
rect 1509 -3170 1543 -3110
rect 3030 -2910 3064 -2848
rect 1940 -2946 1956 -2912
rect 1990 -2946 2006 -2912
rect 2132 -2946 2148 -2912
rect 2182 -2946 2198 -2912
rect 2324 -2946 2340 -2912
rect 2374 -2946 2390 -2912
rect 2516 -2946 2532 -2912
rect 2566 -2946 2582 -2912
rect 2708 -2946 2724 -2912
rect 2758 -2946 2774 -2912
rect 2900 -2946 2916 -2912
rect 2950 -2946 2966 -2912
rect 1956 -3000 1990 -2984
rect 1956 -3096 1990 -3080
rect 2052 -3000 2086 -2984
rect 2052 -3096 2086 -3080
rect 2148 -3000 2182 -2984
rect 2148 -3096 2182 -3080
rect 2244 -3000 2278 -2984
rect 2244 -3096 2278 -3080
rect 2340 -3000 2374 -2984
rect 2340 -3096 2374 -3080
rect 2436 -3000 2470 -2984
rect 2436 -3096 2470 -3080
rect 2532 -3000 2566 -2984
rect 2532 -3096 2566 -3080
rect 2628 -3000 2662 -2984
rect 2628 -3096 2662 -3080
rect 2724 -3000 2758 -2984
rect 2724 -3096 2758 -3080
rect 2820 -3000 2854 -2984
rect 2820 -3096 2854 -3080
rect 2916 -3000 2950 -2984
rect 2916 -3096 2950 -3080
rect 1644 -3168 1660 -3134
rect 1694 -3168 1710 -3134
rect -1256 -3214 -1227 -3180
rect -1193 -3214 -1135 -3180
rect -1101 -3214 -1043 -3180
rect -1009 -3214 -951 -3180
rect -917 -3214 -859 -3180
rect -825 -3214 -767 -3180
rect -733 -3214 -675 -3180
rect -641 -3214 -583 -3180
rect -549 -3214 -491 -3180
rect -457 -3214 -399 -3180
rect -365 -3214 -336 -3180
rect 321 -3204 417 -3170
rect 1447 -3204 1543 -3170
rect 1842 -3170 1876 -3108
rect 3030 -3170 3064 -3110
rect 1842 -3204 1938 -3170
rect 2968 -3204 3064 -3170
rect -2042 -3358 -2008 -3296
rect -3230 -3392 -3134 -3358
rect -2104 -3392 -2008 -3358
rect -687 -3285 -629 -3214
rect -687 -3319 -675 -3285
rect -641 -3319 -629 -3285
rect -687 -3378 -629 -3319
rect -687 -3412 -675 -3378
rect -641 -3412 -629 -3378
rect -687 -3447 -629 -3412
rect -595 -3256 -539 -3214
rect -595 -3290 -573 -3256
rect -595 -3324 -539 -3290
rect -595 -3358 -573 -3324
rect -595 -3392 -539 -3358
rect -595 -3426 -573 -3392
rect -595 -3442 -539 -3426
rect -505 -3256 -439 -3248
rect -505 -3290 -489 -3256
rect -455 -3290 -439 -3256
rect -505 -3324 -439 -3290
rect -505 -3358 -489 -3324
rect -455 -3358 -439 -3324
rect -505 -3392 -439 -3358
rect -505 -3426 -489 -3392
rect -455 -3426 -439 -3392
rect -505 -3444 -439 -3426
rect -405 -3256 -353 -3214
rect -371 -3290 -353 -3256
rect -405 -3324 -353 -3290
rect -371 -3358 -353 -3324
rect -405 -3392 -353 -3358
rect -371 -3426 -353 -3392
rect -405 -3442 -353 -3426
rect 321 -3312 417 -3278
rect 1447 -3312 1543 -3278
rect 321 -3374 355 -3312
rect -3230 -3500 -3134 -3466
rect -2104 -3500 -2008 -3466
rect -3230 -3562 -3196 -3500
rect -2042 -3560 -2008 -3500
rect -593 -3492 -526 -3476
rect -593 -3526 -576 -3492
rect -542 -3526 -526 -3492
rect -593 -3530 -526 -3526
rect -3116 -3590 -3082 -3574
rect -3116 -3686 -3082 -3670
rect -3020 -3590 -2986 -3574
rect -3020 -3686 -2986 -3670
rect -2924 -3590 -2890 -3574
rect -2924 -3686 -2890 -3670
rect -2828 -3590 -2794 -3574
rect -2828 -3686 -2794 -3670
rect -2732 -3590 -2698 -3574
rect -2732 -3686 -2698 -3670
rect -2636 -3590 -2602 -3574
rect -2636 -3686 -2602 -3670
rect -2540 -3590 -2506 -3574
rect -2540 -3686 -2506 -3670
rect -2444 -3590 -2410 -3574
rect -2444 -3686 -2410 -3670
rect -2348 -3590 -2314 -3574
rect -2348 -3686 -2314 -3670
rect -2252 -3590 -2218 -3574
rect -2252 -3686 -2218 -3670
rect -2156 -3590 -2122 -3574
rect -2156 -3686 -2122 -3670
rect -3132 -3758 -3116 -3724
rect -3082 -3758 -3066 -3724
rect -2940 -3758 -2924 -3724
rect -2890 -3758 -2874 -3724
rect -2748 -3758 -2732 -3724
rect -2698 -3758 -2682 -3724
rect -2556 -3758 -2540 -3724
rect -2506 -3758 -2490 -3724
rect -2364 -3758 -2348 -3724
rect -2314 -3758 -2298 -3724
rect -2172 -3758 -2156 -3724
rect -2122 -3758 -2106 -3724
rect -3230 -3822 -3196 -3760
rect -492 -3564 -458 -3444
rect -424 -3487 -357 -3476
rect -424 -3492 -405 -3487
rect -424 -3526 -408 -3492
rect -371 -3521 -357 -3487
rect -374 -3526 -357 -3521
rect -687 -3596 -629 -3579
rect -687 -3630 -675 -3596
rect -641 -3630 -629 -3596
rect -687 -3724 -629 -3630
rect -595 -3580 -533 -3564
rect -595 -3614 -573 -3580
rect -539 -3614 -533 -3580
rect -595 -3648 -533 -3614
rect -595 -3682 -573 -3648
rect -539 -3682 -533 -3648
rect -595 -3724 -533 -3682
rect -492 -3580 -353 -3564
rect -492 -3590 -405 -3580
rect -458 -3614 -405 -3590
rect -371 -3614 -353 -3580
rect -458 -3624 -353 -3614
rect -492 -3648 -353 -3624
rect -492 -3682 -405 -3648
rect -371 -3682 -353 -3648
rect -492 -3690 -353 -3682
rect -704 -3758 -675 -3724
rect -641 -3758 -583 -3724
rect -549 -3758 -491 -3724
rect -457 -3758 -399 -3724
rect -365 -3758 -336 -3724
rect -2042 -3822 -2008 -3760
rect -3230 -3856 -3134 -3822
rect -2104 -3856 -2008 -3822
rect -687 -3852 -629 -3758
rect -687 -3886 -675 -3852
rect -641 -3886 -629 -3852
rect -687 -3903 -629 -3886
rect -548 -3804 -502 -3758
rect 1509 -3374 1543 -3312
rect 435 -3412 469 -3396
rect 435 -3676 469 -3660
rect 531 -3412 565 -3396
rect 531 -3676 565 -3660
rect 627 -3412 661 -3396
rect 627 -3676 661 -3660
rect 723 -3412 757 -3396
rect 723 -3676 757 -3660
rect 819 -3412 853 -3396
rect 819 -3676 853 -3660
rect 915 -3412 949 -3396
rect 915 -3676 949 -3660
rect 1011 -3412 1045 -3396
rect 1011 -3676 1045 -3660
rect 1107 -3412 1141 -3396
rect 1107 -3676 1141 -3660
rect 1203 -3412 1237 -3396
rect 1203 -3676 1237 -3660
rect 1299 -3412 1333 -3396
rect 1299 -3676 1333 -3660
rect 1395 -3412 1429 -3396
rect 1395 -3676 1429 -3660
rect 419 -3754 435 -3720
rect 469 -3754 485 -3720
rect 611 -3754 627 -3720
rect 661 -3754 677 -3720
rect 803 -3754 819 -3720
rect 853 -3754 869 -3720
rect 995 -3754 1011 -3720
rect 1045 -3754 1061 -3720
rect 1187 -3754 1203 -3720
rect 1237 -3754 1253 -3720
rect 1379 -3754 1395 -3720
rect 1429 -3754 1445 -3720
rect -548 -3838 -536 -3804
rect -548 -3872 -502 -3838
rect -548 -3906 -536 -3872
rect -548 -3922 -502 -3906
rect -468 -3804 -402 -3792
rect -468 -3838 -452 -3804
rect -418 -3838 -402 -3804
rect -468 -3872 -402 -3838
rect 321 -3822 355 -3760
rect 1509 -3822 1543 -3760
rect 321 -3856 417 -3822
rect 1447 -3856 1543 -3822
rect 1842 -3312 1938 -3278
rect 2968 -3312 3064 -3278
rect 1842 -3374 1876 -3312
rect 3030 -3374 3064 -3312
rect 1956 -3412 1990 -3396
rect 1956 -3676 1990 -3660
rect 2052 -3412 2086 -3396
rect 2052 -3676 2086 -3660
rect 2148 -3412 2182 -3396
rect 2148 -3676 2182 -3660
rect 2244 -3412 2278 -3396
rect 2244 -3676 2278 -3660
rect 2340 -3412 2374 -3396
rect 2340 -3676 2374 -3660
rect 2436 -3412 2470 -3396
rect 2436 -3676 2470 -3660
rect 2532 -3412 2566 -3396
rect 2532 -3676 2566 -3660
rect 2628 -3412 2662 -3396
rect 2628 -3676 2662 -3660
rect 2724 -3412 2758 -3396
rect 2724 -3676 2758 -3660
rect 2820 -3412 2854 -3396
rect 2820 -3676 2854 -3660
rect 2916 -3412 2950 -3396
rect 2916 -3676 2950 -3660
rect 1940 -3754 1956 -3720
rect 1990 -3754 2006 -3720
rect 2132 -3754 2148 -3720
rect 2182 -3754 2198 -3720
rect 2324 -3754 2340 -3720
rect 2374 -3754 2390 -3720
rect 2516 -3754 2532 -3720
rect 2566 -3754 2582 -3720
rect 2708 -3754 2724 -3720
rect 2758 -3754 2774 -3720
rect 2900 -3754 2916 -3720
rect 2950 -3754 2966 -3720
rect 1842 -3822 1876 -3760
rect 3030 -3822 3064 -3760
rect 1842 -3856 1938 -3822
rect 2968 -3856 3064 -3822
rect -468 -3906 -452 -3872
rect -418 -3906 -402 -3872
rect -468 -3918 -402 -3906
rect -548 -3961 -532 -3956
rect -548 -3995 -539 -3961
rect -498 -3990 -482 -3956
rect -505 -3995 -482 -3990
rect -548 -4004 -482 -3995
rect -687 -4070 -629 -4035
rect -448 -4038 -402 -3918
rect -687 -4104 -675 -4070
rect -641 -4104 -629 -4070
rect -687 -4163 -629 -4104
rect -3230 -4226 -3134 -4192
rect -2104 -4226 -2008 -4192
rect -3230 -4288 -3196 -4226
rect -2042 -4288 -2008 -4226
rect -687 -4197 -675 -4163
rect -641 -4197 -629 -4163
rect -687 -4268 -629 -4197
rect -544 -4056 -502 -4040
rect -544 -4090 -536 -4056
rect -544 -4124 -502 -4090
rect -544 -4158 -536 -4124
rect -544 -4192 -502 -4158
rect -544 -4226 -536 -4192
rect -544 -4268 -502 -4226
rect -468 -4056 -402 -4038
rect -468 -4090 -452 -4056
rect -418 -4090 -402 -4056
rect -468 -4120 -402 -4090
rect -468 -4154 -453 -4120
rect -419 -4124 -402 -4120
rect -468 -4158 -452 -4154
rect -418 -4158 -402 -4124
rect -468 -4192 -402 -4158
rect -468 -4226 -452 -4192
rect -418 -4226 -402 -4192
rect -468 -4234 -402 -4226
rect 321 -4226 417 -4192
rect 1447 -4226 1543 -4192
rect -3132 -4328 -3116 -4294
rect -3082 -4328 -3066 -4294
rect -2940 -4328 -2924 -4294
rect -2890 -4328 -2874 -4294
rect -2748 -4328 -2732 -4294
rect -2698 -4328 -2682 -4294
rect -2556 -4328 -2540 -4294
rect -2506 -4328 -2490 -4294
rect -2364 -4328 -2348 -4294
rect -2314 -4328 -2298 -4294
rect -2172 -4328 -2156 -4294
rect -2122 -4328 -2106 -4294
rect -3116 -4388 -3082 -4372
rect -3116 -4652 -3082 -4636
rect -3020 -4388 -2986 -4372
rect -3020 -4652 -2986 -4636
rect -2924 -4388 -2890 -4372
rect -2924 -4652 -2890 -4636
rect -2828 -4388 -2794 -4372
rect -2828 -4652 -2794 -4636
rect -2732 -4388 -2698 -4372
rect -2732 -4652 -2698 -4636
rect -2636 -4388 -2602 -4372
rect -2636 -4652 -2602 -4636
rect -2540 -4388 -2506 -4372
rect -2540 -4652 -2506 -4636
rect -2444 -4388 -2410 -4372
rect -2444 -4652 -2410 -4636
rect -2348 -4388 -2314 -4372
rect -2348 -4652 -2314 -4636
rect -2252 -4388 -2218 -4372
rect -2252 -4652 -2218 -4636
rect -2156 -4388 -2122 -4372
rect -2156 -4652 -2122 -4636
rect -3230 -4736 -3196 -4674
rect -704 -4302 -675 -4268
rect -641 -4302 -583 -4268
rect -549 -4302 -491 -4268
rect -457 -4302 -399 -4268
rect -365 -4302 -336 -4268
rect 321 -4288 355 -4226
rect -687 -4373 -629 -4302
rect -687 -4407 -675 -4373
rect -641 -4407 -629 -4373
rect -687 -4466 -629 -4407
rect -687 -4500 -675 -4466
rect -641 -4500 -629 -4466
rect -687 -4535 -629 -4500
rect -544 -4344 -502 -4302
rect -544 -4378 -536 -4344
rect -544 -4412 -502 -4378
rect -544 -4446 -536 -4412
rect -544 -4480 -502 -4446
rect -544 -4514 -536 -4480
rect -544 -4530 -502 -4514
rect -468 -4344 -402 -4336
rect -468 -4378 -452 -4344
rect -418 -4378 -402 -4344
rect -468 -4412 -402 -4378
rect -468 -4452 -452 -4412
rect -418 -4452 -402 -4412
rect -468 -4480 -402 -4452
rect -468 -4514 -452 -4480
rect -418 -4514 -402 -4480
rect -468 -4532 -402 -4514
rect -548 -4574 -482 -4566
rect -548 -4608 -540 -4574
rect -506 -4580 -482 -4574
rect -548 -4614 -532 -4608
rect -498 -4614 -482 -4580
rect -548 -4664 -502 -4648
rect -448 -4652 -402 -4532
rect 1509 -4288 1543 -4226
rect 419 -4324 435 -4290
rect 469 -4324 485 -4290
rect 611 -4324 627 -4290
rect 661 -4324 677 -4290
rect 803 -4324 819 -4290
rect 853 -4324 869 -4290
rect 995 -4324 1011 -4290
rect 1045 -4324 1061 -4290
rect 1187 -4324 1203 -4290
rect 1237 -4324 1253 -4290
rect 1379 -4324 1395 -4290
rect 1429 -4324 1445 -4290
rect 435 -4378 469 -4362
rect 435 -4474 469 -4458
rect 531 -4378 565 -4362
rect 531 -4474 565 -4458
rect 627 -4378 661 -4362
rect 627 -4474 661 -4458
rect 723 -4378 757 -4362
rect 723 -4474 757 -4458
rect 819 -4378 853 -4362
rect 819 -4474 853 -4458
rect 915 -4378 949 -4362
rect 915 -4474 949 -4458
rect 1011 -4378 1045 -4362
rect 1011 -4474 1045 -4458
rect 1107 -4378 1141 -4362
rect 1107 -4474 1141 -4458
rect 1203 -4378 1237 -4362
rect 1203 -4474 1237 -4458
rect 1299 -4378 1333 -4362
rect 1299 -4474 1333 -4458
rect 1395 -4378 1429 -4362
rect 1395 -4474 1429 -4458
rect 321 -4548 355 -4486
rect 1842 -4226 1938 -4192
rect 2968 -4226 3064 -4192
rect 1842 -4288 1876 -4226
rect 1616 -4386 1650 -4370
rect 1616 -4478 1650 -4462
rect 1704 -4386 1738 -4370
rect 1704 -4478 1738 -4462
rect 1509 -4548 1543 -4488
rect 3030 -4288 3064 -4226
rect 1940 -4324 1956 -4290
rect 1990 -4324 2006 -4290
rect 2132 -4324 2148 -4290
rect 2182 -4324 2198 -4290
rect 2324 -4324 2340 -4290
rect 2374 -4324 2390 -4290
rect 2516 -4324 2532 -4290
rect 2566 -4324 2582 -4290
rect 2708 -4324 2724 -4290
rect 2758 -4324 2774 -4290
rect 2900 -4324 2916 -4290
rect 2950 -4324 2966 -4290
rect 1956 -4378 1990 -4362
rect 1956 -4474 1990 -4458
rect 2052 -4378 2086 -4362
rect 2052 -4474 2086 -4458
rect 2148 -4378 2182 -4362
rect 2148 -4474 2182 -4458
rect 2244 -4378 2278 -4362
rect 2244 -4474 2278 -4458
rect 2340 -4378 2374 -4362
rect 2340 -4474 2374 -4458
rect 2436 -4378 2470 -4362
rect 2436 -4474 2470 -4458
rect 2532 -4378 2566 -4362
rect 2532 -4474 2566 -4458
rect 2628 -4378 2662 -4362
rect 2628 -4474 2662 -4458
rect 2724 -4378 2758 -4362
rect 2724 -4474 2758 -4458
rect 2820 -4378 2854 -4362
rect 2820 -4474 2854 -4458
rect 2916 -4378 2950 -4362
rect 2916 -4474 2950 -4458
rect 1644 -4546 1660 -4512
rect 1694 -4546 1710 -4512
rect 321 -4582 417 -4548
rect 1447 -4582 1543 -4548
rect 1842 -4548 1876 -4486
rect 3030 -4548 3064 -4488
rect 1842 -4582 1938 -4548
rect 2968 -4582 3064 -4548
rect -2042 -4736 -2008 -4674
rect -3230 -4770 -3134 -4736
rect -2104 -4770 -2008 -4736
rect -687 -4684 -629 -4667
rect -687 -4718 -675 -4684
rect -641 -4718 -629 -4684
rect -687 -4812 -629 -4718
rect -548 -4698 -536 -4664
rect -548 -4732 -502 -4698
rect -548 -4766 -536 -4732
rect -548 -4812 -502 -4766
rect -468 -4664 -402 -4652
rect -468 -4698 -452 -4664
rect -418 -4698 -402 -4664
rect -468 -4732 -402 -4698
rect -468 -4766 -452 -4732
rect -418 -4766 -402 -4732
rect -468 -4778 -402 -4766
rect 321 -4690 417 -4656
rect 1447 -4690 1543 -4656
rect 321 -4752 355 -4690
rect -3230 -4878 -3134 -4844
rect -2104 -4878 -2008 -4844
rect -704 -4846 -675 -4812
rect -641 -4846 -583 -4812
rect -549 -4846 -491 -4812
rect -457 -4846 -399 -4812
rect -365 -4846 -336 -4812
rect -3230 -4940 -3196 -4878
rect -2042 -4938 -2008 -4878
rect -3116 -4968 -3082 -4952
rect -3116 -5064 -3082 -5048
rect -3020 -4968 -2986 -4952
rect -3020 -5064 -2986 -5048
rect -2924 -4968 -2890 -4952
rect -2924 -5064 -2890 -5048
rect -2828 -4968 -2794 -4952
rect -2828 -5064 -2794 -5048
rect -2732 -4968 -2698 -4952
rect -2732 -5064 -2698 -5048
rect -2636 -4968 -2602 -4952
rect -2636 -5064 -2602 -5048
rect -2540 -4968 -2506 -4952
rect -2540 -5064 -2506 -5048
rect -2444 -4968 -2410 -4952
rect -2444 -5064 -2410 -5048
rect -2348 -4968 -2314 -4952
rect -2348 -5064 -2314 -5048
rect -2252 -4968 -2218 -4952
rect -2252 -5064 -2218 -5048
rect -2156 -4968 -2122 -4952
rect -2156 -5064 -2122 -5048
rect -3132 -5136 -3116 -5102
rect -3082 -5136 -3066 -5102
rect -2940 -5136 -2924 -5102
rect -2890 -5136 -2874 -5102
rect -2748 -5136 -2732 -5102
rect -2698 -5136 -2682 -5102
rect -2556 -5136 -2540 -5102
rect -2506 -5136 -2490 -5102
rect -2364 -5136 -2348 -5102
rect -2314 -5136 -2298 -5102
rect -2172 -5136 -2156 -5102
rect -2122 -5136 -2106 -5102
rect -3230 -5200 -3196 -5138
rect -2042 -5200 -2008 -5138
rect -3230 -5234 -3134 -5200
rect -2104 -5234 -2008 -5200
rect 1509 -4752 1543 -4690
rect 435 -4790 469 -4774
rect 435 -5054 469 -5038
rect 531 -4790 565 -4774
rect 531 -5054 565 -5038
rect 627 -4790 661 -4774
rect 627 -5054 661 -5038
rect 723 -4790 757 -4774
rect 723 -5054 757 -5038
rect 819 -4790 853 -4774
rect 819 -5054 853 -5038
rect 915 -4790 949 -4774
rect 915 -5054 949 -5038
rect 1011 -4790 1045 -4774
rect 1011 -5054 1045 -5038
rect 1107 -4790 1141 -4774
rect 1107 -5054 1141 -5038
rect 1203 -4790 1237 -4774
rect 1203 -5054 1237 -5038
rect 1299 -4790 1333 -4774
rect 1299 -5054 1333 -5038
rect 1395 -4790 1429 -4774
rect 1395 -5054 1429 -5038
rect 419 -5132 435 -5098
rect 469 -5132 485 -5098
rect 611 -5132 627 -5098
rect 661 -5132 677 -5098
rect 803 -5132 819 -5098
rect 853 -5132 869 -5098
rect 995 -5132 1011 -5098
rect 1045 -5132 1061 -5098
rect 1187 -5132 1203 -5098
rect 1237 -5132 1253 -5098
rect 1379 -5132 1395 -5098
rect 1429 -5132 1445 -5098
rect 321 -5200 355 -5138
rect 1509 -5200 1543 -5138
rect 321 -5234 417 -5200
rect 1447 -5234 1543 -5200
rect 1842 -4690 1938 -4656
rect 2968 -4690 3064 -4656
rect 1842 -4752 1876 -4690
rect 3030 -4752 3064 -4690
rect 1956 -4790 1990 -4774
rect 1956 -5054 1990 -5038
rect 2052 -4790 2086 -4774
rect 2052 -5054 2086 -5038
rect 2148 -4790 2182 -4774
rect 2148 -5054 2182 -5038
rect 2244 -4790 2278 -4774
rect 2244 -5054 2278 -5038
rect 2340 -4790 2374 -4774
rect 2340 -5054 2374 -5038
rect 2436 -4790 2470 -4774
rect 2436 -5054 2470 -5038
rect 2532 -4790 2566 -4774
rect 2532 -5054 2566 -5038
rect 2628 -4790 2662 -4774
rect 2628 -5054 2662 -5038
rect 2724 -4790 2758 -4774
rect 2724 -5054 2758 -5038
rect 2820 -4790 2854 -4774
rect 2820 -5054 2854 -5038
rect 2916 -4790 2950 -4774
rect 2916 -5054 2950 -5038
rect 1940 -5132 1956 -5098
rect 1990 -5132 2006 -5098
rect 2132 -5132 2148 -5098
rect 2182 -5132 2198 -5098
rect 2324 -5132 2340 -5098
rect 2374 -5132 2390 -5098
rect 2516 -5132 2532 -5098
rect 2566 -5132 2582 -5098
rect 2708 -5132 2724 -5098
rect 2758 -5132 2774 -5098
rect 2900 -5132 2916 -5098
rect 2950 -5132 2966 -5098
rect 1842 -5200 1876 -5138
rect 3030 -5200 3064 -5138
rect 1842 -5234 1938 -5200
rect 2968 -5234 3064 -5200
<< viali >>
rect -3116 -238 -3082 -204
rect -2924 -238 -2890 -204
rect -2732 -238 -2698 -204
rect -2540 -238 -2506 -204
rect -2348 -238 -2314 -204
rect -2156 -238 -2122 -204
rect -3116 -546 -3082 -298
rect -3020 -546 -2986 -298
rect -2924 -546 -2890 -298
rect -2828 -546 -2794 -298
rect -2732 -546 -2698 -298
rect -2636 -546 -2602 -298
rect -2540 -546 -2506 -298
rect -2444 -546 -2410 -298
rect -2348 -546 -2314 -298
rect -2252 -546 -2218 -298
rect -2156 -546 -2122 -298
rect -2042 -584 -2008 -198
rect 435 -234 469 -200
rect 627 -234 661 -200
rect 819 -234 853 -200
rect 1011 -234 1045 -200
rect 1203 -234 1237 -200
rect 1395 -234 1429 -200
rect 435 -368 469 -288
rect 531 -368 565 -288
rect 627 -368 661 -288
rect 723 -368 757 -288
rect 819 -368 853 -288
rect 915 -368 949 -288
rect 1011 -368 1045 -288
rect 1107 -368 1141 -288
rect 1203 -368 1237 -288
rect 1299 -368 1333 -288
rect 1395 -368 1429 -288
rect 1509 -396 1543 -198
rect 1616 -372 1650 -296
rect 1704 -372 1738 -296
rect 1509 -398 1543 -396
rect 1956 -234 1990 -200
rect 2148 -234 2182 -200
rect 2340 -234 2374 -200
rect 2532 -234 2566 -200
rect 2724 -234 2758 -200
rect 2916 -234 2950 -200
rect 1956 -368 1990 -288
rect 2052 -368 2086 -288
rect 2148 -368 2182 -288
rect 2244 -368 2278 -288
rect 2340 -368 2374 -288
rect 2436 -368 2470 -288
rect 2532 -368 2566 -288
rect 2628 -368 2662 -288
rect 2724 -368 2758 -288
rect 2820 -368 2854 -288
rect 2916 -368 2950 -288
rect 1660 -456 1694 -422
rect -951 -494 -917 -460
rect -859 -494 -825 -460
rect -767 -494 -733 -460
rect -675 -494 -641 -460
rect -583 -494 -549 -460
rect -491 -494 -457 -460
rect -399 -494 -365 -460
rect 3030 -396 3064 -198
rect 3030 -398 3064 -396
rect -822 -608 -788 -603
rect -822 -637 -820 -608
rect -820 -637 -788 -608
rect -905 -726 -900 -698
rect -900 -726 -871 -698
rect -905 -732 -871 -726
rect -452 -608 -418 -594
rect -452 -628 -418 -608
rect -538 -726 -532 -700
rect -532 -726 -504 -700
rect -538 -734 -504 -726
rect -2042 -850 -2008 -848
rect -3116 -958 -3082 -878
rect -3020 -958 -2986 -878
rect -2924 -958 -2890 -878
rect -2828 -958 -2794 -878
rect -2732 -958 -2698 -878
rect -2636 -958 -2602 -878
rect -2540 -958 -2506 -878
rect -2444 -958 -2410 -878
rect -2348 -958 -2314 -878
rect -2252 -958 -2218 -878
rect -2156 -958 -2122 -878
rect -3116 -1046 -3082 -1012
rect -2924 -1046 -2890 -1012
rect -2732 -1046 -2698 -1012
rect -2540 -1046 -2506 -1012
rect -2348 -1046 -2314 -1012
rect -2156 -1046 -2122 -1012
rect -2042 -1048 -2008 -850
rect -951 -1038 -917 -1004
rect -859 -1038 -825 -1004
rect -767 -1038 -733 -1004
rect -675 -1038 -641 -1004
rect -583 -1038 -549 -1004
rect -491 -1038 -457 -1004
rect -399 -1038 -365 -1004
rect 435 -948 469 -700
rect 531 -948 565 -700
rect 627 -948 661 -700
rect 723 -948 757 -700
rect 819 -948 853 -700
rect 915 -948 949 -700
rect 1011 -948 1045 -700
rect 1107 -948 1141 -700
rect 1203 -948 1237 -700
rect 1299 -948 1333 -700
rect 1395 -948 1429 -700
rect 435 -1042 469 -1008
rect 627 -1042 661 -1008
rect 819 -1042 853 -1008
rect 1011 -1042 1045 -1008
rect 1203 -1042 1237 -1008
rect 1395 -1042 1429 -1008
rect 1509 -1048 1543 -662
rect 1956 -948 1990 -700
rect 2052 -948 2086 -700
rect 2148 -948 2182 -700
rect 2244 -948 2278 -700
rect 2340 -948 2374 -700
rect 2436 -948 2470 -700
rect 2532 -948 2566 -700
rect 2628 -948 2662 -700
rect 2724 -948 2758 -700
rect 2820 -948 2854 -700
rect 2916 -948 2950 -700
rect 1956 -1042 1990 -1008
rect 2148 -1042 2182 -1008
rect 2340 -1042 2374 -1008
rect 2532 -1042 2566 -1008
rect 2724 -1042 2758 -1008
rect 2916 -1042 2950 -1008
rect 3030 -1048 3064 -662
rect -453 -1216 -419 -1197
rect -453 -1231 -452 -1216
rect -452 -1231 -419 -1216
rect -534 -1316 -500 -1312
rect -534 -1346 -532 -1316
rect -532 -1346 -500 -1316
rect -3116 -1572 -3082 -1538
rect -2924 -1572 -2890 -1538
rect -2732 -1572 -2698 -1538
rect -2540 -1572 -2506 -1538
rect -2348 -1572 -2314 -1538
rect -2156 -1572 -2122 -1538
rect -3116 -1880 -3082 -1632
rect -3020 -1880 -2986 -1632
rect -2924 -1880 -2890 -1632
rect -2828 -1880 -2794 -1632
rect -2732 -1880 -2698 -1632
rect -2636 -1880 -2602 -1632
rect -2540 -1880 -2506 -1632
rect -2444 -1880 -2410 -1632
rect -2348 -1880 -2314 -1632
rect -2252 -1880 -2218 -1632
rect -2156 -1880 -2122 -1632
rect -2042 -1918 -2008 -1532
rect -675 -1582 -641 -1548
rect -583 -1582 -549 -1548
rect -491 -1582 -457 -1548
rect -399 -1582 -365 -1548
rect -469 -1710 -435 -1676
rect 435 -1568 469 -1534
rect 627 -1568 661 -1534
rect 819 -1568 853 -1534
rect 1011 -1568 1045 -1534
rect 1203 -1568 1237 -1534
rect 1395 -1568 1429 -1534
rect 435 -1702 469 -1622
rect 531 -1702 565 -1622
rect 627 -1702 661 -1622
rect 723 -1702 757 -1622
rect 819 -1702 853 -1622
rect 915 -1702 949 -1622
rect 1011 -1702 1045 -1622
rect 1107 -1702 1141 -1622
rect 1203 -1702 1237 -1622
rect 1299 -1702 1333 -1622
rect 1395 -1702 1429 -1622
rect -582 -1814 -576 -1784
rect -576 -1814 -548 -1784
rect -582 -1818 -548 -1814
rect -408 -1814 -374 -1785
rect -408 -1819 -374 -1814
rect 1509 -1730 1543 -1532
rect 1616 -1706 1650 -1630
rect 1704 -1706 1738 -1630
rect 1509 -1732 1543 -1730
rect 1956 -1568 1990 -1534
rect 2148 -1568 2182 -1534
rect 2340 -1568 2374 -1534
rect 2532 -1568 2566 -1534
rect 2724 -1568 2758 -1534
rect 2916 -1568 2950 -1534
rect 1956 -1702 1990 -1622
rect 2052 -1702 2086 -1622
rect 2148 -1702 2182 -1622
rect 2244 -1702 2278 -1622
rect 2340 -1702 2374 -1622
rect 2436 -1702 2470 -1622
rect 2532 -1702 2566 -1622
rect 2628 -1702 2662 -1622
rect 2724 -1702 2758 -1622
rect 2820 -1702 2854 -1622
rect 2916 -1702 2950 -1622
rect 1660 -1790 1694 -1756
rect 3030 -1730 3064 -1532
rect 3030 -1732 3064 -1730
rect -1227 -2126 -1193 -2092
rect -1135 -2126 -1101 -2092
rect -1043 -2126 -1009 -2092
rect -951 -2126 -917 -2092
rect -859 -2126 -825 -2092
rect -767 -2126 -733 -2092
rect -675 -2126 -641 -2092
rect -583 -2126 -549 -2092
rect -491 -2126 -457 -2092
rect -399 -2126 -365 -2092
rect -2042 -2184 -2008 -2182
rect -3116 -2292 -3082 -2212
rect -3020 -2292 -2986 -2212
rect -2924 -2292 -2890 -2212
rect -2828 -2292 -2794 -2212
rect -2732 -2292 -2698 -2212
rect -2636 -2292 -2602 -2212
rect -2540 -2292 -2506 -2212
rect -2444 -2292 -2410 -2212
rect -2348 -2292 -2314 -2212
rect -2252 -2292 -2218 -2212
rect -2156 -2292 -2122 -2212
rect -3116 -2380 -3082 -2346
rect -2924 -2380 -2890 -2346
rect -2732 -2380 -2698 -2346
rect -2540 -2380 -2506 -2346
rect -2348 -2380 -2314 -2346
rect -2156 -2380 -2122 -2346
rect -2042 -2382 -2008 -2184
rect -1004 -2270 -970 -2236
rect -1091 -2404 -1057 -2398
rect -1091 -2432 -1084 -2404
rect -1084 -2432 -1057 -2404
rect -489 -2304 -455 -2270
rect -583 -2404 -549 -2398
rect -583 -2432 -576 -2404
rect -576 -2432 -549 -2404
rect 435 -2282 469 -2034
rect 531 -2282 565 -2034
rect 627 -2282 661 -2034
rect 723 -2282 757 -2034
rect 819 -2282 853 -2034
rect 915 -2282 949 -2034
rect 1011 -2282 1045 -2034
rect 1107 -2282 1141 -2034
rect 1203 -2282 1237 -2034
rect 1299 -2282 1333 -2034
rect 1395 -2282 1429 -2034
rect 435 -2376 469 -2342
rect 627 -2376 661 -2342
rect 819 -2376 853 -2342
rect 1011 -2376 1045 -2342
rect 1203 -2376 1237 -2342
rect 1395 -2376 1429 -2342
rect -402 -2404 -368 -2395
rect -402 -2429 -374 -2404
rect -374 -2429 -368 -2404
rect 1509 -2382 1543 -1996
rect 1956 -2282 1990 -2034
rect 2052 -2282 2086 -2034
rect 2148 -2282 2182 -2034
rect 2244 -2282 2278 -2034
rect 2340 -2282 2374 -2034
rect 2436 -2282 2470 -2034
rect 2532 -2282 2566 -2034
rect 2628 -2282 2662 -2034
rect 2724 -2282 2758 -2034
rect 2820 -2282 2854 -2034
rect 2916 -2282 2950 -2034
rect 1956 -2376 1990 -2342
rect 2148 -2376 2182 -2342
rect 2340 -2376 2374 -2342
rect 2532 -2376 2566 -2342
rect 2724 -2376 2758 -2342
rect 2916 -2376 2950 -2342
rect 3030 -2382 3064 -1996
rect -1227 -2670 -1193 -2636
rect -1135 -2670 -1101 -2636
rect -1043 -2670 -1009 -2636
rect -951 -2670 -917 -2636
rect -859 -2670 -825 -2636
rect -767 -2670 -733 -2636
rect -675 -2670 -641 -2636
rect -583 -2670 -549 -2636
rect -491 -2670 -457 -2636
rect -399 -2670 -365 -2636
rect -3116 -2950 -3082 -2916
rect -2924 -2950 -2890 -2916
rect -2732 -2950 -2698 -2916
rect -2540 -2950 -2506 -2916
rect -2348 -2950 -2314 -2916
rect -2156 -2950 -2122 -2916
rect -3116 -3258 -3082 -3010
rect -3020 -3258 -2986 -3010
rect -2924 -3258 -2890 -3010
rect -2828 -3258 -2794 -3010
rect -2732 -3258 -2698 -3010
rect -2636 -3258 -2602 -3010
rect -2540 -3258 -2506 -3010
rect -2444 -3258 -2410 -3010
rect -2348 -3258 -2314 -3010
rect -2252 -3258 -2218 -3010
rect -2156 -3258 -2122 -3010
rect -2042 -3296 -2008 -2910
rect -1089 -2902 -1084 -2874
rect -1084 -2902 -1055 -2874
rect -1089 -2908 -1055 -2902
rect -994 -2908 -960 -2874
rect -574 -2902 -542 -2874
rect -542 -2902 -540 -2874
rect -574 -2908 -540 -2902
rect -401 -2902 -374 -2875
rect -374 -2902 -367 -2875
rect -401 -2909 -367 -2902
rect -490 -3070 -489 -3036
rect -489 -3070 -456 -3036
rect 435 -2946 469 -2912
rect 627 -2946 661 -2912
rect 819 -2946 853 -2912
rect 1011 -2946 1045 -2912
rect 1203 -2946 1237 -2912
rect 1395 -2946 1429 -2912
rect 435 -3080 469 -3000
rect 531 -3080 565 -3000
rect 627 -3080 661 -3000
rect 723 -3080 757 -3000
rect 819 -3080 853 -3000
rect 915 -3080 949 -3000
rect 1011 -3080 1045 -3000
rect 1107 -3080 1141 -3000
rect 1203 -3080 1237 -3000
rect 1299 -3080 1333 -3000
rect 1395 -3080 1429 -3000
rect 1509 -3108 1543 -2910
rect 1616 -3084 1650 -3008
rect 1704 -3084 1738 -3008
rect 1509 -3110 1543 -3108
rect 1956 -2946 1990 -2912
rect 2148 -2946 2182 -2912
rect 2340 -2946 2374 -2912
rect 2532 -2946 2566 -2912
rect 2724 -2946 2758 -2912
rect 2916 -2946 2950 -2912
rect 1956 -3080 1990 -3000
rect 2052 -3080 2086 -3000
rect 2148 -3080 2182 -3000
rect 2244 -3080 2278 -3000
rect 2340 -3080 2374 -3000
rect 2436 -3080 2470 -3000
rect 2532 -3080 2566 -3000
rect 2628 -3080 2662 -3000
rect 2724 -3080 2758 -3000
rect 2820 -3080 2854 -3000
rect 2916 -3080 2950 -3000
rect 1660 -3168 1694 -3134
rect -1227 -3214 -1193 -3180
rect -1135 -3214 -1101 -3180
rect -1043 -3214 -1009 -3180
rect -951 -3214 -917 -3180
rect -859 -3214 -825 -3180
rect -767 -3214 -733 -3180
rect -675 -3214 -641 -3180
rect -583 -3214 -549 -3180
rect -491 -3214 -457 -3180
rect -399 -3214 -365 -3180
rect 3030 -3108 3064 -2910
rect 3030 -3110 3064 -3108
rect -576 -3526 -542 -3492
rect -2042 -3562 -2008 -3560
rect -3116 -3670 -3082 -3590
rect -3020 -3670 -2986 -3590
rect -2924 -3670 -2890 -3590
rect -2828 -3670 -2794 -3590
rect -2732 -3670 -2698 -3590
rect -2636 -3670 -2602 -3590
rect -2540 -3670 -2506 -3590
rect -2444 -3670 -2410 -3590
rect -2348 -3670 -2314 -3590
rect -2252 -3670 -2218 -3590
rect -2156 -3670 -2122 -3590
rect -3116 -3758 -3082 -3724
rect -2924 -3758 -2890 -3724
rect -2732 -3758 -2698 -3724
rect -2540 -3758 -2506 -3724
rect -2348 -3758 -2314 -3724
rect -2156 -3758 -2122 -3724
rect -2042 -3760 -2008 -3562
rect -405 -3492 -371 -3487
rect -405 -3521 -374 -3492
rect -374 -3521 -371 -3492
rect -492 -3624 -458 -3590
rect -675 -3758 -641 -3724
rect -583 -3758 -549 -3724
rect -491 -3758 -457 -3724
rect -399 -3758 -365 -3724
rect 435 -3660 469 -3412
rect 531 -3660 565 -3412
rect 627 -3660 661 -3412
rect 723 -3660 757 -3412
rect 819 -3660 853 -3412
rect 915 -3660 949 -3412
rect 1011 -3660 1045 -3412
rect 1107 -3660 1141 -3412
rect 1203 -3660 1237 -3412
rect 1299 -3660 1333 -3412
rect 1395 -3660 1429 -3412
rect 435 -3754 469 -3720
rect 627 -3754 661 -3720
rect 819 -3754 853 -3720
rect 1011 -3754 1045 -3720
rect 1203 -3754 1237 -3720
rect 1395 -3754 1429 -3720
rect 1509 -3760 1543 -3374
rect 1956 -3660 1990 -3412
rect 2052 -3660 2086 -3412
rect 2148 -3660 2182 -3412
rect 2244 -3660 2278 -3412
rect 2340 -3660 2374 -3412
rect 2436 -3660 2470 -3412
rect 2532 -3660 2566 -3412
rect 2628 -3660 2662 -3412
rect 2724 -3660 2758 -3412
rect 2820 -3660 2854 -3412
rect 2916 -3660 2950 -3412
rect 1956 -3754 1990 -3720
rect 2148 -3754 2182 -3720
rect 2340 -3754 2374 -3720
rect 2532 -3754 2566 -3720
rect 2724 -3754 2758 -3720
rect 2916 -3754 2950 -3720
rect 3030 -3760 3064 -3374
rect -539 -3990 -532 -3961
rect -532 -3990 -505 -3961
rect -539 -3995 -505 -3990
rect -453 -4124 -419 -4120
rect -453 -4154 -452 -4124
rect -452 -4154 -419 -4124
rect -3116 -4328 -3082 -4294
rect -2924 -4328 -2890 -4294
rect -2732 -4328 -2698 -4294
rect -2540 -4328 -2506 -4294
rect -2348 -4328 -2314 -4294
rect -2156 -4328 -2122 -4294
rect -3116 -4636 -3082 -4388
rect -3020 -4636 -2986 -4388
rect -2924 -4636 -2890 -4388
rect -2828 -4636 -2794 -4388
rect -2732 -4636 -2698 -4388
rect -2636 -4636 -2602 -4388
rect -2540 -4636 -2506 -4388
rect -2444 -4636 -2410 -4388
rect -2348 -4636 -2314 -4388
rect -2252 -4636 -2218 -4388
rect -2156 -4636 -2122 -4388
rect -2042 -4674 -2008 -4288
rect -675 -4302 -641 -4268
rect -583 -4302 -549 -4268
rect -491 -4302 -457 -4268
rect -399 -4302 -365 -4268
rect -452 -4446 -418 -4418
rect -452 -4452 -418 -4446
rect -540 -4580 -506 -4574
rect -540 -4608 -532 -4580
rect -532 -4608 -506 -4580
rect 435 -4324 469 -4290
rect 627 -4324 661 -4290
rect 819 -4324 853 -4290
rect 1011 -4324 1045 -4290
rect 1203 -4324 1237 -4290
rect 1395 -4324 1429 -4290
rect 435 -4458 469 -4378
rect 531 -4458 565 -4378
rect 627 -4458 661 -4378
rect 723 -4458 757 -4378
rect 819 -4458 853 -4378
rect 915 -4458 949 -4378
rect 1011 -4458 1045 -4378
rect 1107 -4458 1141 -4378
rect 1203 -4458 1237 -4378
rect 1299 -4458 1333 -4378
rect 1395 -4458 1429 -4378
rect 1509 -4486 1543 -4288
rect 1616 -4462 1650 -4386
rect 1704 -4462 1738 -4386
rect 1509 -4488 1543 -4486
rect 1956 -4324 1990 -4290
rect 2148 -4324 2182 -4290
rect 2340 -4324 2374 -4290
rect 2532 -4324 2566 -4290
rect 2724 -4324 2758 -4290
rect 2916 -4324 2950 -4290
rect 1956 -4458 1990 -4378
rect 2052 -4458 2086 -4378
rect 2148 -4458 2182 -4378
rect 2244 -4458 2278 -4378
rect 2340 -4458 2374 -4378
rect 2436 -4458 2470 -4378
rect 2532 -4458 2566 -4378
rect 2628 -4458 2662 -4378
rect 2724 -4458 2758 -4378
rect 2820 -4458 2854 -4378
rect 2916 -4458 2950 -4378
rect 1660 -4546 1694 -4512
rect 3030 -4486 3064 -4288
rect 3030 -4488 3064 -4486
rect -675 -4846 -641 -4812
rect -583 -4846 -549 -4812
rect -491 -4846 -457 -4812
rect -399 -4846 -365 -4812
rect -2042 -4940 -2008 -4938
rect -3116 -5048 -3082 -4968
rect -3020 -5048 -2986 -4968
rect -2924 -5048 -2890 -4968
rect -2828 -5048 -2794 -4968
rect -2732 -5048 -2698 -4968
rect -2636 -5048 -2602 -4968
rect -2540 -5048 -2506 -4968
rect -2444 -5048 -2410 -4968
rect -2348 -5048 -2314 -4968
rect -2252 -5048 -2218 -4968
rect -2156 -5048 -2122 -4968
rect -3116 -5136 -3082 -5102
rect -2924 -5136 -2890 -5102
rect -2732 -5136 -2698 -5102
rect -2540 -5136 -2506 -5102
rect -2348 -5136 -2314 -5102
rect -2156 -5136 -2122 -5102
rect -2042 -5138 -2008 -4940
rect 435 -5038 469 -4790
rect 531 -5038 565 -4790
rect 627 -5038 661 -4790
rect 723 -5038 757 -4790
rect 819 -5038 853 -4790
rect 915 -5038 949 -4790
rect 1011 -5038 1045 -4790
rect 1107 -5038 1141 -4790
rect 1203 -5038 1237 -4790
rect 1299 -5038 1333 -4790
rect 1395 -5038 1429 -4790
rect 435 -5132 469 -5098
rect 627 -5132 661 -5098
rect 819 -5132 853 -5098
rect 1011 -5132 1045 -5098
rect 1203 -5132 1237 -5098
rect 1395 -5132 1429 -5098
rect 1509 -5138 1543 -4752
rect 1956 -5038 1990 -4790
rect 2052 -5038 2086 -4790
rect 2148 -5038 2182 -4790
rect 2244 -5038 2278 -4790
rect 2340 -5038 2374 -4790
rect 2436 -5038 2470 -4790
rect 2532 -5038 2566 -4790
rect 2628 -5038 2662 -4790
rect 2724 -5038 2758 -4790
rect 2820 -5038 2854 -4790
rect 2916 -5038 2950 -4790
rect 1956 -5132 1990 -5098
rect 2148 -5132 2182 -5098
rect 2340 -5132 2374 -5098
rect 2532 -5132 2566 -5098
rect 2724 -5132 2758 -5098
rect 2916 -5132 2950 -5098
rect 3030 -5138 3064 -4752
<< metal1 >>
rect -3300 -136 -2218 -102
rect -3429 -246 -3402 -194
rect -3350 -246 -3340 -194
rect -3300 -699 -3266 -136
rect -3135 -246 -3125 -194
rect -3073 -246 -3063 -194
rect -3020 -286 -2986 -136
rect -2942 -246 -2932 -194
rect -2880 -246 -2870 -194
rect -2828 -286 -2794 -136
rect -2751 -246 -2741 -194
rect -2689 -246 -2679 -194
rect -2636 -286 -2602 -136
rect -2559 -246 -2549 -194
rect -2497 -246 -2487 -194
rect -2444 -286 -2410 -136
rect -2367 -246 -2357 -194
rect -2305 -246 -2295 -194
rect -2252 -286 -2218 -136
rect -2175 -246 -2165 -194
rect -2113 -246 -2103 -194
rect -2048 -198 -2002 -66
rect -1597 -121 -1587 -69
rect -1535 -121 -914 -69
rect -862 -121 -852 -69
rect 251 -136 1333 -102
rect -3122 -298 -3076 -286
rect -3122 -546 -3116 -298
rect -3082 -546 -3076 -298
rect -3122 -558 -3076 -546
rect -3026 -298 -2980 -286
rect -3026 -546 -3020 -298
rect -2986 -546 -2980 -298
rect -3026 -558 -2980 -546
rect -2930 -298 -2884 -286
rect -2930 -546 -2924 -298
rect -2890 -546 -2884 -298
rect -2930 -558 -2884 -546
rect -2834 -298 -2788 -286
rect -2834 -546 -2828 -298
rect -2794 -546 -2788 -298
rect -2834 -558 -2788 -546
rect -2738 -298 -2692 -286
rect -2738 -546 -2732 -298
rect -2698 -546 -2692 -298
rect -2738 -558 -2692 -546
rect -2642 -298 -2596 -286
rect -2642 -546 -2636 -298
rect -2602 -546 -2596 -298
rect -2642 -558 -2596 -546
rect -2546 -298 -2500 -286
rect -2546 -546 -2540 -298
rect -2506 -546 -2500 -298
rect -2546 -558 -2500 -546
rect -2450 -298 -2404 -286
rect -2450 -546 -2444 -298
rect -2410 -546 -2404 -298
rect -2450 -558 -2404 -546
rect -2354 -298 -2308 -286
rect -2354 -546 -2348 -298
rect -2314 -546 -2308 -298
rect -2354 -558 -2308 -546
rect -2258 -298 -2212 -286
rect -2258 -546 -2252 -298
rect -2218 -546 -2212 -298
rect -2258 -558 -2212 -546
rect -2162 -298 -2116 -286
rect -2162 -546 -2156 -298
rect -2122 -546 -2116 -298
rect -2162 -558 -2116 -546
rect -3689 -733 -3266 -699
rect -3429 -1053 -3402 -1001
rect -3350 -1053 -3340 -1001
rect -3300 -1110 -3266 -733
rect -3116 -699 -3082 -558
rect -2924 -699 -2890 -558
rect -2732 -699 -2698 -558
rect -2540 -699 -2506 -558
rect -2348 -699 -2314 -558
rect -2156 -699 -2122 -558
rect -2048 -584 -2042 -198
rect -2008 -584 -2002 -198
rect -1952 -246 -1942 -194
rect -1890 -246 -1416 -194
rect -1364 -246 -1354 -194
rect 70 -245 149 -193
rect 201 -245 211 -193
rect -1050 -460 -336 -429
rect -1050 -494 -951 -460
rect -917 -494 -859 -460
rect -825 -494 -767 -460
rect -733 -494 -675 -460
rect -641 -494 -583 -460
rect -549 -494 -491 -460
rect -457 -494 -399 -460
rect -365 -494 -336 -460
rect -1050 -525 -336 -494
rect 251 -513 285 -136
rect 419 -193 485 -188
rect 416 -245 426 -193
rect 478 -245 488 -193
rect 419 -248 485 -245
rect 531 -276 565 -136
rect 611 -193 677 -188
rect 607 -245 617 -193
rect 669 -245 679 -193
rect 611 -248 677 -245
rect 723 -276 757 -136
rect 803 -193 869 -188
rect 799 -245 809 -193
rect 861 -245 871 -193
rect 803 -248 869 -245
rect 915 -276 949 -136
rect 995 -193 1061 -188
rect 991 -245 1001 -193
rect 1053 -245 1063 -193
rect 995 -248 1061 -245
rect 1107 -276 1141 -136
rect 1187 -192 1253 -188
rect 1184 -244 1194 -192
rect 1246 -244 1256 -192
rect 1187 -248 1253 -244
rect 1299 -276 1333 -136
rect 1379 -192 1445 -188
rect 1376 -244 1386 -192
rect 1438 -244 1448 -192
rect 1503 -198 1549 -26
rect 1772 -136 2854 -102
rect 1379 -248 1445 -244
rect 429 -288 475 -276
rect 429 -368 435 -288
rect 469 -368 475 -288
rect 429 -380 475 -368
rect 525 -288 571 -276
rect 525 -368 531 -288
rect 565 -368 571 -288
rect 525 -380 571 -368
rect 621 -288 667 -276
rect 621 -368 627 -288
rect 661 -368 667 -288
rect 621 -380 667 -368
rect 717 -288 763 -276
rect 717 -368 723 -288
rect 757 -368 763 -288
rect 717 -380 763 -368
rect 813 -288 859 -276
rect 813 -368 819 -288
rect 853 -368 859 -288
rect 813 -380 859 -368
rect 909 -288 955 -276
rect 909 -368 915 -288
rect 949 -368 955 -288
rect 909 -380 955 -368
rect 1005 -288 1051 -276
rect 1005 -368 1011 -288
rect 1045 -368 1051 -288
rect 1005 -380 1051 -368
rect 1101 -288 1147 -276
rect 1101 -368 1107 -288
rect 1141 -368 1147 -288
rect 1101 -380 1147 -368
rect 1197 -288 1243 -276
rect 1197 -368 1203 -288
rect 1237 -368 1243 -288
rect 1197 -380 1243 -368
rect 1293 -288 1339 -276
rect 1293 -368 1299 -288
rect 1333 -368 1339 -288
rect 1293 -380 1339 -368
rect 1389 -288 1435 -276
rect 1389 -368 1395 -288
rect 1429 -368 1435 -288
rect 1389 -380 1435 -368
rect -80 -547 285 -513
rect -2048 -596 -2002 -584
rect -1426 -645 -1416 -593
rect -1364 -597 -1354 -593
rect -1364 -603 -776 -597
rect -1364 -637 -822 -603
rect -788 -637 -776 -603
rect -471 -636 -461 -584
rect -409 -636 -399 -584
rect -1364 -643 -776 -637
rect -1364 -645 -1354 -643
rect -3116 -733 -1797 -699
rect -3116 -866 -3082 -733
rect -2924 -866 -2890 -733
rect -2732 -866 -2698 -733
rect -2540 -866 -2506 -733
rect -2348 -866 -2314 -733
rect -2156 -866 -2122 -733
rect -2048 -848 -2002 -836
rect -3122 -878 -3076 -866
rect -3122 -958 -3116 -878
rect -3082 -958 -3076 -878
rect -3122 -970 -3076 -958
rect -3026 -878 -2980 -866
rect -3026 -958 -3020 -878
rect -2986 -958 -2980 -878
rect -3026 -970 -2980 -958
rect -2930 -878 -2884 -866
rect -2930 -958 -2924 -878
rect -2890 -958 -2884 -878
rect -2930 -970 -2884 -958
rect -2834 -878 -2788 -866
rect -2834 -958 -2828 -878
rect -2794 -958 -2788 -878
rect -2834 -970 -2788 -958
rect -2738 -878 -2692 -866
rect -2738 -958 -2732 -878
rect -2698 -958 -2692 -878
rect -2738 -970 -2692 -958
rect -2642 -878 -2596 -866
rect -2642 -958 -2636 -878
rect -2602 -958 -2596 -878
rect -2642 -970 -2596 -958
rect -2546 -878 -2500 -866
rect -2546 -958 -2540 -878
rect -2506 -958 -2500 -878
rect -2546 -970 -2500 -958
rect -2450 -878 -2404 -866
rect -2450 -958 -2444 -878
rect -2410 -958 -2404 -878
rect -2450 -970 -2404 -958
rect -2354 -878 -2308 -866
rect -2354 -958 -2348 -878
rect -2314 -958 -2308 -878
rect -2354 -970 -2308 -958
rect -2258 -878 -2212 -866
rect -2258 -958 -2252 -878
rect -2218 -958 -2212 -878
rect -2258 -970 -2212 -958
rect -2162 -878 -2116 -866
rect -2162 -958 -2156 -878
rect -2122 -958 -2116 -878
rect -2162 -970 -2116 -958
rect -3132 -1001 -3066 -998
rect -3135 -1053 -3125 -1001
rect -3073 -1053 -3063 -1001
rect -3132 -1058 -3066 -1053
rect -3020 -1110 -2986 -970
rect -2940 -1001 -2874 -998
rect -2944 -1053 -2934 -1001
rect -2882 -1053 -2872 -1001
rect -2940 -1058 -2874 -1053
rect -2828 -1110 -2794 -970
rect -2748 -1001 -2682 -998
rect -2752 -1053 -2742 -1001
rect -2690 -1053 -2680 -1001
rect -2748 -1058 -2682 -1053
rect -2636 -1110 -2602 -970
rect -2556 -1001 -2490 -998
rect -2560 -1053 -2550 -1001
rect -2498 -1053 -2488 -1001
rect -2556 -1058 -2490 -1053
rect -2444 -1110 -2410 -970
rect -2364 -1002 -2298 -998
rect -2367 -1054 -2357 -1002
rect -2305 -1054 -2295 -1002
rect -2364 -1058 -2298 -1054
rect -2252 -1110 -2218 -970
rect -2172 -1002 -2106 -998
rect -2175 -1054 -2165 -1002
rect -2113 -1054 -2103 -1002
rect -2048 -1048 -2042 -848
rect -2008 -1048 -2002 -848
rect -1831 -870 -1797 -733
rect -924 -742 -914 -690
rect -862 -742 -852 -690
rect -559 -746 -549 -694
rect -497 -746 -487 -694
rect -80 -870 -46 -547
rect -1831 -904 -46 -870
rect -980 -974 -336 -973
rect -2172 -1058 -2106 -1054
rect -3300 -1144 -2218 -1110
rect -2048 -1180 -2002 -1048
rect -1050 -1004 -336 -974
rect -1050 -1038 -951 -1004
rect -917 -1038 -859 -1004
rect -825 -1038 -767 -1004
rect -733 -1038 -675 -1004
rect -641 -1038 -583 -1004
rect -549 -1038 -491 -1004
rect -457 -1038 -399 -1004
rect -365 -1038 -336 -1004
rect -1050 -1069 -336 -1038
rect 70 -1052 149 -1000
rect 201 -1052 211 -1000
rect -1050 -1070 -951 -1069
rect 251 -1110 285 -547
rect 435 -513 469 -380
rect 627 -513 661 -380
rect 819 -513 853 -380
rect 1011 -513 1045 -380
rect 1203 -513 1237 -380
rect 1395 -513 1429 -380
rect 1503 -398 1509 -198
rect 1543 -285 1549 -198
rect 1643 -245 1670 -193
rect 1722 -245 1732 -193
rect 1610 -285 1656 -284
rect 1543 -296 1656 -285
rect 1543 -372 1616 -296
rect 1650 -372 1656 -296
rect 1543 -384 1656 -372
rect 1698 -285 1744 -284
rect 1772 -285 1806 -136
rect 1940 -193 2006 -188
rect 1937 -245 1947 -193
rect 1999 -245 2009 -193
rect 1940 -248 2006 -245
rect 2052 -276 2086 -136
rect 2132 -193 2198 -188
rect 2128 -245 2138 -193
rect 2190 -245 2200 -193
rect 2132 -248 2198 -245
rect 2244 -276 2278 -136
rect 2324 -193 2390 -188
rect 2320 -245 2330 -193
rect 2382 -245 2392 -193
rect 2324 -248 2390 -245
rect 2436 -276 2470 -136
rect 2516 -193 2582 -188
rect 2512 -245 2522 -193
rect 2574 -245 2584 -193
rect 2516 -248 2582 -245
rect 2628 -276 2662 -136
rect 2708 -192 2774 -188
rect 2705 -244 2715 -192
rect 2767 -244 2777 -192
rect 2708 -248 2774 -244
rect 2820 -276 2854 -136
rect 2900 -192 2966 -188
rect 2897 -244 2907 -192
rect 2959 -244 2969 -192
rect 3024 -198 3070 -26
rect 2900 -248 2966 -244
rect 1698 -296 1806 -285
rect 1698 -372 1704 -296
rect 1738 -372 1806 -296
rect 1698 -384 1806 -372
rect 1950 -288 1996 -276
rect 1950 -368 1956 -288
rect 1990 -368 1996 -288
rect 1950 -380 1996 -368
rect 2046 -288 2092 -276
rect 2046 -368 2052 -288
rect 2086 -368 2092 -288
rect 2046 -380 2092 -368
rect 2142 -288 2188 -276
rect 2142 -368 2148 -288
rect 2182 -368 2188 -288
rect 2142 -380 2188 -368
rect 2238 -288 2284 -276
rect 2238 -368 2244 -288
rect 2278 -368 2284 -288
rect 2238 -380 2284 -368
rect 2334 -288 2380 -276
rect 2334 -368 2340 -288
rect 2374 -368 2380 -288
rect 2334 -380 2380 -368
rect 2430 -288 2476 -276
rect 2430 -368 2436 -288
rect 2470 -368 2476 -288
rect 2430 -380 2476 -368
rect 2526 -288 2572 -276
rect 2526 -368 2532 -288
rect 2566 -368 2572 -288
rect 2526 -380 2572 -368
rect 2622 -288 2668 -276
rect 2622 -368 2628 -288
rect 2662 -368 2668 -288
rect 2622 -380 2668 -368
rect 2718 -288 2764 -276
rect 2718 -368 2724 -288
rect 2758 -368 2764 -288
rect 2718 -380 2764 -368
rect 2814 -288 2860 -276
rect 2814 -368 2820 -288
rect 2854 -368 2860 -288
rect 2814 -380 2860 -368
rect 2910 -288 2956 -276
rect 2910 -368 2916 -288
rect 2950 -368 2956 -288
rect 2910 -380 2956 -368
rect 1543 -385 1649 -384
rect 1703 -385 1806 -384
rect 1543 -398 1549 -385
rect 1503 -410 1549 -398
rect 1648 -422 1706 -416
rect 1648 -423 1660 -422
rect 1694 -423 1706 -422
rect 1640 -475 1650 -423
rect 1702 -475 1712 -423
rect 1772 -513 1806 -385
rect 435 -547 1806 -513
rect 435 -688 469 -547
rect 627 -688 661 -547
rect 819 -688 853 -547
rect 1011 -688 1045 -547
rect 1203 -688 1237 -547
rect 1395 -688 1429 -547
rect 1503 -662 1549 -650
rect 429 -700 475 -688
rect 429 -948 435 -700
rect 469 -948 475 -700
rect 429 -960 475 -948
rect 525 -700 571 -688
rect 525 -948 531 -700
rect 565 -948 571 -700
rect 525 -960 571 -948
rect 621 -700 667 -688
rect 621 -948 627 -700
rect 661 -948 667 -700
rect 621 -960 667 -948
rect 717 -700 763 -688
rect 717 -948 723 -700
rect 757 -948 763 -700
rect 717 -960 763 -948
rect 813 -700 859 -688
rect 813 -948 819 -700
rect 853 -948 859 -700
rect 813 -960 859 -948
rect 909 -700 955 -688
rect 909 -948 915 -700
rect 949 -948 955 -700
rect 909 -960 955 -948
rect 1005 -700 1051 -688
rect 1005 -948 1011 -700
rect 1045 -948 1051 -700
rect 1005 -960 1051 -948
rect 1101 -700 1147 -688
rect 1101 -948 1107 -700
rect 1141 -948 1147 -700
rect 1101 -960 1147 -948
rect 1197 -700 1243 -688
rect 1197 -948 1203 -700
rect 1237 -948 1243 -700
rect 1197 -960 1243 -948
rect 1293 -700 1339 -688
rect 1293 -948 1299 -700
rect 1333 -948 1339 -700
rect 1293 -960 1339 -948
rect 1389 -700 1435 -688
rect 1389 -948 1395 -700
rect 1429 -948 1435 -700
rect 1389 -960 1435 -948
rect 416 -1052 426 -1000
rect 478 -1052 488 -1000
rect 531 -1110 565 -960
rect 609 -1052 619 -1000
rect 671 -1052 681 -1000
rect 723 -1110 757 -960
rect 800 -1052 810 -1000
rect 862 -1052 872 -1000
rect 915 -1110 949 -960
rect 992 -1052 1002 -1000
rect 1054 -1052 1064 -1000
rect 1107 -1110 1141 -960
rect 1184 -1052 1194 -1000
rect 1246 -1052 1256 -1000
rect 1299 -1110 1333 -960
rect 1376 -1052 1386 -1000
rect 1438 -1052 1448 -1000
rect 1503 -1048 1509 -662
rect 1543 -1048 1549 -662
rect 251 -1144 1333 -1110
rect 88 -1191 98 -1188
rect -465 -1197 98 -1191
rect -465 -1231 -453 -1197
rect -419 -1231 98 -1197
rect -465 -1237 98 -1231
rect 88 -1240 98 -1237
rect 150 -1240 160 -1188
rect 1503 -1224 1549 -1048
rect 1643 -1052 1670 -1000
rect 1722 -1052 1732 -1000
rect 1772 -1110 1806 -547
rect 1956 -513 1990 -380
rect 2148 -513 2182 -380
rect 2340 -513 2374 -380
rect 2532 -513 2566 -380
rect 2724 -513 2758 -380
rect 2916 -513 2950 -380
rect 3024 -398 3030 -198
rect 3064 -398 3070 -198
rect 3024 -410 3070 -398
rect 1956 -547 3307 -513
rect 1956 -688 1990 -547
rect 2148 -688 2182 -547
rect 2340 -688 2374 -547
rect 2532 -688 2566 -547
rect 2724 -688 2758 -547
rect 2916 -688 2950 -547
rect 3024 -662 3070 -650
rect 1950 -700 1996 -688
rect 1950 -948 1956 -700
rect 1990 -948 1996 -700
rect 1950 -960 1996 -948
rect 2046 -700 2092 -688
rect 2046 -948 2052 -700
rect 2086 -948 2092 -700
rect 2046 -960 2092 -948
rect 2142 -700 2188 -688
rect 2142 -948 2148 -700
rect 2182 -948 2188 -700
rect 2142 -960 2188 -948
rect 2238 -700 2284 -688
rect 2238 -948 2244 -700
rect 2278 -948 2284 -700
rect 2238 -960 2284 -948
rect 2334 -700 2380 -688
rect 2334 -948 2340 -700
rect 2374 -948 2380 -700
rect 2334 -960 2380 -948
rect 2430 -700 2476 -688
rect 2430 -948 2436 -700
rect 2470 -948 2476 -700
rect 2430 -960 2476 -948
rect 2526 -700 2572 -688
rect 2526 -948 2532 -700
rect 2566 -948 2572 -700
rect 2526 -960 2572 -948
rect 2622 -700 2668 -688
rect 2622 -948 2628 -700
rect 2662 -948 2668 -700
rect 2622 -960 2668 -948
rect 2718 -700 2764 -688
rect 2718 -948 2724 -700
rect 2758 -948 2764 -700
rect 2718 -960 2764 -948
rect 2814 -700 2860 -688
rect 2814 -948 2820 -700
rect 2854 -948 2860 -700
rect 2814 -960 2860 -948
rect 2910 -700 2956 -688
rect 2910 -948 2916 -700
rect 2950 -948 2956 -700
rect 2910 -960 2956 -948
rect 1937 -1052 1947 -1000
rect 1999 -1052 2009 -1000
rect 2052 -1110 2086 -960
rect 2130 -1052 2140 -1000
rect 2192 -1052 2202 -1000
rect 2244 -1110 2278 -960
rect 2321 -1052 2331 -1000
rect 2383 -1052 2393 -1000
rect 2436 -1110 2470 -960
rect 2513 -1052 2523 -1000
rect 2575 -1052 2585 -1000
rect 2628 -1110 2662 -960
rect 2705 -1052 2715 -1000
rect 2767 -1052 2777 -1000
rect 2820 -1110 2854 -960
rect 2897 -1052 2907 -1000
rect 2959 -1052 2969 -1000
rect 3024 -1048 3030 -662
rect 3064 -1048 3070 -662
rect 1772 -1144 2854 -1110
rect 3024 -1224 3070 -1048
rect -549 -1312 -287 -1303
rect -549 -1346 -534 -1312
rect -500 -1346 -287 -1312
rect -549 -1355 -287 -1346
rect -235 -1355 -225 -1303
rect -3300 -1470 -2218 -1436
rect -3429 -1580 -3402 -1528
rect -3350 -1580 -3340 -1528
rect -3300 -2033 -3266 -1470
rect -3135 -1580 -3125 -1528
rect -3073 -1580 -3063 -1528
rect -3020 -1620 -2986 -1470
rect -2942 -1580 -2932 -1528
rect -2880 -1580 -2870 -1528
rect -2828 -1620 -2794 -1470
rect -2751 -1580 -2741 -1528
rect -2689 -1580 -2679 -1528
rect -2636 -1620 -2602 -1470
rect -2559 -1580 -2549 -1528
rect -2497 -1580 -2487 -1528
rect -2444 -1620 -2410 -1470
rect -2367 -1580 -2357 -1528
rect -2305 -1580 -2295 -1528
rect -2252 -1620 -2218 -1470
rect -2175 -1580 -2165 -1528
rect -2113 -1580 -2103 -1528
rect -2048 -1532 -2002 -1400
rect -3122 -1632 -3076 -1620
rect -3122 -1880 -3116 -1632
rect -3082 -1880 -3076 -1632
rect -3122 -1892 -3076 -1880
rect -3026 -1632 -2980 -1620
rect -3026 -1880 -3020 -1632
rect -2986 -1880 -2980 -1632
rect -3026 -1892 -2980 -1880
rect -2930 -1632 -2884 -1620
rect -2930 -1880 -2924 -1632
rect -2890 -1880 -2884 -1632
rect -2930 -1892 -2884 -1880
rect -2834 -1632 -2788 -1620
rect -2834 -1880 -2828 -1632
rect -2794 -1880 -2788 -1632
rect -2834 -1892 -2788 -1880
rect -2738 -1632 -2692 -1620
rect -2738 -1880 -2732 -1632
rect -2698 -1880 -2692 -1632
rect -2738 -1892 -2692 -1880
rect -2642 -1632 -2596 -1620
rect -2642 -1880 -2636 -1632
rect -2602 -1880 -2596 -1632
rect -2642 -1892 -2596 -1880
rect -2546 -1632 -2500 -1620
rect -2546 -1880 -2540 -1632
rect -2506 -1880 -2500 -1632
rect -2546 -1892 -2500 -1880
rect -2450 -1632 -2404 -1620
rect -2450 -1880 -2444 -1632
rect -2410 -1880 -2404 -1632
rect -2450 -1892 -2404 -1880
rect -2354 -1632 -2308 -1620
rect -2354 -1880 -2348 -1632
rect -2314 -1880 -2308 -1632
rect -2354 -1892 -2308 -1880
rect -2258 -1632 -2212 -1620
rect -2258 -1880 -2252 -1632
rect -2218 -1880 -2212 -1632
rect -2258 -1892 -2212 -1880
rect -2162 -1632 -2116 -1620
rect -2162 -1880 -2156 -1632
rect -2122 -1880 -2116 -1632
rect -2162 -1892 -2116 -1880
rect -3690 -2067 -3266 -2033
rect -3429 -2387 -3402 -2335
rect -3350 -2387 -3340 -2335
rect -3300 -2444 -3266 -2067
rect -3116 -2033 -3082 -1892
rect -2924 -2033 -2890 -1892
rect -2732 -2033 -2698 -1892
rect -2540 -2033 -2506 -1892
rect -2348 -2033 -2314 -1892
rect -2156 -2033 -2122 -1892
rect -2048 -1918 -2042 -1532
rect -2008 -1918 -2002 -1532
rect -2048 -1930 -2002 -1918
rect -1852 -1446 -50 -1412
rect -1852 -2033 -1818 -1446
rect -1734 -1580 -1724 -1528
rect -1672 -1580 -1416 -1528
rect -1364 -1580 -1354 -1528
rect -782 -1548 -336 -1517
rect -782 -1582 -675 -1548
rect -641 -1582 -583 -1548
rect -549 -1582 -491 -1548
rect -457 -1582 -399 -1548
rect -365 -1582 -336 -1548
rect -782 -1613 -336 -1582
rect -488 -1721 -478 -1669
rect -426 -1721 -416 -1669
rect -602 -1828 -592 -1776
rect -540 -1828 -530 -1776
rect -426 -1831 -416 -1779
rect -364 -1831 -354 -1779
rect -84 -1847 -50 -1446
rect 251 -1470 1333 -1436
rect 70 -1579 149 -1527
rect 201 -1579 211 -1527
rect 251 -1847 285 -1470
rect 419 -1527 485 -1522
rect 416 -1579 426 -1527
rect 478 -1579 488 -1527
rect 419 -1582 485 -1579
rect 531 -1610 565 -1470
rect 611 -1527 677 -1522
rect 607 -1579 617 -1527
rect 669 -1579 679 -1527
rect 611 -1582 677 -1579
rect 723 -1610 757 -1470
rect 803 -1527 869 -1522
rect 799 -1579 809 -1527
rect 861 -1579 871 -1527
rect 803 -1582 869 -1579
rect 915 -1610 949 -1470
rect 995 -1527 1061 -1522
rect 991 -1579 1001 -1527
rect 1053 -1579 1063 -1527
rect 995 -1582 1061 -1579
rect 1107 -1610 1141 -1470
rect 1187 -1526 1253 -1522
rect 1184 -1578 1194 -1526
rect 1246 -1578 1256 -1526
rect 1187 -1582 1253 -1578
rect 1299 -1610 1333 -1470
rect 1379 -1526 1445 -1522
rect 1376 -1578 1386 -1526
rect 1438 -1578 1448 -1526
rect 1503 -1532 1549 -1360
rect 1772 -1470 2854 -1436
rect 1379 -1582 1445 -1578
rect 429 -1622 475 -1610
rect 429 -1702 435 -1622
rect 469 -1702 475 -1622
rect 429 -1714 475 -1702
rect 525 -1622 571 -1610
rect 525 -1702 531 -1622
rect 565 -1702 571 -1622
rect 525 -1714 571 -1702
rect 621 -1622 667 -1610
rect 621 -1702 627 -1622
rect 661 -1702 667 -1622
rect 621 -1714 667 -1702
rect 717 -1622 763 -1610
rect 717 -1702 723 -1622
rect 757 -1702 763 -1622
rect 717 -1714 763 -1702
rect 813 -1622 859 -1610
rect 813 -1702 819 -1622
rect 853 -1702 859 -1622
rect 813 -1714 859 -1702
rect 909 -1622 955 -1610
rect 909 -1702 915 -1622
rect 949 -1702 955 -1622
rect 909 -1714 955 -1702
rect 1005 -1622 1051 -1610
rect 1005 -1702 1011 -1622
rect 1045 -1702 1051 -1622
rect 1005 -1714 1051 -1702
rect 1101 -1622 1147 -1610
rect 1101 -1702 1107 -1622
rect 1141 -1702 1147 -1622
rect 1101 -1714 1147 -1702
rect 1197 -1622 1243 -1610
rect 1197 -1702 1203 -1622
rect 1237 -1702 1243 -1622
rect 1197 -1714 1243 -1702
rect 1293 -1622 1339 -1610
rect 1293 -1702 1299 -1622
rect 1333 -1702 1339 -1622
rect 1293 -1714 1339 -1702
rect 1389 -1622 1435 -1610
rect 1389 -1702 1395 -1622
rect 1429 -1702 1435 -1622
rect 1389 -1714 1435 -1702
rect -84 -1881 285 -1847
rect -882 -1971 -872 -1919
rect -820 -1971 -416 -1919
rect -364 -1971 -354 -1919
rect -3116 -2067 -1818 -2033
rect -3116 -2200 -3082 -2067
rect -2924 -2200 -2890 -2067
rect -2732 -2200 -2698 -2067
rect -2540 -2200 -2506 -2067
rect -2348 -2200 -2314 -2067
rect -2156 -2200 -2122 -2067
rect -1326 -2092 -336 -2061
rect -1326 -2126 -1227 -2092
rect -1193 -2126 -1135 -2092
rect -1101 -2126 -1043 -2092
rect -1009 -2126 -951 -2092
rect -917 -2126 -859 -2092
rect -825 -2126 -767 -2092
rect -733 -2126 -675 -2092
rect -641 -2126 -583 -2092
rect -549 -2126 -491 -2092
rect -457 -2126 -399 -2092
rect -365 -2126 -336 -2092
rect -1326 -2157 -336 -2126
rect -2048 -2182 -2002 -2170
rect -3122 -2212 -3076 -2200
rect -3122 -2292 -3116 -2212
rect -3082 -2292 -3076 -2212
rect -3122 -2304 -3076 -2292
rect -3026 -2212 -2980 -2200
rect -3026 -2292 -3020 -2212
rect -2986 -2292 -2980 -2212
rect -3026 -2304 -2980 -2292
rect -2930 -2212 -2884 -2200
rect -2930 -2292 -2924 -2212
rect -2890 -2292 -2884 -2212
rect -2930 -2304 -2884 -2292
rect -2834 -2212 -2788 -2200
rect -2834 -2292 -2828 -2212
rect -2794 -2292 -2788 -2212
rect -2834 -2304 -2788 -2292
rect -2738 -2212 -2692 -2200
rect -2738 -2292 -2732 -2212
rect -2698 -2292 -2692 -2212
rect -2738 -2304 -2692 -2292
rect -2642 -2212 -2596 -2200
rect -2642 -2292 -2636 -2212
rect -2602 -2292 -2596 -2212
rect -2642 -2304 -2596 -2292
rect -2546 -2212 -2500 -2200
rect -2546 -2292 -2540 -2212
rect -2506 -2292 -2500 -2212
rect -2546 -2304 -2500 -2292
rect -2450 -2212 -2404 -2200
rect -2450 -2292 -2444 -2212
rect -2410 -2292 -2404 -2212
rect -2450 -2304 -2404 -2292
rect -2354 -2212 -2308 -2200
rect -2354 -2292 -2348 -2212
rect -2314 -2292 -2308 -2212
rect -2354 -2304 -2308 -2292
rect -2258 -2212 -2212 -2200
rect -2258 -2292 -2252 -2212
rect -2218 -2292 -2212 -2212
rect -2258 -2304 -2212 -2292
rect -2162 -2212 -2116 -2200
rect -2162 -2292 -2156 -2212
rect -2122 -2292 -2116 -2212
rect -2162 -2304 -2116 -2292
rect -3132 -2335 -3066 -2332
rect -3135 -2387 -3125 -2335
rect -3073 -2387 -3063 -2335
rect -3132 -2392 -3066 -2387
rect -3020 -2444 -2986 -2304
rect -2940 -2335 -2874 -2332
rect -2944 -2387 -2934 -2335
rect -2882 -2387 -2872 -2335
rect -2940 -2392 -2874 -2387
rect -2828 -2444 -2794 -2304
rect -2748 -2335 -2682 -2332
rect -2752 -2387 -2742 -2335
rect -2690 -2387 -2680 -2335
rect -2748 -2392 -2682 -2387
rect -2636 -2444 -2602 -2304
rect -2556 -2335 -2490 -2332
rect -2560 -2387 -2550 -2335
rect -2498 -2387 -2488 -2335
rect -2556 -2392 -2490 -2387
rect -2444 -2444 -2410 -2304
rect -2364 -2336 -2298 -2332
rect -2367 -2388 -2357 -2336
rect -2305 -2388 -2295 -2336
rect -2364 -2392 -2298 -2388
rect -2252 -2444 -2218 -2304
rect -2172 -2336 -2106 -2332
rect -2175 -2388 -2165 -2336
rect -2113 -2388 -2103 -2336
rect -2048 -2382 -2042 -2182
rect -2008 -2382 -2002 -2182
rect -602 -2230 -592 -2225
rect -1016 -2236 -592 -2230
rect -1016 -2270 -1004 -2236
rect -970 -2270 -592 -2236
rect -1016 -2276 -592 -2270
rect -602 -2277 -592 -2276
rect -540 -2277 -530 -2225
rect -297 -2264 -287 -2261
rect -501 -2270 -287 -2264
rect -501 -2304 -489 -2270
rect -455 -2304 -287 -2270
rect -501 -2310 -287 -2304
rect -297 -2313 -287 -2310
rect -235 -2313 -225 -2261
rect -2172 -2392 -2106 -2388
rect -3300 -2478 -2218 -2444
rect -2048 -2514 -2002 -2382
rect -1111 -2440 -1101 -2388
rect -1049 -2440 -762 -2388
rect -710 -2440 -700 -2388
rect -602 -2442 -592 -2390
rect -540 -2442 -530 -2390
rect -422 -2437 -412 -2385
rect -360 -2437 -350 -2385
rect 70 -2386 149 -2334
rect 201 -2386 211 -2334
rect 251 -2444 285 -1881
rect 435 -1847 469 -1714
rect 627 -1847 661 -1714
rect 819 -1847 853 -1714
rect 1011 -1847 1045 -1714
rect 1203 -1847 1237 -1714
rect 1395 -1847 1429 -1714
rect 1503 -1732 1509 -1532
rect 1543 -1619 1549 -1532
rect 1643 -1579 1670 -1527
rect 1722 -1579 1732 -1527
rect 1610 -1619 1656 -1618
rect 1543 -1630 1656 -1619
rect 1543 -1706 1616 -1630
rect 1650 -1706 1656 -1630
rect 1543 -1718 1656 -1706
rect 1698 -1619 1744 -1618
rect 1772 -1619 1806 -1470
rect 1940 -1527 2006 -1522
rect 1937 -1579 1947 -1527
rect 1999 -1579 2009 -1527
rect 1940 -1582 2006 -1579
rect 2052 -1610 2086 -1470
rect 2132 -1527 2198 -1522
rect 2128 -1579 2138 -1527
rect 2190 -1579 2200 -1527
rect 2132 -1582 2198 -1579
rect 2244 -1610 2278 -1470
rect 2324 -1527 2390 -1522
rect 2320 -1579 2330 -1527
rect 2382 -1579 2392 -1527
rect 2324 -1582 2390 -1579
rect 2436 -1610 2470 -1470
rect 2516 -1527 2582 -1522
rect 2512 -1579 2522 -1527
rect 2574 -1579 2584 -1527
rect 2516 -1582 2582 -1579
rect 2628 -1610 2662 -1470
rect 2708 -1526 2774 -1522
rect 2705 -1578 2715 -1526
rect 2767 -1578 2777 -1526
rect 2708 -1582 2774 -1578
rect 2820 -1610 2854 -1470
rect 2900 -1526 2966 -1522
rect 2897 -1578 2907 -1526
rect 2959 -1578 2969 -1526
rect 3024 -1532 3070 -1360
rect 2900 -1582 2966 -1578
rect 1698 -1630 1806 -1619
rect 1698 -1706 1704 -1630
rect 1738 -1706 1806 -1630
rect 1698 -1718 1806 -1706
rect 1950 -1622 1996 -1610
rect 1950 -1702 1956 -1622
rect 1990 -1702 1996 -1622
rect 1950 -1714 1996 -1702
rect 2046 -1622 2092 -1610
rect 2046 -1702 2052 -1622
rect 2086 -1702 2092 -1622
rect 2046 -1714 2092 -1702
rect 2142 -1622 2188 -1610
rect 2142 -1702 2148 -1622
rect 2182 -1702 2188 -1622
rect 2142 -1714 2188 -1702
rect 2238 -1622 2284 -1610
rect 2238 -1702 2244 -1622
rect 2278 -1702 2284 -1622
rect 2238 -1714 2284 -1702
rect 2334 -1622 2380 -1610
rect 2334 -1702 2340 -1622
rect 2374 -1702 2380 -1622
rect 2334 -1714 2380 -1702
rect 2430 -1622 2476 -1610
rect 2430 -1702 2436 -1622
rect 2470 -1702 2476 -1622
rect 2430 -1714 2476 -1702
rect 2526 -1622 2572 -1610
rect 2526 -1702 2532 -1622
rect 2566 -1702 2572 -1622
rect 2526 -1714 2572 -1702
rect 2622 -1622 2668 -1610
rect 2622 -1702 2628 -1622
rect 2662 -1702 2668 -1622
rect 2622 -1714 2668 -1702
rect 2718 -1622 2764 -1610
rect 2718 -1702 2724 -1622
rect 2758 -1702 2764 -1622
rect 2718 -1714 2764 -1702
rect 2814 -1622 2860 -1610
rect 2814 -1702 2820 -1622
rect 2854 -1702 2860 -1622
rect 2814 -1714 2860 -1702
rect 2910 -1622 2956 -1610
rect 2910 -1702 2916 -1622
rect 2950 -1702 2956 -1622
rect 2910 -1714 2956 -1702
rect 1543 -1719 1649 -1718
rect 1703 -1719 1806 -1718
rect 1543 -1732 1549 -1719
rect 1503 -1744 1549 -1732
rect 1648 -1756 1706 -1750
rect 1648 -1757 1660 -1756
rect 1694 -1757 1706 -1756
rect 1640 -1809 1650 -1757
rect 1702 -1809 1712 -1757
rect 1772 -1847 1806 -1719
rect 435 -1881 1806 -1847
rect 435 -2022 469 -1881
rect 627 -2022 661 -1881
rect 819 -2022 853 -1881
rect 1011 -2022 1045 -1881
rect 1203 -2022 1237 -1881
rect 1395 -2022 1429 -1881
rect 1503 -1996 1549 -1984
rect 429 -2034 475 -2022
rect 429 -2282 435 -2034
rect 469 -2282 475 -2034
rect 429 -2294 475 -2282
rect 525 -2034 571 -2022
rect 525 -2282 531 -2034
rect 565 -2282 571 -2034
rect 525 -2294 571 -2282
rect 621 -2034 667 -2022
rect 621 -2282 627 -2034
rect 661 -2282 667 -2034
rect 621 -2294 667 -2282
rect 717 -2034 763 -2022
rect 717 -2282 723 -2034
rect 757 -2282 763 -2034
rect 717 -2294 763 -2282
rect 813 -2034 859 -2022
rect 813 -2282 819 -2034
rect 853 -2282 859 -2034
rect 813 -2294 859 -2282
rect 909 -2034 955 -2022
rect 909 -2282 915 -2034
rect 949 -2282 955 -2034
rect 909 -2294 955 -2282
rect 1005 -2034 1051 -2022
rect 1005 -2282 1011 -2034
rect 1045 -2282 1051 -2034
rect 1005 -2294 1051 -2282
rect 1101 -2034 1147 -2022
rect 1101 -2282 1107 -2034
rect 1141 -2282 1147 -2034
rect 1101 -2294 1147 -2282
rect 1197 -2034 1243 -2022
rect 1197 -2282 1203 -2034
rect 1237 -2282 1243 -2034
rect 1197 -2294 1243 -2282
rect 1293 -2034 1339 -2022
rect 1293 -2282 1299 -2034
rect 1333 -2282 1339 -2034
rect 1293 -2294 1339 -2282
rect 1389 -2034 1435 -2022
rect 1389 -2282 1395 -2034
rect 1429 -2282 1435 -2034
rect 1389 -2294 1435 -2282
rect 416 -2386 426 -2334
rect 478 -2386 488 -2334
rect 531 -2444 565 -2294
rect 609 -2386 619 -2334
rect 671 -2386 681 -2334
rect 723 -2444 757 -2294
rect 800 -2386 810 -2334
rect 862 -2386 872 -2334
rect 915 -2444 949 -2294
rect 992 -2386 1002 -2334
rect 1054 -2386 1064 -2334
rect 1107 -2444 1141 -2294
rect 1184 -2386 1194 -2334
rect 1246 -2386 1256 -2334
rect 1299 -2444 1333 -2294
rect 1376 -2386 1386 -2334
rect 1438 -2386 1448 -2334
rect 1503 -2382 1509 -1996
rect 1543 -2382 1549 -1996
rect 251 -2478 1333 -2444
rect -1250 -2543 -1240 -2491
rect -1188 -2543 -412 -2491
rect -360 -2543 -350 -2491
rect 1503 -2558 1549 -2382
rect 1643 -2386 1670 -2334
rect 1722 -2386 1732 -2334
rect 1772 -2444 1806 -1881
rect 1956 -1847 1990 -1714
rect 2148 -1847 2182 -1714
rect 2340 -1847 2374 -1714
rect 2532 -1847 2566 -1714
rect 2724 -1847 2758 -1714
rect 2916 -1847 2950 -1714
rect 3024 -1732 3030 -1532
rect 3064 -1732 3070 -1532
rect 3024 -1744 3070 -1732
rect 3273 -1847 3307 -547
rect 1956 -1881 3307 -1847
rect 1956 -2022 1990 -1881
rect 2148 -2022 2182 -1881
rect 2340 -2022 2374 -1881
rect 2532 -2022 2566 -1881
rect 2724 -2022 2758 -1881
rect 2916 -2022 2950 -1881
rect 3024 -1996 3070 -1984
rect 1950 -2034 1996 -2022
rect 1950 -2282 1956 -2034
rect 1990 -2282 1996 -2034
rect 1950 -2294 1996 -2282
rect 2046 -2034 2092 -2022
rect 2046 -2282 2052 -2034
rect 2086 -2282 2092 -2034
rect 2046 -2294 2092 -2282
rect 2142 -2034 2188 -2022
rect 2142 -2282 2148 -2034
rect 2182 -2282 2188 -2034
rect 2142 -2294 2188 -2282
rect 2238 -2034 2284 -2022
rect 2238 -2282 2244 -2034
rect 2278 -2282 2284 -2034
rect 2238 -2294 2284 -2282
rect 2334 -2034 2380 -2022
rect 2334 -2282 2340 -2034
rect 2374 -2282 2380 -2034
rect 2334 -2294 2380 -2282
rect 2430 -2034 2476 -2022
rect 2430 -2282 2436 -2034
rect 2470 -2282 2476 -2034
rect 2430 -2294 2476 -2282
rect 2526 -2034 2572 -2022
rect 2526 -2282 2532 -2034
rect 2566 -2282 2572 -2034
rect 2526 -2294 2572 -2282
rect 2622 -2034 2668 -2022
rect 2622 -2282 2628 -2034
rect 2662 -2282 2668 -2034
rect 2622 -2294 2668 -2282
rect 2718 -2034 2764 -2022
rect 2718 -2282 2724 -2034
rect 2758 -2282 2764 -2034
rect 2718 -2294 2764 -2282
rect 2814 -2034 2860 -2022
rect 2814 -2282 2820 -2034
rect 2854 -2282 2860 -2034
rect 2814 -2294 2860 -2282
rect 2910 -2034 2956 -2022
rect 2910 -2282 2916 -2034
rect 2950 -2282 2956 -2034
rect 2910 -2294 2956 -2282
rect 1937 -2386 1947 -2334
rect 1999 -2386 2009 -2334
rect 2052 -2444 2086 -2294
rect 2130 -2386 2140 -2334
rect 2192 -2386 2202 -2334
rect 2244 -2444 2278 -2294
rect 2321 -2386 2331 -2334
rect 2383 -2386 2393 -2334
rect 2436 -2444 2470 -2294
rect 2513 -2386 2523 -2334
rect 2575 -2386 2585 -2334
rect 2628 -2444 2662 -2294
rect 2705 -2386 2715 -2334
rect 2767 -2386 2777 -2334
rect 2820 -2444 2854 -2294
rect 2897 -2386 2907 -2334
rect 2959 -2386 2969 -2334
rect 3024 -2382 3030 -1996
rect 3064 -2382 3070 -1996
rect 1772 -2478 2854 -2444
rect 3024 -2558 3070 -2382
rect -1326 -2636 -336 -2605
rect -1326 -2670 -1227 -2636
rect -1193 -2670 -1135 -2636
rect -1101 -2670 -1043 -2636
rect -1009 -2670 -951 -2636
rect -917 -2670 -859 -2636
rect -825 -2670 -767 -2636
rect -733 -2670 -675 -2636
rect -641 -2670 -583 -2636
rect -549 -2670 -491 -2636
rect -457 -2670 -399 -2636
rect -365 -2670 -336 -2636
rect -1326 -2701 -336 -2670
rect 3273 -2626 3307 -1881
rect 3273 -2660 3456 -2626
rect -3300 -2848 -2218 -2814
rect -3429 -2958 -3402 -2906
rect -3350 -2958 -3340 -2906
rect -3300 -3411 -3266 -2848
rect -3135 -2958 -3125 -2906
rect -3073 -2958 -3063 -2906
rect -3020 -2998 -2986 -2848
rect -2942 -2958 -2932 -2906
rect -2880 -2958 -2870 -2906
rect -2828 -2998 -2794 -2848
rect -2751 -2958 -2741 -2906
rect -2689 -2958 -2679 -2906
rect -2636 -2998 -2602 -2848
rect -2559 -2958 -2549 -2906
rect -2497 -2958 -2487 -2906
rect -2444 -2998 -2410 -2848
rect -2367 -2958 -2357 -2906
rect -2305 -2958 -2295 -2906
rect -2252 -2998 -2218 -2848
rect -2175 -2958 -2165 -2906
rect -2113 -2958 -2103 -2906
rect -2048 -2910 -2002 -2778
rect -772 -2827 -762 -2775
rect -710 -2827 -412 -2775
rect -360 -2827 -350 -2775
rect 251 -2848 1333 -2814
rect -3122 -3010 -3076 -2998
rect -3122 -3258 -3116 -3010
rect -3082 -3258 -3076 -3010
rect -3122 -3270 -3076 -3258
rect -3026 -3010 -2980 -2998
rect -3026 -3258 -3020 -3010
rect -2986 -3258 -2980 -3010
rect -3026 -3270 -2980 -3258
rect -2930 -3010 -2884 -2998
rect -2930 -3258 -2924 -3010
rect -2890 -3258 -2884 -3010
rect -2930 -3270 -2884 -3258
rect -2834 -3010 -2788 -2998
rect -2834 -3258 -2828 -3010
rect -2794 -3258 -2788 -3010
rect -2834 -3270 -2788 -3258
rect -2738 -3010 -2692 -2998
rect -2738 -3258 -2732 -3010
rect -2698 -3258 -2692 -3010
rect -2738 -3270 -2692 -3258
rect -2642 -3010 -2596 -2998
rect -2642 -3258 -2636 -3010
rect -2602 -3258 -2596 -3010
rect -2642 -3270 -2596 -3258
rect -2546 -3010 -2500 -2998
rect -2546 -3258 -2540 -3010
rect -2506 -3258 -2500 -3010
rect -2546 -3270 -2500 -3258
rect -2450 -3010 -2404 -2998
rect -2450 -3258 -2444 -3010
rect -2410 -3258 -2404 -3010
rect -2450 -3270 -2404 -3258
rect -2354 -3010 -2308 -2998
rect -2354 -3258 -2348 -3010
rect -2314 -3258 -2308 -3010
rect -2354 -3270 -2308 -3258
rect -2258 -3010 -2212 -2998
rect -2258 -3258 -2252 -3010
rect -2218 -3258 -2212 -3010
rect -2258 -3270 -2212 -3258
rect -2162 -3010 -2116 -2998
rect -2162 -3258 -2156 -3010
rect -2122 -3258 -2116 -3010
rect -2162 -3270 -2116 -3258
rect -3690 -3445 -3266 -3411
rect -3429 -3765 -3402 -3713
rect -3350 -3765 -3340 -3713
rect -3300 -3822 -3266 -3445
rect -3116 -3411 -3082 -3270
rect -2924 -3411 -2890 -3270
rect -2732 -3411 -2698 -3270
rect -2540 -3411 -2506 -3270
rect -2348 -3411 -2314 -3270
rect -2156 -3411 -2122 -3270
rect -2048 -3296 -2042 -2910
rect -2008 -3296 -2002 -2910
rect -1936 -2958 -1926 -2906
rect -1874 -2958 -1416 -2906
rect -1364 -2958 -1354 -2906
rect -1108 -2917 -1098 -2865
rect -1046 -2917 -1036 -2865
rect -1002 -2868 -872 -2864
rect -1006 -2874 -872 -2868
rect -1006 -2908 -994 -2874
rect -960 -2908 -872 -2874
rect -1006 -2914 -872 -2908
rect -1002 -2916 -872 -2914
rect -820 -2874 -527 -2864
rect -820 -2908 -574 -2874
rect -540 -2908 -527 -2874
rect -820 -2916 -527 -2908
rect -1002 -2918 -527 -2916
rect -422 -2918 -412 -2866
rect -360 -2918 -350 -2866
rect 70 -2957 149 -2905
rect 201 -2957 211 -2905
rect -246 -3030 -236 -3026
rect -502 -3036 -236 -3030
rect -502 -3070 -490 -3036
rect -456 -3070 -236 -3036
rect -502 -3076 -236 -3070
rect -246 -3078 -236 -3076
rect -184 -3078 -174 -3026
rect -1326 -3180 -336 -3149
rect -1326 -3214 -1227 -3180
rect -1193 -3214 -1135 -3180
rect -1101 -3214 -1043 -3180
rect -1009 -3214 -951 -3180
rect -917 -3214 -859 -3180
rect -825 -3214 -767 -3180
rect -733 -3214 -675 -3180
rect -641 -3214 -583 -3180
rect -549 -3214 -491 -3180
rect -457 -3214 -399 -3180
rect -365 -3214 -336 -3180
rect -1326 -3245 -336 -3214
rect 251 -3225 285 -2848
rect 419 -2905 485 -2900
rect 416 -2957 426 -2905
rect 478 -2957 488 -2905
rect 419 -2960 485 -2957
rect 531 -2988 565 -2848
rect 611 -2905 677 -2900
rect 607 -2957 617 -2905
rect 669 -2957 679 -2905
rect 611 -2960 677 -2957
rect 723 -2988 757 -2848
rect 803 -2905 869 -2900
rect 799 -2957 809 -2905
rect 861 -2957 871 -2905
rect 803 -2960 869 -2957
rect 915 -2988 949 -2848
rect 995 -2905 1061 -2900
rect 991 -2957 1001 -2905
rect 1053 -2957 1063 -2905
rect 995 -2960 1061 -2957
rect 1107 -2988 1141 -2848
rect 1187 -2904 1253 -2900
rect 1184 -2956 1194 -2904
rect 1246 -2956 1256 -2904
rect 1187 -2960 1253 -2956
rect 1299 -2988 1333 -2848
rect 1379 -2904 1445 -2900
rect 1376 -2956 1386 -2904
rect 1438 -2956 1448 -2904
rect 1503 -2910 1549 -2738
rect 1772 -2848 2854 -2814
rect 1379 -2960 1445 -2956
rect 429 -3000 475 -2988
rect 429 -3080 435 -3000
rect 469 -3080 475 -3000
rect 429 -3092 475 -3080
rect 525 -3000 571 -2988
rect 525 -3080 531 -3000
rect 565 -3080 571 -3000
rect 525 -3092 571 -3080
rect 621 -3000 667 -2988
rect 621 -3080 627 -3000
rect 661 -3080 667 -3000
rect 621 -3092 667 -3080
rect 717 -3000 763 -2988
rect 717 -3080 723 -3000
rect 757 -3080 763 -3000
rect 717 -3092 763 -3080
rect 813 -3000 859 -2988
rect 813 -3080 819 -3000
rect 853 -3080 859 -3000
rect 813 -3092 859 -3080
rect 909 -3000 955 -2988
rect 909 -3080 915 -3000
rect 949 -3080 955 -3000
rect 909 -3092 955 -3080
rect 1005 -3000 1051 -2988
rect 1005 -3080 1011 -3000
rect 1045 -3080 1051 -3000
rect 1005 -3092 1051 -3080
rect 1101 -3000 1147 -2988
rect 1101 -3080 1107 -3000
rect 1141 -3080 1147 -3000
rect 1101 -3092 1147 -3080
rect 1197 -3000 1243 -2988
rect 1197 -3080 1203 -3000
rect 1237 -3080 1243 -3000
rect 1197 -3092 1243 -3080
rect 1293 -3000 1339 -2988
rect 1293 -3080 1299 -3000
rect 1333 -3080 1339 -3000
rect 1293 -3092 1339 -3080
rect 1389 -3000 1435 -2988
rect 1389 -3080 1395 -3000
rect 1429 -3080 1435 -3000
rect 1389 -3092 1435 -3080
rect -2048 -3308 -2002 -3296
rect -44 -3259 285 -3225
rect -44 -3308 -10 -3259
rect -1812 -3342 -10 -3308
rect -1812 -3411 -1778 -3342
rect -3116 -3445 -1778 -3411
rect -773 -3445 -762 -3393
rect -710 -3445 -414 -3393
rect -362 -3445 -352 -3393
rect -3116 -3578 -3082 -3445
rect -2924 -3578 -2890 -3445
rect -2732 -3578 -2698 -3445
rect -2540 -3578 -2506 -3445
rect -2348 -3578 -2314 -3445
rect -2156 -3578 -2122 -3445
rect -1251 -3539 -1241 -3485
rect -1187 -3492 -528 -3485
rect -1187 -3526 -576 -3492
rect -542 -3526 -528 -3492
rect -424 -3526 -414 -3474
rect -362 -3526 -352 -3474
rect -1187 -3539 -528 -3526
rect -417 -3527 -359 -3526
rect -2048 -3560 -2002 -3548
rect -3122 -3590 -3076 -3578
rect -3122 -3670 -3116 -3590
rect -3082 -3670 -3076 -3590
rect -3122 -3682 -3076 -3670
rect -3026 -3590 -2980 -3578
rect -3026 -3670 -3020 -3590
rect -2986 -3670 -2980 -3590
rect -3026 -3682 -2980 -3670
rect -2930 -3590 -2884 -3578
rect -2930 -3670 -2924 -3590
rect -2890 -3670 -2884 -3590
rect -2930 -3682 -2884 -3670
rect -2834 -3590 -2788 -3578
rect -2834 -3670 -2828 -3590
rect -2794 -3670 -2788 -3590
rect -2834 -3682 -2788 -3670
rect -2738 -3590 -2692 -3578
rect -2738 -3670 -2732 -3590
rect -2698 -3670 -2692 -3590
rect -2738 -3682 -2692 -3670
rect -2642 -3590 -2596 -3578
rect -2642 -3670 -2636 -3590
rect -2602 -3670 -2596 -3590
rect -2642 -3682 -2596 -3670
rect -2546 -3590 -2500 -3578
rect -2546 -3670 -2540 -3590
rect -2506 -3670 -2500 -3590
rect -2546 -3682 -2500 -3670
rect -2450 -3590 -2404 -3578
rect -2450 -3670 -2444 -3590
rect -2410 -3670 -2404 -3590
rect -2450 -3682 -2404 -3670
rect -2354 -3590 -2308 -3578
rect -2354 -3670 -2348 -3590
rect -2314 -3670 -2308 -3590
rect -2354 -3682 -2308 -3670
rect -2258 -3590 -2212 -3578
rect -2258 -3670 -2252 -3590
rect -2218 -3670 -2212 -3590
rect -2258 -3682 -2212 -3670
rect -2162 -3590 -2116 -3578
rect -2162 -3670 -2156 -3590
rect -2122 -3670 -2116 -3590
rect -2162 -3682 -2116 -3670
rect -3132 -3713 -3066 -3710
rect -3135 -3765 -3125 -3713
rect -3073 -3765 -3063 -3713
rect -3132 -3770 -3066 -3765
rect -3020 -3822 -2986 -3682
rect -2940 -3713 -2874 -3710
rect -2944 -3765 -2934 -3713
rect -2882 -3765 -2872 -3713
rect -2940 -3770 -2874 -3765
rect -2828 -3822 -2794 -3682
rect -2748 -3713 -2682 -3710
rect -2752 -3765 -2742 -3713
rect -2690 -3765 -2680 -3713
rect -2748 -3770 -2682 -3765
rect -2636 -3822 -2602 -3682
rect -2556 -3713 -2490 -3710
rect -2560 -3765 -2550 -3713
rect -2498 -3765 -2488 -3713
rect -2556 -3770 -2490 -3765
rect -2444 -3822 -2410 -3682
rect -2364 -3714 -2298 -3710
rect -2367 -3766 -2357 -3714
rect -2305 -3766 -2295 -3714
rect -2364 -3770 -2298 -3766
rect -2252 -3822 -2218 -3682
rect -2172 -3714 -2106 -3710
rect -2175 -3766 -2165 -3714
rect -2113 -3766 -2103 -3714
rect -2048 -3760 -2042 -3560
rect -2008 -3760 -2002 -3560
rect -510 -3632 -500 -3580
rect -448 -3632 -438 -3580
rect -2172 -3770 -2106 -3766
rect -3300 -3856 -2218 -3822
rect -2048 -3892 -2002 -3760
rect -783 -3724 -336 -3693
rect -783 -3758 -675 -3724
rect -641 -3758 -583 -3724
rect -549 -3758 -491 -3724
rect -457 -3758 -399 -3724
rect -365 -3758 -336 -3724
rect -783 -3789 -336 -3758
rect -245 -3764 -235 -3712
rect -183 -3764 149 -3712
rect 201 -3764 211 -3712
rect 251 -3822 285 -3259
rect 435 -3225 469 -3092
rect 627 -3225 661 -3092
rect 819 -3225 853 -3092
rect 1011 -3225 1045 -3092
rect 1203 -3225 1237 -3092
rect 1395 -3225 1429 -3092
rect 1503 -3110 1509 -2910
rect 1543 -2997 1549 -2910
rect 1643 -2957 1670 -2905
rect 1722 -2957 1732 -2905
rect 1610 -2997 1656 -2996
rect 1543 -3008 1656 -2997
rect 1543 -3084 1616 -3008
rect 1650 -3084 1656 -3008
rect 1543 -3096 1656 -3084
rect 1698 -2997 1744 -2996
rect 1772 -2997 1806 -2848
rect 1940 -2905 2006 -2900
rect 1937 -2957 1947 -2905
rect 1999 -2957 2009 -2905
rect 1940 -2960 2006 -2957
rect 2052 -2988 2086 -2848
rect 2132 -2905 2198 -2900
rect 2128 -2957 2138 -2905
rect 2190 -2957 2200 -2905
rect 2132 -2960 2198 -2957
rect 2244 -2988 2278 -2848
rect 2324 -2905 2390 -2900
rect 2320 -2957 2330 -2905
rect 2382 -2957 2392 -2905
rect 2324 -2960 2390 -2957
rect 2436 -2988 2470 -2848
rect 2516 -2905 2582 -2900
rect 2512 -2957 2522 -2905
rect 2574 -2957 2584 -2905
rect 2516 -2960 2582 -2957
rect 2628 -2988 2662 -2848
rect 2708 -2904 2774 -2900
rect 2705 -2956 2715 -2904
rect 2767 -2956 2777 -2904
rect 2708 -2960 2774 -2956
rect 2820 -2988 2854 -2848
rect 2900 -2904 2966 -2900
rect 2897 -2956 2907 -2904
rect 2959 -2956 2969 -2904
rect 3024 -2910 3070 -2738
rect 2900 -2960 2966 -2956
rect 1698 -3008 1806 -2997
rect 1698 -3084 1704 -3008
rect 1738 -3084 1806 -3008
rect 1698 -3096 1806 -3084
rect 1950 -3000 1996 -2988
rect 1950 -3080 1956 -3000
rect 1990 -3080 1996 -3000
rect 1950 -3092 1996 -3080
rect 2046 -3000 2092 -2988
rect 2046 -3080 2052 -3000
rect 2086 -3080 2092 -3000
rect 2046 -3092 2092 -3080
rect 2142 -3000 2188 -2988
rect 2142 -3080 2148 -3000
rect 2182 -3080 2188 -3000
rect 2142 -3092 2188 -3080
rect 2238 -3000 2284 -2988
rect 2238 -3080 2244 -3000
rect 2278 -3080 2284 -3000
rect 2238 -3092 2284 -3080
rect 2334 -3000 2380 -2988
rect 2334 -3080 2340 -3000
rect 2374 -3080 2380 -3000
rect 2334 -3092 2380 -3080
rect 2430 -3000 2476 -2988
rect 2430 -3080 2436 -3000
rect 2470 -3080 2476 -3000
rect 2430 -3092 2476 -3080
rect 2526 -3000 2572 -2988
rect 2526 -3080 2532 -3000
rect 2566 -3080 2572 -3000
rect 2526 -3092 2572 -3080
rect 2622 -3000 2668 -2988
rect 2622 -3080 2628 -3000
rect 2662 -3080 2668 -3000
rect 2622 -3092 2668 -3080
rect 2718 -3000 2764 -2988
rect 2718 -3080 2724 -3000
rect 2758 -3080 2764 -3000
rect 2718 -3092 2764 -3080
rect 2814 -3000 2860 -2988
rect 2814 -3080 2820 -3000
rect 2854 -3080 2860 -3000
rect 2814 -3092 2860 -3080
rect 2910 -3000 2956 -2988
rect 2910 -3080 2916 -3000
rect 2950 -3080 2956 -3000
rect 2910 -3092 2956 -3080
rect 1543 -3097 1649 -3096
rect 1703 -3097 1806 -3096
rect 1543 -3110 1549 -3097
rect 1503 -3122 1549 -3110
rect 1648 -3134 1706 -3128
rect 1648 -3135 1660 -3134
rect 1694 -3135 1706 -3134
rect 1640 -3187 1650 -3135
rect 1702 -3187 1712 -3135
rect 1772 -3225 1806 -3097
rect 435 -3259 1806 -3225
rect 435 -3400 469 -3259
rect 627 -3400 661 -3259
rect 819 -3400 853 -3259
rect 1011 -3400 1045 -3259
rect 1203 -3400 1237 -3259
rect 1395 -3400 1429 -3259
rect 1503 -3374 1549 -3362
rect 429 -3412 475 -3400
rect 429 -3660 435 -3412
rect 469 -3660 475 -3412
rect 429 -3672 475 -3660
rect 525 -3412 571 -3400
rect 525 -3660 531 -3412
rect 565 -3660 571 -3412
rect 525 -3672 571 -3660
rect 621 -3412 667 -3400
rect 621 -3660 627 -3412
rect 661 -3660 667 -3412
rect 621 -3672 667 -3660
rect 717 -3412 763 -3400
rect 717 -3660 723 -3412
rect 757 -3660 763 -3412
rect 717 -3672 763 -3660
rect 813 -3412 859 -3400
rect 813 -3660 819 -3412
rect 853 -3660 859 -3412
rect 813 -3672 859 -3660
rect 909 -3412 955 -3400
rect 909 -3660 915 -3412
rect 949 -3660 955 -3412
rect 909 -3672 955 -3660
rect 1005 -3412 1051 -3400
rect 1005 -3660 1011 -3412
rect 1045 -3660 1051 -3412
rect 1005 -3672 1051 -3660
rect 1101 -3412 1147 -3400
rect 1101 -3660 1107 -3412
rect 1141 -3660 1147 -3412
rect 1101 -3672 1147 -3660
rect 1197 -3412 1243 -3400
rect 1197 -3660 1203 -3412
rect 1237 -3660 1243 -3412
rect 1197 -3672 1243 -3660
rect 1293 -3412 1339 -3400
rect 1293 -3660 1299 -3412
rect 1333 -3660 1339 -3412
rect 1293 -3672 1339 -3660
rect 1389 -3412 1435 -3400
rect 1389 -3660 1395 -3412
rect 1429 -3660 1435 -3412
rect 1389 -3672 1435 -3660
rect 416 -3764 426 -3712
rect 478 -3764 488 -3712
rect 531 -3822 565 -3672
rect 609 -3764 619 -3712
rect 671 -3764 681 -3712
rect 723 -3822 757 -3672
rect 800 -3764 810 -3712
rect 862 -3764 872 -3712
rect 915 -3822 949 -3672
rect 992 -3764 1002 -3712
rect 1054 -3764 1064 -3712
rect 1107 -3822 1141 -3672
rect 1184 -3764 1194 -3712
rect 1246 -3764 1256 -3712
rect 1299 -3822 1333 -3672
rect 1376 -3764 1386 -3712
rect 1438 -3764 1448 -3712
rect 1503 -3760 1509 -3374
rect 1543 -3760 1549 -3374
rect 251 -3856 1333 -3822
rect 1503 -3936 1549 -3760
rect 1643 -3764 1670 -3712
rect 1722 -3764 1732 -3712
rect 1772 -3822 1806 -3259
rect 1956 -3225 1990 -3092
rect 2148 -3225 2182 -3092
rect 2340 -3225 2374 -3092
rect 2532 -3225 2566 -3092
rect 2724 -3225 2758 -3092
rect 2916 -3225 2950 -3092
rect 3024 -3110 3030 -2910
rect 3064 -3110 3070 -2910
rect 3024 -3122 3070 -3110
rect 3273 -3225 3307 -2660
rect 1956 -3259 3307 -3225
rect 1956 -3400 1990 -3259
rect 2148 -3400 2182 -3259
rect 2340 -3400 2374 -3259
rect 2532 -3400 2566 -3259
rect 2724 -3400 2758 -3259
rect 2916 -3400 2950 -3259
rect 3024 -3374 3070 -3362
rect 1950 -3412 1996 -3400
rect 1950 -3660 1956 -3412
rect 1990 -3660 1996 -3412
rect 1950 -3672 1996 -3660
rect 2046 -3412 2092 -3400
rect 2046 -3660 2052 -3412
rect 2086 -3660 2092 -3412
rect 2046 -3672 2092 -3660
rect 2142 -3412 2188 -3400
rect 2142 -3660 2148 -3412
rect 2182 -3660 2188 -3412
rect 2142 -3672 2188 -3660
rect 2238 -3412 2284 -3400
rect 2238 -3660 2244 -3412
rect 2278 -3660 2284 -3412
rect 2238 -3672 2284 -3660
rect 2334 -3412 2380 -3400
rect 2334 -3660 2340 -3412
rect 2374 -3660 2380 -3412
rect 2334 -3672 2380 -3660
rect 2430 -3412 2476 -3400
rect 2430 -3660 2436 -3412
rect 2470 -3660 2476 -3412
rect 2430 -3672 2476 -3660
rect 2526 -3412 2572 -3400
rect 2526 -3660 2532 -3412
rect 2566 -3660 2572 -3412
rect 2526 -3672 2572 -3660
rect 2622 -3412 2668 -3400
rect 2622 -3660 2628 -3412
rect 2662 -3660 2668 -3412
rect 2622 -3672 2668 -3660
rect 2718 -3412 2764 -3400
rect 2718 -3660 2724 -3412
rect 2758 -3660 2764 -3412
rect 2718 -3672 2764 -3660
rect 2814 -3412 2860 -3400
rect 2814 -3660 2820 -3412
rect 2854 -3660 2860 -3412
rect 2814 -3672 2860 -3660
rect 2910 -3412 2956 -3400
rect 2910 -3660 2916 -3412
rect 2950 -3660 2956 -3412
rect 2910 -3672 2956 -3660
rect 1937 -3764 1947 -3712
rect 1999 -3764 2009 -3712
rect 2052 -3822 2086 -3672
rect 2130 -3764 2140 -3712
rect 2192 -3764 2202 -3712
rect 2244 -3822 2278 -3672
rect 2321 -3764 2331 -3712
rect 2383 -3764 2393 -3712
rect 2436 -3822 2470 -3672
rect 2513 -3764 2523 -3712
rect 2575 -3764 2585 -3712
rect 2628 -3822 2662 -3672
rect 2705 -3764 2715 -3712
rect 2767 -3764 2777 -3712
rect 2820 -3822 2854 -3672
rect 2897 -3764 2907 -3712
rect 2959 -3764 2969 -3712
rect 3024 -3760 3030 -3374
rect 3064 -3760 3070 -3374
rect 1772 -3856 2854 -3822
rect 3024 -3935 3070 -3760
rect -579 -3961 -236 -3951
rect -579 -3995 -539 -3961
rect -505 -3995 -236 -3961
rect -579 -4003 -236 -3995
rect -184 -4003 -173 -3951
rect -91 -4114 -81 -4111
rect -465 -4120 -81 -4114
rect -465 -4154 -453 -4120
rect -419 -4154 -81 -4120
rect -3300 -4226 -2218 -4192
rect -3429 -4336 -3402 -4284
rect -3350 -4336 -3340 -4284
rect -3300 -4789 -3266 -4226
rect -3135 -4336 -3125 -4284
rect -3073 -4336 -3063 -4284
rect -3020 -4376 -2986 -4226
rect -2942 -4336 -2932 -4284
rect -2880 -4336 -2870 -4284
rect -2828 -4376 -2794 -4226
rect -2751 -4336 -2741 -4284
rect -2689 -4336 -2679 -4284
rect -2636 -4376 -2602 -4226
rect -2559 -4336 -2549 -4284
rect -2497 -4336 -2487 -4284
rect -2444 -4376 -2410 -4226
rect -2367 -4336 -2357 -4284
rect -2305 -4336 -2295 -4284
rect -2252 -4376 -2218 -4226
rect -2175 -4336 -2165 -4284
rect -2113 -4336 -2103 -4284
rect -2048 -4288 -2002 -4156
rect -465 -4160 -81 -4154
rect -91 -4163 -81 -4160
rect -29 -4163 -19 -4111
rect 251 -4226 1333 -4192
rect -784 -4268 -336 -4237
rect -3122 -4388 -3076 -4376
rect -3122 -4636 -3116 -4388
rect -3082 -4636 -3076 -4388
rect -3122 -4648 -3076 -4636
rect -3026 -4388 -2980 -4376
rect -3026 -4636 -3020 -4388
rect -2986 -4636 -2980 -4388
rect -3026 -4648 -2980 -4636
rect -2930 -4388 -2884 -4376
rect -2930 -4636 -2924 -4388
rect -2890 -4636 -2884 -4388
rect -2930 -4648 -2884 -4636
rect -2834 -4388 -2788 -4376
rect -2834 -4636 -2828 -4388
rect -2794 -4636 -2788 -4388
rect -2834 -4648 -2788 -4636
rect -2738 -4388 -2692 -4376
rect -2738 -4636 -2732 -4388
rect -2698 -4636 -2692 -4388
rect -2738 -4648 -2692 -4636
rect -2642 -4388 -2596 -4376
rect -2642 -4636 -2636 -4388
rect -2602 -4636 -2596 -4388
rect -2642 -4648 -2596 -4636
rect -2546 -4388 -2500 -4376
rect -2546 -4636 -2540 -4388
rect -2506 -4636 -2500 -4388
rect -2546 -4648 -2500 -4636
rect -2450 -4388 -2404 -4376
rect -2450 -4636 -2444 -4388
rect -2410 -4636 -2404 -4388
rect -2450 -4648 -2404 -4636
rect -2354 -4388 -2308 -4376
rect -2354 -4636 -2348 -4388
rect -2314 -4636 -2308 -4388
rect -2354 -4648 -2308 -4636
rect -2258 -4388 -2212 -4376
rect -2258 -4636 -2252 -4388
rect -2218 -4636 -2212 -4388
rect -2258 -4648 -2212 -4636
rect -2162 -4388 -2116 -4376
rect -2162 -4636 -2156 -4388
rect -2122 -4636 -2116 -4388
rect -2162 -4648 -2116 -4636
rect -3690 -4823 -3266 -4789
rect -3429 -5143 -3402 -5091
rect -3350 -5143 -3340 -5091
rect -3300 -5200 -3266 -4823
rect -3116 -4789 -3082 -4648
rect -2924 -4789 -2890 -4648
rect -2732 -4789 -2698 -4648
rect -2540 -4789 -2506 -4648
rect -2348 -4789 -2314 -4648
rect -2156 -4789 -2122 -4648
rect -2048 -4674 -2042 -4288
rect -2008 -4674 -2002 -4288
rect -1953 -4336 -1943 -4284
rect -1891 -4336 -1416 -4284
rect -1364 -4336 -1354 -4284
rect -784 -4302 -675 -4268
rect -641 -4302 -583 -4268
rect -549 -4302 -491 -4268
rect -457 -4302 -399 -4268
rect -365 -4302 -336 -4268
rect -784 -4333 -336 -4302
rect 70 -4335 149 -4283
rect 201 -4335 211 -4283
rect 82 -4412 92 -4409
rect -464 -4418 92 -4412
rect -464 -4452 -452 -4418
rect -418 -4452 92 -4418
rect -464 -4458 92 -4452
rect 82 -4461 92 -4458
rect 144 -4461 154 -4409
rect -558 -4617 -548 -4565
rect -496 -4617 -486 -4565
rect 251 -4603 285 -4226
rect 419 -4283 485 -4278
rect 416 -4335 426 -4283
rect 478 -4335 488 -4283
rect 419 -4338 485 -4335
rect 531 -4366 565 -4226
rect 611 -4283 677 -4278
rect 607 -4335 617 -4283
rect 669 -4335 679 -4283
rect 611 -4338 677 -4335
rect 723 -4366 757 -4226
rect 803 -4283 869 -4278
rect 799 -4335 809 -4283
rect 861 -4335 871 -4283
rect 803 -4338 869 -4335
rect 915 -4366 949 -4226
rect 995 -4283 1061 -4278
rect 991 -4335 1001 -4283
rect 1053 -4335 1063 -4283
rect 995 -4338 1061 -4335
rect 1107 -4366 1141 -4226
rect 1187 -4282 1253 -4278
rect 1184 -4334 1194 -4282
rect 1246 -4334 1256 -4282
rect 1187 -4338 1253 -4334
rect 1299 -4366 1333 -4226
rect 1379 -4282 1445 -4278
rect 1376 -4334 1386 -4282
rect 1438 -4334 1448 -4282
rect 1503 -4288 1549 -4115
rect 1772 -4226 2854 -4192
rect 1379 -4338 1445 -4334
rect 429 -4378 475 -4366
rect 429 -4458 435 -4378
rect 469 -4458 475 -4378
rect 429 -4470 475 -4458
rect 525 -4378 571 -4366
rect 525 -4458 531 -4378
rect 565 -4458 571 -4378
rect 525 -4470 571 -4458
rect 621 -4378 667 -4366
rect 621 -4458 627 -4378
rect 661 -4458 667 -4378
rect 621 -4470 667 -4458
rect 717 -4378 763 -4366
rect 717 -4458 723 -4378
rect 757 -4458 763 -4378
rect 717 -4470 763 -4458
rect 813 -4378 859 -4366
rect 813 -4458 819 -4378
rect 853 -4458 859 -4378
rect 813 -4470 859 -4458
rect 909 -4378 955 -4366
rect 909 -4458 915 -4378
rect 949 -4458 955 -4378
rect 909 -4470 955 -4458
rect 1005 -4378 1051 -4366
rect 1005 -4458 1011 -4378
rect 1045 -4458 1051 -4378
rect 1005 -4470 1051 -4458
rect 1101 -4378 1147 -4366
rect 1101 -4458 1107 -4378
rect 1141 -4458 1147 -4378
rect 1101 -4470 1147 -4458
rect 1197 -4378 1243 -4366
rect 1197 -4458 1203 -4378
rect 1237 -4458 1243 -4378
rect 1197 -4470 1243 -4458
rect 1293 -4378 1339 -4366
rect 1293 -4458 1299 -4378
rect 1333 -4458 1339 -4378
rect 1293 -4470 1339 -4458
rect 1389 -4378 1435 -4366
rect 1389 -4458 1395 -4378
rect 1429 -4458 1435 -4378
rect 1389 -4470 1435 -4458
rect -48 -4637 285 -4603
rect -48 -4674 -14 -4637
rect -2048 -4686 -2002 -4674
rect -1808 -4708 -14 -4674
rect -1808 -4789 -1774 -4708
rect -3116 -4823 -1774 -4789
rect -774 -4812 -336 -4781
rect -3116 -4956 -3082 -4823
rect -2924 -4956 -2890 -4823
rect -2732 -4956 -2698 -4823
rect -2540 -4956 -2506 -4823
rect -2348 -4956 -2314 -4823
rect -2156 -4956 -2122 -4823
rect -774 -4846 -675 -4812
rect -641 -4846 -583 -4812
rect -549 -4846 -491 -4812
rect -457 -4846 -399 -4812
rect -365 -4846 -336 -4812
rect -774 -4877 -336 -4846
rect -2048 -4938 -2002 -4926
rect -3122 -4968 -3076 -4956
rect -3122 -5048 -3116 -4968
rect -3082 -5048 -3076 -4968
rect -3122 -5060 -3076 -5048
rect -3026 -4968 -2980 -4956
rect -3026 -5048 -3020 -4968
rect -2986 -5048 -2980 -4968
rect -3026 -5060 -2980 -5048
rect -2930 -4968 -2884 -4956
rect -2930 -5048 -2924 -4968
rect -2890 -5048 -2884 -4968
rect -2930 -5060 -2884 -5048
rect -2834 -4968 -2788 -4956
rect -2834 -5048 -2828 -4968
rect -2794 -5048 -2788 -4968
rect -2834 -5060 -2788 -5048
rect -2738 -4968 -2692 -4956
rect -2738 -5048 -2732 -4968
rect -2698 -5048 -2692 -4968
rect -2738 -5060 -2692 -5048
rect -2642 -4968 -2596 -4956
rect -2642 -5048 -2636 -4968
rect -2602 -5048 -2596 -4968
rect -2642 -5060 -2596 -5048
rect -2546 -4968 -2500 -4956
rect -2546 -5048 -2540 -4968
rect -2506 -5048 -2500 -4968
rect -2546 -5060 -2500 -5048
rect -2450 -4968 -2404 -4956
rect -2450 -5048 -2444 -4968
rect -2410 -5048 -2404 -4968
rect -2450 -5060 -2404 -5048
rect -2354 -4968 -2308 -4956
rect -2354 -5048 -2348 -4968
rect -2314 -5048 -2308 -4968
rect -2354 -5060 -2308 -5048
rect -2258 -4968 -2212 -4956
rect -2258 -5048 -2252 -4968
rect -2218 -5048 -2212 -4968
rect -2258 -5060 -2212 -5048
rect -2162 -4968 -2116 -4956
rect -2162 -5048 -2156 -4968
rect -2122 -5048 -2116 -4968
rect -2162 -5060 -2116 -5048
rect -3132 -5091 -3066 -5088
rect -3135 -5143 -3125 -5091
rect -3073 -5143 -3063 -5091
rect -3132 -5148 -3066 -5143
rect -3020 -5200 -2986 -5060
rect -2940 -5091 -2874 -5088
rect -2944 -5143 -2934 -5091
rect -2882 -5143 -2872 -5091
rect -2940 -5148 -2874 -5143
rect -2828 -5200 -2794 -5060
rect -2748 -5091 -2682 -5088
rect -2752 -5143 -2742 -5091
rect -2690 -5143 -2680 -5091
rect -2748 -5148 -2682 -5143
rect -2636 -5200 -2602 -5060
rect -2556 -5091 -2490 -5088
rect -2560 -5143 -2550 -5091
rect -2498 -5143 -2488 -5091
rect -2556 -5148 -2490 -5143
rect -2444 -5200 -2410 -5060
rect -2364 -5092 -2298 -5088
rect -2367 -5144 -2357 -5092
rect -2305 -5144 -2295 -5092
rect -2364 -5148 -2298 -5144
rect -2252 -5200 -2218 -5060
rect -2172 -5092 -2106 -5088
rect -2175 -5144 -2165 -5092
rect -2113 -5144 -2103 -5092
rect -2048 -5138 -2042 -4938
rect -2008 -5138 -2002 -4938
rect -2172 -5148 -2106 -5144
rect -3300 -5234 -2218 -5200
rect -2048 -5270 -2002 -5138
rect 70 -5142 149 -5090
rect 201 -5142 211 -5090
rect 251 -5200 285 -4637
rect 435 -4603 469 -4470
rect 627 -4603 661 -4470
rect 819 -4603 853 -4470
rect 1011 -4603 1045 -4470
rect 1203 -4603 1237 -4470
rect 1395 -4603 1429 -4470
rect 1503 -4488 1509 -4288
rect 1543 -4375 1549 -4288
rect 1643 -4335 1670 -4283
rect 1722 -4335 1732 -4283
rect 1610 -4375 1656 -4374
rect 1543 -4386 1656 -4375
rect 1543 -4462 1616 -4386
rect 1650 -4462 1656 -4386
rect 1543 -4474 1656 -4462
rect 1698 -4375 1744 -4374
rect 1772 -4375 1806 -4226
rect 1940 -4283 2006 -4278
rect 1937 -4335 1947 -4283
rect 1999 -4335 2009 -4283
rect 1940 -4338 2006 -4335
rect 2052 -4366 2086 -4226
rect 2132 -4283 2198 -4278
rect 2128 -4335 2138 -4283
rect 2190 -4335 2200 -4283
rect 2132 -4338 2198 -4335
rect 2244 -4366 2278 -4226
rect 2324 -4283 2390 -4278
rect 2320 -4335 2330 -4283
rect 2382 -4335 2392 -4283
rect 2324 -4338 2390 -4335
rect 2436 -4366 2470 -4226
rect 2516 -4283 2582 -4278
rect 2512 -4335 2522 -4283
rect 2574 -4335 2584 -4283
rect 2516 -4338 2582 -4335
rect 2628 -4366 2662 -4226
rect 2708 -4282 2774 -4278
rect 2705 -4334 2715 -4282
rect 2767 -4334 2777 -4282
rect 2708 -4338 2774 -4334
rect 2820 -4366 2854 -4226
rect 2900 -4282 2966 -4278
rect 2897 -4334 2907 -4282
rect 2959 -4334 2969 -4282
rect 3024 -4288 3070 -4115
rect 2900 -4338 2966 -4334
rect 1698 -4386 1806 -4375
rect 1698 -4462 1704 -4386
rect 1738 -4462 1806 -4386
rect 1698 -4474 1806 -4462
rect 1950 -4378 1996 -4366
rect 1950 -4458 1956 -4378
rect 1990 -4458 1996 -4378
rect 1950 -4470 1996 -4458
rect 2046 -4378 2092 -4366
rect 2046 -4458 2052 -4378
rect 2086 -4458 2092 -4378
rect 2046 -4470 2092 -4458
rect 2142 -4378 2188 -4366
rect 2142 -4458 2148 -4378
rect 2182 -4458 2188 -4378
rect 2142 -4470 2188 -4458
rect 2238 -4378 2284 -4366
rect 2238 -4458 2244 -4378
rect 2278 -4458 2284 -4378
rect 2238 -4470 2284 -4458
rect 2334 -4378 2380 -4366
rect 2334 -4458 2340 -4378
rect 2374 -4458 2380 -4378
rect 2334 -4470 2380 -4458
rect 2430 -4378 2476 -4366
rect 2430 -4458 2436 -4378
rect 2470 -4458 2476 -4378
rect 2430 -4470 2476 -4458
rect 2526 -4378 2572 -4366
rect 2526 -4458 2532 -4378
rect 2566 -4458 2572 -4378
rect 2526 -4470 2572 -4458
rect 2622 -4378 2668 -4366
rect 2622 -4458 2628 -4378
rect 2662 -4458 2668 -4378
rect 2622 -4470 2668 -4458
rect 2718 -4378 2764 -4366
rect 2718 -4458 2724 -4378
rect 2758 -4458 2764 -4378
rect 2718 -4470 2764 -4458
rect 2814 -4378 2860 -4366
rect 2814 -4458 2820 -4378
rect 2854 -4458 2860 -4378
rect 2814 -4470 2860 -4458
rect 2910 -4378 2956 -4366
rect 2910 -4458 2916 -4378
rect 2950 -4458 2956 -4378
rect 2910 -4470 2956 -4458
rect 1543 -4475 1649 -4474
rect 1703 -4475 1806 -4474
rect 1543 -4488 1549 -4475
rect 1503 -4500 1549 -4488
rect 1648 -4512 1706 -4506
rect 1648 -4513 1660 -4512
rect 1694 -4513 1706 -4512
rect 1640 -4565 1650 -4513
rect 1702 -4565 1712 -4513
rect 1772 -4603 1806 -4475
rect 435 -4637 1806 -4603
rect 435 -4778 469 -4637
rect 627 -4778 661 -4637
rect 819 -4778 853 -4637
rect 1011 -4778 1045 -4637
rect 1203 -4778 1237 -4637
rect 1395 -4778 1429 -4637
rect 1503 -4752 1549 -4740
rect 429 -4790 475 -4778
rect 429 -5038 435 -4790
rect 469 -5038 475 -4790
rect 429 -5050 475 -5038
rect 525 -4790 571 -4778
rect 525 -5038 531 -4790
rect 565 -5038 571 -4790
rect 525 -5050 571 -5038
rect 621 -4790 667 -4778
rect 621 -5038 627 -4790
rect 661 -5038 667 -4790
rect 621 -5050 667 -5038
rect 717 -4790 763 -4778
rect 717 -5038 723 -4790
rect 757 -5038 763 -4790
rect 717 -5050 763 -5038
rect 813 -4790 859 -4778
rect 813 -5038 819 -4790
rect 853 -5038 859 -4790
rect 813 -5050 859 -5038
rect 909 -4790 955 -4778
rect 909 -5038 915 -4790
rect 949 -5038 955 -4790
rect 909 -5050 955 -5038
rect 1005 -4790 1051 -4778
rect 1005 -5038 1011 -4790
rect 1045 -5038 1051 -4790
rect 1005 -5050 1051 -5038
rect 1101 -4790 1147 -4778
rect 1101 -5038 1107 -4790
rect 1141 -5038 1147 -4790
rect 1101 -5050 1147 -5038
rect 1197 -4790 1243 -4778
rect 1197 -5038 1203 -4790
rect 1237 -5038 1243 -4790
rect 1197 -5050 1243 -5038
rect 1293 -4790 1339 -4778
rect 1293 -5038 1299 -4790
rect 1333 -5038 1339 -4790
rect 1293 -5050 1339 -5038
rect 1389 -4790 1435 -4778
rect 1389 -5038 1395 -4790
rect 1429 -5038 1435 -4790
rect 1389 -5050 1435 -5038
rect 416 -5142 426 -5090
rect 478 -5142 488 -5090
rect 531 -5200 565 -5050
rect 609 -5142 619 -5090
rect 671 -5142 681 -5090
rect 723 -5200 757 -5050
rect 800 -5142 810 -5090
rect 862 -5142 872 -5090
rect 915 -5200 949 -5050
rect 992 -5142 1002 -5090
rect 1054 -5142 1064 -5090
rect 1107 -5200 1141 -5050
rect 1184 -5142 1194 -5090
rect 1246 -5142 1256 -5090
rect 1299 -5200 1333 -5050
rect 1376 -5142 1386 -5090
rect 1438 -5142 1448 -5090
rect 1503 -5138 1509 -4752
rect 1543 -5138 1549 -4752
rect 251 -5234 1333 -5200
rect 1503 -5314 1549 -5138
rect 1643 -5142 1670 -5090
rect 1722 -5142 1732 -5090
rect 1772 -5200 1806 -4637
rect 1956 -4603 1990 -4470
rect 2148 -4603 2182 -4470
rect 2340 -4603 2374 -4470
rect 2532 -4603 2566 -4470
rect 2724 -4603 2758 -4470
rect 2916 -4603 2950 -4470
rect 3024 -4488 3030 -4288
rect 3064 -4488 3070 -4288
rect 3024 -4500 3070 -4488
rect 3273 -4603 3307 -3259
rect 1956 -4637 3307 -4603
rect 1956 -4778 1990 -4637
rect 2148 -4778 2182 -4637
rect 2340 -4778 2374 -4637
rect 2532 -4778 2566 -4637
rect 2724 -4778 2758 -4637
rect 2916 -4778 2950 -4637
rect 3024 -4752 3070 -4740
rect 1950 -4790 1996 -4778
rect 1950 -5038 1956 -4790
rect 1990 -5038 1996 -4790
rect 1950 -5050 1996 -5038
rect 2046 -4790 2092 -4778
rect 2046 -5038 2052 -4790
rect 2086 -5038 2092 -4790
rect 2046 -5050 2092 -5038
rect 2142 -4790 2188 -4778
rect 2142 -5038 2148 -4790
rect 2182 -5038 2188 -4790
rect 2142 -5050 2188 -5038
rect 2238 -4790 2284 -4778
rect 2238 -5038 2244 -4790
rect 2278 -5038 2284 -4790
rect 2238 -5050 2284 -5038
rect 2334 -4790 2380 -4778
rect 2334 -5038 2340 -4790
rect 2374 -5038 2380 -4790
rect 2334 -5050 2380 -5038
rect 2430 -4790 2476 -4778
rect 2430 -5038 2436 -4790
rect 2470 -5038 2476 -4790
rect 2430 -5050 2476 -5038
rect 2526 -4790 2572 -4778
rect 2526 -5038 2532 -4790
rect 2566 -5038 2572 -4790
rect 2526 -5050 2572 -5038
rect 2622 -4790 2668 -4778
rect 2622 -5038 2628 -4790
rect 2662 -5038 2668 -4790
rect 2622 -5050 2668 -5038
rect 2718 -4790 2764 -4778
rect 2718 -5038 2724 -4790
rect 2758 -5038 2764 -4790
rect 2718 -5050 2764 -5038
rect 2814 -4790 2860 -4778
rect 2814 -5038 2820 -4790
rect 2854 -5038 2860 -4790
rect 2814 -5050 2860 -5038
rect 2910 -4790 2956 -4778
rect 2910 -5038 2916 -4790
rect 2950 -5038 2956 -4790
rect 2910 -5050 2956 -5038
rect 1937 -5142 1947 -5090
rect 1999 -5142 2009 -5090
rect 2052 -5200 2086 -5050
rect 2130 -5142 2140 -5090
rect 2192 -5142 2202 -5090
rect 2244 -5200 2278 -5050
rect 2321 -5142 2331 -5090
rect 2383 -5142 2393 -5090
rect 2436 -5200 2470 -5050
rect 2513 -5142 2523 -5090
rect 2575 -5142 2585 -5090
rect 2628 -5200 2662 -5050
rect 2705 -5142 2715 -5090
rect 2767 -5142 2777 -5090
rect 2820 -5200 2854 -5050
rect 2897 -5142 2907 -5090
rect 2959 -5142 2969 -5090
rect 3024 -5138 3030 -4752
rect 3064 -5138 3070 -4752
rect 1772 -5234 2854 -5200
rect 3024 -5314 3070 -5138
<< via1 >>
rect -3402 -246 -3350 -194
rect -3125 -204 -3073 -194
rect -3125 -238 -3116 -204
rect -3116 -238 -3082 -204
rect -3082 -238 -3073 -204
rect -3125 -246 -3073 -238
rect -2932 -204 -2880 -194
rect -2932 -238 -2924 -204
rect -2924 -238 -2890 -204
rect -2890 -238 -2880 -204
rect -2932 -246 -2880 -238
rect -2741 -204 -2689 -194
rect -2741 -238 -2732 -204
rect -2732 -238 -2698 -204
rect -2698 -238 -2689 -204
rect -2741 -246 -2689 -238
rect -2549 -204 -2497 -194
rect -2549 -238 -2540 -204
rect -2540 -238 -2506 -204
rect -2506 -238 -2497 -204
rect -2549 -246 -2497 -238
rect -2357 -204 -2305 -194
rect -2357 -238 -2348 -204
rect -2348 -238 -2314 -204
rect -2314 -238 -2305 -204
rect -2357 -246 -2305 -238
rect -2165 -204 -2113 -194
rect -2165 -238 -2156 -204
rect -2156 -238 -2122 -204
rect -2122 -238 -2113 -204
rect -2165 -246 -2113 -238
rect -1587 -121 -1535 -69
rect -914 -121 -862 -69
rect -3402 -1053 -3350 -1001
rect -1942 -246 -1890 -194
rect -1416 -246 -1364 -194
rect 149 -245 201 -193
rect 426 -200 478 -193
rect 426 -234 435 -200
rect 435 -234 469 -200
rect 469 -234 478 -200
rect 426 -245 478 -234
rect 617 -200 669 -193
rect 617 -234 627 -200
rect 627 -234 661 -200
rect 661 -234 669 -200
rect 617 -245 669 -234
rect 809 -200 861 -193
rect 809 -234 819 -200
rect 819 -234 853 -200
rect 853 -234 861 -200
rect 809 -245 861 -234
rect 1001 -200 1053 -193
rect 1001 -234 1011 -200
rect 1011 -234 1045 -200
rect 1045 -234 1053 -200
rect 1001 -245 1053 -234
rect 1194 -200 1246 -192
rect 1194 -234 1203 -200
rect 1203 -234 1237 -200
rect 1237 -234 1246 -200
rect 1194 -244 1246 -234
rect 1386 -200 1438 -192
rect 1386 -234 1395 -200
rect 1395 -234 1429 -200
rect 1429 -234 1438 -200
rect 1386 -244 1438 -234
rect -1416 -645 -1364 -593
rect -461 -594 -409 -584
rect -461 -628 -452 -594
rect -452 -628 -418 -594
rect -418 -628 -409 -594
rect -461 -636 -409 -628
rect -3125 -1012 -3073 -1001
rect -3125 -1046 -3116 -1012
rect -3116 -1046 -3082 -1012
rect -3082 -1046 -3073 -1012
rect -3125 -1053 -3073 -1046
rect -2934 -1012 -2882 -1001
rect -2934 -1046 -2924 -1012
rect -2924 -1046 -2890 -1012
rect -2890 -1046 -2882 -1012
rect -2934 -1053 -2882 -1046
rect -2742 -1012 -2690 -1001
rect -2742 -1046 -2732 -1012
rect -2732 -1046 -2698 -1012
rect -2698 -1046 -2690 -1012
rect -2742 -1053 -2690 -1046
rect -2550 -1012 -2498 -1001
rect -2550 -1046 -2540 -1012
rect -2540 -1046 -2506 -1012
rect -2506 -1046 -2498 -1012
rect -2550 -1053 -2498 -1046
rect -2357 -1012 -2305 -1002
rect -2357 -1046 -2348 -1012
rect -2348 -1046 -2314 -1012
rect -2314 -1046 -2305 -1012
rect -2357 -1054 -2305 -1046
rect -2165 -1012 -2113 -1002
rect -2165 -1046 -2156 -1012
rect -2156 -1046 -2122 -1012
rect -2122 -1046 -2113 -1012
rect -2165 -1054 -2113 -1046
rect -914 -698 -862 -690
rect -914 -732 -905 -698
rect -905 -732 -871 -698
rect -871 -732 -862 -698
rect -914 -742 -862 -732
rect -549 -700 -497 -694
rect -549 -734 -538 -700
rect -538 -734 -504 -700
rect -504 -734 -497 -700
rect -549 -746 -497 -734
rect 149 -1052 201 -1000
rect 1670 -245 1722 -193
rect 1947 -200 1999 -193
rect 1947 -234 1956 -200
rect 1956 -234 1990 -200
rect 1990 -234 1999 -200
rect 1947 -245 1999 -234
rect 2138 -200 2190 -193
rect 2138 -234 2148 -200
rect 2148 -234 2182 -200
rect 2182 -234 2190 -200
rect 2138 -245 2190 -234
rect 2330 -200 2382 -193
rect 2330 -234 2340 -200
rect 2340 -234 2374 -200
rect 2374 -234 2382 -200
rect 2330 -245 2382 -234
rect 2522 -200 2574 -193
rect 2522 -234 2532 -200
rect 2532 -234 2566 -200
rect 2566 -234 2574 -200
rect 2522 -245 2574 -234
rect 2715 -200 2767 -192
rect 2715 -234 2724 -200
rect 2724 -234 2758 -200
rect 2758 -234 2767 -200
rect 2715 -244 2767 -234
rect 2907 -200 2959 -192
rect 2907 -234 2916 -200
rect 2916 -234 2950 -200
rect 2950 -234 2959 -200
rect 2907 -244 2959 -234
rect 1650 -456 1660 -423
rect 1660 -456 1694 -423
rect 1694 -456 1702 -423
rect 1650 -475 1702 -456
rect 426 -1008 478 -1000
rect 426 -1042 435 -1008
rect 435 -1042 469 -1008
rect 469 -1042 478 -1008
rect 426 -1052 478 -1042
rect 619 -1008 671 -1000
rect 619 -1042 627 -1008
rect 627 -1042 661 -1008
rect 661 -1042 671 -1008
rect 619 -1052 671 -1042
rect 810 -1008 862 -1000
rect 810 -1042 819 -1008
rect 819 -1042 853 -1008
rect 853 -1042 862 -1008
rect 810 -1052 862 -1042
rect 1002 -1008 1054 -1000
rect 1002 -1042 1011 -1008
rect 1011 -1042 1045 -1008
rect 1045 -1042 1054 -1008
rect 1002 -1052 1054 -1042
rect 1194 -1008 1246 -1000
rect 1194 -1042 1203 -1008
rect 1203 -1042 1237 -1008
rect 1237 -1042 1246 -1008
rect 1194 -1052 1246 -1042
rect 1386 -1008 1438 -1000
rect 1386 -1042 1395 -1008
rect 1395 -1042 1429 -1008
rect 1429 -1042 1438 -1008
rect 1386 -1052 1438 -1042
rect 98 -1240 150 -1188
rect 1670 -1052 1722 -1000
rect 1947 -1008 1999 -1000
rect 1947 -1042 1956 -1008
rect 1956 -1042 1990 -1008
rect 1990 -1042 1999 -1008
rect 1947 -1052 1999 -1042
rect 2140 -1008 2192 -1000
rect 2140 -1042 2148 -1008
rect 2148 -1042 2182 -1008
rect 2182 -1042 2192 -1008
rect 2140 -1052 2192 -1042
rect 2331 -1008 2383 -1000
rect 2331 -1042 2340 -1008
rect 2340 -1042 2374 -1008
rect 2374 -1042 2383 -1008
rect 2331 -1052 2383 -1042
rect 2523 -1008 2575 -1000
rect 2523 -1042 2532 -1008
rect 2532 -1042 2566 -1008
rect 2566 -1042 2575 -1008
rect 2523 -1052 2575 -1042
rect 2715 -1008 2767 -1000
rect 2715 -1042 2724 -1008
rect 2724 -1042 2758 -1008
rect 2758 -1042 2767 -1008
rect 2715 -1052 2767 -1042
rect 2907 -1008 2959 -1000
rect 2907 -1042 2916 -1008
rect 2916 -1042 2950 -1008
rect 2950 -1042 2959 -1008
rect 2907 -1052 2959 -1042
rect -287 -1355 -235 -1303
rect -3402 -1580 -3350 -1528
rect -3125 -1538 -3073 -1528
rect -3125 -1572 -3116 -1538
rect -3116 -1572 -3082 -1538
rect -3082 -1572 -3073 -1538
rect -3125 -1580 -3073 -1572
rect -2932 -1538 -2880 -1528
rect -2932 -1572 -2924 -1538
rect -2924 -1572 -2890 -1538
rect -2890 -1572 -2880 -1538
rect -2932 -1580 -2880 -1572
rect -2741 -1538 -2689 -1528
rect -2741 -1572 -2732 -1538
rect -2732 -1572 -2698 -1538
rect -2698 -1572 -2689 -1538
rect -2741 -1580 -2689 -1572
rect -2549 -1538 -2497 -1528
rect -2549 -1572 -2540 -1538
rect -2540 -1572 -2506 -1538
rect -2506 -1572 -2497 -1538
rect -2549 -1580 -2497 -1572
rect -2357 -1538 -2305 -1528
rect -2357 -1572 -2348 -1538
rect -2348 -1572 -2314 -1538
rect -2314 -1572 -2305 -1538
rect -2357 -1580 -2305 -1572
rect -2165 -1538 -2113 -1528
rect -2165 -1572 -2156 -1538
rect -2156 -1572 -2122 -1538
rect -2122 -1572 -2113 -1538
rect -2165 -1580 -2113 -1572
rect -3402 -2387 -3350 -2335
rect -1724 -1580 -1672 -1528
rect -1416 -1580 -1364 -1528
rect -478 -1676 -426 -1669
rect -478 -1710 -469 -1676
rect -469 -1710 -435 -1676
rect -435 -1710 -426 -1676
rect -478 -1721 -426 -1710
rect -592 -1784 -540 -1776
rect -592 -1818 -582 -1784
rect -582 -1818 -548 -1784
rect -548 -1818 -540 -1784
rect -592 -1828 -540 -1818
rect -416 -1785 -364 -1779
rect -416 -1819 -408 -1785
rect -408 -1819 -374 -1785
rect -374 -1819 -364 -1785
rect -416 -1831 -364 -1819
rect 149 -1579 201 -1527
rect 426 -1534 478 -1527
rect 426 -1568 435 -1534
rect 435 -1568 469 -1534
rect 469 -1568 478 -1534
rect 426 -1579 478 -1568
rect 617 -1534 669 -1527
rect 617 -1568 627 -1534
rect 627 -1568 661 -1534
rect 661 -1568 669 -1534
rect 617 -1579 669 -1568
rect 809 -1534 861 -1527
rect 809 -1568 819 -1534
rect 819 -1568 853 -1534
rect 853 -1568 861 -1534
rect 809 -1579 861 -1568
rect 1001 -1534 1053 -1527
rect 1001 -1568 1011 -1534
rect 1011 -1568 1045 -1534
rect 1045 -1568 1053 -1534
rect 1001 -1579 1053 -1568
rect 1194 -1534 1246 -1526
rect 1194 -1568 1203 -1534
rect 1203 -1568 1237 -1534
rect 1237 -1568 1246 -1534
rect 1194 -1578 1246 -1568
rect 1386 -1534 1438 -1526
rect 1386 -1568 1395 -1534
rect 1395 -1568 1429 -1534
rect 1429 -1568 1438 -1534
rect 1386 -1578 1438 -1568
rect -872 -1971 -820 -1919
rect -416 -1971 -364 -1919
rect -3125 -2346 -3073 -2335
rect -3125 -2380 -3116 -2346
rect -3116 -2380 -3082 -2346
rect -3082 -2380 -3073 -2346
rect -3125 -2387 -3073 -2380
rect -2934 -2346 -2882 -2335
rect -2934 -2380 -2924 -2346
rect -2924 -2380 -2890 -2346
rect -2890 -2380 -2882 -2346
rect -2934 -2387 -2882 -2380
rect -2742 -2346 -2690 -2335
rect -2742 -2380 -2732 -2346
rect -2732 -2380 -2698 -2346
rect -2698 -2380 -2690 -2346
rect -2742 -2387 -2690 -2380
rect -2550 -2346 -2498 -2335
rect -2550 -2380 -2540 -2346
rect -2540 -2380 -2506 -2346
rect -2506 -2380 -2498 -2346
rect -2550 -2387 -2498 -2380
rect -2357 -2346 -2305 -2336
rect -2357 -2380 -2348 -2346
rect -2348 -2380 -2314 -2346
rect -2314 -2380 -2305 -2346
rect -2357 -2388 -2305 -2380
rect -2165 -2346 -2113 -2336
rect -2165 -2380 -2156 -2346
rect -2156 -2380 -2122 -2346
rect -2122 -2380 -2113 -2346
rect -2165 -2388 -2113 -2380
rect -592 -2277 -540 -2225
rect -287 -2313 -235 -2261
rect -1101 -2398 -1049 -2388
rect -1101 -2432 -1091 -2398
rect -1091 -2432 -1057 -2398
rect -1057 -2432 -1049 -2398
rect -1101 -2440 -1049 -2432
rect -762 -2440 -710 -2388
rect -592 -2398 -540 -2390
rect -592 -2432 -583 -2398
rect -583 -2432 -549 -2398
rect -549 -2432 -540 -2398
rect -592 -2442 -540 -2432
rect -412 -2395 -360 -2385
rect -412 -2429 -402 -2395
rect -402 -2429 -368 -2395
rect -368 -2429 -360 -2395
rect -412 -2437 -360 -2429
rect 149 -2386 201 -2334
rect 1670 -1579 1722 -1527
rect 1947 -1534 1999 -1527
rect 1947 -1568 1956 -1534
rect 1956 -1568 1990 -1534
rect 1990 -1568 1999 -1534
rect 1947 -1579 1999 -1568
rect 2138 -1534 2190 -1527
rect 2138 -1568 2148 -1534
rect 2148 -1568 2182 -1534
rect 2182 -1568 2190 -1534
rect 2138 -1579 2190 -1568
rect 2330 -1534 2382 -1527
rect 2330 -1568 2340 -1534
rect 2340 -1568 2374 -1534
rect 2374 -1568 2382 -1534
rect 2330 -1579 2382 -1568
rect 2522 -1534 2574 -1527
rect 2522 -1568 2532 -1534
rect 2532 -1568 2566 -1534
rect 2566 -1568 2574 -1534
rect 2522 -1579 2574 -1568
rect 2715 -1534 2767 -1526
rect 2715 -1568 2724 -1534
rect 2724 -1568 2758 -1534
rect 2758 -1568 2767 -1534
rect 2715 -1578 2767 -1568
rect 2907 -1534 2959 -1526
rect 2907 -1568 2916 -1534
rect 2916 -1568 2950 -1534
rect 2950 -1568 2959 -1534
rect 2907 -1578 2959 -1568
rect 1650 -1790 1660 -1757
rect 1660 -1790 1694 -1757
rect 1694 -1790 1702 -1757
rect 1650 -1809 1702 -1790
rect 426 -2342 478 -2334
rect 426 -2376 435 -2342
rect 435 -2376 469 -2342
rect 469 -2376 478 -2342
rect 426 -2386 478 -2376
rect 619 -2342 671 -2334
rect 619 -2376 627 -2342
rect 627 -2376 661 -2342
rect 661 -2376 671 -2342
rect 619 -2386 671 -2376
rect 810 -2342 862 -2334
rect 810 -2376 819 -2342
rect 819 -2376 853 -2342
rect 853 -2376 862 -2342
rect 810 -2386 862 -2376
rect 1002 -2342 1054 -2334
rect 1002 -2376 1011 -2342
rect 1011 -2376 1045 -2342
rect 1045 -2376 1054 -2342
rect 1002 -2386 1054 -2376
rect 1194 -2342 1246 -2334
rect 1194 -2376 1203 -2342
rect 1203 -2376 1237 -2342
rect 1237 -2376 1246 -2342
rect 1194 -2386 1246 -2376
rect 1386 -2342 1438 -2334
rect 1386 -2376 1395 -2342
rect 1395 -2376 1429 -2342
rect 1429 -2376 1438 -2342
rect 1386 -2386 1438 -2376
rect -1240 -2543 -1188 -2491
rect -412 -2543 -360 -2491
rect 1670 -2386 1722 -2334
rect 1947 -2342 1999 -2334
rect 1947 -2376 1956 -2342
rect 1956 -2376 1990 -2342
rect 1990 -2376 1999 -2342
rect 1947 -2386 1999 -2376
rect 2140 -2342 2192 -2334
rect 2140 -2376 2148 -2342
rect 2148 -2376 2182 -2342
rect 2182 -2376 2192 -2342
rect 2140 -2386 2192 -2376
rect 2331 -2342 2383 -2334
rect 2331 -2376 2340 -2342
rect 2340 -2376 2374 -2342
rect 2374 -2376 2383 -2342
rect 2331 -2386 2383 -2376
rect 2523 -2342 2575 -2334
rect 2523 -2376 2532 -2342
rect 2532 -2376 2566 -2342
rect 2566 -2376 2575 -2342
rect 2523 -2386 2575 -2376
rect 2715 -2342 2767 -2334
rect 2715 -2376 2724 -2342
rect 2724 -2376 2758 -2342
rect 2758 -2376 2767 -2342
rect 2715 -2386 2767 -2376
rect 2907 -2342 2959 -2334
rect 2907 -2376 2916 -2342
rect 2916 -2376 2950 -2342
rect 2950 -2376 2959 -2342
rect 2907 -2386 2959 -2376
rect -3402 -2958 -3350 -2906
rect -3125 -2916 -3073 -2906
rect -3125 -2950 -3116 -2916
rect -3116 -2950 -3082 -2916
rect -3082 -2950 -3073 -2916
rect -3125 -2958 -3073 -2950
rect -2932 -2916 -2880 -2906
rect -2932 -2950 -2924 -2916
rect -2924 -2950 -2890 -2916
rect -2890 -2950 -2880 -2916
rect -2932 -2958 -2880 -2950
rect -2741 -2916 -2689 -2906
rect -2741 -2950 -2732 -2916
rect -2732 -2950 -2698 -2916
rect -2698 -2950 -2689 -2916
rect -2741 -2958 -2689 -2950
rect -2549 -2916 -2497 -2906
rect -2549 -2950 -2540 -2916
rect -2540 -2950 -2506 -2916
rect -2506 -2950 -2497 -2916
rect -2549 -2958 -2497 -2950
rect -2357 -2916 -2305 -2906
rect -2357 -2950 -2348 -2916
rect -2348 -2950 -2314 -2916
rect -2314 -2950 -2305 -2916
rect -2357 -2958 -2305 -2950
rect -2165 -2916 -2113 -2906
rect -2165 -2950 -2156 -2916
rect -2156 -2950 -2122 -2916
rect -2122 -2950 -2113 -2916
rect -2165 -2958 -2113 -2950
rect -762 -2827 -710 -2775
rect -412 -2827 -360 -2775
rect -3402 -3765 -3350 -3713
rect -1926 -2958 -1874 -2906
rect -1416 -2958 -1364 -2906
rect -1098 -2874 -1046 -2865
rect -1098 -2908 -1089 -2874
rect -1089 -2908 -1055 -2874
rect -1055 -2908 -1046 -2874
rect -1098 -2917 -1046 -2908
rect -872 -2916 -820 -2864
rect -412 -2875 -360 -2866
rect -412 -2909 -401 -2875
rect -401 -2909 -367 -2875
rect -367 -2909 -360 -2875
rect -412 -2918 -360 -2909
rect 149 -2957 201 -2905
rect -236 -3078 -184 -3026
rect 426 -2912 478 -2905
rect 426 -2946 435 -2912
rect 435 -2946 469 -2912
rect 469 -2946 478 -2912
rect 426 -2957 478 -2946
rect 617 -2912 669 -2905
rect 617 -2946 627 -2912
rect 627 -2946 661 -2912
rect 661 -2946 669 -2912
rect 617 -2957 669 -2946
rect 809 -2912 861 -2905
rect 809 -2946 819 -2912
rect 819 -2946 853 -2912
rect 853 -2946 861 -2912
rect 809 -2957 861 -2946
rect 1001 -2912 1053 -2905
rect 1001 -2946 1011 -2912
rect 1011 -2946 1045 -2912
rect 1045 -2946 1053 -2912
rect 1001 -2957 1053 -2946
rect 1194 -2912 1246 -2904
rect 1194 -2946 1203 -2912
rect 1203 -2946 1237 -2912
rect 1237 -2946 1246 -2912
rect 1194 -2956 1246 -2946
rect 1386 -2912 1438 -2904
rect 1386 -2946 1395 -2912
rect 1395 -2946 1429 -2912
rect 1429 -2946 1438 -2912
rect 1386 -2956 1438 -2946
rect -762 -3445 -710 -3393
rect -414 -3445 -362 -3393
rect -1241 -3539 -1187 -3485
rect -414 -3487 -362 -3474
rect -414 -3521 -405 -3487
rect -405 -3521 -371 -3487
rect -371 -3521 -362 -3487
rect -414 -3526 -362 -3521
rect -3125 -3724 -3073 -3713
rect -3125 -3758 -3116 -3724
rect -3116 -3758 -3082 -3724
rect -3082 -3758 -3073 -3724
rect -3125 -3765 -3073 -3758
rect -2934 -3724 -2882 -3713
rect -2934 -3758 -2924 -3724
rect -2924 -3758 -2890 -3724
rect -2890 -3758 -2882 -3724
rect -2934 -3765 -2882 -3758
rect -2742 -3724 -2690 -3713
rect -2742 -3758 -2732 -3724
rect -2732 -3758 -2698 -3724
rect -2698 -3758 -2690 -3724
rect -2742 -3765 -2690 -3758
rect -2550 -3724 -2498 -3713
rect -2550 -3758 -2540 -3724
rect -2540 -3758 -2506 -3724
rect -2506 -3758 -2498 -3724
rect -2550 -3765 -2498 -3758
rect -2357 -3724 -2305 -3714
rect -2357 -3758 -2348 -3724
rect -2348 -3758 -2314 -3724
rect -2314 -3758 -2305 -3724
rect -2357 -3766 -2305 -3758
rect -2165 -3724 -2113 -3714
rect -2165 -3758 -2156 -3724
rect -2156 -3758 -2122 -3724
rect -2122 -3758 -2113 -3724
rect -2165 -3766 -2113 -3758
rect -500 -3590 -448 -3580
rect -500 -3624 -492 -3590
rect -492 -3624 -458 -3590
rect -458 -3624 -448 -3590
rect -500 -3632 -448 -3624
rect -235 -3764 -183 -3712
rect 149 -3764 201 -3712
rect 1670 -2957 1722 -2905
rect 1947 -2912 1999 -2905
rect 1947 -2946 1956 -2912
rect 1956 -2946 1990 -2912
rect 1990 -2946 1999 -2912
rect 1947 -2957 1999 -2946
rect 2138 -2912 2190 -2905
rect 2138 -2946 2148 -2912
rect 2148 -2946 2182 -2912
rect 2182 -2946 2190 -2912
rect 2138 -2957 2190 -2946
rect 2330 -2912 2382 -2905
rect 2330 -2946 2340 -2912
rect 2340 -2946 2374 -2912
rect 2374 -2946 2382 -2912
rect 2330 -2957 2382 -2946
rect 2522 -2912 2574 -2905
rect 2522 -2946 2532 -2912
rect 2532 -2946 2566 -2912
rect 2566 -2946 2574 -2912
rect 2522 -2957 2574 -2946
rect 2715 -2912 2767 -2904
rect 2715 -2946 2724 -2912
rect 2724 -2946 2758 -2912
rect 2758 -2946 2767 -2912
rect 2715 -2956 2767 -2946
rect 2907 -2912 2959 -2904
rect 2907 -2946 2916 -2912
rect 2916 -2946 2950 -2912
rect 2950 -2946 2959 -2912
rect 2907 -2956 2959 -2946
rect 1650 -3168 1660 -3135
rect 1660 -3168 1694 -3135
rect 1694 -3168 1702 -3135
rect 1650 -3187 1702 -3168
rect 426 -3720 478 -3712
rect 426 -3754 435 -3720
rect 435 -3754 469 -3720
rect 469 -3754 478 -3720
rect 426 -3764 478 -3754
rect 619 -3720 671 -3712
rect 619 -3754 627 -3720
rect 627 -3754 661 -3720
rect 661 -3754 671 -3720
rect 619 -3764 671 -3754
rect 810 -3720 862 -3712
rect 810 -3754 819 -3720
rect 819 -3754 853 -3720
rect 853 -3754 862 -3720
rect 810 -3764 862 -3754
rect 1002 -3720 1054 -3712
rect 1002 -3754 1011 -3720
rect 1011 -3754 1045 -3720
rect 1045 -3754 1054 -3720
rect 1002 -3764 1054 -3754
rect 1194 -3720 1246 -3712
rect 1194 -3754 1203 -3720
rect 1203 -3754 1237 -3720
rect 1237 -3754 1246 -3720
rect 1194 -3764 1246 -3754
rect 1386 -3720 1438 -3712
rect 1386 -3754 1395 -3720
rect 1395 -3754 1429 -3720
rect 1429 -3754 1438 -3720
rect 1386 -3764 1438 -3754
rect 1670 -3764 1722 -3712
rect 1947 -3720 1999 -3712
rect 1947 -3754 1956 -3720
rect 1956 -3754 1990 -3720
rect 1990 -3754 1999 -3720
rect 1947 -3764 1999 -3754
rect 2140 -3720 2192 -3712
rect 2140 -3754 2148 -3720
rect 2148 -3754 2182 -3720
rect 2182 -3754 2192 -3720
rect 2140 -3764 2192 -3754
rect 2331 -3720 2383 -3712
rect 2331 -3754 2340 -3720
rect 2340 -3754 2374 -3720
rect 2374 -3754 2383 -3720
rect 2331 -3764 2383 -3754
rect 2523 -3720 2575 -3712
rect 2523 -3754 2532 -3720
rect 2532 -3754 2566 -3720
rect 2566 -3754 2575 -3720
rect 2523 -3764 2575 -3754
rect 2715 -3720 2767 -3712
rect 2715 -3754 2724 -3720
rect 2724 -3754 2758 -3720
rect 2758 -3754 2767 -3720
rect 2715 -3764 2767 -3754
rect 2907 -3720 2959 -3712
rect 2907 -3754 2916 -3720
rect 2916 -3754 2950 -3720
rect 2950 -3754 2959 -3720
rect 2907 -3764 2959 -3754
rect -236 -4003 -184 -3951
rect -3402 -4336 -3350 -4284
rect -3125 -4294 -3073 -4284
rect -3125 -4328 -3116 -4294
rect -3116 -4328 -3082 -4294
rect -3082 -4328 -3073 -4294
rect -3125 -4336 -3073 -4328
rect -2932 -4294 -2880 -4284
rect -2932 -4328 -2924 -4294
rect -2924 -4328 -2890 -4294
rect -2890 -4328 -2880 -4294
rect -2932 -4336 -2880 -4328
rect -2741 -4294 -2689 -4284
rect -2741 -4328 -2732 -4294
rect -2732 -4328 -2698 -4294
rect -2698 -4328 -2689 -4294
rect -2741 -4336 -2689 -4328
rect -2549 -4294 -2497 -4284
rect -2549 -4328 -2540 -4294
rect -2540 -4328 -2506 -4294
rect -2506 -4328 -2497 -4294
rect -2549 -4336 -2497 -4328
rect -2357 -4294 -2305 -4284
rect -2357 -4328 -2348 -4294
rect -2348 -4328 -2314 -4294
rect -2314 -4328 -2305 -4294
rect -2357 -4336 -2305 -4328
rect -2165 -4294 -2113 -4284
rect -2165 -4328 -2156 -4294
rect -2156 -4328 -2122 -4294
rect -2122 -4328 -2113 -4294
rect -2165 -4336 -2113 -4328
rect -81 -4163 -29 -4111
rect -3402 -5143 -3350 -5091
rect -1943 -4336 -1891 -4284
rect -1416 -4336 -1364 -4284
rect 149 -4335 201 -4283
rect 92 -4461 144 -4409
rect -548 -4574 -496 -4565
rect -548 -4608 -540 -4574
rect -540 -4608 -506 -4574
rect -506 -4608 -496 -4574
rect -548 -4617 -496 -4608
rect 426 -4290 478 -4283
rect 426 -4324 435 -4290
rect 435 -4324 469 -4290
rect 469 -4324 478 -4290
rect 426 -4335 478 -4324
rect 617 -4290 669 -4283
rect 617 -4324 627 -4290
rect 627 -4324 661 -4290
rect 661 -4324 669 -4290
rect 617 -4335 669 -4324
rect 809 -4290 861 -4283
rect 809 -4324 819 -4290
rect 819 -4324 853 -4290
rect 853 -4324 861 -4290
rect 809 -4335 861 -4324
rect 1001 -4290 1053 -4283
rect 1001 -4324 1011 -4290
rect 1011 -4324 1045 -4290
rect 1045 -4324 1053 -4290
rect 1001 -4335 1053 -4324
rect 1194 -4290 1246 -4282
rect 1194 -4324 1203 -4290
rect 1203 -4324 1237 -4290
rect 1237 -4324 1246 -4290
rect 1194 -4334 1246 -4324
rect 1386 -4290 1438 -4282
rect 1386 -4324 1395 -4290
rect 1395 -4324 1429 -4290
rect 1429 -4324 1438 -4290
rect 1386 -4334 1438 -4324
rect -3125 -5102 -3073 -5091
rect -3125 -5136 -3116 -5102
rect -3116 -5136 -3082 -5102
rect -3082 -5136 -3073 -5102
rect -3125 -5143 -3073 -5136
rect -2934 -5102 -2882 -5091
rect -2934 -5136 -2924 -5102
rect -2924 -5136 -2890 -5102
rect -2890 -5136 -2882 -5102
rect -2934 -5143 -2882 -5136
rect -2742 -5102 -2690 -5091
rect -2742 -5136 -2732 -5102
rect -2732 -5136 -2698 -5102
rect -2698 -5136 -2690 -5102
rect -2742 -5143 -2690 -5136
rect -2550 -5102 -2498 -5091
rect -2550 -5136 -2540 -5102
rect -2540 -5136 -2506 -5102
rect -2506 -5136 -2498 -5102
rect -2550 -5143 -2498 -5136
rect -2357 -5102 -2305 -5092
rect -2357 -5136 -2348 -5102
rect -2348 -5136 -2314 -5102
rect -2314 -5136 -2305 -5102
rect -2357 -5144 -2305 -5136
rect -2165 -5102 -2113 -5092
rect -2165 -5136 -2156 -5102
rect -2156 -5136 -2122 -5102
rect -2122 -5136 -2113 -5102
rect -2165 -5144 -2113 -5136
rect 149 -5142 201 -5090
rect 1670 -4335 1722 -4283
rect 1947 -4290 1999 -4283
rect 1947 -4324 1956 -4290
rect 1956 -4324 1990 -4290
rect 1990 -4324 1999 -4290
rect 1947 -4335 1999 -4324
rect 2138 -4290 2190 -4283
rect 2138 -4324 2148 -4290
rect 2148 -4324 2182 -4290
rect 2182 -4324 2190 -4290
rect 2138 -4335 2190 -4324
rect 2330 -4290 2382 -4283
rect 2330 -4324 2340 -4290
rect 2340 -4324 2374 -4290
rect 2374 -4324 2382 -4290
rect 2330 -4335 2382 -4324
rect 2522 -4290 2574 -4283
rect 2522 -4324 2532 -4290
rect 2532 -4324 2566 -4290
rect 2566 -4324 2574 -4290
rect 2522 -4335 2574 -4324
rect 2715 -4290 2767 -4282
rect 2715 -4324 2724 -4290
rect 2724 -4324 2758 -4290
rect 2758 -4324 2767 -4290
rect 2715 -4334 2767 -4324
rect 2907 -4290 2959 -4282
rect 2907 -4324 2916 -4290
rect 2916 -4324 2950 -4290
rect 2950 -4324 2959 -4290
rect 2907 -4334 2959 -4324
rect 1650 -4546 1660 -4513
rect 1660 -4546 1694 -4513
rect 1694 -4546 1702 -4513
rect 1650 -4565 1702 -4546
rect 426 -5098 478 -5090
rect 426 -5132 435 -5098
rect 435 -5132 469 -5098
rect 469 -5132 478 -5098
rect 426 -5142 478 -5132
rect 619 -5098 671 -5090
rect 619 -5132 627 -5098
rect 627 -5132 661 -5098
rect 661 -5132 671 -5098
rect 619 -5142 671 -5132
rect 810 -5098 862 -5090
rect 810 -5132 819 -5098
rect 819 -5132 853 -5098
rect 853 -5132 862 -5098
rect 810 -5142 862 -5132
rect 1002 -5098 1054 -5090
rect 1002 -5132 1011 -5098
rect 1011 -5132 1045 -5098
rect 1045 -5132 1054 -5098
rect 1002 -5142 1054 -5132
rect 1194 -5098 1246 -5090
rect 1194 -5132 1203 -5098
rect 1203 -5132 1237 -5098
rect 1237 -5132 1246 -5098
rect 1194 -5142 1246 -5132
rect 1386 -5098 1438 -5090
rect 1386 -5132 1395 -5098
rect 1395 -5132 1429 -5098
rect 1429 -5132 1438 -5098
rect 1386 -5142 1438 -5132
rect 1670 -5142 1722 -5090
rect 1947 -5098 1999 -5090
rect 1947 -5132 1956 -5098
rect 1956 -5132 1990 -5098
rect 1990 -5132 1999 -5098
rect 1947 -5142 1999 -5132
rect 2140 -5098 2192 -5090
rect 2140 -5132 2148 -5098
rect 2148 -5132 2182 -5098
rect 2182 -5132 2192 -5098
rect 2140 -5142 2192 -5132
rect 2331 -5098 2383 -5090
rect 2331 -5132 2340 -5098
rect 2340 -5132 2374 -5098
rect 2374 -5132 2383 -5098
rect 2331 -5142 2383 -5132
rect 2523 -5098 2575 -5090
rect 2523 -5132 2532 -5098
rect 2532 -5132 2566 -5098
rect 2566 -5132 2575 -5098
rect 2523 -5142 2575 -5132
rect 2715 -5098 2767 -5090
rect 2715 -5132 2724 -5098
rect 2724 -5132 2758 -5098
rect 2758 -5132 2767 -5098
rect 2715 -5142 2767 -5132
rect 2907 -5098 2959 -5090
rect 2907 -5132 2916 -5098
rect 2916 -5132 2950 -5098
rect 2950 -5132 2959 -5098
rect 2907 -5142 2959 -5132
<< metal2 >>
rect -1587 -69 -1535 148
rect -3402 -194 -3350 -184
rect -3125 -194 -3073 -184
rect -2932 -194 -2880 -184
rect -2741 -194 -2689 -184
rect -2549 -194 -2497 -184
rect -2357 -194 -2305 -184
rect -2165 -194 -2113 -184
rect -1942 -194 -1890 -184
rect -3350 -246 -3125 -194
rect -3073 -246 -2932 -194
rect -2880 -246 -2741 -194
rect -2689 -246 -2549 -194
rect -2497 -246 -2357 -194
rect -2305 -246 -2165 -194
rect -2113 -246 -1942 -194
rect -3402 -256 -3350 -246
rect -3125 -256 -3073 -246
rect -2932 -256 -2880 -246
rect -2741 -256 -2689 -246
rect -2549 -256 -2497 -246
rect -2357 -256 -2305 -246
rect -2165 -256 -2113 -246
rect -1942 -256 -1890 -246
rect -3402 -1001 -3350 -991
rect -3125 -1001 -3073 -991
rect -2934 -1001 -2882 -991
rect -2742 -1001 -2690 -991
rect -2550 -1001 -2498 -991
rect -2357 -1001 -2305 -992
rect -2165 -1001 -2113 -992
rect -1587 -1001 -1535 -121
rect -3350 -1053 -3125 -1001
rect -3073 -1053 -2934 -1001
rect -2882 -1053 -2742 -1001
rect -2690 -1053 -2550 -1001
rect -2498 -1002 -1535 -1001
rect -2498 -1053 -2357 -1002
rect -3402 -1063 -3350 -1053
rect -3125 -1063 -3073 -1053
rect -2934 -1063 -2882 -1053
rect -2742 -1063 -2690 -1053
rect -2550 -1063 -2498 -1053
rect -2305 -1053 -2165 -1002
rect -2357 -1064 -2305 -1054
rect -2113 -1053 -1535 -1002
rect -2165 -1064 -2113 -1054
rect -3402 -1528 -3350 -1518
rect -3125 -1528 -3073 -1518
rect -2932 -1528 -2880 -1518
rect -2741 -1528 -2689 -1518
rect -2549 -1528 -2497 -1518
rect -2357 -1528 -2305 -1518
rect -2165 -1528 -2113 -1518
rect -1724 -1528 -1672 -1518
rect -3350 -1580 -3125 -1528
rect -3073 -1580 -2932 -1528
rect -2880 -1580 -2741 -1528
rect -2689 -1580 -2549 -1528
rect -2497 -1580 -2357 -1528
rect -2305 -1580 -2165 -1528
rect -2113 -1580 -1724 -1528
rect -3402 -1590 -3350 -1580
rect -3125 -1590 -3073 -1580
rect -2932 -1590 -2880 -1580
rect -2741 -1590 -2689 -1580
rect -2549 -1590 -2497 -1580
rect -2357 -1590 -2305 -1580
rect -2165 -1590 -2113 -1580
rect -1724 -1590 -1672 -1580
rect -3402 -2335 -3350 -2325
rect -3125 -2335 -3073 -2325
rect -2934 -2335 -2882 -2325
rect -2742 -2335 -2690 -2325
rect -2550 -2335 -2498 -2325
rect -2357 -2335 -2305 -2326
rect -2165 -2335 -2113 -2326
rect -1587 -2335 -1535 -1053
rect -3350 -2387 -3125 -2335
rect -3073 -2387 -2934 -2335
rect -2882 -2387 -2742 -2335
rect -2690 -2387 -2550 -2335
rect -2498 -2336 -1535 -2335
rect -2498 -2387 -2357 -2336
rect -3402 -2397 -3350 -2387
rect -3125 -2397 -3073 -2387
rect -2934 -2397 -2882 -2387
rect -2742 -2397 -2690 -2387
rect -2550 -2397 -2498 -2387
rect -2305 -2387 -2165 -2336
rect -2357 -2398 -2305 -2388
rect -2113 -2387 -1535 -2336
rect -2165 -2398 -2113 -2388
rect -3402 -2906 -3350 -2896
rect -3125 -2906 -3073 -2896
rect -2932 -2906 -2880 -2896
rect -2741 -2906 -2689 -2896
rect -2549 -2906 -2497 -2896
rect -2357 -2906 -2305 -2896
rect -2165 -2906 -2113 -2896
rect -1926 -2906 -1874 -2896
rect -3350 -2958 -3125 -2906
rect -3073 -2958 -2932 -2906
rect -2880 -2958 -2741 -2906
rect -2689 -2958 -2549 -2906
rect -2497 -2958 -2357 -2906
rect -2305 -2958 -2165 -2906
rect -2113 -2958 -1926 -2906
rect -3402 -2968 -3350 -2958
rect -3125 -2968 -3073 -2958
rect -2932 -2968 -2880 -2958
rect -2741 -2968 -2689 -2958
rect -2549 -2968 -2497 -2958
rect -2357 -2968 -2305 -2958
rect -2165 -2968 -2113 -2958
rect -1926 -2968 -1874 -2958
rect -3402 -3713 -3350 -3703
rect -3125 -3713 -3073 -3703
rect -2934 -3713 -2882 -3703
rect -2742 -3713 -2690 -3703
rect -2550 -3713 -2498 -3703
rect -2357 -3713 -2305 -3704
rect -2165 -3713 -2113 -3704
rect -1587 -3713 -1535 -2387
rect -1416 -194 -1364 -184
rect -1416 -593 -1364 -246
rect -1416 -1528 -1364 -645
rect -1416 -2906 -1364 -1580
rect -3350 -3765 -3125 -3713
rect -3073 -3765 -2934 -3713
rect -2882 -3765 -2742 -3713
rect -2690 -3765 -2550 -3713
rect -2498 -3714 -1532 -3713
rect -2498 -3765 -2357 -3714
rect -3402 -3775 -3350 -3765
rect -3125 -3775 -3073 -3765
rect -2934 -3775 -2882 -3765
rect -2742 -3775 -2690 -3765
rect -2550 -3775 -2498 -3765
rect -2305 -3765 -2165 -3714
rect -2357 -3776 -2305 -3766
rect -2113 -3765 -1532 -3714
rect -2165 -3776 -2113 -3766
rect -3402 -4284 -3350 -4274
rect -3125 -4284 -3073 -4274
rect -2932 -4284 -2880 -4274
rect -2741 -4284 -2689 -4274
rect -2549 -4284 -2497 -4274
rect -2357 -4284 -2305 -4274
rect -2165 -4284 -2113 -4274
rect -1943 -4284 -1891 -4274
rect -3350 -4336 -3125 -4284
rect -3073 -4336 -2932 -4284
rect -2880 -4336 -2741 -4284
rect -2689 -4336 -2549 -4284
rect -2497 -4336 -2357 -4284
rect -2305 -4336 -2165 -4284
rect -2113 -4336 -1943 -4284
rect -3402 -4346 -3350 -4336
rect -3125 -4346 -3073 -4336
rect -2932 -4346 -2880 -4336
rect -2741 -4346 -2689 -4336
rect -2549 -4346 -2497 -4336
rect -2357 -4346 -2305 -4336
rect -2165 -4346 -2113 -4336
rect -1943 -4346 -1891 -4336
rect -3402 -5091 -3350 -5081
rect -3125 -5091 -3073 -5081
rect -2934 -5091 -2882 -5081
rect -2742 -5091 -2690 -5081
rect -2550 -5091 -2498 -5081
rect -2357 -5091 -2305 -5082
rect -2165 -5091 -2113 -5082
rect -1587 -5091 -1535 -3765
rect -1416 -4284 -1364 -2958
rect -1241 -2491 -1187 148
rect -1101 -2388 -1049 148
rect -914 -69 -862 -60
rect -914 -690 -862 -121
rect 149 -193 201 -183
rect 426 -193 478 -183
rect 617 -193 669 -183
rect 809 -193 861 -183
rect 1001 -193 1053 -183
rect 1194 -192 1246 -182
rect -461 -245 149 -193
rect 201 -245 426 -193
rect 478 -245 617 -193
rect 669 -245 809 -193
rect 861 -245 1001 -193
rect 1053 -244 1194 -193
rect 1386 -192 1438 -182
rect 1246 -244 1386 -193
rect 1670 -193 1722 -183
rect 1947 -193 1999 -183
rect 2138 -193 2190 -183
rect 2330 -193 2382 -183
rect 2522 -193 2574 -183
rect 2715 -192 2767 -182
rect 1438 -244 1670 -193
rect 1053 -245 1670 -244
rect 1722 -245 1947 -193
rect 1999 -245 2138 -193
rect 2190 -245 2330 -193
rect 2382 -245 2522 -193
rect 2574 -244 2715 -193
rect 2907 -192 2959 -182
rect 2767 -244 2907 -193
rect 2959 -244 2966 -193
rect 2574 -245 2966 -244
rect -461 -584 -409 -245
rect 149 -255 201 -245
rect 426 -255 478 -245
rect 617 -255 669 -245
rect 809 -255 861 -245
rect 1001 -255 1053 -245
rect 1194 -254 1246 -245
rect 1386 -254 1438 -245
rect 1670 -255 1722 -245
rect 1947 -255 1999 -245
rect 2138 -255 2190 -245
rect 2330 -255 2382 -245
rect 2522 -255 2574 -245
rect 2715 -254 2767 -245
rect 2907 -254 2959 -245
rect -461 -646 -409 -636
rect 1650 -423 1702 -413
rect -914 -752 -862 -742
rect -549 -694 -497 -684
rect -497 -746 -426 -694
rect -549 -756 -426 -746
rect -478 -1000 -426 -756
rect 1650 -990 1702 -475
rect 149 -1000 201 -990
rect 426 -1000 478 -990
rect 619 -1000 671 -990
rect 810 -1000 862 -990
rect 1002 -1000 1054 -990
rect 1194 -1000 1246 -990
rect 1386 -1000 1438 -990
rect 1650 -1000 1722 -990
rect 1947 -1000 1999 -990
rect 2140 -1000 2192 -990
rect 2331 -1000 2383 -990
rect 2523 -1000 2575 -990
rect 2715 -1000 2767 -990
rect 2907 -1000 2959 -990
rect -478 -1052 149 -1000
rect 201 -1052 426 -1000
rect 478 -1052 619 -1000
rect 671 -1052 810 -1000
rect 862 -1052 1002 -1000
rect 1054 -1052 1194 -1000
rect 1246 -1052 1386 -1000
rect 1438 -1052 1670 -1000
rect 1722 -1052 1947 -1000
rect 1999 -1052 2140 -1000
rect 2192 -1052 2331 -1000
rect 2383 -1052 2523 -1000
rect 2575 -1052 2715 -1000
rect 2767 -1052 2907 -1000
rect 2959 -1052 2966 -1000
rect -478 -1669 -426 -1052
rect 149 -1062 201 -1052
rect 426 -1062 478 -1052
rect 619 -1062 671 -1052
rect 810 -1062 862 -1052
rect 1002 -1062 1054 -1052
rect 1194 -1062 1246 -1052
rect 1386 -1062 1438 -1052
rect 1670 -1062 1722 -1052
rect 1947 -1062 1999 -1052
rect 2140 -1062 2192 -1052
rect 2331 -1062 2383 -1052
rect 2523 -1062 2575 -1052
rect 2715 -1062 2767 -1052
rect 2907 -1062 2959 -1052
rect 98 -1188 150 -1178
rect -478 -1731 -426 -1721
rect -287 -1303 -235 -1293
rect -592 -1776 -540 -1766
rect -1101 -2450 -1049 -2440
rect -872 -1919 -820 -1909
rect -1241 -2543 -1240 -2491
rect -1188 -2543 -1187 -2491
rect -1241 -2864 -1187 -2543
rect -1098 -2864 -1046 -2855
rect -872 -2864 -820 -1971
rect -592 -2225 -540 -1828
rect -416 -1779 -364 -1769
rect -416 -1919 -364 -1831
rect -416 -1981 -364 -1971
rect -1241 -2865 -1045 -2864
rect -1241 -2917 -1098 -2865
rect -1046 -2917 -1045 -2865
rect -1241 -2918 -1045 -2917
rect -1241 -3485 -1187 -2918
rect -1098 -2927 -1046 -2918
rect -872 -2926 -820 -2916
rect -762 -2388 -710 -2378
rect -762 -2775 -710 -2440
rect -592 -2390 -540 -2277
rect -287 -2261 -235 -1355
rect 98 -1517 150 -1240
rect 98 -1527 201 -1517
rect 426 -1527 478 -1517
rect 617 -1527 669 -1517
rect 809 -1527 861 -1517
rect 1001 -1527 1053 -1517
rect 1194 -1526 1246 -1516
rect 98 -1579 149 -1527
rect 201 -1579 426 -1527
rect 478 -1579 617 -1527
rect 669 -1579 809 -1527
rect 861 -1579 1001 -1527
rect 1053 -1578 1194 -1527
rect 1386 -1526 1438 -1516
rect 1246 -1578 1386 -1527
rect 1670 -1527 1722 -1517
rect 1947 -1527 1999 -1517
rect 2138 -1527 2190 -1517
rect 2330 -1527 2382 -1517
rect 2522 -1527 2574 -1517
rect 2715 -1526 2767 -1516
rect 1438 -1578 1670 -1527
rect 1053 -1579 1670 -1578
rect 1722 -1579 1947 -1527
rect 1999 -1579 2138 -1527
rect 2190 -1579 2330 -1527
rect 2382 -1579 2522 -1527
rect 2574 -1578 2715 -1527
rect 2907 -1526 2959 -1516
rect 2767 -1578 2907 -1527
rect 2959 -1578 2966 -1527
rect 2574 -1579 2966 -1578
rect 98 -1589 201 -1579
rect 426 -1589 478 -1579
rect 617 -1589 669 -1579
rect 809 -1589 861 -1579
rect 1001 -1589 1053 -1579
rect 1194 -1588 1246 -1579
rect 1386 -1588 1438 -1579
rect 1670 -1589 1722 -1579
rect 1947 -1589 1999 -1579
rect 2138 -1589 2190 -1579
rect 2330 -1589 2382 -1579
rect 2522 -1589 2574 -1579
rect 2715 -1588 2767 -1579
rect 2907 -1588 2959 -1579
rect 1650 -1757 1702 -1747
rect -235 -2313 148 -2261
rect -287 -2323 -235 -2313
rect 96 -2324 148 -2313
rect 1650 -2324 1702 -1809
rect 96 -2334 201 -2324
rect 426 -2334 478 -2324
rect 619 -2334 671 -2324
rect 810 -2334 862 -2324
rect 1002 -2334 1054 -2324
rect 1194 -2334 1246 -2324
rect 1386 -2334 1438 -2324
rect 1650 -2334 1722 -2324
rect 1947 -2334 1999 -2324
rect 2140 -2334 2192 -2324
rect 2331 -2334 2383 -2324
rect 2523 -2334 2575 -2324
rect 2715 -2334 2767 -2324
rect 2907 -2334 2959 -2324
rect -592 -2450 -540 -2442
rect -412 -2385 -360 -2375
rect 96 -2386 149 -2334
rect 201 -2386 426 -2334
rect 478 -2386 619 -2334
rect 671 -2386 810 -2334
rect 862 -2386 1002 -2334
rect 1054 -2386 1194 -2334
rect 1246 -2386 1386 -2334
rect 1438 -2386 1670 -2334
rect 1722 -2386 1947 -2334
rect 1999 -2386 2140 -2334
rect 2192 -2386 2331 -2334
rect 2383 -2386 2523 -2334
rect 2575 -2386 2715 -2334
rect 2767 -2386 2907 -2334
rect 2959 -2386 2966 -2334
rect 96 -2397 201 -2386
rect 426 -2396 478 -2386
rect 619 -2396 671 -2386
rect 810 -2396 862 -2386
rect 1002 -2396 1054 -2386
rect 1194 -2396 1246 -2386
rect 1386 -2396 1438 -2386
rect 1670 -2396 1722 -2386
rect 1947 -2396 1999 -2386
rect 2140 -2396 2192 -2386
rect 2331 -2396 2383 -2386
rect 2523 -2396 2575 -2386
rect 2715 -2396 2767 -2386
rect 2907 -2396 2959 -2386
rect -412 -2491 -360 -2437
rect -412 -2553 -360 -2543
rect -762 -3393 -710 -2827
rect -412 -2775 -360 -2765
rect -412 -2866 -360 -2827
rect 149 -2905 201 -2895
rect 426 -2905 478 -2895
rect 617 -2905 669 -2895
rect 809 -2905 861 -2895
rect 1001 -2905 1053 -2895
rect 1194 -2904 1246 -2894
rect -412 -2928 -360 -2918
rect -81 -2957 149 -2905
rect 201 -2957 426 -2905
rect 478 -2957 617 -2905
rect 669 -2957 809 -2905
rect 861 -2957 1001 -2905
rect 1053 -2956 1194 -2905
rect 1386 -2904 1438 -2894
rect 1246 -2956 1386 -2905
rect 1670 -2905 1722 -2895
rect 1947 -2905 1999 -2895
rect 2138 -2905 2190 -2895
rect 2330 -2905 2382 -2895
rect 2522 -2905 2574 -2895
rect 2715 -2904 2767 -2894
rect 1438 -2956 1670 -2905
rect 1053 -2957 1670 -2956
rect 1722 -2957 1947 -2905
rect 1999 -2957 2138 -2905
rect 2190 -2957 2330 -2905
rect 2382 -2957 2522 -2905
rect 2574 -2956 2715 -2905
rect 2907 -2904 2959 -2894
rect 2767 -2956 2907 -2905
rect 2959 -2956 2966 -2905
rect 2574 -2957 2966 -2956
rect -236 -3026 -184 -3016
rect -762 -3475 -710 -3445
rect -414 -3393 -362 -3383
rect -414 -3474 -362 -3445
rect -414 -3536 -362 -3526
rect -1241 -3549 -1187 -3539
rect -1416 -4346 -1364 -4336
rect -500 -3580 -448 -3570
rect -500 -4555 -448 -3632
rect -236 -3702 -184 -3078
rect -236 -3712 -183 -3702
rect -236 -3764 -235 -3712
rect -236 -3774 -183 -3764
rect -236 -3951 -184 -3774
rect -236 -4013 -184 -4003
rect -81 -4111 -29 -2957
rect 149 -2967 201 -2957
rect 426 -2967 478 -2957
rect 617 -2967 669 -2957
rect 809 -2967 861 -2957
rect 1001 -2967 1053 -2957
rect 1194 -2966 1246 -2957
rect 1386 -2966 1438 -2957
rect 1670 -2967 1722 -2957
rect 1947 -2967 1999 -2957
rect 2138 -2967 2190 -2957
rect 2330 -2967 2382 -2957
rect 2522 -2967 2574 -2957
rect 2715 -2966 2767 -2957
rect 2907 -2966 2959 -2957
rect 1650 -3135 1702 -3125
rect 1650 -3702 1702 -3187
rect 149 -3712 201 -3702
rect 426 -3712 478 -3702
rect 619 -3712 671 -3702
rect 810 -3712 862 -3702
rect 1002 -3712 1054 -3702
rect 1194 -3712 1246 -3702
rect 1386 -3712 1438 -3702
rect 1650 -3712 1722 -3702
rect 1947 -3712 1999 -3702
rect 2140 -3712 2192 -3702
rect 2331 -3712 2383 -3702
rect 2523 -3712 2575 -3702
rect 2715 -3712 2767 -3702
rect 2907 -3712 2959 -3702
rect 201 -3764 426 -3712
rect 478 -3764 619 -3712
rect 671 -3764 810 -3712
rect 862 -3764 1002 -3712
rect 1054 -3764 1194 -3712
rect 1246 -3764 1386 -3712
rect 1438 -3764 1670 -3712
rect 1722 -3764 1947 -3712
rect 1999 -3764 2140 -3712
rect 2192 -3764 2331 -3712
rect 2383 -3764 2523 -3712
rect 2575 -3764 2715 -3712
rect 2767 -3764 2907 -3712
rect 2959 -3764 2966 -3712
rect 149 -3774 201 -3764
rect 426 -3774 478 -3764
rect 619 -3774 671 -3764
rect 810 -3774 862 -3764
rect 1002 -3774 1054 -3764
rect 1194 -3774 1246 -3764
rect 1386 -3774 1438 -3764
rect 1670 -3774 1722 -3764
rect 1947 -3774 1999 -3764
rect 2140 -3774 2192 -3764
rect 2331 -3774 2383 -3764
rect 2523 -3774 2575 -3764
rect 2715 -3774 2767 -3764
rect 2907 -3774 2959 -3764
rect -81 -4173 -29 -4163
rect 92 -4283 201 -4273
rect 426 -4283 478 -4273
rect 617 -4283 669 -4273
rect 809 -4283 861 -4273
rect 1001 -4283 1053 -4273
rect 1194 -4282 1246 -4272
rect 92 -4335 149 -4283
rect 201 -4335 426 -4283
rect 478 -4335 617 -4283
rect 669 -4335 809 -4283
rect 861 -4335 1001 -4283
rect 1053 -4334 1194 -4283
rect 1386 -4282 1438 -4272
rect 1246 -4334 1386 -4283
rect 1670 -4283 1722 -4273
rect 1947 -4283 1999 -4273
rect 2138 -4283 2190 -4273
rect 2330 -4283 2382 -4273
rect 2522 -4283 2574 -4273
rect 2715 -4282 2767 -4272
rect 1438 -4334 1670 -4283
rect 1053 -4335 1670 -4334
rect 1722 -4335 1947 -4283
rect 1999 -4335 2138 -4283
rect 2190 -4335 2330 -4283
rect 2382 -4335 2522 -4283
rect 2574 -4334 2715 -4283
rect 2907 -4282 2959 -4272
rect 2767 -4334 2907 -4283
rect 2959 -4334 2966 -4283
rect 2574 -4335 2966 -4334
rect 92 -4345 201 -4335
rect 426 -4345 478 -4335
rect 617 -4345 669 -4335
rect 809 -4345 861 -4335
rect 1001 -4345 1053 -4335
rect 1194 -4344 1246 -4335
rect 1386 -4344 1438 -4335
rect 1670 -4345 1722 -4335
rect 1947 -4345 1999 -4335
rect 2138 -4345 2190 -4335
rect 2330 -4345 2382 -4335
rect 2522 -4345 2574 -4335
rect 2715 -4344 2767 -4335
rect 2907 -4344 2959 -4335
rect 92 -4409 144 -4345
rect 92 -4471 144 -4461
rect -548 -4565 -448 -4555
rect -496 -4617 -448 -4565
rect -548 -4627 -448 -4617
rect -3350 -5143 -3125 -5091
rect -3073 -5143 -2934 -5091
rect -2882 -5143 -2742 -5091
rect -2690 -5143 -2550 -5091
rect -2498 -5092 -1535 -5091
rect -2498 -5143 -2357 -5092
rect -3402 -5153 -3350 -5143
rect -3125 -5153 -3073 -5143
rect -2934 -5153 -2882 -5143
rect -2742 -5153 -2690 -5143
rect -2550 -5153 -2498 -5143
rect -2305 -5143 -2165 -5092
rect -2357 -5154 -2305 -5144
rect -2113 -5143 -1535 -5092
rect -500 -5089 -448 -4627
rect 1650 -4513 1702 -4503
rect 1650 -5080 1702 -4565
rect 149 -5089 201 -5080
rect -500 -5090 203 -5089
rect 426 -5090 478 -5080
rect 619 -5090 671 -5080
rect 810 -5090 862 -5080
rect 1002 -5090 1054 -5080
rect 1194 -5090 1246 -5080
rect 1386 -5090 1438 -5080
rect 1650 -5090 1722 -5080
rect 1947 -5090 1999 -5080
rect 2140 -5090 2192 -5080
rect 2331 -5090 2383 -5080
rect 2523 -5090 2575 -5080
rect 2715 -5090 2767 -5080
rect 2907 -5090 2959 -5080
rect -500 -5141 149 -5090
rect -2165 -5154 -2113 -5144
rect -1587 -5148 -1535 -5143
rect 201 -5142 426 -5090
rect 478 -5142 619 -5090
rect 671 -5142 810 -5090
rect 862 -5142 1002 -5090
rect 1054 -5142 1194 -5090
rect 1246 -5142 1386 -5090
rect 1438 -5142 1670 -5090
rect 1722 -5142 1947 -5090
rect 1999 -5142 2140 -5090
rect 2192 -5142 2331 -5090
rect 2383 -5142 2523 -5090
rect 2575 -5142 2715 -5090
rect 2767 -5142 2907 -5090
rect 2959 -5142 2966 -5090
rect 149 -5152 201 -5142
rect 426 -5152 478 -5142
rect 619 -5152 671 -5142
rect 810 -5152 862 -5142
rect 1002 -5152 1054 -5142
rect 1194 -5152 1246 -5142
rect 1386 -5152 1438 -5142
rect 1670 -5152 1722 -5142
rect 1947 -5152 1999 -5142
rect 2140 -5152 2192 -5142
rect 2331 -5152 2383 -5142
rect 2523 -5152 2575 -5142
rect 2715 -5152 2767 -5142
rect 2907 -5152 2959 -5142
<< labels >>
flabel metal1 -3682 -716 -3682 -716 1 FreeSans 400 0 0 0 in0
port 4 n
flabel metal1 -3684 -2051 -3684 -2051 1 FreeSans 400 0 0 0 in1
port 5 n
flabel metal1 -3682 -3429 -3682 -3429 1 FreeSans 400 0 0 0 in2
port 6 n
flabel metal1 -3683 -4808 -3683 -4808 1 FreeSans 400 0 0 0 in3
port 7 n
flabel metal1 1525 -1212 1525 -1212 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 3046 -1214 3046 -1214 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 1527 -1369 1527 -1369 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 3048 -1371 3048 -1371 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 1527 -2546 1527 -2546 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 3048 -2550 3048 -2550 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 3048 -2746 3048 -2746 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 1527 -2744 1527 -2744 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 1525 -3926 1525 -3926 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 3049 -3925 3049 -3925 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 1525 -4130 1525 -4130 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 3049 -4128 3049 -4128 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 1523 -5306 1523 -5306 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 3045 -5302 3045 -5302 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 3438 -2641 3438 -2641 1 FreeSans 400 0 0 0 out
port 8 n
flabel metal2 -1562 128 -1562 128 1 FreeSans 400 0 0 0 en
port 1 n
flabel metal2 -1216 128 -1216 128 1 FreeSans 400 0 0 0 s1
port 2 n
flabel metal2 -1073 128 -1073 128 1 FreeSans 400 0 0 0 s0
port 3 n
flabel metal1 -1030 -478 -1030 -478 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -1037 -1022 -1037 -1022 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -752 -1566 -752 -1566 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -1314 -2113 -1314 -2113 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -1303 -2653 -1303 -2653 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -1315 -3203 -1315 -3203 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -767 -3742 -767 -3742 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -769 -4286 -769 -4286 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -748 -4830 -748 -4830 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -2025 -77 -2025 -77 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -2025 -1170 -2025 -1170 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -2025 -1408 -2025 -1408 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -2025 -2505 -2025 -2505 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -2025 -2787 -2025 -2787 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -2025 -3884 -2025 -3884 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 -2028 -4172 -2028 -4172 1 FreeSans 400 0 0 0 VDD
port 9 n power bidirectional
flabel metal1 -2026 -5260 -2026 -5260 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 1528 -56 1528 -56 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel metal1 3048 -56 3048 -56 1 FreeSans 400 0 0 0 VSS
port 10 n power bidirectional
flabel locali -448 -4064 -414 -4030 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_5/Y
flabel locali -448 -3996 -414 -3962 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_5/Y
flabel locali -540 -3996 -506 -3962 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_5/A
flabel nwell -583 -4302 -549 -4268 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VPB
flabel pwell -583 -3758 -549 -3724 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VNB
flabel metal1 -583 -3758 -549 -3724 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VGND
flabel metal1 -583 -4302 -549 -4268 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_5/VPWR
rlabel comment -612 -3741 -612 -3741 2 sky130_fd_sc_hd__inv_1_5/inv_1
rlabel metal1 -612 -3789 -336 -3693 5 sky130_fd_sc_hd__inv_1_5/VGND
rlabel metal1 -612 -4333 -336 -4237 5 sky130_fd_sc_hd__inv_1_5/VPWR
flabel locali -448 -4540 -414 -4506 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_6/Y
flabel locali -448 -4608 -414 -4574 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_6/Y
flabel locali -540 -4608 -506 -4574 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_6/A
flabel nwell -583 -4302 -549 -4268 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VPB
flabel pwell -583 -4846 -549 -4812 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VNB
flabel metal1 -583 -4846 -549 -4812 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VGND
flabel metal1 -583 -4302 -549 -4268 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_6/VPWR
rlabel comment -612 -4829 -612 -4829 4 sky130_fd_sc_hd__inv_1_6/inv_1
rlabel metal1 -612 -4877 -336 -4781 1 sky130_fd_sc_hd__inv_1_6/VGND
rlabel metal1 -612 -4333 -336 -4237 1 sky130_fd_sc_hd__inv_1_6/VPWR
flabel metal1 -687 -4294 -634 -4265 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VPWR
flabel metal1 -684 -3761 -633 -3723 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VGND
rlabel comment -612 -3741 -612 -3741 8 sky130_fd_sc_hd__tapvpwrvgnd_1_6/tapvpwrvgnd_1
rlabel metal1 -704 -3789 -612 -3693 5 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VGND
rlabel metal1 -704 -4333 -612 -4237 5 sky130_fd_sc_hd__tapvpwrvgnd_1_6/VPWR
flabel metal1 -682 -4305 -629 -4276 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VPWR
flabel metal1 -683 -4847 -632 -4809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VGND
rlabel comment -704 -4829 -704 -4829 4 sky130_fd_sc_hd__tapvpwrvgnd_1_7/tapvpwrvgnd_1
rlabel metal1 -704 -4877 -612 -4781 1 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VGND
rlabel metal1 -704 -4333 -612 -4237 1 sky130_fd_sc_hd__tapvpwrvgnd_1_7/VPWR
flabel metal1 -3424 -4310 -3424 -4310 3 FreeSans 400 0 0 0 transmission_gate_3/en_b
flabel metal1 -3425 -4806 -3425 -4806 3 FreeSans 400 0 0 0 transmission_gate_3/in
flabel metal1 -3425 -5117 -3425 -5117 3 FreeSans 400 0 0 0 transmission_gate_3/en
flabel metal1 -1934 -4807 -1934 -4807 7 FreeSans 400 0 0 0 transmission_gate_3/out
flabel metal1 -2025 -4161 -2025 -4161 5 FreeSans 400 0 0 0 transmission_gate_3/VDD
flabel metal1 -2025 -5267 -2025 -5267 1 FreeSans 400 0 0 0 transmission_gate_3/VSS
flabel metal1 1526 -5305 1526 -5305 5 FreeSans 400 0 0 0 switch_5t_3/VDD
flabel metal1 1526 -4123 1526 -4123 5 FreeSans 400 0 0 0 switch_5t_3/VSS
flabel metal1 80 -5115 80 -5115 5 FreeSans 400 0 0 0 switch_5t_3/en_b
flabel metal1 78 -4309 78 -4309 5 FreeSans 400 0 0 0 switch_5t_3/en
flabel metal1 79 -4620 79 -4620 5 FreeSans 400 0 0 0 switch_5t_3/in
flabel metal1 3174 -4619 3174 -4619 7 FreeSans 400 0 0 0 switch_5t_3/out
flabel metal1 3047 -5306 3047 -5306 5 FreeSans 400 0 0 0 switch_5t_3/VDD
flabel metal1 3047 -4124 3047 -4124 5 FreeSans 400 0 0 0 switch_5t_3/VSS
flabel metal1 1648 -5116 1648 -5116 3 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_1/en_b
flabel metal1 1647 -4620 1647 -4620 3 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_1/in
flabel metal1 1647 -4309 1647 -4309 3 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_1/en
flabel metal1 3138 -4619 3138 -4619 7 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_1/out
flabel metal1 3047 -5265 3047 -5265 1 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_1/VDD
flabel metal1 3047 -4159 3047 -4159 5 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_1/VSS
flabel metal1 127 -5116 127 -5116 3 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_0/en_b
flabel metal1 126 -4620 126 -4620 3 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_0/in
flabel metal1 126 -4309 126 -4309 3 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_0/en
flabel metal1 1617 -4619 1617 -4619 7 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_0/out
flabel metal1 1526 -5265 1526 -5265 1 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_0/VDD
flabel metal1 1526 -4159 1526 -4159 5 FreeSans 400 0 0 0 switch_5t_3/transmission_gate_0/VSS
flabel metal1 -777 -2671 -724 -2639 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VGND
flabel metal1 -777 -3214 -725 -3183 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VPWR
flabel nwell -766 -3206 -732 -3188 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VPB
flabel pwell -767 -2665 -735 -2643 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_0/VNB
rlabel comment -704 -2653 -704 -2653 8 sky130_fd_sc_hd__fill_2_0/fill_2
rlabel metal1 -888 -2701 -704 -2605 5 sky130_fd_sc_hd__fill_2_0/VGND
rlabel metal1 -888 -3245 -704 -3149 5 sky130_fd_sc_hd__fill_2_0/VPWR
flabel locali -1000 -2976 -966 -2942 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -1000 -2908 -966 -2874 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/Y
flabel locali -1092 -2908 -1058 -2874 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_0/A
flabel nwell -1135 -3214 -1101 -3180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPB
flabel pwell -1135 -2670 -1101 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VNB
flabel metal1 -1135 -2670 -1101 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VGND
flabel metal1 -1135 -3214 -1101 -3180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_0/VPWR
rlabel comment -1164 -2653 -1164 -2653 2 sky130_fd_sc_hd__inv_1_0/inv_1
rlabel metal1 -1164 -2701 -888 -2605 5 sky130_fd_sc_hd__inv_1_0/VGND
rlabel metal1 -1164 -3245 -888 -3149 5 sky130_fd_sc_hd__inv_1_0/VPWR
flabel locali -492 -3656 -458 -3622 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali -492 -3588 -458 -3554 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali -492 -3520 -458 -3486 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/Y
flabel locali -584 -3520 -550 -3486 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/B
flabel locali -400 -3520 -366 -3486 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_0/A
flabel nwell -584 -3214 -550 -3180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPB
flabel pwell -584 -3758 -550 -3724 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VNB
flabel metal1 -584 -3758 -550 -3724 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VGND
flabel metal1 -584 -3214 -550 -3180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_0/VPWR
rlabel comment -612 -3741 -612 -3741 4 sky130_fd_sc_hd__nand2_1_0/nand2_1
rlabel metal1 -612 -3789 -336 -3693 1 sky130_fd_sc_hd__nand2_1_0/VGND
rlabel metal1 -612 -3245 -336 -3149 1 sky130_fd_sc_hd__nand2_1_0/VPWR
flabel locali -492 -2772 -458 -2738 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali -492 -2840 -458 -2806 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali -492 -2908 -458 -2874 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/Y
flabel locali -584 -2908 -550 -2874 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/B
flabel locali -400 -2908 -366 -2874 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_1/A
flabel nwell -584 -3214 -550 -3180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VPB
flabel pwell -584 -2670 -550 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VNB
flabel metal1 -584 -2670 -550 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VGND
flabel metal1 -584 -3214 -550 -3180 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_1/VPWR
rlabel comment -612 -2653 -612 -2653 2 sky130_fd_sc_hd__nand2_1_1/nand2_1
rlabel metal1 -612 -2701 -336 -2605 5 sky130_fd_sc_hd__nand2_1_1/VGND
rlabel metal1 -612 -3245 -336 -3149 5 sky130_fd_sc_hd__nand2_1_1/VPWR
flabel metal1 -1239 -3206 -1186 -3177 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -1236 -2673 -1185 -2635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel comment -1164 -2653 -1164 -2653 8 sky130_fd_sc_hd__tapvpwrvgnd_1_0/tapvpwrvgnd_1
rlabel metal1 -1256 -2701 -1164 -2605 5 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VGND
rlabel metal1 -1256 -3245 -1164 -3149 5 sky130_fd_sc_hd__tapvpwrvgnd_1_0/VPWR
flabel metal1 -682 -3217 -629 -3188 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 -683 -3759 -632 -3721 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel comment -704 -3741 -704 -3741 4 sky130_fd_sc_hd__tapvpwrvgnd_1_3/tapvpwrvgnd_1
rlabel metal1 -704 -3789 -612 -3693 1 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VGND
rlabel metal1 -704 -3245 -612 -3149 1 sky130_fd_sc_hd__tapvpwrvgnd_1_3/VPWR
flabel metal1 -687 -3206 -634 -3177 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VPWR
flabel metal1 -684 -2673 -633 -2635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VGND
rlabel comment -612 -2653 -612 -2653 8 sky130_fd_sc_hd__tapvpwrvgnd_1_8/tapvpwrvgnd_1
rlabel metal1 -704 -2701 -612 -2605 5 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VGND
rlabel metal1 -704 -3245 -612 -3149 5 sky130_fd_sc_hd__tapvpwrvgnd_1_8/VPWR
flabel metal1 -3424 -2932 -3424 -2932 3 FreeSans 400 0 0 0 transmission_gate_2/en_b
flabel metal1 -3425 -3428 -3425 -3428 3 FreeSans 400 0 0 0 transmission_gate_2/in
flabel metal1 -3425 -3739 -3425 -3739 3 FreeSans 400 0 0 0 transmission_gate_2/en
flabel metal1 -1934 -3429 -1934 -3429 7 FreeSans 400 0 0 0 transmission_gate_2/out
flabel metal1 -2025 -2783 -2025 -2783 5 FreeSans 400 0 0 0 transmission_gate_2/VDD
flabel metal1 -2025 -3889 -2025 -3889 1 FreeSans 400 0 0 0 transmission_gate_2/VSS
flabel metal1 1526 -3927 1526 -3927 5 FreeSans 400 0 0 0 switch_5t_2/VDD
flabel metal1 1526 -2745 1526 -2745 5 FreeSans 400 0 0 0 switch_5t_2/VSS
flabel metal1 80 -3737 80 -3737 5 FreeSans 400 0 0 0 switch_5t_2/en_b
flabel metal1 78 -2931 78 -2931 5 FreeSans 400 0 0 0 switch_5t_2/en
flabel metal1 79 -3242 79 -3242 5 FreeSans 400 0 0 0 switch_5t_2/in
flabel metal1 3174 -3241 3174 -3241 7 FreeSans 400 0 0 0 switch_5t_2/out
flabel metal1 3047 -3928 3047 -3928 5 FreeSans 400 0 0 0 switch_5t_2/VDD
flabel metal1 3047 -2746 3047 -2746 5 FreeSans 400 0 0 0 switch_5t_2/VSS
flabel metal1 1648 -3738 1648 -3738 3 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_1/en_b
flabel metal1 1647 -3242 1647 -3242 3 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_1/in
flabel metal1 1647 -2931 1647 -2931 3 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_1/en
flabel metal1 3138 -3241 3138 -3241 7 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_1/out
flabel metal1 3047 -3887 3047 -3887 1 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_1/VDD
flabel metal1 3047 -2781 3047 -2781 5 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_1/VSS
flabel metal1 127 -3738 127 -3738 3 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_0/en_b
flabel metal1 126 -3242 126 -3242 3 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_0/in
flabel metal1 126 -2931 126 -2931 3 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_0/en
flabel metal1 1617 -3241 1617 -3241 7 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_0/out
flabel metal1 1526 -3887 1526 -3887 1 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_0/VDD
flabel metal1 1526 -2781 1526 -2781 5 FreeSans 400 0 0 0 switch_5t_2/transmission_gate_0/VSS
flabel metal1 -868 -2667 -815 -2635 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VGND
flabel metal1 -867 -2123 -815 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VPWR
flabel nwell -860 -2118 -826 -2100 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VPB
flabel pwell -857 -2663 -825 -2641 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__fill_2_1/VNB
rlabel comment -888 -2653 -888 -2653 4 sky130_fd_sc_hd__fill_2_1/fill_2
rlabel metal1 -888 -2701 -704 -2605 1 sky130_fd_sc_hd__fill_2_1/VGND
rlabel metal1 -888 -2157 -704 -2061 1 sky130_fd_sc_hd__fill_2_1/VPWR
flabel locali -1000 -2364 -966 -2330 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali -1000 -2432 -966 -2398 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/Y
flabel locali -1092 -2432 -1058 -2398 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_1/A
flabel nwell -1135 -2126 -1101 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPB
flabel pwell -1135 -2670 -1101 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VNB
flabel metal1 -1135 -2670 -1101 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VGND
flabel metal1 -1135 -2126 -1101 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_1/VPWR
rlabel comment -1164 -2653 -1164 -2653 4 sky130_fd_sc_hd__inv_1_1/inv_1
rlabel metal1 -1164 -2701 -888 -2605 1 sky130_fd_sc_hd__inv_1_1/VGND
rlabel metal1 -1164 -2157 -888 -2061 1 sky130_fd_sc_hd__inv_1_1/VPWR
flabel locali -492 -2568 -458 -2534 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/Y
flabel locali -492 -2500 -458 -2466 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/Y
flabel locali -492 -2432 -458 -2398 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/Y
flabel locali -584 -2432 -550 -2398 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/B
flabel locali -400 -2432 -366 -2398 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_2/A
flabel nwell -584 -2126 -550 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VPB
flabel pwell -584 -2670 -550 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VNB
flabel metal1 -584 -2670 -550 -2636 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VGND
flabel metal1 -584 -2126 -550 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_2/VPWR
rlabel comment -612 -2653 -612 -2653 4 sky130_fd_sc_hd__nand2_1_2/nand2_1
rlabel metal1 -612 -2701 -336 -2605 1 sky130_fd_sc_hd__nand2_1_2/VGND
rlabel metal1 -612 -2157 -336 -2061 1 sky130_fd_sc_hd__nand2_1_2/VPWR
flabel locali -492 -1684 -458 -1650 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/Y
flabel locali -492 -1752 -458 -1718 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/Y
flabel locali -492 -1820 -458 -1786 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/Y
flabel locali -584 -1820 -550 -1786 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/B
flabel locali -400 -1820 -366 -1786 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__nand2_1_3/A
flabel nwell -584 -2126 -550 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VPB
flabel pwell -584 -1582 -550 -1548 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VNB
flabel metal1 -584 -1582 -550 -1548 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VGND
flabel metal1 -584 -2126 -550 -2092 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__nand2_1_3/VPWR
rlabel comment -612 -1565 -612 -1565 2 sky130_fd_sc_hd__nand2_1_3/nand2_1
rlabel metal1 -612 -1613 -336 -1517 5 sky130_fd_sc_hd__nand2_1_3/VGND
rlabel metal1 -612 -2157 -336 -2061 5 sky130_fd_sc_hd__nand2_1_3/VPWR
flabel metal1 -1234 -2129 -1181 -2100 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -1235 -2671 -1184 -2633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel comment -1256 -2653 -1256 -2653 4 sky130_fd_sc_hd__tapvpwrvgnd_1_1/tapvpwrvgnd_1
rlabel metal1 -1256 -2701 -1164 -2605 1 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VGND
rlabel metal1 -1256 -2157 -1164 -2061 1 sky130_fd_sc_hd__tapvpwrvgnd_1_1/VPWR
flabel metal1 -687 -2118 -634 -2089 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 -684 -1585 -633 -1547 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel comment -612 -1565 -612 -1565 8 sky130_fd_sc_hd__tapvpwrvgnd_1_2/tapvpwrvgnd_1
rlabel metal1 -704 -1613 -612 -1517 5 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VGND
rlabel metal1 -704 -2157 -612 -2061 5 sky130_fd_sc_hd__tapvpwrvgnd_1_2/VPWR
flabel metal1 -682 -2129 -629 -2100 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VPWR
flabel metal1 -683 -2671 -632 -2633 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VGND
rlabel comment -704 -2653 -704 -2653 4 sky130_fd_sc_hd__tapvpwrvgnd_1_9/tapvpwrvgnd_1
rlabel metal1 -704 -2701 -612 -2605 1 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VGND
rlabel metal1 -704 -2157 -612 -2061 1 sky130_fd_sc_hd__tapvpwrvgnd_1_9/VPWR
flabel metal1 -3424 -1554 -3424 -1554 3 FreeSans 400 0 0 0 transmission_gate_1/en_b
flabel metal1 -3425 -2050 -3425 -2050 3 FreeSans 400 0 0 0 transmission_gate_1/in
flabel metal1 -3425 -2361 -3425 -2361 3 FreeSans 400 0 0 0 transmission_gate_1/en
flabel metal1 -1934 -2051 -1934 -2051 7 FreeSans 400 0 0 0 transmission_gate_1/out
flabel metal1 -2025 -1405 -2025 -1405 5 FreeSans 400 0 0 0 transmission_gate_1/VDD
flabel metal1 -2025 -2511 -2025 -2511 1 FreeSans 400 0 0 0 transmission_gate_1/VSS
flabel metal1 1526 -2549 1526 -2549 5 FreeSans 400 0 0 0 switch_5t_0/VDD
flabel metal1 1526 -1367 1526 -1367 5 FreeSans 400 0 0 0 switch_5t_0/VSS
flabel metal1 80 -2359 80 -2359 5 FreeSans 400 0 0 0 switch_5t_0/en_b
flabel metal1 78 -1553 78 -1553 5 FreeSans 400 0 0 0 switch_5t_0/en
flabel metal1 79 -1864 79 -1864 5 FreeSans 400 0 0 0 switch_5t_0/in
flabel metal1 3174 -1863 3174 -1863 7 FreeSans 400 0 0 0 switch_5t_0/out
flabel metal1 3047 -2550 3047 -2550 5 FreeSans 400 0 0 0 switch_5t_0/VDD
flabel metal1 3047 -1368 3047 -1368 5 FreeSans 400 0 0 0 switch_5t_0/VSS
flabel metal1 1648 -2360 1648 -2360 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/en_b
flabel metal1 1647 -1864 1647 -1864 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/in
flabel metal1 1647 -1553 1647 -1553 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/en
flabel metal1 3138 -1863 3138 -1863 7 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/out
flabel metal1 3047 -2509 3047 -2509 1 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/VDD
flabel metal1 3047 -1403 3047 -1403 5 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_1/VSS
flabel metal1 127 -2360 127 -2360 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/en_b
flabel metal1 126 -1864 126 -1864 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/in
flabel metal1 126 -1553 126 -1553 3 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/en
flabel metal1 1617 -1863 1617 -1863 7 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/out
flabel metal1 1526 -2509 1526 -2509 1 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/VDD
flabel metal1 1526 -1403 1526 -1403 5 FreeSans 400 0 0 0 switch_5t_0/transmission_gate_0/VSS
flabel locali -448 -1276 -414 -1242 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/Y
flabel locali -448 -1344 -414 -1310 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/Y
flabel locali -540 -1344 -506 -1310 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_3/A
flabel nwell -583 -1038 -549 -1004 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VPB
flabel pwell -583 -1582 -549 -1548 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VNB
flabel metal1 -583 -1582 -549 -1548 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VGND
flabel metal1 -583 -1038 -549 -1004 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_3/VPWR
rlabel comment -612 -1565 -612 -1565 4 sky130_fd_sc_hd__inv_1_3/inv_1
rlabel metal1 -612 -1613 -336 -1517 1 sky130_fd_sc_hd__inv_1_3/VGND
rlabel metal1 -612 -1069 -336 -973 1 sky130_fd_sc_hd__inv_1_3/VPWR
flabel locali -448 -800 -414 -766 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_4/Y
flabel locali -448 -732 -414 -698 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_4/Y
flabel locali -540 -732 -506 -698 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_4/A
flabel nwell -583 -1038 -549 -1004 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VPB
flabel pwell -583 -494 -549 -460 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VNB
flabel metal1 -583 -494 -549 -460 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VGND
flabel metal1 -583 -1038 -549 -1004 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_4/VPWR
rlabel comment -612 -477 -612 -477 2 sky130_fd_sc_hd__inv_1_4/inv_1
rlabel metal1 -612 -525 -336 -429 5 sky130_fd_sc_hd__inv_1_4/VGND
rlabel metal1 -612 -1069 -336 -973 5 sky130_fd_sc_hd__inv_1_4/VPWR
flabel locali -816 -800 -782 -766 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_8/Y
flabel locali -816 -732 -782 -698 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_8/Y
flabel locali -908 -732 -874 -698 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_1_8/A
flabel nwell -951 -1038 -917 -1004 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VPB
flabel pwell -951 -494 -917 -460 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VNB
flabel metal1 -951 -494 -917 -460 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VGND
flabel metal1 -951 -1038 -917 -1004 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_1_8/VPWR
rlabel comment -980 -477 -980 -477 2 sky130_fd_sc_hd__inv_1_8/inv_1
rlabel metal1 -980 -525 -704 -429 5 sky130_fd_sc_hd__inv_1_8/VGND
rlabel metal1 -980 -1069 -704 -973 5 sky130_fd_sc_hd__inv_1_8/VPWR
flabel metal1 -682 -1041 -629 -1012 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR
flabel metal1 -683 -1583 -632 -1545 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VGND
rlabel comment -704 -1565 -704 -1565 4 sky130_fd_sc_hd__tapvpwrvgnd_1_4/tapvpwrvgnd_1
rlabel metal1 -704 -1613 -612 -1517 1 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VGND
rlabel metal1 -704 -1069 -612 -973 1 sky130_fd_sc_hd__tapvpwrvgnd_1_4/VPWR
flabel metal1 -687 -1030 -634 -1001 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VPWR
flabel metal1 -684 -497 -633 -459 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VGND
rlabel comment -612 -477 -612 -477 8 sky130_fd_sc_hd__tapvpwrvgnd_1_5/tapvpwrvgnd_1
rlabel metal1 -704 -525 -612 -429 5 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VGND
rlabel metal1 -704 -1069 -612 -973 5 sky130_fd_sc_hd__tapvpwrvgnd_1_5/VPWR
flabel metal1 -3424 -220 -3424 -220 3 FreeSans 400 0 0 0 transmission_gate_0/en_b
flabel metal1 -3425 -716 -3425 -716 3 FreeSans 400 0 0 0 transmission_gate_0/in
flabel metal1 -3425 -1027 -3425 -1027 3 FreeSans 400 0 0 0 transmission_gate_0/en
flabel metal1 -1934 -717 -1934 -717 7 FreeSans 400 0 0 0 transmission_gate_0/out
flabel metal1 -2025 -71 -2025 -71 5 FreeSans 400 0 0 0 transmission_gate_0/VDD
flabel metal1 -2025 -1177 -2025 -1177 1 FreeSans 400 0 0 0 transmission_gate_0/VSS
flabel metal1 1526 -1215 1526 -1215 5 FreeSans 400 0 0 0 switch_5t_1/VDD
flabel metal1 1526 -33 1526 -33 5 FreeSans 400 0 0 0 switch_5t_1/VSS
flabel metal1 80 -1025 80 -1025 5 FreeSans 400 0 0 0 switch_5t_1/en_b
flabel metal1 78 -219 78 -219 5 FreeSans 400 0 0 0 switch_5t_1/en
flabel metal1 79 -530 79 -530 5 FreeSans 400 0 0 0 switch_5t_1/in
flabel metal1 3174 -529 3174 -529 7 FreeSans 400 0 0 0 switch_5t_1/out
flabel metal1 3047 -1216 3047 -1216 5 FreeSans 400 0 0 0 switch_5t_1/VDD
flabel metal1 3047 -34 3047 -34 5 FreeSans 400 0 0 0 switch_5t_1/VSS
flabel metal1 1648 -1026 1648 -1026 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/en_b
flabel metal1 1647 -530 1647 -530 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/in
flabel metal1 1647 -219 1647 -219 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/en
flabel metal1 3138 -529 3138 -529 7 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/out
flabel metal1 3047 -1175 3047 -1175 1 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/VDD
flabel metal1 3047 -69 3047 -69 5 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_1/VSS
flabel metal1 127 -1026 127 -1026 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/en_b
flabel metal1 126 -530 126 -530 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/in
flabel metal1 126 -219 126 -219 3 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/en
flabel metal1 1617 -529 1617 -529 7 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/out
flabel metal1 1526 -1175 1526 -1175 1 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/VDD
flabel metal1 1526 -69 1526 -69 5 FreeSans 400 0 0 0 switch_5t_1/transmission_gate_0/VSS
<< end >>
