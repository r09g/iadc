magic
tech sky130A
magscale 1 2
timestamp 1655456512
<< error_p >>
rect 337 466 395 472
rect 757 466 815 472
rect 1177 466 1235 472
rect 1597 466 1655 472
rect 2017 466 2075 472
rect 2437 466 2495 472
rect 2857 466 2915 472
rect 3277 466 3335 472
rect 3697 466 3755 472
rect 4117 466 4175 472
rect 4537 466 4595 472
rect 4957 466 5015 472
rect 5377 466 5435 472
rect 5797 466 5855 472
rect 6217 466 6275 472
rect 6637 466 6695 472
rect 7057 466 7115 472
rect 7477 466 7535 472
rect 7897 466 7955 472
rect 8317 466 8375 472
rect 337 432 349 466
rect 757 432 769 466
rect 1177 432 1189 466
rect 1597 432 1609 466
rect 2017 432 2029 466
rect 2437 432 2449 466
rect 2857 432 2869 466
rect 3277 432 3289 466
rect 3697 432 3709 466
rect 4117 432 4129 466
rect 4537 432 4549 466
rect 4957 432 4969 466
rect 5377 432 5389 466
rect 5797 432 5809 466
rect 6217 432 6229 466
rect 6637 432 6649 466
rect 7057 432 7069 466
rect 7477 432 7489 466
rect 7897 432 7909 466
rect 8317 432 8329 466
rect 337 426 395 432
rect 757 426 815 432
rect 1177 426 1235 432
rect 1597 426 1655 432
rect 2017 426 2075 432
rect 2437 426 2495 432
rect 2857 426 2915 432
rect 3277 426 3335 432
rect 3697 426 3755 432
rect 4117 426 4175 432
rect 4537 426 4595 432
rect 4957 426 5015 432
rect 5377 426 5435 432
rect 5797 426 5855 432
rect 6217 426 6275 432
rect 6637 426 6695 432
rect 7057 426 7115 432
rect 7477 426 7535 432
rect 7897 426 7955 432
rect 8317 426 8375 432
rect 547 138 605 144
rect 967 138 1025 144
rect 1387 138 1445 144
rect 1807 138 1865 144
rect 2227 138 2285 144
rect 2647 138 2705 144
rect 3067 138 3125 144
rect 3487 138 3545 144
rect 3907 138 3965 144
rect 4327 138 4385 144
rect 4747 138 4805 144
rect 5167 138 5225 144
rect 5587 138 5645 144
rect 6007 138 6065 144
rect 6427 138 6485 144
rect 6847 138 6905 144
rect 7267 138 7325 144
rect 7687 138 7745 144
rect 8107 138 8165 144
rect 8527 138 8585 144
rect 547 104 559 138
rect 967 104 979 138
rect 1387 104 1399 138
rect 1807 104 1819 138
rect 2227 104 2239 138
rect 2647 104 2659 138
rect 3067 104 3079 138
rect 3487 104 3499 138
rect 3907 104 3919 138
rect 4327 104 4339 138
rect 4747 104 4759 138
rect 5167 104 5179 138
rect 5587 104 5599 138
rect 6007 104 6019 138
rect 6427 104 6439 138
rect 6847 104 6859 138
rect 7267 104 7279 138
rect 7687 104 7699 138
rect 8107 104 8119 138
rect 8527 104 8539 138
rect 547 98 605 104
rect 967 98 1025 104
rect 1387 98 1445 104
rect 1807 98 1865 104
rect 2227 98 2285 104
rect 2647 98 2705 104
rect 3067 98 3125 104
rect 3487 98 3545 104
rect 3907 98 3965 104
rect 4327 98 4385 104
rect 4747 98 4805 104
rect 5167 98 5225 104
rect 5587 98 5645 104
rect 6007 98 6065 104
rect 6427 98 6485 104
rect 6847 98 6905 104
rect 7267 98 7325 104
rect 7687 98 7745 104
rect 8107 98 8165 104
rect 8527 98 8585 104
rect 339 -66 397 -60
rect 759 -66 817 -60
rect 1179 -66 1237 -60
rect 1599 -66 1657 -60
rect 2019 -66 2077 -60
rect 2439 -66 2497 -60
rect 2859 -66 2917 -60
rect 3279 -66 3337 -60
rect 3699 -66 3757 -60
rect 4119 -66 4177 -60
rect 4539 -66 4597 -60
rect 4959 -66 5017 -60
rect 5379 -66 5437 -60
rect 5799 -66 5857 -60
rect 6219 -66 6277 -60
rect 6639 -66 6697 -60
rect 7059 -66 7117 -60
rect 7479 -66 7537 -60
rect 7899 -66 7957 -60
rect 8319 -66 8377 -60
rect 339 -100 351 -66
rect 759 -100 771 -66
rect 1179 -100 1191 -66
rect 1599 -100 1611 -66
rect 2019 -100 2031 -66
rect 2439 -100 2451 -66
rect 2859 -100 2871 -66
rect 3279 -100 3291 -66
rect 3699 -100 3711 -66
rect 4119 -100 4131 -66
rect 4539 -100 4551 -66
rect 4959 -100 4971 -66
rect 5379 -100 5391 -66
rect 5799 -100 5811 -66
rect 6219 -100 6231 -66
rect 6639 -100 6651 -66
rect 7059 -100 7071 -66
rect 7479 -100 7491 -66
rect 7899 -100 7911 -66
rect 8319 -100 8331 -66
rect 339 -106 397 -100
rect 759 -106 817 -100
rect 1179 -106 1237 -100
rect 1599 -106 1657 -100
rect 2019 -106 2077 -100
rect 2439 -106 2497 -100
rect 2859 -106 2917 -100
rect 3279 -106 3337 -100
rect 3699 -106 3757 -100
rect 4119 -106 4177 -100
rect 4539 -106 4597 -100
rect 4959 -106 5017 -100
rect 5379 -106 5437 -100
rect 5799 -106 5857 -100
rect 6219 -106 6277 -100
rect 6639 -106 6697 -100
rect 7059 -106 7117 -100
rect 7479 -106 7537 -100
rect 7899 -106 7957 -100
rect 8319 -106 8377 -100
rect 549 -395 607 -389
rect 969 -395 1027 -389
rect 1389 -395 1447 -389
rect 1809 -395 1867 -389
rect 2229 -395 2287 -389
rect 2649 -395 2707 -389
rect 3069 -395 3127 -389
rect 3489 -395 3547 -389
rect 3909 -395 3967 -389
rect 4329 -395 4387 -389
rect 4749 -395 4807 -389
rect 5169 -395 5227 -389
rect 5589 -395 5647 -389
rect 6009 -395 6067 -389
rect 6429 -395 6487 -389
rect 6849 -395 6907 -389
rect 7269 -395 7327 -389
rect 7689 -395 7747 -389
rect 8109 -395 8167 -389
rect 8529 -395 8587 -389
rect 549 -429 561 -395
rect 969 -429 981 -395
rect 1389 -429 1401 -395
rect 1809 -429 1821 -395
rect 2229 -429 2241 -395
rect 2649 -429 2661 -395
rect 3069 -429 3081 -395
rect 3489 -429 3501 -395
rect 3909 -429 3921 -395
rect 4329 -429 4341 -395
rect 4749 -429 4761 -395
rect 5169 -429 5181 -395
rect 5589 -429 5601 -395
rect 6009 -429 6021 -395
rect 6429 -429 6441 -395
rect 6849 -429 6861 -395
rect 7269 -429 7281 -395
rect 7689 -429 7701 -395
rect 8109 -429 8121 -395
rect 8529 -429 8541 -395
rect 549 -435 607 -429
rect 969 -435 1027 -429
rect 1389 -435 1447 -429
rect 1809 -435 1867 -429
rect 2229 -435 2287 -429
rect 2649 -435 2707 -429
rect 3069 -435 3127 -429
rect 3489 -435 3547 -429
rect 3909 -435 3967 -429
rect 4329 -435 4387 -429
rect 4749 -435 4807 -429
rect 5169 -435 5227 -429
rect 5589 -435 5647 -429
rect 6009 -435 6067 -429
rect 6429 -435 6487 -429
rect 6849 -435 6907 -429
rect 7269 -435 7327 -429
rect 7689 -435 7747 -429
rect 8109 -435 8167 -429
rect 8529 -435 8587 -429
use sky130_fd_pr__pfet_01v8_VCQUSW  sky130_fd_pr__pfet_01v8_VCQUSW_0
timestamp 1655456512
transform 1 0 4461 0 1 285
box -4520 -852 4520 319
<< end >>
