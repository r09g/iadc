magic
tech sky130A
timestamp 1654734873
<< nwell >>
rect -32 751 1777 1548
<< pwell >>
rect -17 -32 1762 726
<< mvnmos >>
rect 97 97 147 597
rect 176 97 226 597
rect 255 97 305 597
rect 334 97 384 597
rect 413 97 463 597
rect 492 97 542 597
rect 571 97 621 597
rect 650 97 700 597
rect 729 97 779 597
rect 808 97 858 597
rect 887 97 937 597
rect 966 97 1016 597
rect 1045 97 1095 597
rect 1124 97 1174 597
rect 1203 97 1253 597
rect 1282 97 1332 597
rect 1361 97 1411 597
rect 1440 97 1490 597
rect 1519 97 1569 597
rect 1598 97 1648 597
<< mvpmos >>
rect 97 899 147 1399
rect 176 899 226 1399
rect 255 899 305 1399
rect 334 899 384 1399
rect 413 899 463 1399
rect 492 899 542 1399
rect 571 899 621 1399
rect 650 899 700 1399
rect 729 899 779 1399
rect 808 899 858 1399
rect 887 899 937 1399
rect 966 899 1016 1399
rect 1045 899 1095 1399
rect 1124 899 1174 1399
rect 1203 899 1253 1399
rect 1282 899 1332 1399
rect 1361 899 1411 1399
rect 1440 899 1490 1399
rect 1519 899 1569 1399
rect 1598 899 1648 1399
<< mvndiff >>
rect 68 591 97 597
rect 68 103 74 591
rect 91 103 97 591
rect 68 97 97 103
rect 147 591 176 597
rect 147 103 153 591
rect 170 103 176 591
rect 147 97 176 103
rect 226 591 255 597
rect 226 103 232 591
rect 249 103 255 591
rect 226 97 255 103
rect 305 591 334 597
rect 305 103 311 591
rect 328 103 334 591
rect 305 97 334 103
rect 384 591 413 597
rect 384 103 390 591
rect 407 103 413 591
rect 384 97 413 103
rect 463 591 492 597
rect 463 103 469 591
rect 486 103 492 591
rect 463 97 492 103
rect 542 591 571 597
rect 542 103 548 591
rect 565 103 571 591
rect 542 97 571 103
rect 621 591 650 597
rect 621 103 627 591
rect 644 103 650 591
rect 621 97 650 103
rect 700 591 729 597
rect 700 103 706 591
rect 723 103 729 591
rect 700 97 729 103
rect 779 591 808 597
rect 779 103 785 591
rect 802 103 808 591
rect 779 97 808 103
rect 858 591 887 597
rect 858 103 864 591
rect 881 103 887 591
rect 858 97 887 103
rect 937 591 966 597
rect 937 103 943 591
rect 960 103 966 591
rect 937 97 966 103
rect 1016 591 1045 597
rect 1016 103 1022 591
rect 1039 103 1045 591
rect 1016 97 1045 103
rect 1095 591 1124 597
rect 1095 103 1101 591
rect 1118 103 1124 591
rect 1095 97 1124 103
rect 1174 591 1203 597
rect 1174 103 1180 591
rect 1197 103 1203 591
rect 1174 97 1203 103
rect 1253 591 1282 597
rect 1253 103 1259 591
rect 1276 103 1282 591
rect 1253 97 1282 103
rect 1332 591 1361 597
rect 1332 103 1338 591
rect 1355 103 1361 591
rect 1332 97 1361 103
rect 1411 591 1440 597
rect 1411 103 1417 591
rect 1434 103 1440 591
rect 1411 97 1440 103
rect 1490 591 1519 597
rect 1490 103 1496 591
rect 1513 103 1519 591
rect 1490 97 1519 103
rect 1569 591 1598 597
rect 1569 103 1575 591
rect 1592 103 1598 591
rect 1569 97 1598 103
rect 1648 591 1677 597
rect 1648 103 1654 591
rect 1671 103 1677 591
rect 1648 97 1677 103
<< mvpdiff >>
rect 68 1393 97 1399
rect 68 905 74 1393
rect 91 905 97 1393
rect 68 899 97 905
rect 147 1393 176 1399
rect 147 905 153 1393
rect 170 905 176 1393
rect 147 899 176 905
rect 226 1393 255 1399
rect 226 905 232 1393
rect 249 905 255 1393
rect 226 899 255 905
rect 305 1393 334 1399
rect 305 905 311 1393
rect 328 905 334 1393
rect 305 899 334 905
rect 384 1393 413 1399
rect 384 905 390 1393
rect 407 905 413 1393
rect 384 899 413 905
rect 463 1393 492 1399
rect 463 905 469 1393
rect 486 905 492 1393
rect 463 899 492 905
rect 542 1393 571 1399
rect 542 905 548 1393
rect 565 905 571 1393
rect 542 899 571 905
rect 621 1393 650 1399
rect 621 905 627 1393
rect 644 905 650 1393
rect 621 899 650 905
rect 700 1393 729 1399
rect 700 905 706 1393
rect 723 905 729 1393
rect 700 899 729 905
rect 779 1393 808 1399
rect 779 905 785 1393
rect 802 905 808 1393
rect 779 899 808 905
rect 858 1393 887 1399
rect 858 905 864 1393
rect 881 905 887 1393
rect 858 899 887 905
rect 937 1393 966 1399
rect 937 905 943 1393
rect 960 905 966 1393
rect 937 899 966 905
rect 1016 1393 1045 1399
rect 1016 905 1022 1393
rect 1039 905 1045 1393
rect 1016 899 1045 905
rect 1095 1393 1124 1399
rect 1095 905 1101 1393
rect 1118 905 1124 1393
rect 1095 899 1124 905
rect 1174 1393 1203 1399
rect 1174 905 1180 1393
rect 1197 905 1203 1393
rect 1174 899 1203 905
rect 1253 1393 1282 1399
rect 1253 905 1259 1393
rect 1276 905 1282 1393
rect 1253 899 1282 905
rect 1332 1393 1361 1399
rect 1332 905 1338 1393
rect 1355 905 1361 1393
rect 1332 899 1361 905
rect 1411 1393 1440 1399
rect 1411 905 1417 1393
rect 1434 905 1440 1393
rect 1411 899 1440 905
rect 1490 1393 1519 1399
rect 1490 905 1496 1393
rect 1513 905 1519 1393
rect 1490 899 1519 905
rect 1569 1393 1598 1399
rect 1569 905 1575 1393
rect 1592 905 1598 1393
rect 1569 899 1598 905
rect 1648 1393 1677 1399
rect 1648 905 1654 1393
rect 1671 905 1677 1393
rect 1648 899 1677 905
<< mvndiffc >>
rect 74 103 91 591
rect 153 103 170 591
rect 232 103 249 591
rect 311 103 328 591
rect 390 103 407 591
rect 469 103 486 591
rect 548 103 565 591
rect 627 103 644 591
rect 706 103 723 591
rect 785 103 802 591
rect 864 103 881 591
rect 943 103 960 591
rect 1022 103 1039 591
rect 1101 103 1118 591
rect 1180 103 1197 591
rect 1259 103 1276 591
rect 1338 103 1355 591
rect 1417 103 1434 591
rect 1496 103 1513 591
rect 1575 103 1592 591
rect 1654 103 1671 591
<< mvpdiffc >>
rect 74 905 91 1393
rect 153 905 170 1393
rect 232 905 249 1393
rect 311 905 328 1393
rect 390 905 407 1393
rect 469 905 486 1393
rect 548 905 565 1393
rect 627 905 644 1393
rect 706 905 723 1393
rect 785 905 802 1393
rect 864 905 881 1393
rect 943 905 960 1393
rect 1022 905 1039 1393
rect 1101 905 1118 1393
rect 1180 905 1197 1393
rect 1259 905 1276 1393
rect 1338 905 1355 1393
rect 1417 905 1434 1393
rect 1496 905 1513 1393
rect 1575 905 1592 1393
rect 1654 905 1671 1393
<< mvpsubdiff >>
rect 1 702 1744 708
rect 1 685 55 702
rect 1690 685 1744 702
rect 1 679 1744 685
rect 1 654 30 679
rect 1 40 7 654
rect 24 40 30 654
rect 1715 654 1744 679
rect 1 15 30 40
rect 1715 40 1721 654
rect 1738 40 1744 654
rect 1715 15 1744 40
rect 1 9 1744 15
rect 1 -8 55 9
rect 1690 -8 1744 9
rect 1 -14 1744 -8
<< mvnsubdiff >>
rect 1 1509 1744 1515
rect 1 1492 55 1509
rect 1690 1492 1744 1509
rect 1 1486 1744 1492
rect 1 1461 30 1486
rect 1 838 7 1461
rect 24 838 30 1461
rect 1715 1461 1744 1486
rect 1 813 30 838
rect 1715 838 1721 1461
rect 1738 838 1744 1461
rect 1715 813 1744 838
rect 1 807 1744 813
rect 1 790 55 807
rect 1690 790 1744 807
rect 1 784 1744 790
<< mvpsubdiffcont >>
rect 55 685 1690 702
rect 7 40 24 654
rect 1721 40 1738 654
rect 55 -8 1690 9
<< mvnsubdiffcont >>
rect 55 1492 1690 1509
rect 7 838 24 1461
rect 1721 838 1738 1461
rect 55 790 1690 807
<< poly >>
rect 97 1440 147 1448
rect 97 1423 105 1440
rect 139 1423 147 1440
rect 97 1399 147 1423
rect 176 1440 226 1448
rect 176 1423 184 1440
rect 218 1423 226 1440
rect 176 1399 226 1423
rect 255 1440 305 1448
rect 255 1423 263 1440
rect 297 1423 305 1440
rect 255 1399 305 1423
rect 334 1440 384 1448
rect 334 1423 342 1440
rect 376 1423 384 1440
rect 334 1399 384 1423
rect 413 1440 463 1448
rect 413 1423 421 1440
rect 455 1423 463 1440
rect 413 1399 463 1423
rect 492 1440 542 1448
rect 492 1423 500 1440
rect 534 1423 542 1440
rect 492 1399 542 1423
rect 571 1440 621 1448
rect 571 1423 579 1440
rect 613 1423 621 1440
rect 571 1399 621 1423
rect 650 1440 700 1448
rect 650 1423 658 1440
rect 692 1423 700 1440
rect 650 1399 700 1423
rect 729 1440 779 1448
rect 729 1423 737 1440
rect 771 1423 779 1440
rect 729 1399 779 1423
rect 808 1440 858 1448
rect 808 1423 816 1440
rect 850 1423 858 1440
rect 808 1399 858 1423
rect 887 1440 937 1448
rect 887 1423 895 1440
rect 929 1423 937 1440
rect 887 1399 937 1423
rect 966 1440 1016 1448
rect 966 1423 974 1440
rect 1008 1423 1016 1440
rect 966 1399 1016 1423
rect 1045 1440 1095 1448
rect 1045 1423 1053 1440
rect 1087 1423 1095 1440
rect 1045 1399 1095 1423
rect 1124 1440 1174 1448
rect 1124 1423 1132 1440
rect 1166 1423 1174 1440
rect 1124 1399 1174 1423
rect 1203 1440 1253 1448
rect 1203 1423 1211 1440
rect 1245 1423 1253 1440
rect 1203 1399 1253 1423
rect 1282 1440 1332 1448
rect 1282 1423 1290 1440
rect 1324 1423 1332 1440
rect 1282 1399 1332 1423
rect 1361 1440 1411 1448
rect 1361 1423 1369 1440
rect 1403 1423 1411 1440
rect 1361 1399 1411 1423
rect 1440 1440 1490 1448
rect 1440 1423 1448 1440
rect 1482 1423 1490 1440
rect 1440 1399 1490 1423
rect 1519 1440 1569 1448
rect 1519 1423 1527 1440
rect 1561 1423 1569 1440
rect 1519 1399 1569 1423
rect 1598 1440 1648 1448
rect 1598 1423 1606 1440
rect 1640 1423 1648 1440
rect 1598 1399 1648 1423
rect 97 876 147 899
rect 97 859 105 876
rect 139 859 147 876
rect 97 851 147 859
rect 176 876 226 899
rect 176 859 184 876
rect 218 859 226 876
rect 176 851 226 859
rect 255 876 305 899
rect 255 859 263 876
rect 297 859 305 876
rect 255 851 305 859
rect 334 876 384 899
rect 334 859 342 876
rect 376 859 384 876
rect 334 851 384 859
rect 413 876 463 899
rect 413 859 421 876
rect 455 859 463 876
rect 413 851 463 859
rect 492 876 542 899
rect 492 859 500 876
rect 534 859 542 876
rect 492 851 542 859
rect 571 876 621 899
rect 571 859 579 876
rect 613 859 621 876
rect 571 851 621 859
rect 650 876 700 899
rect 650 859 658 876
rect 692 859 700 876
rect 650 851 700 859
rect 729 876 779 899
rect 729 859 737 876
rect 771 859 779 876
rect 729 851 779 859
rect 808 876 858 899
rect 808 859 816 876
rect 850 859 858 876
rect 808 851 858 859
rect 887 876 937 899
rect 887 859 895 876
rect 929 859 937 876
rect 887 851 937 859
rect 966 876 1016 899
rect 966 859 974 876
rect 1008 859 1016 876
rect 966 851 1016 859
rect 1045 876 1095 899
rect 1045 859 1053 876
rect 1087 859 1095 876
rect 1045 851 1095 859
rect 1124 876 1174 899
rect 1124 859 1132 876
rect 1166 859 1174 876
rect 1124 851 1174 859
rect 1203 876 1253 899
rect 1203 859 1211 876
rect 1245 859 1253 876
rect 1203 851 1253 859
rect 1282 876 1332 899
rect 1282 859 1290 876
rect 1324 859 1332 876
rect 1282 851 1332 859
rect 1361 876 1411 899
rect 1361 859 1369 876
rect 1403 859 1411 876
rect 1361 851 1411 859
rect 1440 876 1490 899
rect 1440 859 1448 876
rect 1482 859 1490 876
rect 1440 851 1490 859
rect 1519 876 1569 899
rect 1519 859 1527 876
rect 1561 859 1569 876
rect 1519 851 1569 859
rect 1598 876 1648 899
rect 1598 859 1606 876
rect 1640 859 1648 876
rect 1598 851 1648 859
rect 97 633 147 641
rect 97 616 105 633
rect 139 616 147 633
rect 97 597 147 616
rect 176 633 226 641
rect 176 616 184 633
rect 218 616 226 633
rect 176 597 226 616
rect 255 633 305 641
rect 255 616 263 633
rect 297 616 305 633
rect 255 597 305 616
rect 334 633 384 641
rect 334 616 342 633
rect 376 616 384 633
rect 334 597 384 616
rect 413 633 463 641
rect 413 616 421 633
rect 455 616 463 633
rect 413 597 463 616
rect 492 633 542 641
rect 492 616 500 633
rect 534 616 542 633
rect 492 597 542 616
rect 571 633 621 641
rect 571 616 579 633
rect 613 616 621 633
rect 571 597 621 616
rect 650 633 700 641
rect 650 616 658 633
rect 692 616 700 633
rect 650 597 700 616
rect 729 633 779 641
rect 729 616 737 633
rect 771 616 779 633
rect 729 597 779 616
rect 808 633 858 641
rect 808 616 816 633
rect 850 616 858 633
rect 808 597 858 616
rect 887 633 937 641
rect 887 616 895 633
rect 929 616 937 633
rect 887 597 937 616
rect 966 633 1016 641
rect 966 616 974 633
rect 1008 616 1016 633
rect 966 597 1016 616
rect 1045 633 1095 641
rect 1045 616 1053 633
rect 1087 616 1095 633
rect 1045 597 1095 616
rect 1124 633 1174 641
rect 1124 616 1132 633
rect 1166 616 1174 633
rect 1124 597 1174 616
rect 1203 633 1253 641
rect 1203 616 1211 633
rect 1245 616 1253 633
rect 1203 597 1253 616
rect 1282 633 1332 641
rect 1282 616 1290 633
rect 1324 616 1332 633
rect 1282 597 1332 616
rect 1361 633 1411 641
rect 1361 616 1369 633
rect 1403 616 1411 633
rect 1361 597 1411 616
rect 1440 633 1490 641
rect 1440 616 1448 633
rect 1482 616 1490 633
rect 1440 597 1490 616
rect 1519 633 1569 641
rect 1519 616 1527 633
rect 1561 616 1569 633
rect 1519 597 1569 616
rect 1598 633 1648 641
rect 1598 616 1606 633
rect 1640 616 1648 633
rect 1598 597 1648 616
rect 97 78 147 97
rect 97 61 105 78
rect 139 61 147 78
rect 97 53 147 61
rect 176 78 226 97
rect 176 61 184 78
rect 218 61 226 78
rect 176 53 226 61
rect 255 78 305 97
rect 255 61 263 78
rect 297 61 305 78
rect 255 53 305 61
rect 334 78 384 97
rect 334 61 342 78
rect 376 61 384 78
rect 334 53 384 61
rect 413 78 463 97
rect 413 61 421 78
rect 455 61 463 78
rect 413 53 463 61
rect 492 78 542 97
rect 492 61 500 78
rect 534 61 542 78
rect 492 53 542 61
rect 571 78 621 97
rect 571 61 579 78
rect 613 61 621 78
rect 571 53 621 61
rect 650 78 700 97
rect 650 61 658 78
rect 692 61 700 78
rect 650 53 700 61
rect 729 78 779 97
rect 729 61 737 78
rect 771 61 779 78
rect 729 53 779 61
rect 808 78 858 97
rect 808 61 816 78
rect 850 61 858 78
rect 808 53 858 61
rect 887 78 937 97
rect 887 61 895 78
rect 929 61 937 78
rect 887 53 937 61
rect 966 78 1016 97
rect 966 61 974 78
rect 1008 61 1016 78
rect 966 53 1016 61
rect 1045 78 1095 97
rect 1045 61 1053 78
rect 1087 61 1095 78
rect 1045 53 1095 61
rect 1124 78 1174 97
rect 1124 61 1132 78
rect 1166 61 1174 78
rect 1124 53 1174 61
rect 1203 78 1253 97
rect 1203 61 1211 78
rect 1245 61 1253 78
rect 1203 53 1253 61
rect 1282 78 1332 97
rect 1282 61 1290 78
rect 1324 61 1332 78
rect 1282 53 1332 61
rect 1361 78 1411 97
rect 1361 61 1369 78
rect 1403 61 1411 78
rect 1361 53 1411 61
rect 1440 78 1490 97
rect 1440 61 1448 78
rect 1482 61 1490 78
rect 1440 53 1490 61
rect 1519 78 1569 97
rect 1519 61 1527 78
rect 1561 61 1569 78
rect 1519 53 1569 61
rect 1598 78 1648 97
rect 1598 61 1606 78
rect 1640 61 1648 78
rect 1598 53 1648 61
<< polycont >>
rect 105 1423 139 1440
rect 184 1423 218 1440
rect 263 1423 297 1440
rect 342 1423 376 1440
rect 421 1423 455 1440
rect 500 1423 534 1440
rect 579 1423 613 1440
rect 658 1423 692 1440
rect 737 1423 771 1440
rect 816 1423 850 1440
rect 895 1423 929 1440
rect 974 1423 1008 1440
rect 1053 1423 1087 1440
rect 1132 1423 1166 1440
rect 1211 1423 1245 1440
rect 1290 1423 1324 1440
rect 1369 1423 1403 1440
rect 1448 1423 1482 1440
rect 1527 1423 1561 1440
rect 1606 1423 1640 1440
rect 105 859 139 876
rect 184 859 218 876
rect 263 859 297 876
rect 342 859 376 876
rect 421 859 455 876
rect 500 859 534 876
rect 579 859 613 876
rect 658 859 692 876
rect 737 859 771 876
rect 816 859 850 876
rect 895 859 929 876
rect 974 859 1008 876
rect 1053 859 1087 876
rect 1132 859 1166 876
rect 1211 859 1245 876
rect 1290 859 1324 876
rect 1369 859 1403 876
rect 1448 859 1482 876
rect 1527 859 1561 876
rect 1606 859 1640 876
rect 105 616 139 633
rect 184 616 218 633
rect 263 616 297 633
rect 342 616 376 633
rect 421 616 455 633
rect 500 616 534 633
rect 579 616 613 633
rect 658 616 692 633
rect 737 616 771 633
rect 816 616 850 633
rect 895 616 929 633
rect 974 616 1008 633
rect 1053 616 1087 633
rect 1132 616 1166 633
rect 1211 616 1245 633
rect 1290 616 1324 633
rect 1369 616 1403 633
rect 1448 616 1482 633
rect 1527 616 1561 633
rect 1606 616 1640 633
rect 105 61 139 78
rect 184 61 218 78
rect 263 61 297 78
rect 342 61 376 78
rect 421 61 455 78
rect 500 61 534 78
rect 579 61 613 78
rect 658 61 692 78
rect 737 61 771 78
rect 816 61 850 78
rect 895 61 929 78
rect 974 61 1008 78
rect 1053 61 1087 78
rect 1132 61 1166 78
rect 1211 61 1245 78
rect 1290 61 1324 78
rect 1369 61 1403 78
rect 1448 61 1482 78
rect 1527 61 1561 78
rect 1606 61 1640 78
<< locali >>
rect 7 1492 55 1509
rect 1690 1492 1738 1509
rect 7 1461 24 1492
rect 1721 1461 1738 1492
rect 97 1423 105 1440
rect 139 1423 147 1440
rect 176 1423 184 1440
rect 218 1423 226 1440
rect 255 1423 263 1440
rect 297 1423 305 1440
rect 334 1423 342 1440
rect 376 1423 384 1440
rect 413 1423 421 1440
rect 455 1423 463 1440
rect 492 1423 500 1440
rect 534 1423 542 1440
rect 571 1423 579 1440
rect 613 1423 621 1440
rect 650 1423 658 1440
rect 692 1423 700 1440
rect 729 1423 737 1440
rect 771 1423 779 1440
rect 808 1423 816 1440
rect 850 1423 858 1440
rect 887 1423 895 1440
rect 929 1423 937 1440
rect 966 1423 974 1440
rect 1008 1423 1016 1440
rect 1045 1423 1053 1440
rect 1087 1423 1095 1440
rect 1124 1423 1132 1440
rect 1166 1423 1174 1440
rect 1203 1423 1211 1440
rect 1245 1423 1253 1440
rect 1282 1423 1290 1440
rect 1324 1423 1332 1440
rect 1361 1423 1369 1440
rect 1403 1423 1411 1440
rect 1440 1423 1448 1440
rect 1482 1423 1490 1440
rect 1519 1423 1527 1440
rect 1561 1423 1569 1440
rect 1598 1423 1606 1440
rect 1640 1423 1648 1440
rect 74 1393 91 1401
rect 74 897 91 905
rect 153 1393 170 1401
rect 153 897 170 905
rect 232 1393 249 1401
rect 232 897 249 905
rect 311 1393 328 1401
rect 311 897 328 905
rect 390 1393 407 1401
rect 390 897 407 905
rect 469 1393 486 1401
rect 469 897 486 905
rect 548 1393 565 1401
rect 548 897 565 905
rect 627 1393 644 1401
rect 627 897 644 905
rect 706 1393 723 1401
rect 706 897 723 905
rect 785 1393 802 1401
rect 785 897 802 905
rect 864 1393 881 1401
rect 864 897 881 905
rect 943 1393 960 1401
rect 943 897 960 905
rect 1022 1393 1039 1401
rect 1022 897 1039 905
rect 1101 1393 1118 1401
rect 1101 897 1118 905
rect 1180 1393 1197 1401
rect 1180 897 1197 905
rect 1259 1393 1276 1401
rect 1259 897 1276 905
rect 1338 1393 1355 1401
rect 1338 897 1355 905
rect 1417 1393 1434 1401
rect 1417 897 1434 905
rect 1496 1393 1513 1401
rect 1496 897 1513 905
rect 1575 1393 1592 1401
rect 1575 897 1592 905
rect 1654 1393 1671 1401
rect 1654 897 1671 905
rect 97 859 105 876
rect 139 859 147 876
rect 176 859 184 876
rect 218 859 226 876
rect 255 859 263 876
rect 297 859 305 876
rect 334 859 342 876
rect 376 859 384 876
rect 413 859 421 876
rect 455 859 463 876
rect 492 859 500 876
rect 534 859 542 876
rect 571 859 579 876
rect 613 859 621 876
rect 650 859 658 876
rect 692 859 700 876
rect 729 859 737 876
rect 771 859 779 876
rect 808 859 816 876
rect 850 859 858 876
rect 887 859 895 876
rect 929 859 937 876
rect 966 859 974 876
rect 1008 859 1016 876
rect 1045 859 1053 876
rect 1087 859 1095 876
rect 1124 859 1132 876
rect 1166 859 1174 876
rect 1203 859 1211 876
rect 1245 859 1253 876
rect 1282 859 1290 876
rect 1324 859 1332 876
rect 1361 859 1369 876
rect 1403 859 1411 876
rect 1440 859 1448 876
rect 1482 859 1490 876
rect 1519 859 1527 876
rect 1561 859 1569 876
rect 1598 859 1606 876
rect 1640 859 1648 876
rect 7 807 24 838
rect 1721 807 1738 838
rect 7 790 55 807
rect 1690 790 1738 807
rect 7 685 55 702
rect 1690 685 1738 702
rect 7 654 24 685
rect 1721 654 1738 685
rect 97 616 105 633
rect 139 616 147 633
rect 176 616 184 633
rect 218 616 226 633
rect 255 616 263 633
rect 297 616 305 633
rect 334 616 342 633
rect 376 616 384 633
rect 413 616 421 633
rect 455 616 463 633
rect 492 616 500 633
rect 534 616 542 633
rect 571 616 579 633
rect 613 616 621 633
rect 650 616 658 633
rect 692 616 700 633
rect 729 616 737 633
rect 771 616 779 633
rect 808 616 816 633
rect 850 616 858 633
rect 887 616 895 633
rect 929 616 937 633
rect 966 616 974 633
rect 1008 616 1016 633
rect 1045 616 1053 633
rect 1087 616 1095 633
rect 1124 616 1132 633
rect 1166 616 1174 633
rect 1203 616 1211 633
rect 1245 616 1253 633
rect 1282 616 1290 633
rect 1324 616 1332 633
rect 1361 616 1369 633
rect 1403 616 1411 633
rect 1440 616 1448 633
rect 1482 616 1490 633
rect 1519 616 1527 633
rect 1561 616 1569 633
rect 1598 616 1606 633
rect 1640 616 1648 633
rect 74 591 91 599
rect 74 95 91 103
rect 153 591 170 599
rect 153 95 170 103
rect 232 591 249 599
rect 232 95 249 103
rect 311 591 328 599
rect 311 95 328 103
rect 390 591 407 599
rect 390 95 407 103
rect 469 591 486 599
rect 469 95 486 103
rect 548 591 565 599
rect 548 95 565 103
rect 627 591 644 599
rect 627 95 644 103
rect 706 591 723 599
rect 706 95 723 103
rect 785 591 802 599
rect 785 95 802 103
rect 864 591 881 599
rect 864 95 881 103
rect 943 591 960 599
rect 943 95 960 103
rect 1022 591 1039 599
rect 1022 95 1039 103
rect 1101 591 1118 599
rect 1101 95 1118 103
rect 1180 591 1197 599
rect 1180 95 1197 103
rect 1259 591 1276 599
rect 1259 95 1276 103
rect 1338 591 1355 599
rect 1338 95 1355 103
rect 1417 591 1434 599
rect 1417 95 1434 103
rect 1496 591 1513 599
rect 1496 95 1513 103
rect 1575 591 1592 599
rect 1575 95 1592 103
rect 1654 591 1671 599
rect 1654 95 1671 103
rect 97 61 105 78
rect 139 61 147 78
rect 176 61 184 78
rect 218 61 226 78
rect 255 61 263 78
rect 297 61 305 78
rect 334 61 342 78
rect 376 61 384 78
rect 413 61 421 78
rect 455 61 463 78
rect 492 61 500 78
rect 534 61 542 78
rect 571 61 579 78
rect 613 61 621 78
rect 650 61 658 78
rect 692 61 700 78
rect 729 61 737 78
rect 771 61 779 78
rect 808 61 816 78
rect 850 61 858 78
rect 887 61 895 78
rect 929 61 937 78
rect 966 61 974 78
rect 1008 61 1016 78
rect 1045 61 1053 78
rect 1087 61 1095 78
rect 1124 61 1132 78
rect 1166 61 1174 78
rect 1203 61 1211 78
rect 1245 61 1253 78
rect 1282 61 1290 78
rect 1324 61 1332 78
rect 1361 61 1369 78
rect 1403 61 1411 78
rect 1440 61 1448 78
rect 1482 61 1490 78
rect 1519 61 1527 78
rect 1561 61 1569 78
rect 1598 61 1606 78
rect 1640 61 1648 78
rect 7 9 24 40
rect 1721 9 1738 40
rect 7 -8 55 9
rect 1690 -8 1738 9
<< viali >>
rect 55 1492 1690 1509
rect 7 838 24 1461
rect 113 1423 130 1440
rect 192 1423 209 1440
rect 271 1423 288 1440
rect 350 1423 367 1440
rect 429 1423 446 1440
rect 508 1423 525 1440
rect 587 1423 604 1440
rect 666 1423 683 1440
rect 745 1423 762 1440
rect 824 1423 841 1440
rect 904 1423 921 1440
rect 983 1423 1000 1440
rect 1062 1423 1079 1440
rect 1141 1423 1158 1440
rect 1220 1423 1237 1440
rect 1299 1423 1316 1440
rect 1378 1423 1395 1440
rect 1457 1423 1474 1440
rect 1536 1423 1553 1440
rect 1615 1423 1632 1440
rect 74 905 91 1393
rect 153 905 170 1393
rect 232 905 249 1393
rect 311 905 328 1393
rect 390 905 407 1393
rect 469 905 486 1393
rect 548 905 565 1393
rect 627 905 644 1393
rect 706 905 723 1393
rect 785 905 802 1393
rect 864 905 881 1393
rect 943 905 960 1393
rect 1022 905 1039 1393
rect 1101 905 1118 1393
rect 1180 905 1197 1393
rect 1259 905 1276 1393
rect 1338 905 1355 1393
rect 1417 905 1434 1393
rect 1496 905 1513 1393
rect 1575 905 1592 1393
rect 1654 905 1671 1393
rect 113 859 130 876
rect 192 859 209 876
rect 271 859 288 876
rect 350 859 367 876
rect 429 859 446 876
rect 508 859 525 876
rect 587 859 604 876
rect 666 859 683 876
rect 745 859 762 876
rect 824 859 841 876
rect 904 859 921 876
rect 983 859 1000 876
rect 1062 859 1079 876
rect 1141 859 1158 876
rect 1220 859 1237 876
rect 1299 859 1316 876
rect 1378 859 1395 876
rect 1457 859 1474 876
rect 1536 859 1553 876
rect 1615 859 1632 876
rect 1721 838 1738 1461
rect 7 40 24 654
rect 113 616 130 633
rect 192 616 209 633
rect 271 616 288 633
rect 350 616 367 633
rect 429 616 446 633
rect 508 616 525 633
rect 587 616 604 633
rect 666 616 683 633
rect 745 616 762 633
rect 824 616 841 633
rect 904 616 921 633
rect 983 616 1000 633
rect 1062 616 1079 633
rect 1141 616 1158 633
rect 1220 616 1237 633
rect 1299 616 1316 633
rect 1378 616 1395 633
rect 1457 616 1474 633
rect 1536 616 1553 633
rect 1615 616 1632 633
rect 74 103 91 591
rect 153 103 170 591
rect 232 103 249 591
rect 311 103 328 591
rect 390 103 407 591
rect 469 103 486 591
rect 548 103 565 591
rect 627 103 644 591
rect 706 103 723 591
rect 785 103 802 591
rect 864 103 881 591
rect 943 103 960 591
rect 1022 103 1039 591
rect 1101 103 1118 591
rect 1180 103 1197 591
rect 1259 103 1276 591
rect 1338 103 1355 591
rect 1417 103 1434 591
rect 1496 103 1513 591
rect 1575 103 1592 591
rect 1654 103 1671 591
rect 113 61 130 78
rect 192 61 209 78
rect 271 61 288 78
rect 350 61 367 78
rect 429 61 446 78
rect 508 61 525 78
rect 587 61 604 78
rect 666 61 683 78
rect 745 61 762 78
rect 824 61 841 78
rect 904 61 921 78
rect 983 61 1000 78
rect 1062 61 1079 78
rect 1141 61 1158 78
rect 1220 61 1237 78
rect 1299 61 1316 78
rect 1378 61 1395 78
rect 1457 61 1474 78
rect 1536 61 1553 78
rect 1615 61 1632 78
rect 1721 40 1738 654
rect 55 -8 1690 9
<< metal1 >>
rect 4 1509 1741 1512
rect 4 1492 55 1509
rect 1690 1492 1741 1509
rect 4 1461 1741 1492
rect 4 838 7 1461
rect 24 1440 1721 1461
rect 24 1423 113 1440
rect 130 1423 192 1440
rect 209 1423 271 1440
rect 288 1423 350 1440
rect 367 1423 429 1440
rect 446 1423 508 1440
rect 525 1423 587 1440
rect 604 1423 666 1440
rect 683 1423 745 1440
rect 762 1423 824 1440
rect 841 1423 904 1440
rect 921 1423 983 1440
rect 1000 1423 1062 1440
rect 1079 1423 1141 1440
rect 1158 1423 1220 1440
rect 1237 1423 1299 1440
rect 1316 1423 1378 1440
rect 1395 1423 1457 1440
rect 1474 1423 1536 1440
rect 1553 1423 1615 1440
rect 1632 1423 1721 1440
rect 24 1420 1721 1423
rect 24 879 30 1420
rect 71 1393 94 1420
rect 150 1393 173 1399
rect 229 1393 252 1420
rect 308 1393 331 1399
rect 387 1393 410 1420
rect 466 1393 489 1399
rect 545 1393 568 1420
rect 624 1393 647 1399
rect 703 1393 726 1420
rect 782 1393 805 1399
rect 861 1393 884 1420
rect 940 1393 963 1399
rect 1019 1393 1042 1420
rect 1098 1393 1121 1399
rect 1177 1393 1200 1420
rect 1256 1393 1279 1399
rect 1335 1393 1358 1420
rect 1414 1393 1437 1399
rect 1493 1393 1516 1420
rect 1572 1393 1595 1399
rect 1651 1393 1674 1420
rect 71 905 74 1393
rect 91 905 94 1393
rect 143 905 148 1393
rect 174 905 179 1393
rect 229 905 232 1393
rect 249 905 252 1393
rect 301 905 306 1393
rect 332 905 337 1393
rect 387 905 390 1393
rect 407 905 410 1393
rect 459 905 464 1393
rect 490 905 495 1393
rect 545 905 548 1393
rect 565 905 568 1393
rect 617 905 622 1393
rect 648 905 653 1393
rect 703 905 706 1393
rect 723 905 726 1393
rect 775 905 780 1393
rect 806 905 811 1393
rect 861 905 864 1393
rect 881 905 884 1393
rect 933 905 938 1393
rect 964 905 969 1393
rect 1019 905 1022 1393
rect 1039 905 1042 1393
rect 1091 905 1096 1393
rect 1122 905 1127 1393
rect 1177 905 1180 1393
rect 1197 905 1200 1393
rect 1249 905 1254 1393
rect 1280 905 1285 1393
rect 1335 905 1338 1393
rect 1355 905 1358 1393
rect 1407 905 1412 1393
rect 1438 905 1443 1393
rect 1493 905 1496 1393
rect 1513 905 1516 1393
rect 1565 905 1570 1393
rect 1596 905 1601 1393
rect 1651 905 1654 1393
rect 1671 905 1674 1393
rect 71 879 94 905
rect 150 899 173 905
rect 229 899 252 905
rect 308 899 331 905
rect 387 899 410 905
rect 466 899 489 905
rect 545 899 568 905
rect 624 899 647 905
rect 703 899 726 905
rect 782 899 805 905
rect 861 899 884 905
rect 940 899 963 905
rect 1019 899 1042 905
rect 1098 899 1121 905
rect 1177 899 1200 905
rect 1256 899 1279 905
rect 1335 899 1358 905
rect 1414 899 1437 905
rect 1493 899 1516 905
rect 1572 899 1595 905
rect 1651 879 1674 905
rect 1715 879 1721 1420
rect 24 876 1721 879
rect 24 859 113 876
rect 130 859 192 876
rect 209 859 271 876
rect 288 859 350 876
rect 367 859 429 876
rect 446 859 508 876
rect 525 859 587 876
rect 604 859 666 876
rect 683 859 745 876
rect 762 859 824 876
rect 841 859 904 876
rect 921 859 983 876
rect 1000 859 1062 876
rect 1079 859 1141 876
rect 1158 859 1220 876
rect 1237 859 1299 876
rect 1316 859 1378 876
rect 1395 859 1457 876
rect 1474 859 1536 876
rect 1553 859 1615 876
rect 1632 859 1721 876
rect 24 856 1721 859
rect 24 838 27 856
rect 4 832 27 838
rect 1718 838 1721 856
rect 1738 838 1741 1461
rect 1718 832 1741 838
rect -32 772 1777 778
rect -32 720 148 772
rect 174 720 306 772
rect 332 720 464 772
rect 490 720 622 772
rect 648 720 780 772
rect 806 720 938 772
rect 964 720 1096 772
rect 1122 720 1254 772
rect 1280 720 1412 772
rect 1438 720 1570 772
rect 1596 720 1777 772
rect -32 714 1777 720
rect 4 654 27 660
rect 4 40 7 654
rect 24 636 27 654
rect 1718 654 1741 660
rect 1718 636 1721 654
rect 24 633 1721 636
rect 24 616 113 633
rect 130 616 192 633
rect 209 616 271 633
rect 288 616 350 633
rect 367 616 429 633
rect 446 616 508 633
rect 525 616 587 633
rect 604 616 666 633
rect 683 616 745 633
rect 762 616 824 633
rect 841 616 904 633
rect 921 616 983 633
rect 1000 616 1062 633
rect 1079 616 1141 633
rect 1158 616 1220 633
rect 1237 616 1299 633
rect 1316 616 1378 633
rect 1395 616 1457 633
rect 1474 616 1536 633
rect 1553 616 1615 633
rect 1632 616 1721 633
rect 24 613 1721 616
rect 24 81 27 613
rect 71 591 94 597
rect 150 591 173 597
rect 229 591 252 597
rect 308 591 331 597
rect 387 591 410 597
rect 466 591 489 597
rect 545 591 568 597
rect 624 591 647 597
rect 703 591 726 597
rect 782 591 805 597
rect 861 591 884 597
rect 940 591 963 597
rect 1019 591 1042 597
rect 1098 591 1121 597
rect 1177 591 1200 597
rect 1256 591 1279 597
rect 1335 591 1358 597
rect 1414 591 1437 597
rect 1493 591 1516 597
rect 1572 591 1595 597
rect 1651 591 1674 613
rect 71 103 74 591
rect 91 103 94 591
rect 143 103 148 591
rect 174 103 179 591
rect 229 103 232 591
rect 249 103 252 591
rect 301 103 306 591
rect 332 103 337 591
rect 387 103 390 591
rect 407 103 410 591
rect 459 103 464 591
rect 490 103 495 591
rect 545 103 548 591
rect 565 103 568 591
rect 617 103 622 591
rect 648 103 653 591
rect 703 103 706 591
rect 723 103 726 591
rect 775 103 780 591
rect 806 103 811 591
rect 861 103 864 591
rect 881 103 884 591
rect 933 103 938 591
rect 964 103 969 591
rect 1019 103 1022 591
rect 1039 103 1042 591
rect 1091 103 1096 591
rect 1122 103 1127 591
rect 1177 103 1180 591
rect 1197 103 1200 591
rect 1249 103 1254 591
rect 1280 103 1285 591
rect 1335 103 1338 591
rect 1355 103 1358 591
rect 1407 103 1412 591
rect 1438 103 1443 591
rect 1493 103 1496 591
rect 1513 103 1516 591
rect 1565 103 1570 591
rect 1596 103 1601 591
rect 1651 103 1654 591
rect 1671 103 1674 591
rect 71 81 94 103
rect 150 97 173 103
rect 229 81 252 103
rect 308 97 331 103
rect 387 81 410 103
rect 466 97 489 103
rect 545 81 568 103
rect 624 97 647 103
rect 703 81 726 103
rect 782 97 805 103
rect 861 81 884 103
rect 940 97 963 103
rect 1019 81 1042 103
rect 1098 97 1121 103
rect 1177 81 1200 103
rect 1256 97 1279 103
rect 1335 81 1358 103
rect 1414 97 1437 103
rect 1493 81 1516 103
rect 1572 97 1595 103
rect 1651 81 1674 103
rect 1718 81 1721 613
rect 24 78 1721 81
rect 24 61 113 78
rect 130 61 192 78
rect 209 61 271 78
rect 288 61 350 78
rect 367 61 429 78
rect 446 61 508 78
rect 525 61 587 78
rect 604 61 666 78
rect 683 61 745 78
rect 762 61 824 78
rect 841 61 904 78
rect 921 61 983 78
rect 1000 61 1062 78
rect 1079 61 1141 78
rect 1158 61 1220 78
rect 1237 61 1299 78
rect 1316 61 1378 78
rect 1395 61 1457 78
rect 1474 61 1536 78
rect 1553 61 1615 78
rect 1632 61 1721 78
rect 24 40 1721 61
rect 1738 40 1741 654
rect 4 9 1741 40
rect 4 -8 55 9
rect 1690 -8 1741 9
rect 4 -11 1741 -8
<< via1 >>
rect 148 905 153 1393
rect 153 905 170 1393
rect 170 905 174 1393
rect 306 905 311 1393
rect 311 905 328 1393
rect 328 905 332 1393
rect 464 905 469 1393
rect 469 905 486 1393
rect 486 905 490 1393
rect 622 905 627 1393
rect 627 905 644 1393
rect 644 905 648 1393
rect 780 905 785 1393
rect 785 905 802 1393
rect 802 905 806 1393
rect 938 905 943 1393
rect 943 905 960 1393
rect 960 905 964 1393
rect 1096 905 1101 1393
rect 1101 905 1118 1393
rect 1118 905 1122 1393
rect 1254 905 1259 1393
rect 1259 905 1276 1393
rect 1276 905 1280 1393
rect 1412 905 1417 1393
rect 1417 905 1434 1393
rect 1434 905 1438 1393
rect 1570 905 1575 1393
rect 1575 905 1592 1393
rect 1592 905 1596 1393
rect 148 720 174 772
rect 306 720 332 772
rect 464 720 490 772
rect 622 720 648 772
rect 780 720 806 772
rect 938 720 964 772
rect 1096 720 1122 772
rect 1254 720 1280 772
rect 1412 720 1438 772
rect 1570 720 1596 772
rect 148 103 153 591
rect 153 103 170 591
rect 170 103 174 591
rect 306 103 311 591
rect 311 103 328 591
rect 328 103 332 591
rect 464 103 469 591
rect 469 103 486 591
rect 486 103 490 591
rect 622 103 627 591
rect 627 103 644 591
rect 644 103 648 591
rect 780 103 785 591
rect 785 103 802 591
rect 802 103 806 591
rect 938 103 943 591
rect 943 103 960 591
rect 960 103 964 591
rect 1096 103 1101 591
rect 1101 103 1118 591
rect 1118 103 1122 591
rect 1254 103 1259 591
rect 1259 103 1276 591
rect 1276 103 1280 591
rect 1412 103 1417 591
rect 1417 103 1434 591
rect 1434 103 1438 591
rect 1570 103 1575 591
rect 1575 103 1592 591
rect 1592 103 1596 591
<< metal2 >>
rect 148 1393 174 1398
rect 148 772 174 905
rect 148 591 174 720
rect 148 98 174 103
rect 306 1393 332 1398
rect 306 772 332 905
rect 306 591 332 720
rect 306 98 332 103
rect 464 1393 490 1398
rect 464 772 490 905
rect 464 591 490 720
rect 464 98 490 103
rect 622 1393 648 1398
rect 622 772 648 905
rect 622 591 648 720
rect 622 98 648 103
rect 780 1393 806 1398
rect 780 772 806 905
rect 780 591 806 720
rect 780 98 806 103
rect 938 1393 964 1398
rect 938 772 964 905
rect 938 591 964 720
rect 938 98 964 103
rect 1096 1393 1122 1398
rect 1096 772 1122 905
rect 1096 591 1122 720
rect 1096 98 1122 103
rect 1254 1393 1280 1398
rect 1254 772 1280 905
rect 1254 591 1280 720
rect 1254 98 1280 103
rect 1412 1393 1438 1398
rect 1412 772 1438 905
rect 1412 591 1438 720
rect 1412 98 1438 103
rect 1570 1393 1596 1398
rect 1570 772 1596 905
rect 1570 591 1596 720
rect 1570 98 1596 103
<< labels >>
flabel metal1 -26 744 -26 744 1 FreeSans 200 0 0 0 esd
port 1 n
flabel metal1 15 1464 15 1464 1 FreeSans 200 0 0 0 VDD
port 2 n power bidirectional
flabel metal1 15 36 15 36 1 FreeSans 200 0 0 0 VSS
port 3 n power bidirectional
<< end >>
