magic
tech sky130A
magscale 1 2
timestamp 1652749834
<< metal1 >>
rect -133 934 0 986
rect -300 438 -238 490
rect -186 438 -176 490
rect -298 -38 -236 14
rect -184 -38 -174 14
rect -133 -326 -81 934
rect -10 438 0 490
rect 52 438 62 490
rect 1465 447 1524 481
rect 1368 281 1378 333
rect 1430 281 1440 333
rect -31 14 21 179
rect -41 -38 -31 14
rect 21 -38 31 14
rect -31 -218 21 -38
rect -313 -378 -81 -326
rect -300 -715 -238 -663
rect -186 -715 -176 -663
rect -133 -973 -81 -378
rect -17 -715 -7 -663
rect 45 -715 55 -663
rect 1490 -671 1524 447
rect 1559 281 1569 333
rect 1621 281 1631 333
rect 1483 -705 1524 -671
rect 1578 -820 1612 281
rect 1381 -854 1612 -820
rect -133 -1025 -6 -973
<< via1 >>
rect -238 438 -186 490
rect -236 -38 -184 14
rect 0 438 52 490
rect 1378 281 1430 333
rect -31 -38 21 14
rect -238 -715 -186 -663
rect -7 -715 45 -663
rect 1569 281 1621 333
<< metal2 >>
rect -238 490 -186 500
rect 0 490 52 500
rect -186 438 0 490
rect -238 428 -186 438
rect 0 428 52 438
rect 1378 333 1430 343
rect 1569 333 1621 343
rect 1430 281 1569 333
rect 1378 271 1430 281
rect 1569 271 1621 281
rect -236 14 -184 24
rect -31 14 21 24
rect -184 -38 -31 14
rect -236 -48 -184 -38
rect -31 -48 21 -38
rect -238 -663 -186 -653
rect -7 -663 45 -653
rect -186 -715 -7 -663
rect -238 -725 -186 -715
rect -7 -725 45 -715
use transmission_gate  transmission_gate_0 ~/EE372/incremental_delta_sigma_adc/design/analog_modulator/layout/transmission_gate
timestamp 1652661863
transform 1 0 216 0 1 51
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1652661863
transform 1 0 210 0 1 -1101
box -216 -51 1283 1063
<< end >>
