magic
tech sky130A
magscale 1 2
timestamp 1655484843
<< error_p >>
rect -1531 581 -1473 587
rect -1373 581 -1315 587
rect -1215 581 -1157 587
rect -1057 581 -999 587
rect -899 581 -841 587
rect -741 581 -683 587
rect -583 581 -525 587
rect -425 581 -367 587
rect -267 581 -209 587
rect -109 581 -51 587
rect 51 581 109 587
rect 209 581 267 587
rect 367 581 425 587
rect 525 581 583 587
rect 683 581 741 587
rect 841 581 899 587
rect 999 581 1057 587
rect 1157 581 1215 587
rect 1315 581 1373 587
rect 1473 581 1531 587
rect -1531 547 -1519 581
rect -1373 547 -1361 581
rect -1215 547 -1203 581
rect -1057 547 -1045 581
rect -899 547 -887 581
rect -741 547 -729 581
rect -583 547 -571 581
rect -425 547 -413 581
rect -267 547 -255 581
rect -109 547 -97 581
rect 51 547 63 581
rect 209 547 221 581
rect 367 547 379 581
rect 525 547 537 581
rect 683 547 695 581
rect 841 547 853 581
rect 999 547 1011 581
rect 1157 547 1169 581
rect 1315 547 1327 581
rect 1473 547 1485 581
rect -1531 541 -1473 547
rect -1373 541 -1315 547
rect -1215 541 -1157 547
rect -1057 541 -999 547
rect -899 541 -841 547
rect -741 541 -683 547
rect -583 541 -525 547
rect -425 541 -367 547
rect -267 541 -209 547
rect -109 541 -51 547
rect 51 541 109 547
rect 209 541 267 547
rect 367 541 425 547
rect 525 541 583 547
rect 683 541 741 547
rect 841 541 899 547
rect 999 541 1057 547
rect 1157 541 1215 547
rect 1315 541 1373 547
rect 1473 541 1531 547
rect -1531 -547 -1473 -541
rect -1373 -547 -1315 -541
rect -1215 -547 -1157 -541
rect -1057 -547 -999 -541
rect -899 -547 -841 -541
rect -741 -547 -683 -541
rect -583 -547 -525 -541
rect -425 -547 -367 -541
rect -267 -547 -209 -541
rect -109 -547 -51 -541
rect 51 -547 109 -541
rect 209 -547 267 -541
rect 367 -547 425 -541
rect 525 -547 583 -541
rect 683 -547 741 -541
rect 841 -547 899 -541
rect 999 -547 1057 -541
rect 1157 -547 1215 -541
rect 1315 -547 1373 -541
rect 1473 -547 1531 -541
rect -1531 -581 -1519 -547
rect -1373 -581 -1361 -547
rect -1215 -581 -1203 -547
rect -1057 -581 -1045 -547
rect -899 -581 -887 -547
rect -741 -581 -729 -547
rect -583 -581 -571 -547
rect -425 -581 -413 -547
rect -267 -581 -255 -547
rect -109 -581 -97 -547
rect 51 -581 63 -547
rect 209 -581 221 -547
rect 367 -581 379 -547
rect 525 -581 537 -547
rect 683 -581 695 -547
rect 841 -581 853 -547
rect 999 -581 1011 -547
rect 1157 -581 1169 -547
rect 1315 -581 1327 -547
rect 1473 -581 1485 -547
rect -1531 -587 -1473 -581
rect -1373 -587 -1315 -581
rect -1215 -587 -1157 -581
rect -1057 -587 -999 -581
rect -899 -587 -841 -581
rect -741 -587 -683 -581
rect -583 -587 -525 -581
rect -425 -587 -367 -581
rect -267 -587 -209 -581
rect -109 -587 -51 -581
rect 51 -587 109 -581
rect 209 -587 267 -581
rect 367 -587 425 -581
rect 525 -587 583 -581
rect 683 -587 741 -581
rect 841 -587 899 -581
rect 999 -587 1057 -581
rect 1157 -587 1215 -581
rect 1315 -587 1373 -581
rect 1473 -587 1531 -581
<< nwell >>
rect -1809 -797 1809 797
<< mvpmos >>
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
<< mvpdiff >>
rect -1609 488 -1551 500
rect -1609 -488 -1597 488
rect -1563 -488 -1551 488
rect -1609 -500 -1551 -488
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
rect 1551 488 1609 500
rect 1551 -488 1563 488
rect 1597 -488 1609 488
rect 1551 -500 1609 -488
<< mvpdiffc >>
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
<< mvnsubdiff >>
rect -1743 719 1743 731
rect -1743 685 -1635 719
rect 1635 685 1743 719
rect -1743 673 1743 685
rect -1743 623 -1685 673
rect -1743 -623 -1731 623
rect -1697 -623 -1685 623
rect 1685 623 1743 673
rect -1743 -673 -1685 -623
rect 1685 -623 1697 623
rect 1731 -623 1743 623
rect 1685 -673 1743 -623
rect -1743 -685 1743 -673
rect -1743 -719 -1635 -685
rect 1635 -719 1743 -685
rect -1743 -731 1743 -719
<< mvnsubdiffcont >>
rect -1635 685 1635 719
rect -1731 -623 -1697 623
rect 1697 -623 1731 623
rect -1635 -719 1635 -685
<< poly >>
rect -1551 581 -1451 597
rect -1551 547 -1535 581
rect -1467 547 -1451 581
rect -1551 500 -1451 547
rect -1393 581 -1293 597
rect -1393 547 -1377 581
rect -1309 547 -1293 581
rect -1393 500 -1293 547
rect -1235 581 -1135 597
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1235 500 -1135 547
rect -1077 581 -977 597
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -1077 500 -977 547
rect -919 581 -819 597
rect -919 547 -903 581
rect -835 547 -819 581
rect -919 500 -819 547
rect -761 581 -661 597
rect -761 547 -745 581
rect -677 547 -661 581
rect -761 500 -661 547
rect -603 581 -503 597
rect -603 547 -587 581
rect -519 547 -503 581
rect -603 500 -503 547
rect -445 581 -345 597
rect -445 547 -429 581
rect -361 547 -345 581
rect -445 500 -345 547
rect -287 581 -187 597
rect -287 547 -271 581
rect -203 547 -187 581
rect -287 500 -187 547
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 500 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 500 129 547
rect 187 581 287 597
rect 187 547 203 581
rect 271 547 287 581
rect 187 500 287 547
rect 345 581 445 597
rect 345 547 361 581
rect 429 547 445 581
rect 345 500 445 547
rect 503 581 603 597
rect 503 547 519 581
rect 587 547 603 581
rect 503 500 603 547
rect 661 581 761 597
rect 661 547 677 581
rect 745 547 761 581
rect 661 500 761 547
rect 819 581 919 597
rect 819 547 835 581
rect 903 547 919 581
rect 819 500 919 547
rect 977 581 1077 597
rect 977 547 993 581
rect 1061 547 1077 581
rect 977 500 1077 547
rect 1135 581 1235 597
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1135 500 1235 547
rect 1293 581 1393 597
rect 1293 547 1309 581
rect 1377 547 1393 581
rect 1293 500 1393 547
rect 1451 581 1551 597
rect 1451 547 1467 581
rect 1535 547 1551 581
rect 1451 500 1551 547
rect -1551 -547 -1451 -500
rect -1551 -581 -1535 -547
rect -1467 -581 -1451 -547
rect -1551 -597 -1451 -581
rect -1393 -547 -1293 -500
rect -1393 -581 -1377 -547
rect -1309 -581 -1293 -547
rect -1393 -597 -1293 -581
rect -1235 -547 -1135 -500
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1235 -597 -1135 -581
rect -1077 -547 -977 -500
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -1077 -597 -977 -581
rect -919 -547 -819 -500
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -919 -597 -819 -581
rect -761 -547 -661 -500
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -761 -597 -661 -581
rect -603 -547 -503 -500
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -603 -597 -503 -581
rect -445 -547 -345 -500
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -445 -597 -345 -581
rect -287 -547 -187 -500
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -500
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -500
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -500
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 187 -597 287 -581
rect 345 -547 445 -500
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 345 -597 445 -581
rect 503 -547 603 -500
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 503 -597 603 -581
rect 661 -547 761 -500
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 661 -597 761 -581
rect 819 -547 919 -500
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 819 -597 919 -581
rect 977 -547 1077 -500
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 977 -597 1077 -581
rect 1135 -547 1235 -500
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1135 -597 1235 -581
rect 1293 -547 1393 -500
rect 1293 -581 1309 -547
rect 1377 -581 1393 -547
rect 1293 -597 1393 -581
rect 1451 -547 1551 -500
rect 1451 -581 1467 -547
rect 1535 -581 1551 -547
rect 1451 -597 1551 -581
<< polycont >>
rect -1535 547 -1467 581
rect -1377 547 -1309 581
rect -1219 547 -1151 581
rect -1061 547 -993 581
rect -903 547 -835 581
rect -745 547 -677 581
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect 677 547 745 581
rect 835 547 903 581
rect 993 547 1061 581
rect 1151 547 1219 581
rect 1309 547 1377 581
rect 1467 547 1535 581
rect -1535 -581 -1467 -547
rect -1377 -581 -1309 -547
rect -1219 -581 -1151 -547
rect -1061 -581 -993 -547
rect -903 -581 -835 -547
rect -745 -581 -677 -547
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
rect 677 -581 745 -547
rect 835 -581 903 -547
rect 993 -581 1061 -547
rect 1151 -581 1219 -547
rect 1309 -581 1377 -547
rect 1467 -581 1535 -547
<< locali >>
rect -1731 685 -1635 719
rect 1635 685 1731 719
rect -1731 623 -1697 685
rect 1697 623 1731 685
rect -1551 547 -1535 581
rect -1467 547 -1451 581
rect -1393 547 -1377 581
rect -1309 547 -1293 581
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -919 547 -903 581
rect -835 547 -819 581
rect -761 547 -745 581
rect -677 547 -661 581
rect -603 547 -587 581
rect -519 547 -503 581
rect -445 547 -429 581
rect -361 547 -345 581
rect -287 547 -271 581
rect -203 547 -187 581
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect 187 547 203 581
rect 271 547 287 581
rect 345 547 361 581
rect 429 547 445 581
rect 503 547 519 581
rect 587 547 603 581
rect 661 547 677 581
rect 745 547 761 581
rect 819 547 835 581
rect 903 547 919 581
rect 977 547 993 581
rect 1061 547 1077 581
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1293 547 1309 581
rect 1377 547 1393 581
rect 1451 547 1467 581
rect 1535 547 1551 581
rect -1597 488 -1563 504
rect -1597 -504 -1563 -488
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect 1563 488 1597 504
rect 1563 -504 1597 -488
rect -1551 -581 -1535 -547
rect -1467 -581 -1451 -547
rect -1393 -581 -1377 -547
rect -1309 -581 -1293 -547
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1293 -581 1309 -547
rect 1377 -581 1393 -547
rect 1451 -581 1467 -547
rect 1535 -581 1551 -547
rect -1731 -685 -1697 -623
rect 1697 -685 1731 -623
rect -1731 -719 -1635 -685
rect 1635 -719 1731 -685
<< viali >>
rect -1519 547 -1485 581
rect -1361 547 -1327 581
rect -1203 547 -1169 581
rect -1045 547 -1011 581
rect -887 547 -853 581
rect -729 547 -695 581
rect -571 547 -537 581
rect -413 547 -379 581
rect -255 547 -221 581
rect -97 547 -63 581
rect 63 547 97 581
rect 221 547 255 581
rect 379 547 413 581
rect 537 547 571 581
rect 695 547 729 581
rect 853 547 887 581
rect 1011 547 1045 581
rect 1169 547 1203 581
rect 1327 547 1361 581
rect 1485 547 1519 581
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
rect -1519 -581 -1485 -547
rect -1361 -581 -1327 -547
rect -1203 -581 -1169 -547
rect -1045 -581 -1011 -547
rect -887 -581 -853 -547
rect -729 -581 -695 -547
rect -571 -581 -537 -547
rect -413 -581 -379 -547
rect -255 -581 -221 -547
rect -97 -581 -63 -547
rect 63 -581 97 -547
rect 221 -581 255 -547
rect 379 -581 413 -547
rect 537 -581 571 -547
rect 695 -581 729 -547
rect 853 -581 887 -547
rect 1011 -581 1045 -547
rect 1169 -581 1203 -547
rect 1327 -581 1361 -547
rect 1485 -581 1519 -547
<< metal1 >>
rect -1531 581 -1473 587
rect -1531 547 -1519 581
rect -1485 547 -1473 581
rect -1531 541 -1473 547
rect -1373 581 -1315 587
rect -1373 547 -1361 581
rect -1327 547 -1315 581
rect -1373 541 -1315 547
rect -1215 581 -1157 587
rect -1215 547 -1203 581
rect -1169 547 -1157 581
rect -1215 541 -1157 547
rect -1057 581 -999 587
rect -1057 547 -1045 581
rect -1011 547 -999 581
rect -1057 541 -999 547
rect -899 581 -841 587
rect -899 547 -887 581
rect -853 547 -841 581
rect -899 541 -841 547
rect -741 581 -683 587
rect -741 547 -729 581
rect -695 547 -683 581
rect -741 541 -683 547
rect -583 581 -525 587
rect -583 547 -571 581
rect -537 547 -525 581
rect -583 541 -525 547
rect -425 581 -367 587
rect -425 547 -413 581
rect -379 547 -367 581
rect -425 541 -367 547
rect -267 581 -209 587
rect -267 547 -255 581
rect -221 547 -209 581
rect -267 541 -209 547
rect -109 581 -51 587
rect -109 547 -97 581
rect -63 547 -51 581
rect -109 541 -51 547
rect 51 581 109 587
rect 51 547 63 581
rect 97 547 109 581
rect 51 541 109 547
rect 209 581 267 587
rect 209 547 221 581
rect 255 547 267 581
rect 209 541 267 547
rect 367 581 425 587
rect 367 547 379 581
rect 413 547 425 581
rect 367 541 425 547
rect 525 581 583 587
rect 525 547 537 581
rect 571 547 583 581
rect 525 541 583 547
rect 683 581 741 587
rect 683 547 695 581
rect 729 547 741 581
rect 683 541 741 547
rect 841 581 899 587
rect 841 547 853 581
rect 887 547 899 581
rect 841 541 899 547
rect 999 581 1057 587
rect 999 547 1011 581
rect 1045 547 1057 581
rect 999 541 1057 547
rect 1157 581 1215 587
rect 1157 547 1169 581
rect 1203 547 1215 581
rect 1157 541 1215 547
rect 1315 581 1373 587
rect 1315 547 1327 581
rect 1361 547 1373 581
rect 1315 541 1373 547
rect 1473 581 1531 587
rect 1473 547 1485 581
rect 1519 547 1531 581
rect 1473 541 1531 547
rect -1603 488 -1557 500
rect -1603 -488 -1597 488
rect -1563 -488 -1557 488
rect -1603 -500 -1557 -488
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect 1557 488 1603 500
rect 1557 -488 1563 488
rect 1597 -488 1603 488
rect 1557 -500 1603 -488
rect -1531 -547 -1473 -541
rect -1531 -581 -1519 -547
rect -1485 -581 -1473 -547
rect -1531 -587 -1473 -581
rect -1373 -547 -1315 -541
rect -1373 -581 -1361 -547
rect -1327 -581 -1315 -547
rect -1373 -587 -1315 -581
rect -1215 -547 -1157 -541
rect -1215 -581 -1203 -547
rect -1169 -581 -1157 -547
rect -1215 -587 -1157 -581
rect -1057 -547 -999 -541
rect -1057 -581 -1045 -547
rect -1011 -581 -999 -547
rect -1057 -587 -999 -581
rect -899 -547 -841 -541
rect -899 -581 -887 -547
rect -853 -581 -841 -547
rect -899 -587 -841 -581
rect -741 -547 -683 -541
rect -741 -581 -729 -547
rect -695 -581 -683 -547
rect -741 -587 -683 -581
rect -583 -547 -525 -541
rect -583 -581 -571 -547
rect -537 -581 -525 -547
rect -583 -587 -525 -581
rect -425 -547 -367 -541
rect -425 -581 -413 -547
rect -379 -581 -367 -547
rect -425 -587 -367 -581
rect -267 -547 -209 -541
rect -267 -581 -255 -547
rect -221 -581 -209 -547
rect -267 -587 -209 -581
rect -109 -547 -51 -541
rect -109 -581 -97 -547
rect -63 -581 -51 -547
rect -109 -587 -51 -581
rect 51 -547 109 -541
rect 51 -581 63 -547
rect 97 -581 109 -547
rect 51 -587 109 -581
rect 209 -547 267 -541
rect 209 -581 221 -547
rect 255 -581 267 -547
rect 209 -587 267 -581
rect 367 -547 425 -541
rect 367 -581 379 -547
rect 413 -581 425 -547
rect 367 -587 425 -581
rect 525 -547 583 -541
rect 525 -581 537 -547
rect 571 -581 583 -547
rect 525 -587 583 -581
rect 683 -547 741 -541
rect 683 -581 695 -547
rect 729 -581 741 -547
rect 683 -587 741 -581
rect 841 -547 899 -541
rect 841 -581 853 -547
rect 887 -581 899 -547
rect 841 -587 899 -581
rect 999 -547 1057 -541
rect 999 -581 1011 -547
rect 1045 -581 1057 -547
rect 999 -587 1057 -581
rect 1157 -547 1215 -541
rect 1157 -581 1169 -547
rect 1203 -581 1215 -547
rect 1157 -587 1215 -581
rect 1315 -547 1373 -541
rect 1315 -581 1327 -547
rect 1361 -581 1373 -547
rect 1315 -587 1373 -581
rect 1473 -547 1531 -541
rect 1473 -581 1485 -547
rect 1519 -581 1531 -547
rect 1473 -587 1531 -581
<< properties >>
string FIXED_BBOX -1714 -702 1714 702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
