magic
tech sky130A
magscale 1 2
timestamp 1654656593
<< nwell >>
rect 599 4730 7350 6437
<< pwell >>
rect -428 -610 8353 4694
<< psubdiff >>
rect 8274 4649 8323 4650
rect 3135 4600 3281 4649
rect 8057 4600 8323 4649
rect 3135 4534 3184 4600
rect 3135 -541 3184 -462
rect 8274 4517 8323 4600
rect 8274 -541 8323 -498
rect 3135 -590 3275 -541
rect 8165 -590 8323 -541
<< nsubdiff >>
rect 664 6346 769 6380
rect 7174 6346 7283 6380
rect 664 6308 698 6346
rect 664 4802 698 4872
rect 7249 6281 7283 6346
rect 7249 4802 7283 4914
rect 664 4768 784 4802
rect 7177 4768 7283 4802
<< psubdiffcont >>
rect 3281 4600 8057 4649
rect 3135 -462 3184 4534
rect 8274 -498 8323 4517
rect 3275 -590 8165 -541
<< nsubdiffcont >>
rect 769 6346 7174 6380
rect 664 4872 698 6308
rect 7249 4914 7283 6281
rect 784 4768 7177 4802
<< locali >>
rect -430 6380 8656 6436
rect -430 6346 769 6380
rect 7174 6346 8656 6380
rect -430 6308 8656 6346
rect 972 4942 1100 6308
rect 2521 4942 2649 6308
rect 3177 4943 3305 6308
rect 4717 4936 4845 6308
rect 5369 4945 5497 6308
rect 6910 4942 7038 6308
rect 7249 6281 7283 6308
rect 664 4802 698 4872
rect 7249 4802 7283 4914
rect 664 4768 784 4802
rect 7177 4768 7283 4802
rect 8274 4649 8323 4650
rect -378 -462 -250 4625
rect 115 2099 243 2109
rect 115 17 309 2099
rect 2259 2091 2387 2112
rect 2259 17 2445 2091
rect 115 -17 264 17
rect 2292 -17 2445 17
rect 115 -462 309 -17
rect 495 -462 2119 -17
rect 2259 -462 2445 -17
rect 2625 -462 2753 4617
rect 3135 4600 3281 4649
rect 8057 4600 8323 4649
rect 3135 4534 3184 4600
rect 3184 2863 3281 4534
rect 8154 4517 8203 4600
rect 3184 2735 3806 2863
rect 3184 -462 3281 2735
rect 8066 2863 8203 4517
rect 4510 2735 8203 2863
rect 3565 -11 3693 10
rect 3565 -98 3579 -11
rect 3672 -98 3693 -11
rect 3565 -462 3693 -98
rect 4984 0 5112 19
rect 4984 -87 5001 0
rect 5094 -87 5112 0
rect 4984 -462 5112 -87
rect 5234 -462 5362 2735
rect 5874 21 6002 2735
rect 8066 1888 8203 2735
rect 7946 1751 8203 1888
rect 8066 1371 8203 1751
rect 7955 1234 8203 1371
rect 8066 885 8203 1234
rect 7945 748 8203 885
rect 8066 383 8203 748
rect 7931 246 8203 383
rect 8066 21 8203 246
rect 5874 3 8203 21
rect 5874 -94 6259 3
rect 6362 2 8203 3
rect 6362 -94 7429 2
rect 5874 -95 7429 -94
rect 7532 -95 8203 2
rect 5874 -107 8203 -95
rect 5874 -462 6002 -107
rect 8066 -462 8203 -107
rect 8274 4517 8323 4600
rect -430 -482 8274 -462
rect -430 -484 7430 -482
rect -430 -489 5006 -484
rect -430 -541 3579 -489
rect 3672 -541 5006 -489
rect 5099 -488 7430 -484
rect 5099 -541 6269 -488
rect 6362 -541 7430 -488
rect 7523 -498 8274 -482
rect 8323 -498 8656 -462
rect 7523 -541 8656 -498
rect -430 -590 3275 -541
rect 8165 -590 8656 -541
<< viali >>
rect 769 6346 7174 6380
rect -72 4393 -38 4427
rect 284 4393 318 4427
rect 640 4393 674 4427
rect 996 4393 1030 4427
rect 1352 4393 1386 4427
rect 1708 4393 1742 4427
rect 2064 4393 2098 4427
rect 2420 4393 2454 4427
rect 106 4171 140 4205
rect 462 4171 496 4205
rect 818 4171 852 4205
rect 1174 4171 1208 4205
rect 1530 4171 1564 4205
rect 1886 4171 1920 4205
rect 2242 4171 2276 4205
rect -72 3895 -38 3929
rect 284 3895 318 3929
rect 640 3895 674 3929
rect 996 3895 1030 3929
rect 1352 3895 1386 3929
rect 1708 3895 1742 3929
rect 2064 3895 2098 3929
rect 2420 3895 2454 3929
rect 106 3673 140 3707
rect 462 3673 496 3707
rect 818 3673 852 3707
rect 1174 3673 1208 3707
rect 1530 3673 1564 3707
rect 1886 3673 1920 3707
rect 2242 3673 2276 3707
rect -72 3397 -38 3431
rect 284 3397 318 3431
rect 640 3397 674 3431
rect 996 3397 1030 3431
rect 1352 3397 1386 3431
rect 1708 3397 1742 3431
rect 2064 3397 2098 3431
rect 2420 3397 2454 3431
rect 106 3175 140 3209
rect 462 3175 496 3209
rect 818 3175 852 3209
rect 1174 3175 1208 3209
rect 1530 3175 1564 3209
rect 1886 3175 1920 3209
rect 2242 3175 2276 3209
rect -72 2899 -38 2933
rect 284 2899 318 2933
rect 640 2899 674 2933
rect 996 2899 1030 2933
rect 1352 2899 1386 2933
rect 1708 2899 1742 2933
rect 2064 2899 2098 2933
rect 2420 2899 2454 2933
rect 106 2677 140 2711
rect 462 2677 496 2711
rect 818 2677 852 2711
rect 1174 2677 1208 2711
rect 1530 2677 1564 2711
rect 1886 2677 1920 2711
rect 2242 2677 2276 2711
rect -223 2491 2588 2525
rect 460 1885 494 1919
rect 816 1885 850 1919
rect 1172 1885 1206 1919
rect 1528 1885 1562 1919
rect 1884 1885 1918 1919
rect 638 1663 672 1697
rect 994 1663 1028 1697
rect 1350 1663 1384 1697
rect 1706 1663 1740 1697
rect 2062 1663 2096 1697
rect 460 1387 494 1421
rect 816 1387 850 1421
rect 1172 1387 1206 1421
rect 1528 1387 1562 1421
rect 1884 1387 1918 1421
rect 638 1165 672 1199
rect 994 1165 1028 1199
rect 1350 1165 1384 1199
rect 1706 1165 1740 1199
rect 2062 1165 2096 1199
rect 460 859 494 893
rect 816 859 850 893
rect 1172 859 1206 893
rect 1528 859 1562 893
rect 1884 859 1918 893
rect 638 697 672 731
rect 994 697 1028 731
rect 1350 697 1384 731
rect 1706 697 1740 731
rect 2062 697 2096 731
rect 460 361 494 395
rect 816 361 850 395
rect 1172 361 1206 395
rect 1528 361 1562 395
rect 1884 361 1918 395
rect 638 199 672 233
rect 994 199 1028 233
rect 1350 199 1384 233
rect 1706 199 1740 233
rect 2062 199 2096 233
rect 264 -17 2292 17
rect 3429 4402 3463 4436
rect 3785 4402 3819 4436
rect 4141 4402 4175 4436
rect 4497 4402 4531 4436
rect 4853 4402 4887 4436
rect 5209 4402 5243 4436
rect 5565 4402 5599 4436
rect 5921 4402 5955 4436
rect 6277 4402 6311 4436
rect 6633 4402 6667 4436
rect 6989 4402 7023 4436
rect 7345 4402 7379 4436
rect 7701 4402 7735 4436
rect 3607 4180 3641 4214
rect 3963 4180 3997 4214
rect 4319 4180 4353 4214
rect 4675 4180 4709 4214
rect 5031 4180 5065 4214
rect 5387 4180 5421 4214
rect 5743 4180 5777 4214
rect 6099 4180 6133 4214
rect 6455 4180 6489 4214
rect 6811 4180 6845 4214
rect 7167 4180 7201 4214
rect 7523 4180 7557 4214
rect 7879 4180 7913 4214
rect 3429 3902 3463 3936
rect 3785 3902 3819 3936
rect 4141 3902 4175 3936
rect 4497 3902 4531 3936
rect 4853 3902 4887 3936
rect 5209 3902 5243 3936
rect 5565 3902 5599 3936
rect 5921 3902 5955 3936
rect 6277 3902 6311 3936
rect 6633 3902 6667 3936
rect 6989 3902 7023 3936
rect 7345 3902 7379 3936
rect 7701 3902 7735 3936
rect 3607 3680 3641 3714
rect 3963 3680 3997 3714
rect 4319 3680 4353 3714
rect 4675 3680 4709 3714
rect 5031 3680 5065 3714
rect 5387 3680 5421 3714
rect 5743 3680 5777 3714
rect 6099 3680 6133 3714
rect 6455 3680 6489 3714
rect 6811 3680 6845 3714
rect 7167 3680 7201 3714
rect 7523 3680 7557 3714
rect 7879 3680 7913 3714
rect 3965 2836 3999 2932
rect 4143 2676 4177 2793
rect 4321 2676 4355 2932
rect 3433 1959 3467 1993
rect 3789 1959 3823 1993
rect 4145 1959 4179 1993
rect 4501 1959 4535 1993
rect 4857 1959 4891 1993
rect 3611 1737 3645 1771
rect 3967 1737 4001 1771
rect 4323 1737 4357 1771
rect 4679 1737 4713 1771
rect 5035 1737 5069 1771
rect 3433 1459 3467 1493
rect 3789 1459 3823 1493
rect 4145 1459 4179 1493
rect 4501 1459 4535 1493
rect 4857 1459 4891 1493
rect 3611 1237 3645 1271
rect 3967 1237 4001 1271
rect 4323 1237 4357 1271
rect 4679 1237 4713 1271
rect 5035 1237 5069 1271
rect 3433 899 3467 933
rect 3789 899 3823 933
rect 4145 899 4179 933
rect 4501 899 4535 933
rect 4857 899 4891 933
rect 3611 677 3645 711
rect 3967 677 4001 711
rect 4323 677 4357 711
rect 4679 677 4713 711
rect 5035 677 5069 711
rect 3433 399 3467 433
rect 3789 399 3823 433
rect 4145 399 4179 433
rect 4501 399 4535 433
rect 4857 399 4891 433
rect 3611 177 3645 211
rect 3967 177 4001 211
rect 4323 177 4357 211
rect 4679 177 4713 211
rect 5035 177 5069 211
rect 3579 -98 3672 -11
rect 5001 -87 5094 0
rect 6259 -94 6362 3
rect 7429 -95 7532 2
rect 3579 -541 3672 -489
rect 5006 -541 5099 -484
rect 6269 -541 6362 -488
rect 7430 -541 7523 -482
rect 3275 -590 8165 -541
<< metal1 >>
rect -256 6380 8656 6436
rect -256 6346 769 6380
rect 7174 6346 8656 6380
rect -256 6308 8656 6346
rect 1442 6228 2190 6308
rect 1443 6193 2190 6228
rect 1243 5997 1253 6055
rect 1311 5997 1321 6055
rect 1443 6053 1478 6193
rect 1599 5997 1609 6055
rect 1667 5997 1677 6055
rect 1798 6041 1833 6193
rect 1955 5997 1965 6055
rect 2023 5997 2033 6055
rect 2155 6045 2190 6193
rect 3642 6192 4390 6308
rect 2311 5997 2321 6055
rect 2379 5997 2389 6055
rect 3443 5997 3453 6055
rect 3511 5997 3521 6055
rect 3642 6051 3677 6192
rect 3799 5997 3809 6055
rect 3867 5997 3877 6055
rect 3998 6038 4033 6192
rect 4155 5997 4165 6055
rect 4223 5997 4233 6055
rect 4355 6026 4390 6192
rect 5843 6202 6591 6308
rect 4510 5997 4520 6055
rect 4578 5997 4588 6055
rect 5643 5997 5653 6055
rect 5711 5997 5721 6055
rect 5843 6053 5878 6202
rect 5999 5997 6009 6055
rect 6067 5997 6077 6055
rect 6199 6039 6234 6202
rect 6355 5997 6365 6055
rect 6423 5997 6433 6055
rect 6555 6039 6590 6202
rect 6711 5997 6721 6055
rect 6779 5997 6789 6055
rect 1421 5799 1431 5857
rect 1489 5799 1499 5857
rect 1777 5799 1787 5857
rect 1845 5799 1855 5857
rect 2133 5799 2143 5857
rect 2201 5799 2211 5857
rect 3621 5799 3631 5857
rect 3689 5799 3699 5857
rect 3977 5798 3987 5856
rect 4045 5798 4055 5856
rect 4333 5799 4343 5857
rect 4401 5799 4411 5857
rect 5821 5799 5831 5857
rect 5889 5799 5899 5857
rect 6177 5799 6187 5857
rect 6245 5799 6255 5857
rect 6533 5799 6543 5857
rect 6601 5799 6611 5857
rect 1332 5688 1342 5746
rect 1400 5740 1410 5746
rect 6199 5740 6234 5741
rect 1400 5706 2273 5740
rect 3583 5706 4459 5740
rect 5786 5706 6662 5740
rect 1400 5688 1410 5706
rect 1798 5617 1915 5706
rect 3956 5617 4073 5706
rect 6158 5617 6275 5706
rect 1798 5500 8372 5617
rect 1169 5230 1179 5288
rect 1310 5230 1320 5288
rect 1598 5230 1608 5288
rect 1666 5230 1676 5288
rect 1954 5230 1964 5288
rect 2022 5230 2032 5288
rect 2309 5230 2319 5288
rect 2377 5230 2387 5288
rect 3442 5230 3452 5288
rect 3510 5230 3520 5288
rect 3798 5230 3808 5288
rect 3866 5230 3876 5288
rect 4154 5230 4164 5288
rect 4222 5230 4232 5288
rect 4510 5230 4520 5288
rect 4578 5230 4588 5288
rect 5642 5230 5652 5288
rect 5710 5230 5720 5288
rect 5998 5230 6008 5288
rect 6066 5230 6076 5288
rect 6354 5230 6364 5288
rect 6422 5230 6432 5288
rect 6710 5230 6720 5288
rect 6778 5230 6788 5288
rect 1420 5032 1430 5090
rect 1488 5032 1498 5090
rect 1776 5032 1786 5090
rect 1844 5032 1854 5090
rect 2131 5032 2141 5090
rect 2199 5032 2209 5090
rect 3620 5032 3630 5090
rect 3688 5032 3698 5090
rect 3976 5032 3986 5090
rect 4044 5032 4054 5090
rect 4331 5032 4341 5090
rect 4399 5032 4409 5090
rect 5821 5032 5831 5090
rect 5889 5032 5899 5090
rect 6176 5032 6186 5090
rect 6244 5032 6254 5090
rect 6532 5032 6542 5090
rect 6600 5032 6610 5090
rect 2220 4973 2230 4979
rect 1332 4939 2230 4973
rect 1798 4851 1915 4939
rect 2220 4921 2230 4939
rect 2288 4921 2298 4979
rect 3532 4939 4498 4973
rect 5732 4939 6778 4973
rect 3949 4851 4066 4939
rect 6156 4851 6273 4939
rect 1798 4734 8372 4851
rect -378 2569 -250 4625
rect 1116 4511 1164 4530
rect -95 4504 1164 4511
rect -95 4495 451 4504
rect -95 4411 -84 4495
rect -26 4427 451 4495
rect -94 4375 -84 4411
rect -26 4393 284 4427
rect 318 4415 451 4427
rect 509 4427 1164 4504
rect 509 4415 640 4427
rect 318 4393 640 4415
rect 674 4393 996 4427
rect 1030 4393 1164 4427
rect -26 4390 1164 4393
rect 1310 4511 1320 4530
rect 1310 4499 2475 4511
rect 1310 4427 1874 4499
rect 1310 4393 1352 4427
rect 1386 4393 1708 4427
rect 1742 4410 1874 4427
rect 1932 4495 2475 4499
rect 1932 4427 2408 4495
rect 1932 4410 2064 4427
rect 1742 4393 2064 4410
rect 2098 4393 2408 4427
rect 1310 4390 2408 4393
rect -26 4387 2408 4390
rect -26 4375 -16 4387
rect 2398 4375 2408 4387
rect 2466 4375 2476 4495
rect 84 4165 94 4223
rect 152 4211 162 4223
rect 794 4211 804 4224
rect 152 4205 804 4211
rect 862 4211 872 4224
rect 1508 4211 1518 4220
rect 862 4205 1518 4211
rect 1576 4211 1586 4220
rect 2220 4211 2230 4223
rect 1576 4205 2230 4211
rect 152 4171 462 4205
rect 496 4171 804 4205
rect 862 4171 1174 4205
rect 1208 4171 1518 4205
rect 1576 4171 1886 4205
rect 1920 4171 2230 4205
rect 152 4166 804 4171
rect 862 4166 1518 4171
rect 152 4165 1518 4166
rect 1508 4162 1518 4165
rect 1576 4165 2230 4171
rect 2288 4165 2298 4223
rect 1576 4162 1586 4165
rect -95 4119 2473 4122
rect -95 4112 1163 4119
rect -95 4105 450 4112
rect -95 3910 -84 4105
rect -26 3929 450 4105
rect -94 3877 -84 3910
rect -26 3895 284 3929
rect 318 3904 450 3929
rect 508 3929 1163 4112
rect 508 3904 640 3929
rect 318 3895 640 3904
rect 674 3895 996 3929
rect 1030 3911 1163 3929
rect 1221 4114 2473 4119
rect 1221 4108 2407 4114
rect 1221 3929 1873 4108
rect 1221 3911 1352 3929
rect 1030 3895 1352 3911
rect 1386 3895 1708 3929
rect 1742 3900 1873 3929
rect 1931 3929 2407 4108
rect 2465 3935 2475 4114
rect 1931 3900 2064 3929
rect 1742 3895 2064 3900
rect 2098 3906 2407 3929
rect 2098 3895 2408 3906
rect -26 3889 2408 3895
rect -26 3877 -16 3889
rect 2398 3877 2408 3889
rect 2466 3877 2476 3935
rect 84 3667 94 3725
rect 152 3713 162 3725
rect 795 3713 805 3723
rect 152 3707 805 3713
rect 863 3713 873 3723
rect 1508 3713 1518 3720
rect 863 3707 1518 3713
rect 1576 3713 1586 3720
rect 2220 3713 2230 3725
rect 1576 3707 2230 3713
rect 152 3673 462 3707
rect 496 3673 805 3707
rect 863 3673 1174 3707
rect 1208 3673 1518 3707
rect 1576 3673 1886 3707
rect 1920 3673 2230 3707
rect 152 3667 805 3673
rect 795 3665 805 3667
rect 863 3667 1518 3673
rect 863 3665 873 3667
rect 1508 3662 1518 3667
rect 1576 3667 2230 3673
rect 2288 3667 2298 3725
rect 1576 3662 1586 3667
rect -94 3619 2474 3623
rect -94 3607 450 3619
rect -94 3437 -83 3607
rect -94 3379 -84 3437
rect -25 3431 450 3607
rect -25 3399 284 3431
rect -26 3397 284 3399
rect 318 3411 450 3431
rect 508 3613 2474 3619
rect 508 3612 2408 3613
rect 508 3431 1161 3612
rect 508 3411 640 3431
rect 318 3397 640 3411
rect 674 3397 996 3431
rect 1030 3404 1161 3431
rect 1219 3431 1874 3612
rect 1219 3404 1352 3431
rect 1030 3397 1352 3404
rect 1386 3397 1708 3431
rect 1742 3404 1874 3431
rect 1932 3431 2408 3612
rect 1932 3404 2064 3431
rect 1742 3397 2064 3404
rect 2098 3397 2408 3431
rect -26 3391 2408 3397
rect -26 3379 -16 3391
rect 2398 3379 2408 3391
rect 2466 3379 2476 3613
rect 84 3169 94 3227
rect 152 3215 162 3227
rect 799 3215 809 3230
rect 152 3209 809 3215
rect 867 3215 877 3230
rect 1508 3215 1518 3226
rect 867 3209 1518 3215
rect 1576 3215 1586 3226
rect 2220 3215 2230 3227
rect 1576 3209 2230 3215
rect 152 3175 462 3209
rect 496 3175 809 3209
rect 867 3175 1174 3209
rect 1208 3175 1518 3209
rect 1576 3175 1886 3209
rect 1920 3175 2230 3209
rect 152 3172 809 3175
rect 867 3172 1518 3175
rect 152 3169 1518 3172
rect 1508 3168 1518 3169
rect 1576 3169 2230 3175
rect 2288 3169 2298 3227
rect 1576 3168 1586 3169
rect -94 2881 -84 3125
rect -26 3095 8 3125
rect 60 3115 2408 3125
rect 60 3112 1875 3115
rect 60 3110 1163 3112
rect 60 3109 450 3110
rect 23 3095 450 3109
rect -26 3016 450 3095
rect -26 2985 8 3016
rect 11 2985 450 3016
rect -26 2933 450 2985
rect -26 2899 284 2933
rect 318 2902 450 2933
rect 508 2933 1163 3110
rect 508 2902 640 2933
rect 318 2899 640 2902
rect 674 2899 996 2933
rect 1030 2904 1163 2933
rect 1221 2933 1875 3112
rect 1221 2904 1352 2933
rect 1030 2899 1352 2904
rect 1386 2899 1708 2933
rect 1742 2907 1875 2933
rect 1933 2933 2408 3115
rect 1933 2907 2064 2933
rect 1742 2899 2064 2907
rect 2098 2899 2408 2933
rect -26 2893 2408 2899
rect -26 2881 -16 2893
rect 2398 2881 2408 2893
rect 2466 2881 2476 3125
rect 84 2671 94 2729
rect 152 2717 162 2729
rect 438 2717 448 2727
rect 152 2671 448 2717
rect 506 2717 516 2727
rect 794 2717 804 2726
rect 438 2669 448 2671
rect 506 2671 804 2717
rect 862 2717 872 2726
rect 1150 2717 1160 2729
rect 506 2669 516 2671
rect 794 2668 804 2671
rect 862 2671 1160 2717
rect 1218 2717 1228 2729
rect 1507 2717 1517 2728
rect 1218 2671 1517 2717
rect 1575 2717 1585 2728
rect 1863 2717 1873 2728
rect 862 2668 872 2671
rect 1507 2670 1517 2671
rect 1575 2671 1873 2717
rect 1931 2717 1941 2728
rect 2220 2717 2230 2729
rect 1575 2670 1585 2671
rect 1863 2670 1873 2671
rect 1931 2671 2230 2717
rect 2288 2671 2298 2729
rect 1931 2670 1941 2671
rect -386 2441 -378 2543
rect 2625 2543 2753 4617
rect 3429 4446 7850 4520
rect 3383 4329 3393 4446
rect 3510 4442 7850 4446
rect 3510 4436 5553 4442
rect 5611 4436 7689 4442
rect 3510 4402 3785 4436
rect 3819 4402 4141 4436
rect 4175 4402 4497 4436
rect 4531 4402 4853 4436
rect 4887 4402 5209 4436
rect 5243 4402 5553 4436
rect 5611 4402 5921 4436
rect 5955 4402 6277 4436
rect 6311 4402 6633 4436
rect 6667 4402 6989 4436
rect 7023 4402 7345 4436
rect 7379 4402 7689 4436
rect 3510 4384 5553 4402
rect 5611 4384 7689 4402
rect 7747 4384 7850 4442
rect 3510 4380 7850 4384
rect 3510 4374 7757 4380
rect 3510 4329 3520 4374
rect 3585 4232 7935 4259
rect 3585 4174 3595 4232
rect 3653 4214 5731 4232
rect 5789 4214 7867 4232
rect 3653 4180 3963 4214
rect 3997 4180 4319 4214
rect 4353 4180 4675 4214
rect 4709 4180 5031 4214
rect 5065 4180 5387 4214
rect 5421 4180 5731 4214
rect 5789 4180 6099 4214
rect 6133 4180 6455 4214
rect 6489 4180 6811 4214
rect 6845 4180 7167 4214
rect 7201 4180 7523 4214
rect 7557 4180 7867 4214
rect 3653 4174 5731 4180
rect 5789 4174 7867 4180
rect 7925 4174 7935 4232
rect 3428 4105 7843 4131
rect 3428 4019 7845 4105
rect 3428 3942 7843 4019
rect 3382 3825 3392 3942
rect 3509 3936 5553 3942
rect 5611 3936 7689 3942
rect 3509 3902 3785 3936
rect 3819 3902 4141 3936
rect 4175 3902 4497 3936
rect 4531 3902 4853 3936
rect 4887 3902 5209 3936
rect 5243 3902 5553 3936
rect 5611 3902 5921 3936
rect 5955 3902 6277 3936
rect 6311 3902 6633 3936
rect 6667 3902 6989 3936
rect 7023 3902 7345 3936
rect 7379 3902 7689 3936
rect 3509 3884 5553 3902
rect 5611 3884 7689 3902
rect 7747 3884 7843 3942
rect 3509 3861 7843 3884
rect 3509 3825 3519 3861
rect 3585 3674 3595 3732
rect 3653 3720 3663 3732
rect 3879 3720 3889 3776
rect 3653 3675 3889 3720
rect 4011 3720 4021 3776
rect 5721 3720 5731 3732
rect 4011 3714 5731 3720
rect 5789 3720 5799 3732
rect 7857 3720 7867 3732
rect 5789 3714 7867 3720
rect 4011 3680 4319 3714
rect 4353 3680 4675 3714
rect 4709 3680 5031 3714
rect 5065 3680 5387 3714
rect 5421 3680 5731 3714
rect 5789 3680 6099 3714
rect 6133 3680 6455 3714
rect 6489 3680 6811 3714
rect 6845 3680 7167 3714
rect 7201 3680 7523 3714
rect 7557 3680 7867 3714
rect 3653 3674 3953 3675
rect 4011 3674 5731 3680
rect 5789 3674 7867 3680
rect 7925 3674 7935 3732
rect 4094 3630 4255 3636
rect 3551 3596 4131 3630
rect 4094 3590 4131 3596
rect 4121 3572 4131 3590
rect 4189 3596 7809 3630
rect 4189 3590 4255 3596
rect 4189 3572 4199 3590
rect 3879 3396 3889 3514
rect 4011 3397 8403 3514
rect 4011 3396 4021 3397
rect 4121 3022 4131 3040
rect 4089 3016 4131 3022
rect 3879 2982 4131 3016
rect 4189 3022 4199 3040
rect 4189 3016 4257 3022
rect 4189 2982 4442 3016
rect 4089 2976 4257 2982
rect 3959 2939 4005 2944
rect 3879 2822 3889 2939
rect 4010 2938 4020 2939
rect 4315 2938 4361 2944
rect 4011 2932 4373 2938
rect 4011 2919 4321 2932
rect 4355 2919 4373 2932
rect 4011 2882 4309 2919
rect 4011 2880 4026 2882
rect 4291 2881 4309 2882
rect 4010 2822 4026 2880
rect 4121 2668 4131 2805
rect 4189 2668 4199 2805
rect 4121 2664 4199 2668
rect 4299 2667 4309 2881
rect 4367 2667 4377 2919
rect 4315 2664 4361 2667
rect -250 2525 2753 2543
rect -250 2491 -223 2525
rect 2588 2491 2753 2525
rect -250 2441 2753 2491
rect 153 1969 2030 2003
rect 153 1607 281 1969
rect 794 1925 804 1928
rect 438 1867 448 1925
rect 506 1879 804 1925
rect 862 1925 872 1928
rect 1507 1925 1517 1926
rect 506 1867 516 1879
rect 794 1870 804 1879
rect 862 1879 1160 1925
rect 862 1870 872 1879
rect 1150 1867 1160 1879
rect 1218 1879 1517 1925
rect 1575 1925 1585 1926
rect 1218 1867 1228 1879
rect 1507 1868 1517 1879
rect 1575 1879 1872 1925
rect 1575 1868 1585 1879
rect 1862 1867 1872 1879
rect 1930 1867 1940 1925
rect 616 1657 626 1715
rect 684 1703 694 1715
rect 1328 1703 1338 1710
rect 684 1697 1338 1703
rect 1396 1703 1406 1710
rect 2040 1703 2050 1715
rect 1396 1697 2050 1703
rect 684 1663 994 1697
rect 1028 1663 1338 1697
rect 1396 1663 1706 1697
rect 1740 1663 2050 1697
rect 684 1657 1338 1663
rect 1328 1652 1338 1657
rect 1396 1657 2050 1663
rect 2108 1657 2118 1715
rect 1396 1652 1406 1657
rect 580 1607 2003 1613
rect 153 1479 2038 1607
rect 153 1109 281 1479
rect 557 1471 1980 1479
rect 1149 1427 1159 1430
rect 438 1369 448 1427
rect 506 1381 804 1427
rect 506 1369 516 1381
rect 794 1369 804 1381
rect 862 1381 1159 1427
rect 1217 1427 1227 1430
rect 1507 1427 1517 1429
rect 862 1369 872 1381
rect 1149 1372 1159 1381
rect 1217 1381 1517 1427
rect 1575 1427 1585 1429
rect 1217 1372 1227 1381
rect 1507 1371 1517 1381
rect 1575 1381 1872 1427
rect 1575 1371 1585 1381
rect 1862 1369 1872 1381
rect 1930 1369 1940 1427
rect 616 1160 626 1218
rect 684 1205 694 1218
rect 1328 1205 1338 1216
rect 684 1199 1338 1205
rect 1396 1205 1406 1216
rect 2040 1205 2050 1216
rect 1396 1199 2050 1205
rect 684 1165 994 1199
rect 1028 1165 1338 1199
rect 1396 1165 1706 1199
rect 1740 1165 2050 1199
rect 684 1160 1338 1165
rect 626 1159 1338 1160
rect 1328 1158 1338 1159
rect 1396 1159 2050 1165
rect 1396 1158 1406 1159
rect 2040 1158 2050 1159
rect 2108 1158 2118 1216
rect 592 1109 2015 1115
rect 153 981 2038 1109
rect 153 609 281 981
rect 460 973 1994 981
rect 460 899 494 973
rect 816 899 850 973
rect 1172 907 1206 973
rect 1150 899 1160 907
rect 438 841 448 899
rect 506 893 1160 899
rect 1218 899 1228 907
rect 1528 899 1562 973
rect 1884 899 1918 973
rect 1218 893 1872 899
rect 506 859 816 893
rect 850 859 1160 893
rect 1218 859 1528 893
rect 1562 859 1872 893
rect 506 853 1160 859
rect 506 841 516 853
rect 1150 849 1160 853
rect 1218 853 1872 859
rect 1218 849 1228 853
rect 1862 841 1872 853
rect 1930 841 1940 899
rect 616 691 626 749
rect 684 737 694 749
rect 1329 737 1339 748
rect 684 731 1339 737
rect 1397 737 1407 748
rect 2040 737 2050 748
rect 1397 731 2050 737
rect 684 697 994 731
rect 1028 697 1339 731
rect 1397 697 1706 731
rect 1740 697 2050 731
rect 684 691 1339 697
rect 1329 690 1339 691
rect 1397 691 2050 697
rect 1397 690 1407 691
rect 2040 690 2050 691
rect 2108 690 2118 748
rect 445 609 2006 617
rect -100 481 2032 609
rect 153 119 281 481
rect 445 475 2004 481
rect 460 401 494 475
rect 816 401 850 475
rect 1172 409 1206 475
rect 1150 401 1160 409
rect 438 343 448 401
rect 506 395 1160 401
rect 1218 401 1228 409
rect 1528 401 1562 475
rect 1884 401 1918 475
rect 1218 395 1872 401
rect 506 361 816 395
rect 850 361 1160 395
rect 1218 361 1528 395
rect 1562 361 1872 395
rect 506 355 1160 361
rect 506 343 516 355
rect 1150 351 1160 355
rect 1218 355 1872 361
rect 1218 351 1228 355
rect 1862 343 1872 355
rect 1930 343 1940 401
rect 616 193 626 251
rect 684 239 694 251
rect 972 239 982 247
rect 684 193 982 239
rect 1040 239 1050 247
rect 1328 239 1338 244
rect 972 189 982 193
rect 1040 193 1338 239
rect 1396 239 1406 244
rect 1684 239 1694 246
rect 1040 189 1050 193
rect 1328 186 1338 193
rect 1396 193 1694 239
rect 1752 239 1762 246
rect 2040 239 2050 251
rect 1396 186 1406 193
rect 1684 188 1694 193
rect 1752 193 2050 239
rect 2108 193 2118 251
rect 1752 188 1762 193
rect 153 85 2028 119
rect 616 24 626 28
rect 495 23 626 24
rect 252 17 626 23
rect 684 23 694 28
rect 972 23 982 29
rect 684 17 982 23
rect 1040 23 1050 29
rect 1328 23 1338 31
rect 1040 17 1338 23
rect 1396 23 1406 31
rect 1684 23 1694 28
rect 1396 17 1694 23
rect 1752 23 1762 28
rect 2040 23 2050 29
rect 1752 17 2050 23
rect 2108 23 2118 29
rect 2108 17 2304 23
rect 252 -17 264 17
rect 2292 -17 2304 17
rect 252 -23 626 -17
rect 495 -30 626 -23
rect 684 -29 982 -17
rect 1040 -27 1338 -17
rect 1396 -27 1694 -17
rect 1040 -29 1694 -27
rect 684 -30 1694 -29
rect 1752 -29 2050 -17
rect 2108 -23 2304 -17
rect 2108 -29 2119 -23
rect 1752 -30 2119 -29
rect 495 -462 2119 -30
rect 2625 -462 2753 2441
rect 6710 2428 6720 2486
rect 6778 2428 6788 2486
rect 4277 2077 4311 2101
rect 3548 2043 4311 2077
rect 4369 2077 4403 2101
rect 4369 2043 4961 2077
rect 6720 2011 6778 2428
rect 3411 1941 3421 1999
rect 3479 1993 4106 1999
rect 4221 1997 4903 1999
rect 4221 1993 4845 1997
rect 3479 1959 3789 1993
rect 3823 1959 4106 1993
rect 4221 1959 4501 1993
rect 4535 1959 4845 1993
rect 3479 1953 4106 1959
rect 3479 1941 3489 1953
rect 4096 1903 4106 1953
rect 4221 1953 4845 1959
rect 4221 1903 4231 1953
rect 4835 1939 4845 1953
rect 4903 1939 4913 1997
rect 6293 1977 6945 2011
rect 7021 1977 7589 2011
rect 6293 1927 6327 1977
rect 7461 1927 7495 1977
rect 6271 1869 6281 1927
rect 6339 1869 6349 1927
rect 6563 1869 6573 1927
rect 6631 1869 6641 1927
rect 6855 1869 6865 1927
rect 6923 1869 6933 1927
rect 7147 1869 7157 1927
rect 7215 1869 7225 1927
rect 7439 1869 7449 1927
rect 7507 1869 7517 1927
rect 3589 1731 3599 1789
rect 3657 1777 3667 1789
rect 5013 1777 5023 1789
rect 3657 1771 5023 1777
rect 3657 1737 3967 1771
rect 4001 1737 4323 1771
rect 4357 1737 4679 1771
rect 4713 1737 5023 1771
rect 3657 1731 5023 1737
rect 5081 1731 5091 1789
rect 4919 1687 5001 1688
rect 3560 1672 5001 1687
rect 3560 1658 4280 1672
rect 3501 1653 4280 1658
rect 3501 1577 3577 1653
rect 4270 1577 4280 1653
rect 3501 1573 4280 1577
rect 3555 1555 4280 1573
rect 4398 1653 5001 1672
rect 4398 1577 4408 1653
rect 4919 1577 5001 1653
rect 4398 1555 5001 1577
rect 3555 1543 5001 1555
rect 4835 1499 4845 1504
rect 3411 1441 3421 1499
rect 3479 1493 4044 1499
rect 3479 1459 3789 1493
rect 3823 1459 4044 1493
rect 3479 1453 4044 1459
rect 3479 1441 3489 1453
rect 4034 1441 4044 1453
rect 4102 1493 4400 1499
rect 4102 1459 4145 1493
rect 4179 1459 4400 1493
rect 4102 1453 4400 1459
rect 4102 1441 4112 1453
rect 4390 1441 4400 1453
rect 4458 1493 4845 1499
rect 4458 1459 4501 1493
rect 4535 1459 4845 1493
rect 4458 1453 4845 1459
rect 4458 1441 4468 1453
rect 4835 1446 4845 1453
rect 4903 1446 4913 1504
rect 6382 1479 6416 1615
rect 6471 1426 6505 1682
rect 6674 1482 6708 1618
rect 6763 1422 6797 1678
rect 6966 1483 7000 1619
rect 7055 1417 7089 1673
rect 7259 1483 7293 1619
rect 7347 1428 7381 1684
rect 7550 1483 7584 1619
rect 7639 1420 7673 1676
rect 3589 1231 3599 1289
rect 3657 1277 3667 1289
rect 3767 1277 3777 1289
rect 3657 1231 3777 1277
rect 3835 1277 3845 1289
rect 4658 1277 4668 1290
rect 3835 1271 4668 1277
rect 4726 1277 4736 1290
rect 5013 1277 5023 1289
rect 3835 1237 3967 1271
rect 4001 1237 4323 1271
rect 4357 1237 4668 1271
rect 3835 1232 4668 1237
rect 4726 1232 5023 1277
rect 3835 1231 5023 1232
rect 5081 1231 5091 1289
rect 3498 1145 5005 1193
rect 4034 1017 4044 1035
rect 3546 983 4044 1017
rect 4034 977 4044 983
rect 4102 1017 4112 1035
rect 4390 1017 4400 1035
rect 4102 983 4400 1017
rect 4102 977 4112 983
rect 4390 977 4400 983
rect 4458 1017 4468 1035
rect 4458 983 4959 1017
rect 4458 977 4468 983
rect 3411 881 3421 939
rect 3479 893 3777 939
rect 3835 933 4667 939
rect 3835 899 4145 933
rect 4179 899 4501 933
rect 4535 899 4667 933
rect 3479 881 3489 893
rect 3767 881 3777 893
rect 3835 893 4667 899
rect 3835 881 3845 893
rect 4657 881 4667 893
rect 4725 893 4845 939
rect 4725 881 4735 893
rect 4835 881 4845 893
rect 4903 881 4913 939
rect 6293 922 6327 1178
rect 6383 983 6417 1119
rect 6585 923 6619 1179
rect 6674 985 6708 1121
rect 6877 922 6911 1178
rect 6966 983 7000 1119
rect 7169 923 7203 1179
rect 7258 985 7292 1121
rect 7461 921 7495 1177
rect 7550 983 7584 1119
rect 3589 671 3599 729
rect 3657 717 3667 729
rect 5013 717 5023 729
rect 3657 711 5023 717
rect 3657 677 3967 711
rect 4001 677 4323 711
rect 4357 677 4679 711
rect 4713 677 5023 711
rect 3657 671 5023 677
rect 5081 671 5091 729
rect 3565 601 4978 627
rect 3565 593 5001 601
rect 3501 517 3577 593
rect 4925 517 5001 593
rect 3501 516 5001 517
rect 3501 508 4970 516
rect 3557 483 4970 508
rect 6383 486 6417 622
rect 3411 381 3421 439
rect 3479 433 4845 439
rect 3479 399 3789 433
rect 3823 399 4145 433
rect 4179 399 4501 433
rect 4535 399 4845 433
rect 3479 393 4845 399
rect 3479 381 3489 393
rect 4835 381 4845 393
rect 4903 381 4913 439
rect 6471 422 6505 678
rect 6673 486 6707 622
rect 6763 422 6797 678
rect 6965 487 6999 623
rect 7055 433 7089 689
rect 7259 486 7293 622
rect 7347 423 7381 679
rect 7551 485 7585 621
rect 7639 427 7673 683
rect 3589 171 3599 229
rect 3657 217 3667 229
rect 5013 217 5023 229
rect 3657 211 5023 217
rect 3657 177 3967 211
rect 4001 177 4323 211
rect 4357 177 4679 211
rect 4713 177 5023 211
rect 3657 171 5023 177
rect 5081 171 5091 229
rect 6271 177 6281 235
rect 6339 177 6349 235
rect 6563 177 6573 235
rect 6631 177 6641 235
rect 6855 177 6865 235
rect 6923 177 6933 235
rect 7147 177 7157 235
rect 7215 177 7225 235
rect 7439 177 7449 235
rect 7507 177 7517 235
rect 4212 127 4222 128
rect 3547 93 4222 127
rect 4212 70 4222 93
rect 4280 127 4290 128
rect 4280 93 4960 127
rect 6425 93 7576 127
rect 4280 70 4290 93
rect 4989 0 5106 6
rect 3567 -11 3684 -5
rect 3567 -98 3579 -11
rect 3672 -98 3684 -11
rect 4989 -87 5001 0
rect 5094 -87 5106 0
rect 4989 -93 5106 -87
rect 6247 3 6374 9
rect 3567 -104 3684 -98
rect 6247 -94 6259 3
rect 6362 -94 6374 3
rect 6247 -100 6374 -94
rect 7417 2 7544 8
rect 7417 -95 7429 2
rect 7532 -95 7544 2
rect 7417 -101 7544 -95
rect 4212 -231 8604 -201
rect 4212 -289 4222 -231
rect 4280 -289 8604 -231
rect 4212 -318 8604 -289
rect -430 -463 8656 -462
rect -430 -590 -378 -463
rect -384 -591 -378 -590
rect -250 -482 8656 -463
rect -250 -484 7430 -482
rect -250 -489 5006 -484
rect -250 -541 3579 -489
rect -250 -590 3275 -541
rect 3672 -541 5006 -489
rect 5099 -488 7430 -484
rect 5099 -541 6269 -488
rect 6362 -541 7430 -488
rect 7523 -541 8656 -482
rect 8165 -590 8656 -541
rect -250 -591 -244 -590
rect 3263 -596 8177 -590
<< via1 >>
rect 1253 5997 1311 6055
rect 1609 5997 1667 6055
rect 1965 5997 2023 6055
rect 2321 5997 2379 6055
rect 3453 5997 3511 6055
rect 3809 5997 3867 6055
rect 4165 5997 4223 6055
rect 4520 5997 4578 6055
rect 5653 5997 5711 6055
rect 6009 5997 6067 6055
rect 6365 5997 6423 6055
rect 6721 5997 6779 6055
rect 1431 5799 1489 5857
rect 1787 5799 1845 5857
rect 2143 5799 2201 5857
rect 3631 5799 3689 5857
rect 3987 5798 4045 5856
rect 4343 5799 4401 5857
rect 5831 5799 5889 5857
rect 6187 5799 6245 5857
rect 6543 5799 6601 5857
rect 1342 5688 1400 5746
rect 1179 5230 1310 5288
rect 1608 5230 1666 5288
rect 1964 5230 2022 5288
rect 2319 5230 2377 5288
rect 3452 5230 3510 5288
rect 3808 5230 3866 5288
rect 4164 5230 4222 5288
rect 4520 5230 4578 5288
rect 5652 5230 5710 5288
rect 6008 5230 6066 5288
rect 6364 5230 6422 5288
rect 6720 5230 6778 5288
rect 1430 5032 1488 5090
rect 1786 5032 1844 5090
rect 2141 5032 2199 5090
rect 3630 5032 3688 5090
rect 3986 5032 4044 5090
rect 4341 5032 4399 5090
rect 5831 5032 5889 5090
rect 6186 5032 6244 5090
rect 6542 5032 6600 5090
rect 2230 4921 2288 4979
rect -84 4427 -26 4495
rect -84 4393 -72 4427
rect -72 4393 -38 4427
rect -38 4393 -26 4427
rect 451 4415 509 4504
rect -84 4375 -26 4393
rect 1164 4390 1310 4530
rect 1874 4410 1932 4499
rect 2408 4427 2466 4495
rect 2408 4393 2420 4427
rect 2420 4393 2454 4427
rect 2454 4393 2466 4427
rect 2408 4375 2466 4393
rect 94 4205 152 4223
rect 804 4205 862 4224
rect 1518 4205 1576 4220
rect 2230 4205 2288 4223
rect 94 4171 106 4205
rect 106 4171 140 4205
rect 140 4171 152 4205
rect 804 4171 818 4205
rect 818 4171 852 4205
rect 852 4171 862 4205
rect 1518 4171 1530 4205
rect 1530 4171 1564 4205
rect 1564 4171 1576 4205
rect 2230 4171 2242 4205
rect 2242 4171 2276 4205
rect 2276 4171 2288 4205
rect 94 4165 152 4171
rect 804 4166 862 4171
rect 1518 4162 1576 4171
rect 2230 4165 2288 4171
rect -84 3929 -26 4105
rect -84 3895 -72 3929
rect -72 3895 -38 3929
rect -38 3895 -26 3929
rect 450 3904 508 4112
rect 1163 3911 1221 4119
rect 1873 3900 1931 4108
rect 2407 3935 2465 4114
rect 2407 3929 2466 3935
rect 2407 3906 2420 3929
rect 2408 3895 2420 3906
rect 2420 3895 2454 3929
rect 2454 3895 2466 3929
rect -84 3877 -26 3895
rect 2408 3877 2466 3895
rect 94 3707 152 3725
rect 805 3707 863 3723
rect 1518 3707 1576 3720
rect 2230 3707 2288 3725
rect 94 3673 106 3707
rect 106 3673 140 3707
rect 140 3673 152 3707
rect 805 3673 818 3707
rect 818 3673 852 3707
rect 852 3673 863 3707
rect 1518 3673 1530 3707
rect 1530 3673 1564 3707
rect 1564 3673 1576 3707
rect 2230 3673 2242 3707
rect 2242 3673 2276 3707
rect 2276 3673 2288 3707
rect 94 3667 152 3673
rect 805 3665 863 3673
rect 1518 3662 1576 3673
rect 2230 3667 2288 3673
rect -83 3437 -25 3607
rect -84 3431 -25 3437
rect -84 3397 -72 3431
rect -72 3397 -38 3431
rect -38 3399 -25 3431
rect -38 3397 -26 3399
rect 450 3411 508 3619
rect 1161 3404 1219 3612
rect 1874 3404 1932 3612
rect 2408 3431 2466 3613
rect 2408 3397 2420 3431
rect 2420 3397 2454 3431
rect 2454 3397 2466 3431
rect -84 3379 -26 3397
rect 2408 3379 2466 3397
rect 94 3209 152 3227
rect 809 3209 867 3230
rect 1518 3209 1576 3226
rect 2230 3209 2288 3227
rect 94 3175 106 3209
rect 106 3175 140 3209
rect 140 3175 152 3209
rect 809 3175 818 3209
rect 818 3175 852 3209
rect 852 3175 867 3209
rect 1518 3175 1530 3209
rect 1530 3175 1564 3209
rect 1564 3175 1576 3209
rect 2230 3175 2242 3209
rect 2242 3175 2276 3209
rect 2276 3175 2288 3209
rect 94 3169 152 3175
rect 809 3172 867 3175
rect 1518 3168 1576 3175
rect 2230 3169 2288 3175
rect -84 2933 -26 3125
rect -84 2899 -72 2933
rect -72 2899 -38 2933
rect -38 2899 -26 2933
rect 450 2902 508 3110
rect 1163 2904 1221 3112
rect 1875 2907 1933 3115
rect 2408 2933 2466 3125
rect 2408 2899 2420 2933
rect 2420 2899 2454 2933
rect 2454 2899 2466 2933
rect -84 2881 -26 2899
rect 2408 2881 2466 2899
rect 94 2711 152 2729
rect 94 2677 106 2711
rect 106 2677 140 2711
rect 140 2677 152 2711
rect 94 2671 152 2677
rect 448 2711 506 2727
rect 448 2677 462 2711
rect 462 2677 496 2711
rect 496 2677 506 2711
rect 448 2669 506 2677
rect 804 2711 862 2726
rect 804 2677 818 2711
rect 818 2677 852 2711
rect 852 2677 862 2711
rect 804 2668 862 2677
rect 1160 2711 1218 2729
rect 1160 2677 1174 2711
rect 1174 2677 1208 2711
rect 1208 2677 1218 2711
rect 1160 2671 1218 2677
rect 1517 2711 1575 2728
rect 1517 2677 1530 2711
rect 1530 2677 1564 2711
rect 1564 2677 1575 2711
rect 1517 2670 1575 2677
rect 1873 2711 1931 2728
rect 1873 2677 1886 2711
rect 1886 2677 1920 2711
rect 1920 2677 1931 2711
rect 1873 2670 1931 2677
rect 2230 2711 2288 2729
rect 2230 2677 2242 2711
rect 2242 2677 2276 2711
rect 2276 2677 2288 2711
rect 2230 2671 2288 2677
rect -378 2441 -250 2569
rect 3393 4436 3510 4446
rect 5553 4436 5611 4442
rect 7689 4436 7747 4442
rect 3393 4402 3429 4436
rect 3429 4402 3463 4436
rect 3463 4402 3510 4436
rect 5553 4402 5565 4436
rect 5565 4402 5599 4436
rect 5599 4402 5611 4436
rect 7689 4402 7701 4436
rect 7701 4402 7735 4436
rect 7735 4402 7747 4436
rect 3393 4329 3510 4402
rect 5553 4384 5611 4402
rect 7689 4384 7747 4402
rect 3595 4214 3653 4232
rect 5731 4214 5789 4232
rect 7867 4214 7925 4232
rect 3595 4180 3607 4214
rect 3607 4180 3641 4214
rect 3641 4180 3653 4214
rect 5731 4180 5743 4214
rect 5743 4180 5777 4214
rect 5777 4180 5789 4214
rect 7867 4180 7879 4214
rect 7879 4180 7913 4214
rect 7913 4180 7925 4214
rect 3595 4174 3653 4180
rect 5731 4174 5789 4180
rect 7867 4174 7925 4180
rect 3392 3936 3509 3942
rect 5553 3936 5611 3942
rect 7689 3936 7747 3942
rect 3392 3902 3429 3936
rect 3429 3902 3463 3936
rect 3463 3902 3509 3936
rect 5553 3902 5565 3936
rect 5565 3902 5599 3936
rect 5599 3902 5611 3936
rect 7689 3902 7701 3936
rect 7701 3902 7735 3936
rect 7735 3902 7747 3936
rect 3392 3825 3509 3902
rect 5553 3884 5611 3902
rect 7689 3884 7747 3902
rect 3595 3714 3653 3732
rect 3595 3680 3607 3714
rect 3607 3680 3641 3714
rect 3641 3680 3653 3714
rect 3595 3674 3653 3680
rect 3889 3714 4011 3776
rect 5731 3714 5789 3732
rect 7867 3714 7925 3732
rect 3889 3680 3963 3714
rect 3963 3680 3997 3714
rect 3997 3680 4011 3714
rect 5731 3680 5743 3714
rect 5743 3680 5777 3714
rect 5777 3680 5789 3714
rect 7867 3680 7879 3714
rect 7879 3680 7913 3714
rect 7913 3680 7925 3714
rect 3889 3675 4011 3680
rect 3953 3674 4011 3675
rect 5731 3674 5789 3680
rect 7867 3674 7925 3680
rect 4131 3572 4189 3630
rect 3889 3396 4011 3514
rect 4131 2982 4189 3040
rect 3889 2938 4010 2939
rect 3889 2932 4011 2938
rect 3889 2836 3965 2932
rect 3965 2836 3999 2932
rect 3999 2880 4011 2932
rect 3999 2836 4010 2880
rect 3889 2822 4010 2836
rect 4131 2793 4189 2805
rect 4131 2676 4143 2793
rect 4143 2676 4177 2793
rect 4177 2676 4189 2793
rect 4131 2668 4189 2676
rect 4309 2676 4321 2919
rect 4321 2676 4355 2919
rect 4355 2676 4367 2919
rect 4309 2667 4367 2676
rect 448 1919 506 1925
rect 448 1885 460 1919
rect 460 1885 494 1919
rect 494 1885 506 1919
rect 448 1867 506 1885
rect 804 1919 862 1928
rect 804 1885 816 1919
rect 816 1885 850 1919
rect 850 1885 862 1919
rect 804 1870 862 1885
rect 1160 1919 1218 1925
rect 1160 1885 1172 1919
rect 1172 1885 1206 1919
rect 1206 1885 1218 1919
rect 1160 1867 1218 1885
rect 1517 1919 1575 1926
rect 1517 1885 1528 1919
rect 1528 1885 1562 1919
rect 1562 1885 1575 1919
rect 1517 1868 1575 1885
rect 1872 1919 1930 1925
rect 1872 1885 1884 1919
rect 1884 1885 1918 1919
rect 1918 1885 1930 1919
rect 1872 1867 1930 1885
rect 626 1697 684 1715
rect 1338 1697 1396 1710
rect 2050 1697 2108 1715
rect 626 1663 638 1697
rect 638 1663 672 1697
rect 672 1663 684 1697
rect 1338 1663 1350 1697
rect 1350 1663 1384 1697
rect 1384 1663 1396 1697
rect 2050 1663 2062 1697
rect 2062 1663 2096 1697
rect 2096 1663 2108 1697
rect 626 1657 684 1663
rect 1338 1652 1396 1663
rect 2050 1657 2108 1663
rect 448 1421 506 1427
rect 448 1387 460 1421
rect 460 1387 494 1421
rect 494 1387 506 1421
rect 448 1369 506 1387
rect 804 1421 862 1427
rect 804 1387 816 1421
rect 816 1387 850 1421
rect 850 1387 862 1421
rect 804 1369 862 1387
rect 1159 1421 1217 1430
rect 1159 1387 1172 1421
rect 1172 1387 1206 1421
rect 1206 1387 1217 1421
rect 1159 1372 1217 1387
rect 1517 1421 1575 1429
rect 1517 1387 1528 1421
rect 1528 1387 1562 1421
rect 1562 1387 1575 1421
rect 1517 1371 1575 1387
rect 1872 1421 1930 1427
rect 1872 1387 1884 1421
rect 1884 1387 1918 1421
rect 1918 1387 1930 1421
rect 1872 1369 1930 1387
rect 626 1199 684 1218
rect 1338 1199 1396 1216
rect 2050 1199 2108 1216
rect 626 1165 638 1199
rect 638 1165 672 1199
rect 672 1165 684 1199
rect 1338 1165 1350 1199
rect 1350 1165 1384 1199
rect 1384 1165 1396 1199
rect 2050 1165 2062 1199
rect 2062 1165 2096 1199
rect 2096 1165 2108 1199
rect 626 1160 684 1165
rect 1338 1158 1396 1165
rect 2050 1158 2108 1165
rect 448 893 506 899
rect 1160 893 1218 907
rect 1872 893 1930 899
rect 448 859 460 893
rect 460 859 494 893
rect 494 859 506 893
rect 1160 859 1172 893
rect 1172 859 1206 893
rect 1206 859 1218 893
rect 1872 859 1884 893
rect 1884 859 1918 893
rect 1918 859 1930 893
rect 448 841 506 859
rect 1160 849 1218 859
rect 1872 841 1930 859
rect 626 731 684 749
rect 1339 731 1397 748
rect 2050 731 2108 748
rect 626 697 638 731
rect 638 697 672 731
rect 672 697 684 731
rect 1339 697 1350 731
rect 1350 697 1384 731
rect 1384 697 1397 731
rect 2050 697 2062 731
rect 2062 697 2096 731
rect 2096 697 2108 731
rect 626 691 684 697
rect 1339 690 1397 697
rect 2050 690 2108 697
rect 448 395 506 401
rect 1160 395 1218 409
rect 1872 395 1930 401
rect 448 361 460 395
rect 460 361 494 395
rect 494 361 506 395
rect 1160 361 1172 395
rect 1172 361 1206 395
rect 1206 361 1218 395
rect 1872 361 1884 395
rect 1884 361 1918 395
rect 1918 361 1930 395
rect 448 343 506 361
rect 1160 351 1218 361
rect 1872 343 1930 361
rect 626 233 684 251
rect 626 199 638 233
rect 638 199 672 233
rect 672 199 684 233
rect 626 193 684 199
rect 982 233 1040 247
rect 982 199 994 233
rect 994 199 1028 233
rect 1028 199 1040 233
rect 982 189 1040 199
rect 1338 233 1396 244
rect 1338 199 1350 233
rect 1350 199 1384 233
rect 1384 199 1396 233
rect 1338 186 1396 199
rect 1694 233 1752 246
rect 1694 199 1706 233
rect 1706 199 1740 233
rect 1740 199 1752 233
rect 1694 188 1752 199
rect 2050 233 2108 251
rect 2050 199 2062 233
rect 2062 199 2096 233
rect 2096 199 2108 233
rect 2050 193 2108 199
rect 626 17 684 28
rect 982 17 1040 29
rect 1338 17 1396 31
rect 1694 17 1752 28
rect 2050 17 2108 29
rect 626 -17 684 17
rect 982 -17 1040 17
rect 1338 -17 1396 17
rect 1694 -17 1752 17
rect 2050 -17 2108 17
rect 626 -30 684 -17
rect 982 -29 1040 -17
rect 1338 -27 1396 -17
rect 1694 -30 1752 -17
rect 2050 -29 2108 -17
rect 6720 2428 6778 2486
rect 4311 2043 4369 2101
rect 3421 1993 3479 1999
rect 4106 1993 4221 1999
rect 4845 1993 4903 1997
rect 3421 1959 3433 1993
rect 3433 1959 3467 1993
rect 3467 1959 3479 1993
rect 4106 1959 4145 1993
rect 4145 1959 4179 1993
rect 4179 1959 4221 1993
rect 4845 1959 4857 1993
rect 4857 1959 4891 1993
rect 4891 1959 4903 1993
rect 3421 1941 3479 1959
rect 4106 1903 4221 1959
rect 4845 1939 4903 1959
rect 6281 1869 6339 1927
rect 6573 1869 6631 1927
rect 6865 1869 6923 1927
rect 7157 1869 7215 1927
rect 7449 1869 7507 1927
rect 3599 1771 3657 1789
rect 5023 1771 5081 1789
rect 3599 1737 3611 1771
rect 3611 1737 3645 1771
rect 3645 1737 3657 1771
rect 5023 1737 5035 1771
rect 5035 1737 5069 1771
rect 5069 1737 5081 1771
rect 3599 1731 3657 1737
rect 5023 1731 5081 1737
rect 4280 1555 4398 1672
rect 3421 1493 3479 1499
rect 3421 1459 3433 1493
rect 3433 1459 3467 1493
rect 3467 1459 3479 1493
rect 3421 1441 3479 1459
rect 4044 1441 4102 1499
rect 4400 1441 4458 1499
rect 4845 1493 4903 1504
rect 4845 1459 4857 1493
rect 4857 1459 4891 1493
rect 4891 1459 4903 1493
rect 4845 1446 4903 1459
rect 3599 1271 3657 1289
rect 3599 1237 3611 1271
rect 3611 1237 3645 1271
rect 3645 1237 3657 1271
rect 3599 1231 3657 1237
rect 3777 1231 3835 1289
rect 4668 1271 4726 1290
rect 4668 1237 4679 1271
rect 4679 1237 4713 1271
rect 4713 1237 4726 1271
rect 4668 1232 4726 1237
rect 5023 1271 5081 1289
rect 5023 1237 5035 1271
rect 5035 1237 5069 1271
rect 5069 1237 5081 1271
rect 5023 1231 5081 1237
rect 4044 977 4102 1035
rect 4400 977 4458 1035
rect 3421 933 3479 939
rect 3421 899 3433 933
rect 3433 899 3467 933
rect 3467 899 3479 933
rect 3421 881 3479 899
rect 3777 933 3835 939
rect 3777 899 3789 933
rect 3789 899 3823 933
rect 3823 899 3835 933
rect 3777 881 3835 899
rect 4667 881 4725 939
rect 4845 933 4903 939
rect 4845 899 4857 933
rect 4857 899 4891 933
rect 4891 899 4903 933
rect 4845 881 4903 899
rect 3599 711 3657 729
rect 5023 711 5081 729
rect 3599 677 3611 711
rect 3611 677 3645 711
rect 3645 677 3657 711
rect 5023 677 5035 711
rect 5035 677 5069 711
rect 5069 677 5081 711
rect 3599 671 3657 677
rect 5023 671 5081 677
rect 3421 433 3479 439
rect 4845 433 4903 439
rect 3421 399 3433 433
rect 3433 399 3467 433
rect 3467 399 3479 433
rect 4845 399 4857 433
rect 4857 399 4891 433
rect 4891 399 4903 433
rect 3421 381 3479 399
rect 4845 381 4903 399
rect 3599 211 3657 229
rect 5023 211 5081 229
rect 3599 177 3611 211
rect 3611 177 3645 211
rect 3645 177 3657 211
rect 5023 177 5035 211
rect 5035 177 5069 211
rect 5069 177 5081 211
rect 3599 171 3657 177
rect 5023 171 5081 177
rect 6281 177 6339 235
rect 6573 177 6631 235
rect 6865 177 6923 235
rect 7157 177 7215 235
rect 7449 177 7507 235
rect 4222 70 4280 128
rect 3579 -98 3672 -11
rect 5001 -87 5094 0
rect 6259 -94 6362 3
rect 7429 -95 7532 2
rect 4222 -289 4280 -231
rect -378 -591 -250 -463
rect 3579 -576 3672 -489
rect 5006 -571 5099 -484
rect 6269 -575 6362 -488
rect 7430 -569 7523 -482
<< metal2 >>
rect 1253 6055 1311 6065
rect 1609 6055 1667 6065
rect 1965 6055 2023 6065
rect 2321 6055 2379 6065
rect 3453 6055 3511 6065
rect 3809 6055 3867 6065
rect 4165 6055 4223 6065
rect 4520 6055 4578 6065
rect 5653 6055 5711 6065
rect 6009 6055 6067 6065
rect 6365 6055 6423 6065
rect 6721 6055 6779 6065
rect 1311 5997 1609 6055
rect 1667 5997 1965 6055
rect 2023 5997 2321 6055
rect 2379 5997 2567 6055
rect 1253 5957 2567 5997
rect 3452 5997 3453 6055
rect 3511 5997 3809 6055
rect 3867 5997 4165 6055
rect 4223 5997 4520 6055
rect 4578 5997 4748 6055
rect 3452 5957 4748 5997
rect 1431 5857 1489 5867
rect 1787 5857 1845 5867
rect 2143 5857 2201 5867
rect 1489 5799 1787 5857
rect 1845 5799 2143 5857
rect 1431 5789 1489 5799
rect 1787 5789 1845 5799
rect 2143 5789 2201 5799
rect 1342 5746 1400 5756
rect 1179 5288 1310 5298
rect 1342 5288 1400 5688
rect 1608 5288 1666 5298
rect 1964 5288 2022 5298
rect 2319 5288 2377 5298
rect 1310 5230 1608 5288
rect 1666 5230 1964 5288
rect 2022 5230 2319 5288
rect 1179 4540 1310 5230
rect 1608 5220 1666 5230
rect 1964 5220 2022 5230
rect 2319 5220 2377 5230
rect 2441 5120 2567 5957
rect 3631 5857 3689 5867
rect 3987 5857 4045 5866
rect 4343 5857 4401 5867
rect 3689 5856 4343 5857
rect 3689 5799 3987 5856
rect 3631 5789 3689 5799
rect 4045 5799 4343 5856
rect 3987 5788 4045 5798
rect 4343 5789 4401 5799
rect 1430 5090 2567 5120
rect 1488 5032 1786 5090
rect 1844 5032 2141 5090
rect 2199 5032 2567 5090
rect 1430 5022 2567 5032
rect 3393 5298 4577 5319
rect 3393 5288 4578 5298
rect 3393 5230 3452 5288
rect 3510 5230 3808 5288
rect 3866 5230 4164 5288
rect 4222 5230 4520 5288
rect 3393 5221 4578 5230
rect 1164 4530 1310 4540
rect -84 4495 -26 4505
rect 451 4504 509 4514
rect -84 4105 -26 4375
rect 450 4415 451 4498
rect 450 4405 509 4415
rect -84 3617 -26 3877
rect 94 4223 152 4233
rect 94 3725 152 4165
rect -84 3607 -25 3617
rect -84 3437 -83 3607
rect -26 3389 -25 3399
rect -84 3125 -26 3379
rect -84 2871 -26 2881
rect 94 3227 152 3667
rect 94 2729 152 3169
rect 450 4112 508 4405
rect 1163 4390 1164 4502
rect 2230 4979 2288 4989
rect 1163 4380 1310 4390
rect 1874 4499 1932 4509
rect 450 3619 508 3904
rect 450 3110 508 3411
rect 450 2892 508 2902
rect 804 4224 862 4234
rect 804 3733 862 4166
rect 1163 4119 1221 4380
rect 804 3723 863 3733
rect 804 3665 805 3723
rect 804 3655 863 3665
rect 804 3240 862 3655
rect 1163 3622 1221 3911
rect 1161 3612 1221 3622
rect 1219 3404 1221 3612
rect 1161 3394 1221 3404
rect 804 3230 867 3240
rect 804 3172 809 3230
rect 804 3162 867 3172
rect 94 2661 152 2671
rect 448 2727 506 2737
rect -390 2569 -239 2581
rect -390 2441 -378 2569
rect -250 2441 -239 2569
rect -390 2431 -239 2441
rect -378 -463 -250 2431
rect 448 1925 506 2669
rect 448 1427 506 1867
rect 804 2726 862 3162
rect 1163 3112 1221 3394
rect 1163 2894 1221 2904
rect 1517 4230 1575 4232
rect 1517 4220 1576 4230
rect 1517 4162 1518 4220
rect 1517 4152 1576 4162
rect 1517 3730 1575 4152
rect 1874 4118 1932 4410
rect 1873 4108 1932 4118
rect 1931 3900 1932 4108
rect 1873 3890 1932 3900
rect 1517 3720 1576 3730
rect 1517 3662 1518 3720
rect 1517 3652 1576 3662
rect 1517 3236 1575 3652
rect 1874 3612 1932 3890
rect 1517 3226 1576 3236
rect 1517 3168 1518 3226
rect 1517 3158 1576 3168
rect 804 1928 862 2668
rect 448 1359 506 1369
rect 626 1715 684 1725
rect 626 1218 684 1657
rect 804 1427 862 1870
rect 1160 2729 1218 2739
rect 1160 1925 1218 2671
rect 1160 1440 1218 1867
rect 1517 2728 1575 3158
rect 1874 3125 1932 3404
rect 2230 4223 2288 4921
rect 2230 3725 2288 4165
rect 2408 4495 2466 4505
rect 2408 4124 2466 4375
rect 2407 4114 2466 4124
rect 2465 3935 2466 4114
rect 3393 4446 3510 5221
rect 3808 5220 3866 5221
rect 4164 5220 4222 5221
rect 4520 5220 4578 5221
rect 4641 5127 4748 5957
rect 3619 5090 4748 5127
rect 3619 5032 3630 5090
rect 3688 5032 3986 5090
rect 4044 5032 4341 5090
rect 4399 5032 4748 5090
rect 5532 5997 5653 6055
rect 5711 5997 6009 6055
rect 6067 5997 6365 6055
rect 6423 5997 6721 6055
rect 5532 5090 5590 5997
rect 5653 5987 5711 5997
rect 6009 5987 6067 5997
rect 6365 5987 6423 5997
rect 6721 5987 6779 5997
rect 5831 5857 5889 5867
rect 6187 5857 6245 5867
rect 6543 5857 6601 5867
rect 5889 5799 6187 5857
rect 6245 5799 6543 5857
rect 5831 5789 5889 5799
rect 6187 5789 6245 5799
rect 6543 5789 6601 5799
rect 5652 5288 5710 5298
rect 6008 5288 6066 5298
rect 6364 5288 6422 5298
rect 6720 5288 6778 5298
rect 5710 5230 6008 5288
rect 6066 5230 6364 5288
rect 6422 5230 6720 5288
rect 5652 5220 5710 5230
rect 6008 5220 6066 5230
rect 6364 5220 6422 5230
rect 5831 5090 5889 5100
rect 6186 5090 6244 5100
rect 6542 5090 6600 5100
rect 5532 5032 5831 5090
rect 5889 5032 6186 5090
rect 6244 5032 6542 5090
rect 3619 5029 4748 5032
rect 3630 5022 3688 5029
rect 3986 5022 4044 5029
rect 4341 5022 4399 5029
rect 5831 5022 5889 5032
rect 6186 5022 6244 5032
rect 6542 5022 6600 5032
rect 6720 4839 6778 5230
rect 6720 4771 6778 4781
rect 3393 3952 3510 4329
rect 5553 4442 5611 4452
rect 2407 3896 2408 3906
rect 2230 3227 2288 3667
rect 1874 3115 1933 3125
rect 1874 3069 1875 3115
rect 1875 2897 1933 2907
rect 1873 2728 1931 2738
rect 1517 1926 1575 2670
rect 804 1359 862 1369
rect 1159 1430 1218 1440
rect 1217 1372 1218 1430
rect 1159 1362 1218 1372
rect 1338 1710 1396 1720
rect 448 899 506 909
rect 448 401 506 841
rect 448 333 506 343
rect 626 749 684 1160
rect 1338 1216 1396 1652
rect 1517 1429 1575 1868
rect 1517 1361 1575 1371
rect 1872 2670 1873 2724
rect 1872 2660 1931 2670
rect 2230 2729 2288 3169
rect 2408 3613 2466 3877
rect 3392 3942 3510 3952
rect 3509 3833 3510 3942
rect 3595 4232 3653 4242
rect 3392 3815 3509 3825
rect 3595 3732 3653 4174
rect 5553 3942 5611 4384
rect 7689 4442 7747 4452
rect 5553 3874 5611 3884
rect 5731 4232 5789 4242
rect 3595 3664 3653 3674
rect 3889 3776 4011 3786
rect 3889 3674 3953 3675
rect 2408 3125 2466 3379
rect 2408 2871 2466 2881
rect 3889 3514 4011 3674
rect 5731 3732 5789 4174
rect 7689 3942 7747 4384
rect 7689 3874 7747 3884
rect 7867 4232 7925 4242
rect 5731 3664 5789 3674
rect 7867 3732 7925 4174
rect 7867 3664 7925 3674
rect 3889 2939 4011 3396
rect 4131 3630 4189 3640
rect 4131 3040 4189 3572
rect 4131 2972 4189 2982
rect 4010 2938 4011 2939
rect 4010 2870 4011 2880
rect 4309 2919 4367 2929
rect 3889 2812 4010 2822
rect 2230 2661 2288 2671
rect 4106 2805 4208 2815
rect 4106 2668 4131 2805
rect 4189 2668 4208 2805
rect 1872 1925 1930 2660
rect 4106 2009 4208 2668
rect 4367 2667 4369 2723
rect 4309 2657 4369 2667
rect 4311 2101 4369 2657
rect 6720 2486 6778 2496
rect 6720 2418 6778 2428
rect 1872 1427 1930 1867
rect 3421 1999 3479 2009
rect 1872 1359 1930 1369
rect 2050 1715 2108 1725
rect 626 251 684 691
rect 1160 907 1218 917
rect 1160 409 1218 849
rect 1160 341 1218 351
rect 1338 758 1396 1158
rect 2050 1216 2108 1657
rect 3421 1499 3479 1941
rect 4106 1999 4221 2009
rect 4106 1893 4221 1903
rect 3421 1431 3479 1441
rect 3599 1789 3657 1799
rect 3599 1289 3657 1731
rect 4311 1682 4369 2043
rect 4845 1997 4903 2007
rect 4280 1672 4398 1682
rect 4280 1545 4398 1555
rect 4044 1499 4102 1509
rect 3599 1221 3657 1231
rect 3777 1289 3835 1299
rect 1872 899 1930 909
rect 1338 748 1397 758
rect 1338 690 1339 748
rect 1338 680 1397 690
rect 626 28 684 193
rect 626 -40 684 -30
rect 982 247 1040 257
rect 982 29 1040 189
rect 982 -39 1040 -29
rect 1338 244 1396 680
rect 1872 401 1930 841
rect 1872 333 1930 343
rect 2050 748 2108 1158
rect 1338 31 1396 186
rect 1338 -37 1396 -27
rect 1694 246 1752 256
rect 1694 28 1752 188
rect 1694 -40 1752 -30
rect 2050 251 2108 690
rect 3421 939 3479 949
rect 3421 439 3479 881
rect 3777 939 3835 1231
rect 4044 1035 4102 1441
rect 4044 967 4102 977
rect 4400 1499 4458 1509
rect 4400 1035 4458 1441
rect 4845 1504 4903 1939
rect 6281 1927 6339 1937
rect 6573 1927 6631 1937
rect 6865 1927 6923 1937
rect 7157 1927 7215 1937
rect 7449 1927 7507 1937
rect 6339 1869 6573 1927
rect 6631 1869 6865 1927
rect 6923 1869 7157 1927
rect 7215 1869 7449 1927
rect 6281 1859 6339 1869
rect 6573 1859 6631 1869
rect 6865 1859 6923 1869
rect 7157 1859 7215 1869
rect 7449 1859 7507 1869
rect 4845 1436 4903 1446
rect 5023 1789 5081 1799
rect 4668 1290 4726 1300
rect 4400 967 4458 977
rect 4667 1232 4668 1269
rect 4667 1222 4726 1232
rect 5023 1289 5081 1731
rect 3777 871 3835 881
rect 4667 939 4725 1222
rect 5023 1221 5081 1231
rect 4667 871 4725 881
rect 4845 939 4903 949
rect 3421 371 3479 381
rect 3599 729 3657 739
rect 2050 29 2108 193
rect 3599 229 3657 671
rect 4845 439 4903 881
rect 4845 371 4903 381
rect 5023 729 5081 739
rect 3599 -1 3657 171
rect 5023 229 5081 671
rect 4222 128 4280 138
rect 2050 -39 2108 -29
rect 3579 -11 3672 -1
rect 3579 -108 3672 -98
rect 3599 -479 3657 -108
rect 4222 -231 4280 70
rect 5023 10 5081 171
rect 6281 235 6339 245
rect 6573 235 6631 245
rect 6865 235 6923 245
rect 7157 235 7215 245
rect 7449 235 7507 245
rect 6339 177 6573 235
rect 6631 177 6865 235
rect 6923 177 7157 235
rect 7215 177 7449 235
rect 7507 177 7508 190
rect 6281 13 6339 177
rect 6573 167 6631 177
rect 6865 167 6923 177
rect 7157 167 7215 177
rect 7449 167 7508 177
rect 5001 0 5094 10
rect 5001 -97 5094 -87
rect 6259 3 6362 13
rect 7450 12 7508 167
rect 4222 -299 4280 -289
rect 5023 -474 5081 -97
rect 6259 -104 6362 -94
rect 7429 2 7532 12
rect 3579 -489 3672 -479
rect 3579 -586 3672 -576
rect 5006 -484 5099 -474
rect 6281 -478 6339 -104
rect 7429 -105 7532 -95
rect 7450 -472 7508 -105
rect 5006 -581 5099 -571
rect 6269 -488 6362 -478
rect 6269 -585 6362 -575
rect 7430 -482 7523 -472
rect 7430 -579 7523 -569
rect -378 -597 -250 -591
<< via2 >>
rect 6720 4781 6778 4839
rect 6720 2428 6778 2486
<< metal3 >>
rect 6710 4839 6788 4844
rect 6710 4781 6720 4839
rect 6778 4781 6788 4839
rect 6710 2486 6788 4781
rect 6710 2428 6720 2486
rect 6778 2428 6788 2486
rect 6710 2419 6788 2428
use sky130_fd_pr__nfet_01v8_6RUDQZ  sky130_fd_pr__nfet_01v8_6RUDQZ_0
timestamp 1654656593
transform 1 0 4251 0 1 305
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_6RUDQZ  sky130_fd_pr__nfet_01v8_6RUDQZ_1
timestamp 1654656593
transform 1 0 4251 0 1 805
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_6RUDQZ  sky130_fd_pr__nfet_01v8_6RUDQZ_2
timestamp 1654656593
transform 1 0 4251 0 1 1365
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_6RUDQZ  sky130_fd_pr__nfet_01v8_6RUDQZ_3
timestamp 1654656593
transform 1 0 4251 0 1 1865
box -1008 -228 1008 228
use sky130_fd_pr__nfet_01v8_EL6FQZ  sky130_fd_pr__nfet_01v8_EL6FQZ_0
timestamp 1654656593
transform 1 0 5671 0 1 3808
box -2432 -228 2432 228
use sky130_fd_pr__nfet_01v8_EL6FQZ  sky130_fd_pr__nfet_01v8_EL6FQZ_1
timestamp 1654656593
transform 1 0 5671 0 1 4308
box -2432 -228 2432 228
use sky130_fd_pr__nfet_01v8_EZNTQN  sky130_fd_pr__nfet_01v8_EZNTQN_0
timestamp 1654656593
transform 1 0 1278 0 1 1044
box -1146 -1097 1146 1097
use sky130_fd_pr__nfet_01v8_LJREPQ  sky130_fd_pr__nfet_01v8_LJREPQ_0
timestamp 1654656593
transform 1 0 4160 0 1 2804
box -385 -228 385 228
use sky130_fd_pr__nfet_01v8_SD55Q9  sky130_fd_pr__nfet_01v8_SD55Q9_0
timestamp 1654656593
transform 1 0 6983 0 1 1052
box -994 -975 994 975
use sky130_fd_pr__nfet_01v8_lvt_28TRYY  sky130_fd_pr__nfet_01v8_lvt_28TRYY_0
timestamp 1654656593
transform 1 0 1191 0 1 3552
box -1591 -1097 1591 1097
use sky130_fd_pr__pfet_01v8_JJWXCM  sky130_fd_pr__pfet_01v8_JJWXCM_0
timestamp 1654656593
transform 1 0 1815 0 1 5160
box -777 -240 777 240
use sky130_fd_pr__pfet_01v8_JJWXCM  sky130_fd_pr__pfet_01v8_JJWXCM_1
timestamp 1654656593
transform 1 0 4015 0 1 5160
box -777 -240 777 240
use sky130_fd_pr__pfet_01v8_JJWXCM  sky130_fd_pr__pfet_01v8_JJWXCM_2
timestamp 1654656593
transform 1 0 6215 0 1 5160
box -777 -240 777 240
use sky130_fd_pr__pfet_01v8_lvt_SAWXCM  sky130_fd_pr__pfet_01v8_lvt_SAWXCM_0
timestamp 1654656593
transform 1 0 1816 0 1 5927
box -777 -240 777 240
use sky130_fd_pr__pfet_01v8_lvt_SAWXCM  sky130_fd_pr__pfet_01v8_lvt_SAWXCM_1
timestamp 1654656593
transform 1 0 4016 0 1 5927
box -777 -240 777 240
use sky130_fd_pr__pfet_01v8_lvt_SAWXCM  sky130_fd_pr__pfet_01v8_lvt_SAWXCM_2
timestamp 1654656593
transform 1 0 6216 0 1 5927
box -777 -240 777 240
<< labels >>
flabel metal2 1283 4772 1283 4772 1 FreeSans 800 0 0 0 bias_b
port 2 n
flabel metal3 6749 2677 6749 2677 1 FreeSans 800 0 0 0 bias_e
port 5 n
flabel metal2 1190 2273 1190 2273 1 FreeSans 800 0 0 0 bias_c
port 3 n
flabel metal1 -43 535 -43 535 1 FreeSans 800 0 0 0 i_bias
port 6 n
flabel metal1 8289 3446 8289 3446 1 FreeSans 800 0 0 0 bias_d
port 4 n
flabel metal1 8556 -250 8556 -250 1 FreeSans 800 0 0 0 bias_a
port 1 n
flabel locali -301 -525 -301 -525 1 FreeSans 800 0 0 0 VSS
port 8 n ground bidirectional
flabel locali -390 6367 -390 6367 1 FreeSans 800 0 0 0 VDD
port 7 n power bidirectional
<< end >>
