magic
tech sky130A
magscale 1 2
timestamp 1654674269
<< nwell >>
rect -1311 -241 1311 241
<< pmoslvt >>
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
<< pdiff >>
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
<< pdiffc >>
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
<< poly >>
rect -1199 221 -1115 237
rect -1199 205 -1183 221
rect -1217 187 -1183 205
rect -1131 205 -1115 221
rect -1021 221 -937 237
rect -1021 205 -1005 221
rect -1131 187 -1097 205
rect -1217 140 -1097 187
rect -1039 187 -1005 205
rect -953 205 -937 221
rect -843 221 -759 237
rect -843 205 -827 221
rect -953 187 -919 205
rect -1039 140 -919 187
rect -861 187 -827 205
rect -775 205 -759 221
rect -665 221 -581 237
rect -665 205 -649 221
rect -775 187 -741 205
rect -861 140 -741 187
rect -683 187 -649 205
rect -597 205 -581 221
rect -487 221 -403 237
rect -487 205 -471 221
rect -597 187 -563 205
rect -683 140 -563 187
rect -505 187 -471 205
rect -419 205 -403 221
rect -309 221 -225 237
rect -309 205 -293 221
rect -419 187 -385 205
rect -505 140 -385 187
rect -327 187 -293 205
rect -241 205 -225 221
rect -131 221 -47 237
rect -131 205 -115 221
rect -241 187 -207 205
rect -327 140 -207 187
rect -149 187 -115 205
rect -63 205 -47 221
rect 47 221 131 237
rect 47 205 63 221
rect -63 187 -29 205
rect -149 140 -29 187
rect 29 187 63 205
rect 115 205 131 221
rect 225 221 309 237
rect 225 205 241 221
rect 115 187 149 205
rect 29 140 149 187
rect 207 187 241 205
rect 293 205 309 221
rect 403 221 487 237
rect 403 205 419 221
rect 293 187 327 205
rect 207 140 327 187
rect 385 187 419 205
rect 471 205 487 221
rect 581 221 665 237
rect 581 205 597 221
rect 471 187 505 205
rect 385 140 505 187
rect 563 187 597 205
rect 649 205 665 221
rect 759 221 843 237
rect 759 205 775 221
rect 649 187 683 205
rect 563 140 683 187
rect 741 187 775 205
rect 827 205 843 221
rect 937 221 1021 237
rect 937 205 953 221
rect 827 187 861 205
rect 741 140 861 187
rect 919 187 953 205
rect 1005 205 1021 221
rect 1115 221 1199 237
rect 1115 205 1131 221
rect 1005 187 1039 205
rect 919 140 1039 187
rect 1097 187 1131 205
rect 1183 205 1199 221
rect 1183 187 1217 205
rect 1097 140 1217 187
rect -1217 -187 -1097 -140
rect -1217 -205 -1183 -187
rect -1199 -221 -1183 -205
rect -1131 -205 -1097 -187
rect -1039 -187 -919 -140
rect -1039 -205 -1005 -187
rect -1131 -221 -1115 -205
rect -1199 -237 -1115 -221
rect -1021 -221 -1005 -205
rect -953 -205 -919 -187
rect -861 -187 -741 -140
rect -861 -205 -827 -187
rect -953 -221 -937 -205
rect -1021 -237 -937 -221
rect -843 -221 -827 -205
rect -775 -205 -741 -187
rect -683 -187 -563 -140
rect -683 -205 -649 -187
rect -775 -221 -759 -205
rect -843 -237 -759 -221
rect -665 -221 -649 -205
rect -597 -205 -563 -187
rect -505 -187 -385 -140
rect -505 -205 -471 -187
rect -597 -221 -581 -205
rect -665 -237 -581 -221
rect -487 -221 -471 -205
rect -419 -205 -385 -187
rect -327 -187 -207 -140
rect -327 -205 -293 -187
rect -419 -221 -403 -205
rect -487 -237 -403 -221
rect -309 -221 -293 -205
rect -241 -205 -207 -187
rect -149 -187 -29 -140
rect -149 -205 -115 -187
rect -241 -221 -225 -205
rect -309 -237 -225 -221
rect -131 -221 -115 -205
rect -63 -205 -29 -187
rect 29 -187 149 -140
rect 29 -205 63 -187
rect -63 -221 -47 -205
rect -131 -237 -47 -221
rect 47 -221 63 -205
rect 115 -205 149 -187
rect 207 -187 327 -140
rect 207 -205 241 -187
rect 115 -221 131 -205
rect 47 -237 131 -221
rect 225 -221 241 -205
rect 293 -205 327 -187
rect 385 -187 505 -140
rect 385 -205 419 -187
rect 293 -221 309 -205
rect 225 -237 309 -221
rect 403 -221 419 -205
rect 471 -205 505 -187
rect 563 -187 683 -140
rect 563 -205 597 -187
rect 471 -221 487 -205
rect 403 -237 487 -221
rect 581 -221 597 -205
rect 649 -205 683 -187
rect 741 -187 861 -140
rect 741 -205 775 -187
rect 649 -221 665 -205
rect 581 -237 665 -221
rect 759 -221 775 -205
rect 827 -205 861 -187
rect 919 -187 1039 -140
rect 919 -205 953 -187
rect 827 -221 843 -205
rect 759 -237 843 -221
rect 937 -221 953 -205
rect 1005 -205 1039 -187
rect 1097 -187 1217 -140
rect 1097 -205 1131 -187
rect 1005 -221 1021 -205
rect 937 -237 1021 -221
rect 1115 -221 1131 -205
rect 1183 -205 1217 -187
rect 1183 -221 1199 -205
rect 1115 -237 1199 -221
<< polycont >>
rect -1183 187 -1131 221
rect -1005 187 -953 221
rect -827 187 -775 221
rect -649 187 -597 221
rect -471 187 -419 221
rect -293 187 -241 221
rect -115 187 -63 221
rect 63 187 115 221
rect 241 187 293 221
rect 419 187 471 221
rect 597 187 649 221
rect 775 187 827 221
rect 953 187 1005 221
rect 1131 187 1183 221
rect -1183 -221 -1131 -187
rect -1005 -221 -953 -187
rect -827 -221 -775 -187
rect -649 -221 -597 -187
rect -471 -221 -419 -187
rect -293 -221 -241 -187
rect -115 -221 -63 -187
rect 63 -221 115 -187
rect 241 -221 293 -187
rect 419 -221 471 -187
rect 597 -221 649 -187
rect 775 -221 827 -187
rect 953 -221 1005 -187
rect 1131 -221 1183 -187
<< locali >>
rect -1263 187 -1183 221
rect -1131 187 -1115 221
rect -1021 187 -1005 221
rect -953 187 -937 221
rect -843 187 -827 221
rect -775 187 -759 221
rect -665 187 -649 221
rect -597 187 -581 221
rect -487 187 -471 221
rect -419 187 -403 221
rect -309 187 -293 221
rect -241 187 -225 221
rect -131 187 -115 221
rect -63 187 -47 221
rect 47 187 63 221
rect 115 187 131 221
rect 225 187 241 221
rect 293 187 309 221
rect 403 187 419 221
rect 471 187 487 221
rect 581 187 597 221
rect 649 187 665 221
rect 759 187 775 221
rect 827 187 843 221
rect 937 187 953 221
rect 1005 187 1021 221
rect 1115 187 1131 221
rect 1183 187 1263 221
rect -1263 128 -1229 187
rect -1263 -187 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 187
rect 1229 -187 1263 -128
rect -1263 -221 -1183 -187
rect -1131 -221 -1115 -187
rect -1021 -221 -1005 -187
rect -953 -221 -937 -187
rect -843 -221 -827 -187
rect -775 -221 -759 -187
rect -665 -221 -649 -187
rect -597 -221 -581 -187
rect -487 -221 -471 -187
rect -419 -221 -403 -187
rect -309 -221 -293 -187
rect -241 -221 -225 -187
rect -131 -221 -115 -187
rect -63 -221 -47 -187
rect 47 -221 63 -187
rect 115 -221 131 -187
rect 225 -221 241 -187
rect 293 -221 309 -187
rect 403 -221 419 -187
rect 471 -221 487 -187
rect 581 -221 597 -187
rect 649 -221 665 -187
rect 759 -221 775 -187
rect 827 -221 843 -187
rect 937 -221 953 -187
rect 1005 -221 1021 -187
rect 1115 -221 1131 -187
rect 1183 -221 1263 -187
<< viali >>
rect -1005 187 -953 221
rect -827 187 -775 221
rect -649 187 -597 221
rect -471 187 -419 221
rect -293 187 -241 221
rect -115 187 -63 221
rect 63 187 115 221
rect 241 187 293 221
rect 419 187 471 221
rect 597 187 649 221
rect 775 187 827 221
rect 953 187 1005 221
rect -1005 -221 -953 -187
rect -827 -221 -775 -187
rect -649 -221 -597 -187
rect -471 -221 -419 -187
rect -293 -221 -241 -187
rect -115 -221 -63 -187
rect 63 -221 115 -187
rect 241 -221 293 -187
rect 419 -221 471 -187
rect 597 -221 649 -187
rect 775 -221 827 -187
rect 953 -221 1005 -187
<< metal1 >>
rect -1017 221 -941 227
rect -1017 187 -1005 221
rect -953 187 -941 221
rect -1017 181 -941 187
rect -839 221 -763 227
rect -839 187 -827 221
rect -775 187 -763 221
rect -839 181 -763 187
rect -661 221 -585 227
rect -661 187 -649 221
rect -597 187 -585 221
rect -661 181 -585 187
rect -483 221 -407 227
rect -483 187 -471 221
rect -419 187 -407 221
rect -483 181 -407 187
rect -305 221 -229 227
rect -305 187 -293 221
rect -241 187 -229 221
rect -305 181 -229 187
rect -127 221 -51 227
rect -127 187 -115 221
rect -63 187 -51 221
rect -127 181 -51 187
rect 51 221 127 227
rect 51 187 63 221
rect 115 187 127 221
rect 51 181 127 187
rect 229 221 305 227
rect 229 187 241 221
rect 293 187 305 221
rect 229 181 305 187
rect 407 221 483 227
rect 407 187 419 221
rect 471 187 483 221
rect 407 181 483 187
rect 585 221 661 227
rect 585 187 597 221
rect 649 187 661 221
rect 585 181 661 187
rect 763 221 839 227
rect 763 187 775 221
rect 827 187 839 221
rect 763 181 839 187
rect 941 221 1017 227
rect 941 187 953 221
rect 1005 187 1017 221
rect 941 181 1017 187
rect -1017 -187 -941 -181
rect -1017 -221 -1005 -187
rect -953 -221 -941 -187
rect -1017 -227 -941 -221
rect -839 -187 -763 -181
rect -839 -221 -827 -187
rect -775 -221 -763 -187
rect -839 -227 -763 -221
rect -661 -187 -585 -181
rect -661 -221 -649 -187
rect -597 -221 -585 -187
rect -661 -227 -585 -221
rect -483 -187 -407 -181
rect -483 -221 -471 -187
rect -419 -221 -407 -187
rect -483 -227 -407 -221
rect -305 -187 -229 -181
rect -305 -221 -293 -187
rect -241 -221 -229 -187
rect -305 -227 -229 -221
rect -127 -187 -51 -181
rect -127 -221 -115 -187
rect -63 -221 -51 -187
rect -127 -227 -51 -221
rect 51 -187 127 -181
rect 51 -221 63 -187
rect 115 -221 127 -187
rect 51 -227 127 -221
rect 229 -187 305 -181
rect 229 -221 241 -187
rect 293 -221 305 -187
rect 229 -227 305 -221
rect 407 -187 483 -181
rect 407 -221 419 -187
rect 471 -221 483 -187
rect 407 -227 483 -221
rect 585 -187 661 -181
rect 585 -221 597 -187
rect 649 -221 661 -187
rect 585 -227 661 -221
rect 763 -187 839 -181
rect 763 -221 775 -187
rect 827 -221 839 -187
rect 763 -227 839 -221
rect 941 -187 1017 -181
rect 941 -221 953 -187
rect 1005 -221 1017 -187
rect 941 -227 1017 -221
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 14 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
