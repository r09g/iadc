* NGSPICE file created from ota_w_test_v2.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_YVTR7C a_n207_n140# a_n1039_n205# a_29_n205# a_327_n140#
+ a_n683_n205# a_n1275_n140# a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_1097_n205#
+ a_n505_n205# a_n741_n140# a_563_n205# a_861_n140# w_n1311_n241# a_919_n205# a_n327_n205#
+ a_n563_n140# a_385_n205# a_683_n140# a_n919_n140# a_n149_n205# a_1039_n140# a_n385_n140#
+ a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_327_n140# a_207_n205# a_149_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_149_n140# a_29_n205# a_n29_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_861_n140# a_741_n205# a_683_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_n140# a_n327_n205# a_n385_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1097_n205# a_1097_n205# a_1039_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n741_n140# a_n861_n205# a_n919_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n1097_n140# a_n1275_n140# a_n1275_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_683_n140# a_563_n205# a_505_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1039_n140# a_919_n205# a_861_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n29_n140# a_n149_n205# a_n207_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n563_n140# a_n683_n205# a_n741_n140# w_n1311_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_505_n140# a_n563_n140# 0.01fF
C1 a_919_n205# a_1097_n205# 0.07fF
C2 a_n29_n140# a_149_n140# 0.06fF
C3 a_29_n205# a_n505_n205# 0.02fF
C4 a_n327_n205# a_n683_n205# 0.03fF
C5 a_683_n140# a_n207_n140# 0.01fF
C6 a_385_n205# a_n683_n205# 0.01fF
C7 a_n29_n140# a_861_n140# 0.01fF
C8 a_149_n140# a_683_n140# 0.02fF
C9 a_1097_n205# a_n385_n140# 0.01fF
C10 a_563_n205# a_1097_n205# 0.01fF
C11 a_741_n205# a_919_n205# 0.10fF
C12 a_207_n205# a_n149_n205# 0.03fF
C13 a_207_n205# a_n861_n205# 0.01fF
C14 a_385_n205# a_n327_n205# 0.01fF
C15 a_n1097_n140# w_n1311_n241# 0.02fF
C16 a_327_n140# a_n919_n140# 0.01fF
C17 a_149_n140# a_n207_n140# 0.03fF
C18 a_683_n140# a_861_n140# 0.06fF
C19 a_207_n205# a_n1039_n205# 0.01fF
C20 a_563_n205# a_741_n205# 0.10fF
C21 a_919_n205# a_29_n205# 0.01fF
C22 a_n149_n205# a_n683_n205# 0.02fF
C23 a_n1097_n140# a_n1275_n140# 0.06fF
C24 a_n861_n205# a_n683_n205# 0.10fF
C25 a_861_n140# a_n207_n140# 0.01fF
C26 a_207_n205# w_n1311_n241# 0.18fF
C27 a_n1039_n205# a_n683_n205# 0.03fF
C28 a_n29_n140# w_n1311_n241# 0.02fF
C29 a_149_n140# a_861_n140# 0.01fF
C30 a_n149_n205# a_n327_n205# 0.10fF
C31 a_741_n205# a_1097_n205# 0.02fF
C32 a_563_n205# a_29_n205# 0.02fF
C33 a_327_n140# a_n385_n140# 0.01fF
C34 a_385_n205# a_n149_n205# 0.02fF
C35 a_n327_n205# a_n861_n205# 0.02fF
C36 a_n919_n140# a_n741_n140# 0.06fF
C37 a_n1097_n140# a_n563_n140# 0.02fF
C38 a_n29_n140# a_1039_n140# 0.01fF
C39 a_385_n205# a_n861_n205# 0.01fF
C40 a_207_n205# a_n1275_n140# 0.00fF
C41 a_n327_n205# a_n1039_n205# 0.01fF
C42 a_n683_n205# w_n1311_n241# 0.20fF
C43 a_505_n140# a_n919_n140# 0.01fF
C44 a_n29_n140# a_n1275_n140# 0.01fF
C45 a_683_n140# w_n1311_n241# 0.02fF
C46 a_385_n205# a_n1039_n205# 0.01fF
C47 a_1097_n205# a_29_n205# 0.01fF
C48 a_1039_n140# a_683_n140# 0.03fF
C49 a_1097_n205# a_327_n140# 0.01fF
C50 a_n327_n205# w_n1311_n241# 0.20fF
C51 a_n1275_n140# a_n683_n205# 0.01fF
C52 a_n207_n140# w_n1311_n241# 0.02fF
C53 a_n29_n140# a_n563_n140# 0.02fF
C54 a_385_n205# w_n1311_n241# 0.17fF
C55 a_n741_n140# a_n385_n140# 0.03fF
C56 a_149_n140# w_n1311_n241# 0.02fF
C57 a_n149_n205# a_n861_n205# 0.01fF
C58 a_1039_n140# a_n207_n140# 0.01fF
C59 a_741_n205# a_29_n205# 0.01fF
C60 a_505_n140# a_n385_n140# 0.01fF
C61 a_n149_n205# a_n1039_n205# 0.01fF
C62 a_n1275_n140# a_n327_n205# 0.01fF
C63 a_149_n140# a_1039_n140# 0.01fF
C64 a_n1275_n140# a_n207_n140# 0.01fF
C65 a_n563_n140# a_683_n140# 0.01fF
C66 a_385_n205# a_n1275_n140# 0.00fF
C67 a_n1039_n205# a_n861_n205# 0.10fF
C68 a_149_n140# a_n1275_n140# 0.01fF
C69 a_861_n140# w_n1311_n241# 0.01fF
C70 a_n149_n205# w_n1311_n241# 0.19fF
C71 a_1039_n140# a_861_n140# 0.06fF
C72 a_1097_n205# a_505_n140# 0.01fF
C73 a_n563_n140# a_n207_n140# 0.03fF
C74 a_n861_n205# w_n1311_n241# 0.20fF
C75 a_149_n140# a_n563_n140# 0.01fF
C76 a_n1039_n205# w_n1311_n241# 0.20fF
C77 a_n149_n205# a_n1275_n140# 0.01fF
C78 a_n1097_n140# a_n919_n140# 0.06fF
C79 a_207_n205# a_n505_n205# 0.01fF
C80 a_n1275_n140# a_n861_n205# 0.02fF
C81 a_n563_n140# a_861_n140# 0.01fF
C82 a_n1275_n140# a_n1039_n205# 0.07fF
C83 a_327_n140# a_n741_n140# 0.01fF
C84 a_1039_n140# w_n1311_n241# 0.01fF
C85 a_n505_n205# a_n683_n205# 0.10fF
C86 a_327_n140# a_505_n140# 0.06fF
C87 a_n29_n140# a_n919_n140# 0.01fF
C88 a_n1275_n140# w_n1311_n241# 0.33fF
C89 a_n1097_n140# a_n385_n140# 0.01fF
C90 a_207_n205# a_919_n205# 0.01fF
C91 a_n505_n205# a_n327_n205# 0.10fF
C92 a_385_n205# a_n505_n205# 0.01fF
C93 a_n919_n140# a_683_n140# 0.01fF
C94 a_n563_n140# w_n1311_n241# 0.02fF
C95 a_919_n205# a_n683_n205# 0.01fF
C96 a_563_n205# a_207_n205# 0.03fF
C97 a_n563_n140# a_1039_n140# 0.01fF
C98 a_n29_n140# a_n385_n140# 0.03fF
C99 a_505_n140# a_n741_n140# 0.01fF
C100 a_n919_n140# a_n207_n140# 0.01fF
C101 a_n563_n140# a_n1275_n140# 0.01fF
C102 a_149_n140# a_n919_n140# 0.01fF
C103 a_919_n205# a_n327_n205# 0.01fF
C104 a_n149_n205# a_n505_n205# 0.03fF
C105 a_683_n140# a_n385_n140# 0.01fF
C106 a_563_n205# a_n683_n205# 0.01fF
C107 a_207_n205# a_1097_n205# 0.01fF
C108 a_385_n205# a_919_n205# 0.02fF
C109 a_n505_n205# a_n861_n205# 0.03fF
C110 a_1097_n205# a_n29_n140# 0.01fF
C111 a_n505_n205# a_n1039_n205# 0.02fF
C112 a_563_n205# a_n327_n205# 0.01fF
C113 a_n385_n140# a_n207_n140# 0.06fF
C114 a_563_n205# a_385_n205# 0.10fF
C115 a_741_n205# a_207_n205# 0.02fF
C116 a_1097_n205# a_683_n140# 0.02fF
C117 a_327_n140# a_n1097_n140# 0.01fF
C118 a_149_n140# a_n385_n140# 0.02fF
C119 a_n505_n205# w_n1311_n241# 0.20fF
C120 a_919_n205# a_n149_n205# 0.01fF
C121 a_1097_n205# a_n327_n205# 0.00fF
C122 a_1097_n205# a_n207_n140# 0.01fF
C123 a_861_n140# a_n385_n140# 0.01fF
C124 a_741_n205# a_n683_n205# 0.01fF
C125 a_385_n205# a_1097_n205# 0.01fF
C126 a_207_n205# a_29_n205# 0.10fF
C127 a_1097_n205# a_149_n140# 0.01fF
C128 a_n1275_n140# a_n505_n205# 0.01fF
C129 a_n29_n140# a_327_n140# 0.03fF
C130 a_563_n205# a_n149_n205# 0.01fF
C131 a_n919_n140# w_n1311_n241# 0.02fF
C132 a_n1097_n140# a_n741_n140# 0.03fF
C133 a_741_n205# a_n327_n205# 0.01fF
C134 a_563_n205# a_n861_n205# 0.01fF
C135 a_919_n205# w_n1311_n241# 0.14fF
C136 a_741_n205# a_385_n205# 0.03fF
C137 a_1097_n205# a_861_n140# 0.03fF
C138 a_505_n140# a_n1097_n140# 0.01fF
C139 a_29_n205# a_n683_n205# 0.01fF
C140 a_563_n205# a_n1039_n205# 0.01fF
C141 a_327_n140# a_683_n140# 0.03fF
C142 a_n919_n140# a_n1275_n140# 0.03fF
C143 a_1097_n205# a_n149_n205# 0.00fF
C144 a_29_n205# a_n327_n205# 0.03fF
C145 a_n385_n140# w_n1311_n241# 0.02fF
C146 a_563_n205# w_n1311_n241# 0.16fF
C147 a_n29_n140# a_n741_n140# 0.01fF
C148 a_327_n140# a_n207_n140# 0.02fF
C149 a_385_n205# a_29_n205# 0.03fF
C150 a_n919_n140# a_n563_n140# 0.03fF
C151 a_n29_n140# a_505_n140# 0.02fF
C152 a_149_n140# a_327_n140# 0.06fF
C153 a_1039_n140# a_n385_n140# 0.01fF
C154 a_741_n205# a_n149_n205# 0.01fF
C155 a_n1275_n140# a_n385_n140# 0.01fF
C156 a_741_n205# a_n861_n205# 0.01fF
C157 a_n741_n140# a_683_n140# 0.01fF
C158 a_1097_n205# w_n1311_n241# 0.28fF
C159 a_327_n140# a_861_n140# 0.02fF
C160 a_505_n140# a_683_n140# 0.06fF
C161 a_1097_n205# a_1039_n140# 0.06fF
C162 a_n149_n205# a_29_n205# 0.10fF
C163 a_n741_n140# a_n207_n140# 0.02fF
C164 a_n563_n140# a_n385_n140# 0.06fF
C165 a_29_n205# a_n861_n205# 0.01fF
C166 a_149_n140# a_n741_n140# 0.01fF
C167 a_741_n205# w_n1311_n241# 0.15fF
C168 a_505_n140# a_n207_n140# 0.01fF
C169 a_29_n205# a_n1039_n205# 0.01fF
C170 a_149_n140# a_505_n140# 0.03fF
C171 a_n741_n140# a_861_n140# 0.01fF
C172 a_29_n205# w_n1311_n241# 0.19fF
C173 a_327_n140# w_n1311_n241# 0.02fF
C174 a_505_n140# a_861_n140# 0.03fF
C175 a_919_n205# a_n505_n205# 0.01fF
C176 a_327_n140# a_1039_n140# 0.01fF
C177 a_n29_n140# a_n1097_n140# 0.01fF
C178 a_29_n205# a_n1275_n140# 0.00fF
C179 a_327_n140# a_n1275_n140# 0.01fF
C180 a_563_n205# a_n505_n205# 0.01fF
C181 a_n741_n140# w_n1311_n241# 0.02fF
C182 a_327_n140# a_n563_n140# 0.01fF
C183 a_505_n140# w_n1311_n241# 0.02fF
C184 a_1097_n205# a_n505_n205# 0.00fF
C185 a_n919_n140# a_n385_n140# 0.02fF
C186 a_n1097_n140# a_n207_n140# 0.01fF
C187 a_n741_n140# a_n1275_n140# 0.02fF
C188 a_505_n140# a_1039_n140# 0.02fF
C189 a_207_n205# a_n683_n205# 0.01fF
C190 a_149_n140# a_n1097_n140# 0.01fF
C191 a_n29_n140# a_683_n140# 0.01fF
C192 a_563_n205# a_919_n205# 0.03fF
C193 a_n741_n140# a_n563_n140# 0.06fF
C194 a_741_n205# a_n505_n205# 0.01fF
C195 a_207_n205# a_n327_n205# 0.02fF
C196 a_207_n205# a_385_n205# 0.10fF
C197 a_n29_n140# a_n207_n140# 0.06fF
C198 w_n1311_n241# VSUBS 3.79fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AKSJZW a_n149_n195# a_n207_n140# a_207_n195# a_327_n140#
+ a_n1275_n140# a_n861_n195# a_n29_n140# a_149_n140# a_n1097_n140# a_n1039_n195# a_29_n195#
+ a_n683_n195# a_n741_n140# a_741_n195# a_861_n140# a_1097_n195# a_n563_n140# a_n505_n195#
+ a_563_n195# a_683_n140# a_n919_n140# a_919_n195# a_1039_n140# a_n385_n140# a_n327_n195#
+ a_385_n195# a_505_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n195# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n195# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n195# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n195# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_327_n140# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_861_n140# a_741_n195# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n207_n140# a_n327_n195# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_1097_n195# a_1097_n195# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n195# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1275_n140# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n195# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n195# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_29_n195# a_n683_n195# 0.01fF
C1 a_1039_n140# a_149_n140# 0.01fF
C2 a_n327_n195# a_385_n195# 0.01fF
C3 a_327_n140# a_1097_n195# 0.01fF
C4 a_n741_n140# a_n919_n140# 0.06fF
C5 a_n1097_n140# a_n919_n140# 0.06fF
C6 a_n1039_n195# a_563_n195# 0.01fF
C7 a_n29_n140# a_n1275_n140# 0.01fF
C8 a_n385_n140# a_861_n140# 0.01fF
C9 a_n207_n140# a_n741_n140# 0.02fF
C10 a_n207_n140# a_n1097_n140# 0.01fF
C11 a_n563_n140# a_n1097_n140# 0.02fF
C12 a_n563_n140# a_n741_n140# 0.06fF
C13 a_207_n195# a_385_n195# 0.10fF
C14 a_n861_n195# a_385_n195# 0.01fF
C15 a_505_n140# a_1097_n195# 0.01fF
C16 a_n327_n195# a_919_n195# 0.01fF
C17 a_563_n195# a_1097_n195# 0.01fF
C18 a_n1097_n140# a_149_n140# 0.01fF
C19 a_n741_n140# a_149_n140# 0.01fF
C20 a_741_n195# a_563_n195# 0.10fF
C21 a_n505_n195# a_563_n195# 0.01fF
C22 a_n149_n195# a_n1039_n195# 0.01fF
C23 a_385_n195# a_n1275_n140# 0.00fF
C24 a_683_n140# a_1097_n195# 0.02fF
C25 a_207_n195# a_919_n195# 0.01fF
C26 a_327_n140# a_n919_n140# 0.01fF
C27 a_n1039_n195# a_n683_n195# 0.03fF
C28 a_29_n195# a_n1039_n195# 0.01fF
C29 a_n207_n140# a_327_n140# 0.02fF
C30 a_n149_n195# a_1097_n195# 0.00fF
C31 a_327_n140# a_n563_n140# 0.01fF
C32 a_n149_n195# a_741_n195# 0.01fF
C33 a_n29_n140# a_1039_n140# 0.01fF
C34 a_n149_n195# a_n505_n195# 0.03fF
C35 a_505_n140# a_n919_n140# 0.01fF
C36 a_505_n140# a_n207_n140# 0.01fF
C37 a_327_n140# a_149_n140# 0.06fF
C38 a_29_n195# a_1097_n195# 0.01fF
C39 a_505_n140# a_n563_n140# 0.01fF
C40 a_741_n195# a_n683_n195# 0.01fF
C41 a_29_n195# a_741_n195# 0.01fF
C42 a_n1097_n140# a_n1275_n140# 0.06fF
C43 a_n741_n140# a_n1275_n140# 0.02fF
C44 a_1097_n195# a_861_n140# 0.03fF
C45 a_n505_n195# a_n683_n195# 0.10fF
C46 a_n385_n140# a_1097_n195# 0.01fF
C47 a_29_n195# a_n505_n195# 0.02fF
C48 a_683_n140# a_n919_n140# 0.01fF
C49 a_505_n140# a_149_n140# 0.03fF
C50 a_n207_n140# a_683_n140# 0.01fF
C51 a_n29_n140# a_n1097_n140# 0.01fF
C52 a_n741_n140# a_n29_n140# 0.01fF
C53 a_n563_n140# a_683_n140# 0.01fF
C54 a_n327_n195# a_563_n195# 0.01fF
C55 a_385_n195# a_919_n195# 0.02fF
C56 a_683_n140# a_149_n140# 0.02fF
C57 a_327_n140# a_n1275_n140# 0.01fF
C58 a_207_n195# a_563_n195# 0.03fF
C59 a_n385_n140# a_n919_n140# 0.02fF
C60 a_n207_n140# a_861_n140# 0.01fF
C61 a_n861_n195# a_563_n195# 0.01fF
C62 a_n207_n140# a_n385_n140# 0.06fF
C63 a_n563_n140# a_861_n140# 0.01fF
C64 a_n563_n140# a_n385_n140# 0.06fF
C65 a_n149_n195# a_n327_n195# 0.10fF
C66 a_327_n140# a_n29_n140# 0.03fF
C67 a_n1039_n195# a_n505_n195# 0.02fF
C68 a_861_n140# a_149_n140# 0.01fF
C69 a_n385_n140# a_149_n140# 0.02fF
C70 a_n327_n195# a_n683_n195# 0.03fF
C71 a_29_n195# a_n327_n195# 0.03fF
C72 a_207_n195# a_n149_n195# 0.03fF
C73 a_741_n195# a_1097_n195# 0.02fF
C74 a_505_n140# a_n29_n140# 0.02fF
C75 a_n149_n195# a_n861_n195# 0.01fF
C76 a_n505_n195# a_1097_n195# 0.00fF
C77 a_741_n195# a_n505_n195# 0.01fF
C78 a_n741_n140# a_n1097_n140# 0.03fF
C79 a_207_n195# a_n683_n195# 0.01fF
C80 a_29_n195# a_207_n195# 0.10fF
C81 a_n149_n195# a_n1275_n140# 0.01fF
C82 a_n861_n195# a_n683_n195# 0.10fF
C83 a_29_n195# a_n861_n195# 0.01fF
C84 a_683_n140# a_n29_n140# 0.01fF
C85 a_327_n140# a_1039_n140# 0.01fF
C86 a_385_n195# a_563_n195# 0.10fF
C87 a_n1275_n140# a_n683_n195# 0.01fF
C88 a_29_n195# a_n1275_n140# 0.00fF
C89 a_505_n140# a_1039_n140# 0.02fF
C90 a_n385_n140# a_n1275_n140# 0.01fF
C91 a_n207_n140# a_1097_n195# 0.01fF
C92 a_327_n140# a_n1097_n140# 0.01fF
C93 a_327_n140# a_n741_n140# 0.01fF
C94 a_n1039_n195# a_n327_n195# 0.01fF
C95 a_n29_n140# a_861_n140# 0.01fF
C96 a_n385_n140# a_n29_n140# 0.03fF
C97 a_563_n195# a_919_n195# 0.03fF
C98 a_683_n140# a_1039_n140# 0.03fF
C99 a_n149_n195# a_385_n195# 0.02fF
C100 a_1097_n195# a_149_n140# 0.01fF
C101 a_505_n140# a_n1097_n140# 0.01fF
C102 a_505_n140# a_n741_n140# 0.01fF
C103 a_207_n195# a_n1039_n195# 0.01fF
C104 a_n327_n195# a_1097_n195# 0.00fF
C105 a_n861_n195# a_n1039_n195# 0.10fF
C106 a_385_n195# a_n683_n195# 0.01fF
C107 a_n327_n195# a_741_n195# 0.01fF
C108 a_29_n195# a_385_n195# 0.03fF
C109 a_n327_n195# a_n505_n195# 0.10fF
C110 a_n149_n195# a_919_n195# 0.01fF
C111 a_n207_n140# a_n919_n140# 0.01fF
C112 a_n741_n140# a_683_n140# 0.01fF
C113 a_n1039_n195# a_n1275_n140# 0.06fF
C114 a_n563_n140# a_n919_n140# 0.03fF
C115 a_207_n195# a_1097_n195# 0.01fF
C116 a_1039_n140# a_861_n140# 0.06fF
C117 a_n207_n140# a_n563_n140# 0.03fF
C118 a_n385_n140# a_1039_n140# 0.01fF
C119 a_207_n195# a_741_n195# 0.02fF
C120 a_n861_n195# a_741_n195# 0.01fF
C121 a_207_n195# a_n505_n195# 0.01fF
C122 a_n683_n195# a_919_n195# 0.01fF
C123 a_29_n195# a_919_n195# 0.01fF
C124 a_n861_n195# a_n505_n195# 0.03fF
C125 a_149_n140# a_n919_n140# 0.01fF
C126 a_n207_n140# a_149_n140# 0.03fF
C127 a_n563_n140# a_149_n140# 0.01fF
C128 a_505_n140# a_327_n140# 0.06fF
C129 a_n505_n195# a_n1275_n140# 0.01fF
C130 a_n741_n140# a_861_n140# 0.01fF
C131 a_n385_n140# a_n741_n140# 0.03fF
C132 a_n385_n140# a_n1097_n140# 0.01fF
C133 a_n29_n140# a_1097_n195# 0.01fF
C134 a_327_n140# a_683_n140# 0.03fF
C135 a_n1039_n195# a_385_n195# 0.01fF
C136 a_505_n140# a_683_n140# 0.06fF
C137 a_385_n195# a_1097_n195# 0.01fF
C138 a_n1275_n140# a_n919_n140# 0.03fF
C139 a_741_n195# a_385_n195# 0.03fF
C140 a_n207_n140# a_n1275_n140# 0.01fF
C141 a_n563_n140# a_n1275_n140# 0.01fF
C142 a_385_n195# a_n505_n195# 0.01fF
C143 a_1097_n195# a_1039_n140# 0.06fF
C144 a_n149_n195# a_563_n195# 0.01fF
C145 a_327_n140# a_861_n140# 0.02fF
C146 a_207_n195# a_n327_n195# 0.02fF
C147 a_327_n140# a_n385_n140# 0.01fF
C148 a_n29_n140# a_n919_n140# 0.01fF
C149 a_n861_n195# a_n327_n195# 0.02fF
C150 a_n207_n140# a_n29_n140# 0.06fF
C151 a_n1275_n140# a_149_n140# 0.01fF
C152 a_n563_n140# a_n29_n140# 0.02fF
C153 a_1097_n195# a_919_n195# 0.06fF
C154 a_563_n195# a_n683_n195# 0.01fF
C155 a_29_n195# a_563_n195# 0.02fF
C156 a_741_n195# a_919_n195# 0.10fF
C157 a_505_n140# a_861_n140# 0.03fF
C158 a_n327_n195# a_n1275_n140# 0.01fF
C159 a_n505_n195# a_919_n195# 0.01fF
C160 a_505_n140# a_n385_n140# 0.01fF
C161 a_n29_n140# a_149_n140# 0.06fF
C162 a_207_n195# a_n861_n195# 0.01fF
C163 a_683_n140# a_861_n140# 0.06fF
C164 a_n385_n140# a_683_n140# 0.01fF
C165 a_207_n195# a_n1275_n140# 0.00fF
C166 a_n861_n195# a_n1275_n140# 0.02fF
C167 a_n149_n195# a_n683_n195# 0.02fF
C168 a_n207_n140# a_1039_n140# 0.01fF
C169 a_29_n195# a_n149_n195# 0.10fF
C170 a_n563_n140# a_1039_n140# 0.01fF
C171 a_1039_n140# VSUBS 0.01fF
C172 a_861_n140# VSUBS 0.01fF
C173 a_683_n140# VSUBS 0.02fF
C174 a_505_n140# VSUBS 0.02fF
C175 a_327_n140# VSUBS 0.02fF
C176 a_149_n140# VSUBS 0.02fF
C177 a_n29_n140# VSUBS 0.02fF
C178 a_n207_n140# VSUBS 0.02fF
C179 a_n385_n140# VSUBS 0.02fF
C180 a_n563_n140# VSUBS 0.02fF
C181 a_n741_n140# VSUBS 0.02fF
C182 a_n919_n140# VSUBS 0.02fF
C183 a_n1097_n140# VSUBS 0.02fF
C184 a_1097_n195# VSUBS 0.31fF
C185 a_919_n195# VSUBS 0.19fF
C186 a_741_n195# VSUBS 0.20fF
C187 a_563_n195# VSUBS 0.21fF
C188 a_385_n195# VSUBS 0.22fF
C189 a_207_n195# VSUBS 0.23fF
C190 a_29_n195# VSUBS 0.23fF
C191 a_n149_n195# VSUBS 0.24fF
C192 a_n327_n195# VSUBS 0.24fF
C193 a_n505_n195# VSUBS 0.24fF
C194 a_n683_n195# VSUBS 0.24fF
C195 a_n861_n195# VSUBS 0.24fF
C196 a_n1039_n195# VSUBS 0.24fF
C197 a_n1275_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_K7HVMB a_664_n120# a_n608_n120# a_n86_n120# a_72_n208#
+ a_240_n120# a_n184_n120# a_n562_142# a_n510_n120# a_28_n120# a_n298_n120# a_126_n120#
+ a_452_n120# a_n396_n120# a_284_142# a_n138_142# a_550_n120# a_496_n208# a_338_n120#
+ a_n350_n208# a_n820_n120# VSUBS
X0 a_n820_n120# a_n820_n120# a_n820_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X1 a_n510_n120# a_n562_142# a_n608_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X2 a_664_n120# a_664_n120# a_664_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=6.96e+11p pd=5.96e+06u as=0p ps=0u w=1.2e+06u l=200000u
X3 a_n298_n120# a_n350_n208# a_n396_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X4 a_550_n120# a_496_n208# a_452_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X5 a_126_n120# a_72_n208# a_28_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X6 a_n86_n120# a_n138_142# a_n184_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
X7 a_338_n120# a_284_142# a_240_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
C0 a_n86_n120# a_338_n120# 0.02fF
C1 a_126_n120# a_n298_n120# 0.02fF
C2 a_n350_n208# a_496_n208# 0.01fF
C3 a_550_n120# a_n396_n120# 0.01fF
C4 a_n184_n120# a_n298_n120# 0.09fF
C5 a_452_n120# a_n298_n120# 0.01fF
C6 a_550_n120# a_n820_n120# 0.01fF
C7 a_126_n120# a_n608_n120# 0.01fF
C8 a_n138_142# a_496_n208# 0.00fF
C9 a_664_n120# a_284_142# 0.01fF
C10 a_n510_n120# a_n396_n120# 0.09fF
C11 a_240_n120# a_n396_n120# 0.01fF
C12 a_28_n120# a_550_n120# 0.01fF
C13 a_126_n120# a_664_n120# 0.03fF
C14 a_n820_n120# a_496_n208# 0.00fF
C15 a_n184_n120# a_n608_n120# 0.02fF
C16 a_452_n120# a_n608_n120# 0.01fF
C17 a_n510_n120# a_n820_n120# 0.06fF
C18 a_n820_n120# a_240_n120# 0.01fF
C19 a_550_n120# a_338_n120# 0.04fF
C20 a_n86_n120# a_550_n120# 0.01fF
C21 a_n184_n120# a_664_n120# 0.02fF
C22 a_28_n120# a_n510_n120# 0.01fF
C23 a_452_n120# a_664_n120# 0.06fF
C24 a_28_n120# a_240_n120# 0.04fF
C25 a_n350_n208# a_284_142# 0.00fF
C26 a_n510_n120# a_338_n120# 0.01fF
C27 a_n86_n120# a_n510_n120# 0.02fF
C28 a_496_n208# a_n562_142# 0.00fF
C29 a_240_n120# a_338_n120# 0.11fF
C30 a_n86_n120# a_240_n120# 0.02fF
C31 a_n510_n120# a_n562_142# 0.00fF
C32 a_n138_142# a_284_142# 0.01fF
C33 a_72_n208# a_664_n120# 0.00fF
C34 a_126_n120# a_n396_n120# 0.01fF
C35 a_n298_n120# a_n608_n120# 0.03fF
C36 a_n820_n120# a_284_142# 0.00fF
C37 a_n298_n120# a_664_n120# 0.01fF
C38 a_126_n120# a_n820_n120# 0.02fF
C39 a_n184_n120# a_n396_n120# 0.04fF
C40 a_452_n120# a_n396_n120# 0.01fF
C41 a_28_n120# a_126_n120# 0.11fF
C42 a_550_n120# a_n510_n120# 0.01fF
C43 a_n350_n208# a_72_n208# 0.01fF
C44 a_550_n120# a_240_n120# 0.03fF
C45 a_n184_n120# a_n820_n120# 0.03fF
C46 a_452_n120# a_n820_n120# 0.01fF
C47 a_n562_142# a_284_142# 0.01fF
C48 a_664_n120# a_n608_n120# 0.01fF
C49 a_126_n120# a_338_n120# 0.04fF
C50 a_n86_n120# a_126_n120# 0.04fF
C51 a_n184_n120# a_28_n120# 0.04fF
C52 a_n138_142# a_72_n208# 0.01fF
C53 a_28_n120# a_452_n120# 0.02fF
C54 a_n510_n120# a_240_n120# 0.01fF
C55 a_n350_n208# a_n298_n120# 0.00fF
C56 a_n184_n120# a_338_n120# 0.01fF
C57 a_n86_n120# a_n184_n120# 0.11fF
C58 a_452_n120# a_338_n120# 0.09fF
C59 a_n86_n120# a_452_n120# 0.01fF
C60 a_n820_n120# a_72_n208# 0.00fF
C61 a_n298_n120# a_n396_n120# 0.11fF
C62 a_28_n120# a_72_n208# 0.00fF
C63 a_n298_n120# a_n820_n120# 0.03fF
C64 a_n350_n208# a_664_n120# 0.00fF
C65 a_550_n120# a_126_n120# 0.02fF
C66 a_72_n208# a_n562_142# 0.00fF
C67 a_n396_n120# a_n608_n120# 0.04fF
C68 a_28_n120# a_n298_n120# 0.02fF
C69 a_496_n208# a_284_142# 0.01fF
C70 a_240_n120# a_284_142# 0.00fF
C71 a_n138_142# a_664_n120# 0.00fF
C72 a_664_n120# a_n396_n120# 0.01fF
C73 a_n184_n120# a_550_n120# 0.01fF
C74 a_n820_n120# a_n608_n120# 0.13fF
C75 a_452_n120# a_550_n120# 0.11fF
C76 a_n298_n120# a_338_n120# 0.01fF
C77 a_126_n120# a_n510_n120# 0.01fF
C78 a_n86_n120# a_n298_n120# 0.04fF
C79 a_126_n120# a_240_n120# 0.09fF
C80 a_28_n120# a_n608_n120# 0.01fF
C81 a_n820_n120# a_664_n120# 0.02fF
C82 a_452_n120# a_496_n208# 0.00fF
C83 a_n184_n120# a_n510_n120# 0.02fF
C84 a_452_n120# a_n510_n120# 0.01fF
C85 a_n184_n120# a_240_n120# 0.02fF
C86 a_28_n120# a_664_n120# 0.02fF
C87 a_338_n120# a_n608_n120# 0.01fF
C88 a_452_n120# a_240_n120# 0.04fF
C89 a_n86_n120# a_n608_n120# 0.01fF
C90 a_n138_142# a_n350_n208# 0.01fF
C91 a_664_n120# a_338_n120# 0.04fF
C92 a_n86_n120# a_664_n120# 0.02fF
C93 a_664_n120# a_n562_142# 0.00fF
C94 a_72_n208# a_496_n208# 0.01fF
C95 a_n350_n208# a_n820_n120# 0.01fF
C96 a_550_n120# a_n298_n120# 0.01fF
C97 a_n138_142# a_n820_n120# 0.00fF
C98 a_n820_n120# a_n396_n120# 0.04fF
C99 a_n510_n120# a_n298_n120# 0.04fF
C100 a_550_n120# a_n608_n120# 0.01fF
C101 a_n298_n120# a_240_n120# 0.01fF
C102 a_28_n120# a_n396_n120# 0.02fF
C103 a_n350_n208# a_n562_142# 0.01fF
C104 a_n184_n120# a_126_n120# 0.03fF
C105 a_452_n120# a_126_n120# 0.02fF
C106 a_550_n120# a_664_n120# 0.13fF
C107 a_n86_n120# a_n138_142# 0.00fF
C108 a_28_n120# a_n820_n120# 0.02fF
C109 a_n396_n120# a_338_n120# 0.01fF
C110 a_n86_n120# a_n396_n120# 0.03fF
C111 a_n510_n120# a_n608_n120# 0.11fF
C112 a_n138_142# a_n562_142# 0.01fF
C113 a_240_n120# a_n608_n120# 0.01fF
C114 a_72_n208# a_284_142# 0.01fF
C115 a_n184_n120# a_452_n120# 0.01fF
C116 a_664_n120# a_496_n208# 0.01fF
C117 a_n820_n120# a_338_n120# 0.01fF
C118 a_n510_n120# a_664_n120# 0.01fF
C119 a_n86_n120# a_n820_n120# 0.02fF
C120 a_240_n120# a_664_n120# 0.03fF
C121 a_n820_n120# a_n562_142# 0.01fF
C122 a_28_n120# a_338_n120# 0.03fF
C123 a_n86_n120# a_28_n120# 0.09fF
C124 a_550_n120# VSUBS 0.01fF
C125 a_452_n120# VSUBS 0.01fF
C126 a_338_n120# VSUBS 0.01fF
C127 a_240_n120# VSUBS 0.01fF
C128 a_126_n120# VSUBS 0.02fF
C129 a_28_n120# VSUBS 0.01fF
C130 a_n86_n120# VSUBS 0.01fF
C131 a_n184_n120# VSUBS 0.02fF
C132 a_n298_n120# VSUBS 0.02fF
C133 a_n396_n120# VSUBS 0.02fF
C134 a_n510_n120# VSUBS 0.02fF
C135 a_n608_n120# VSUBS 0.02fF
C136 a_496_n208# VSUBS 0.11fF
C137 a_664_n120# VSUBS 0.17fF
C138 a_72_n208# VSUBS 0.10fF
C139 a_284_142# VSUBS 0.10fF
C140 a_n350_n208# VSUBS 0.12fF
C141 a_n138_142# VSUBS 0.11fF
C142 a_n820_n120# VSUBS 0.20fF
C143 a_n562_142# VSUBS 0.14fF
.ends

.subckt sky130_fd_pr__nfet_01v8_S6RQQZ a_n149_n194# a_n207_n140# a_207_n194# a_1453_n194#
+ a_n1217_n194# a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140#
+ a_n1097_n140# a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194#
+ a_861_n140# a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140#
+ a_n919_n140# a_919_n194# a_n1631_n140# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194#
+ a_n1395_n194# a_505_n140# a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n1453_n140# a_n1631_n140# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1453_n194# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n327_n194# a_n1039_n194# 0.01fF
C1 a_n683_n194# a_29_n194# 0.01fF
C2 a_1217_n140# a_327_n140# 0.01fF
C3 a_n1631_n140# a_n29_n140# 0.01fF
C4 a_1395_n140# a_861_n140# 0.02fF
C5 a_n563_n140# a_n1631_n140# 0.01fF
C6 a_n385_n140# a_n1631_n140# 0.01fF
C7 a_1453_n194# a_741_n194# 0.01fF
C8 a_n207_n140# a_n29_n140# 0.06fF
C9 a_n1395_n194# a_207_n194# 0.01fF
C10 a_149_n140# a_n1097_n140# 0.01fF
C11 a_n563_n140# a_n207_n140# 0.03fF
C12 a_1453_n194# a_385_n194# 0.01fF
C13 a_n385_n140# a_n207_n140# 0.06fF
C14 a_1275_n194# a_563_n194# 0.01fF
C15 a_n149_n194# a_29_n194# 0.10fF
C16 a_n1217_n194# a_29_n194# 0.01fF
C17 a_n683_n194# a_563_n194# 0.01fF
C18 a_1217_n140# a_149_n140# 0.01fF
C19 a_207_n194# a_741_n194# 0.02fF
C20 a_919_n194# a_1275_n194# 0.03fF
C21 a_385_n194# a_207_n194# 0.10fF
C22 a_n683_n194# a_n1631_n140# 0.01fF
C23 a_n861_n194# a_207_n194# 0.01fF
C24 a_n505_n194# a_n1395_n194# 0.01fF
C25 a_1395_n140# a_1039_n140# 0.03fF
C26 a_n683_n194# a_919_n194# 0.01fF
C27 a_n149_n194# a_563_n194# 0.01fF
C28 a_505_n140# a_n29_n140# 0.02fF
C29 a_861_n140# a_n207_n140# 0.01fF
C30 a_n563_n140# a_505_n140# 0.01fF
C31 a_29_n194# a_1097_n194# 0.01fF
C32 a_1453_n194# a_n29_n140# 0.01fF
C33 a_n1395_n194# a_n1039_n194# 0.03fF
C34 a_n149_n194# a_n1631_n140# 0.00fF
C35 a_n327_n194# a_n1395_n194# 0.01fF
C36 a_n385_n140# a_505_n140# 0.01fF
C37 a_n1217_n194# a_n1631_n140# 0.02fF
C38 a_n505_n194# a_741_n194# 0.01fF
C39 a_n149_n194# a_919_n194# 0.01fF
C40 a_n505_n194# a_385_n194# 0.01fF
C41 a_n505_n194# a_n861_n194# 0.03fF
C42 a_n1453_n140# a_n29_n140# 0.01fF
C43 a_n1453_n140# a_n563_n140# 0.01fF
C44 a_1453_n194# a_1275_n194# 0.06fF
C45 a_n327_n194# a_741_n194# 0.01fF
C46 a_n741_n140# a_n29_n140# 0.01fF
C47 a_n1453_n140# a_n385_n140# 0.01fF
C48 a_385_n194# a_n1039_n194# 0.01fF
C49 a_n327_n194# a_385_n194# 0.01fF
C50 a_n563_n140# a_n741_n140# 0.06fF
C51 a_1097_n194# a_563_n194# 0.02fF
C52 a_n861_n194# a_n1039_n194# 0.10fF
C53 a_n385_n140# a_n741_n140# 0.03fF
C54 a_n327_n194# a_n861_n194# 0.02fF
C55 a_683_n140# a_n29_n140# 0.01fF
C56 a_1039_n140# a_n207_n140# 0.01fF
C57 a_n563_n140# a_683_n140# 0.01fF
C58 a_n1275_n140# a_n29_n140# 0.01fF
C59 a_n385_n140# a_683_n140# 0.01fF
C60 a_861_n140# a_505_n140# 0.03fF
C61 a_n563_n140# a_n1275_n140# 0.01fF
C62 a_1097_n194# a_919_n194# 0.10fF
C63 a_207_n194# a_1275_n194# 0.01fF
C64 a_861_n140# a_1453_n194# 0.01fF
C65 a_n385_n140# a_n1275_n140# 0.01fF
C66 a_327_n140# a_n29_n140# 0.03fF
C67 a_n563_n140# a_327_n140# 0.01fF
C68 a_n149_n194# a_1453_n194# 0.00fF
C69 a_n683_n194# a_207_n194# 0.01fF
C70 a_n385_n140# a_327_n140# 0.01fF
C71 a_29_n194# a_563_n194# 0.02fF
C72 a_29_n194# a_n1631_n140# 0.00fF
C73 a_861_n140# a_n741_n140# 0.01fF
C74 a_1395_n140# a_n207_n140# 0.01fF
C75 a_29_n194# a_919_n194# 0.01fF
C76 a_n1097_n140# a_n29_n140# 0.01fF
C77 a_n149_n194# a_207_n194# 0.03fF
C78 a_n919_n140# a_n1631_n140# 0.01fF
C79 a_149_n140# a_n29_n140# 0.06fF
C80 a_861_n140# a_683_n140# 0.06fF
C81 a_1039_n140# a_505_n140# 0.02fF
C82 a_n563_n140# a_n1097_n140# 0.02fF
C83 a_n1217_n194# a_207_n194# 0.01fF
C84 a_n563_n140# a_149_n140# 0.01fF
C85 a_1039_n140# a_1453_n194# 0.02fF
C86 a_n385_n140# a_n1097_n140# 0.01fF
C87 a_n207_n140# a_n919_n140# 0.01fF
C88 a_n385_n140# a_149_n140# 0.02fF
C89 a_n505_n194# a_n683_n194# 0.10fF
C90 a_1453_n194# a_1097_n194# 0.02fF
C91 a_n1395_n194# a_n861_n194# 0.02fF
C92 a_n327_n194# a_1275_n194# 0.01fF
C93 a_861_n140# a_327_n140# 0.02fF
C94 a_1217_n140# a_n29_n140# 0.01fF
C95 a_919_n194# a_563_n194# 0.03fF
C96 a_1217_n140# a_n385_n140# 0.01fF
C97 a_n683_n194# a_n1039_n194# 0.03fF
C98 a_n327_n194# a_n683_n194# 0.03fF
C99 a_n149_n194# a_n505_n194# 0.03fF
C100 a_385_n194# a_741_n194# 0.03fF
C101 a_n207_n140# a_n1631_n140# 0.01fF
C102 a_n505_n194# a_n1217_n194# 0.01fF
C103 a_1395_n140# a_505_n140# 0.01fF
C104 a_n861_n194# a_741_n194# 0.01fF
C105 a_1097_n194# a_207_n194# 0.01fF
C106 a_1395_n140# a_1453_n194# 0.06fF
C107 a_1039_n140# a_683_n140# 0.03fF
C108 a_385_n194# a_n861_n194# 0.01fF
C109 a_1453_n194# a_29_n194# 0.00fF
C110 a_861_n140# a_149_n140# 0.01fF
C111 a_n149_n194# a_n1039_n194# 0.01fF
C112 a_n327_n194# a_n149_n194# 0.10fF
C113 a_n1217_n194# a_n1039_n194# 0.10fF
C114 a_505_n140# a_n919_n140# 0.01fF
C115 a_n327_n194# a_n1217_n194# 0.01fF
C116 a_1039_n140# a_327_n140# 0.01fF
C117 a_1217_n140# a_861_n140# 0.03fF
C118 a_29_n194# a_207_n194# 0.10fF
C119 a_n505_n194# a_1097_n194# 0.01fF
C120 a_1453_n194# a_563_n194# 0.01fF
C121 a_1395_n140# a_683_n140# 0.01fF
C122 a_n1453_n140# a_n919_n140# 0.02fF
C123 a_n919_n140# a_n741_n140# 0.06fF
C124 a_1039_n140# a_149_n140# 0.01fF
C125 a_n207_n140# a_505_n140# 0.01fF
C126 a_n327_n194# a_1097_n194# 0.01fF
C127 a_1453_n194# a_919_n194# 0.01fF
C128 a_n1395_n194# a_n683_n194# 0.01fF
C129 a_1395_n140# a_327_n140# 0.01fF
C130 a_683_n140# a_n919_n140# 0.01fF
C131 a_207_n194# a_563_n194# 0.03fF
C132 a_n1275_n140# a_n919_n140# 0.03fF
C133 a_n505_n194# a_29_n194# 0.02fF
C134 a_741_n194# a_1275_n194# 0.02fF
C135 a_n1453_n140# a_n1631_n140# 0.06fF
C136 a_1217_n140# a_1039_n140# 0.06fF
C137 a_385_n194# a_1275_n194# 0.01fF
C138 a_n1631_n140# a_n741_n140# 0.01fF
C139 a_n919_n140# a_327_n140# 0.01fF
C140 a_n1453_n140# a_n207_n140# 0.01fF
C141 a_919_n194# a_207_n194# 0.01fF
C142 a_n149_n194# a_n1395_n194# 0.01fF
C143 a_n683_n194# a_741_n194# 0.01fF
C144 a_n207_n140# a_n741_n140# 0.02fF
C145 a_n1217_n194# a_n1395_n194# 0.10fF
C146 a_29_n194# a_n1039_n194# 0.01fF
C147 a_n683_n194# a_385_n194# 0.01fF
C148 a_n327_n194# a_29_n194# 0.03fF
C149 a_1395_n140# a_149_n140# 0.01fF
C150 a_n683_n194# a_n861_n194# 0.10fF
C151 a_n1275_n140# a_n1631_n140# 0.03fF
C152 a_n207_n140# a_683_n140# 0.01fF
C153 a_n505_n194# a_563_n194# 0.01fF
C154 a_n563_n140# a_n29_n140# 0.02fF
C155 a_n207_n140# a_n1275_n140# 0.01fF
C156 a_n385_n140# a_n29_n140# 0.03fF
C157 a_n149_n194# a_741_n194# 0.01fF
C158 a_1453_n194# a_505_n140# 0.01fF
C159 a_n919_n140# a_n1097_n140# 0.06fF
C160 a_n563_n140# a_n385_n140# 0.06fF
C161 a_n505_n194# a_n1631_n140# 0.01fF
C162 a_149_n140# a_n919_n140# 0.01fF
C163 a_1217_n140# a_1395_n140# 0.06fF
C164 a_n149_n194# a_385_n194# 0.02fF
C165 a_n1217_n194# a_385_n194# 0.01fF
C166 a_n207_n140# a_327_n140# 0.02fF
C167 a_n149_n194# a_n861_n194# 0.01fF
C168 a_n505_n194# a_919_n194# 0.01fF
C169 a_n1039_n194# a_563_n194# 0.01fF
C170 a_n327_n194# a_563_n194# 0.01fF
C171 a_n1217_n194# a_n861_n194# 0.03fF
C172 a_n1631_n140# a_n1039_n194# 0.01fF
C173 a_n327_n194# a_n1631_n140# 0.00fF
C174 a_505_n140# a_n741_n140# 0.01fF
C175 a_1453_n194# a_207_n194# 0.00fF
C176 a_n1631_n140# a_n1097_n140# 0.02fF
C177 a_n327_n194# a_919_n194# 0.01fF
C178 a_n207_n140# a_n1097_n140# 0.01fF
C179 a_505_n140# a_683_n140# 0.06fF
C180 a_149_n140# a_n207_n140# 0.03fF
C181 a_1097_n194# a_741_n194# 0.03fF
C182 a_861_n140# a_n29_n140# 0.01fF
C183 a_1453_n194# a_683_n140# 0.01fF
C184 a_861_n140# a_n563_n140# 0.01fF
C185 a_385_n194# a_1097_n194# 0.01fF
C186 a_861_n140# a_n385_n140# 0.01fF
C187 a_n1395_n194# a_29_n194# 0.01fF
C188 a_n1453_n140# a_n741_n140# 0.01fF
C189 a_505_n140# a_327_n140# 0.06fF
C190 a_1217_n140# a_n207_n140# 0.01fF
C191 a_1453_n194# a_327_n140# 0.01fF
C192 a_n1453_n140# a_n1275_n140# 0.06fF
C193 a_683_n140# a_n741_n140# 0.01fF
C194 a_29_n194# a_741_n194# 0.01fF
C195 a_n1275_n140# a_n741_n140# 0.02fF
C196 a_385_n194# a_29_n194# 0.03fF
C197 a_n149_n194# a_1275_n194# 0.01fF
C198 a_29_n194# a_n861_n194# 0.01fF
C199 a_1039_n140# a_n29_n140# 0.01fF
C200 a_1039_n140# a_n563_n140# 0.01fF
C201 a_505_n140# a_n1097_n140# 0.01fF
C202 a_n505_n194# a_207_n194# 0.01fF
C203 a_327_n140# a_n741_n140# 0.01fF
C204 a_149_n140# a_505_n140# 0.03fF
C205 a_1039_n140# a_n385_n140# 0.01fF
C206 a_n1395_n194# a_n1631_n140# 0.06fF
C207 a_n149_n194# a_n683_n194# 0.02fF
C208 a_1453_n194# a_149_n140# 0.01fF
C209 a_n1217_n194# a_n683_n194# 0.02fF
C210 a_683_n140# a_327_n140# 0.03fF
C211 a_741_n194# a_563_n194# 0.10fF
C212 a_n1275_n140# a_327_n140# 0.01fF
C213 a_207_n194# a_n1039_n194# 0.01fF
C214 a_1217_n140# a_505_n140# 0.01fF
C215 a_n327_n194# a_207_n194# 0.02fF
C216 a_385_n194# a_563_n194# 0.10fF
C217 a_n1453_n140# a_n1097_n140# 0.03fF
C218 a_1217_n140# a_1453_n194# 0.03fF
C219 a_n861_n194# a_563_n194# 0.01fF
C220 a_n1453_n140# a_149_n140# 0.01fF
C221 a_n1097_n140# a_n741_n140# 0.03fF
C222 a_1097_n194# a_1275_n194# 0.10fF
C223 a_n149_n194# a_n1217_n194# 0.01fF
C224 a_149_n140# a_n741_n140# 0.01fF
C225 a_1395_n140# a_n29_n140# 0.01fF
C226 a_919_n194# a_741_n194# 0.10fF
C227 a_n861_n194# a_n1631_n140# 0.01fF
C228 a_385_n194# a_919_n194# 0.02fF
C229 a_149_n140# a_683_n140# 0.02fF
C230 a_861_n140# a_1039_n140# 0.06fF
C231 a_n1275_n140# a_n1097_n140# 0.06fF
C232 a_149_n140# a_n1275_n140# 0.01fF
C233 a_n919_n140# a_n29_n140# 0.01fF
C234 a_n505_n194# a_n1039_n194# 0.02fF
C235 a_n563_n140# a_n919_n140# 0.03fF
C236 a_n327_n194# a_n505_n194# 0.10fF
C237 a_n385_n140# a_n919_n140# 0.02fF
C238 a_327_n140# a_n1097_n140# 0.01fF
C239 a_149_n140# a_327_n140# 0.06fF
C240 a_1217_n140# a_683_n140# 0.02fF
C241 a_29_n194# a_1275_n194# 0.01fF
C242 a_n149_n194# a_1097_n194# 0.01fF
C243 a_1395_n140# VSUBS 0.01fF
C244 a_1217_n140# VSUBS 0.01fF
C245 a_1039_n140# VSUBS 0.02fF
C246 a_861_n140# VSUBS 0.02fF
C247 a_683_n140# VSUBS 0.02fF
C248 a_505_n140# VSUBS 0.02fF
C249 a_327_n140# VSUBS 0.02fF
C250 a_149_n140# VSUBS 0.02fF
C251 a_n29_n140# VSUBS 0.02fF
C252 a_n207_n140# VSUBS 0.02fF
C253 a_n385_n140# VSUBS 0.02fF
C254 a_n563_n140# VSUBS 0.02fF
C255 a_n741_n140# VSUBS 0.02fF
C256 a_n919_n140# VSUBS 0.02fF
C257 a_n1097_n140# VSUBS 0.02fF
C258 a_n1275_n140# VSUBS 0.02fF
C259 a_n1453_n140# VSUBS 0.02fF
C260 a_1453_n194# VSUBS 0.31fF
C261 a_1275_n194# VSUBS 0.19fF
C262 a_1097_n194# VSUBS 0.20fF
C263 a_919_n194# VSUBS 0.21fF
C264 a_741_n194# VSUBS 0.22fF
C265 a_563_n194# VSUBS 0.23fF
C266 a_385_n194# VSUBS 0.23fF
C267 a_207_n194# VSUBS 0.24fF
C268 a_29_n194# VSUBS 0.24fF
C269 a_n149_n194# VSUBS 0.24fF
C270 a_n327_n194# VSUBS 0.24fF
C271 a_n505_n194# VSUBS 0.24fF
C272 a_n683_n194# VSUBS 0.24fF
C273 a_n861_n194# VSUBS 0.24fF
C274 a_n1039_n194# VSUBS 0.24fF
C275 a_n1217_n194# VSUBS 0.24fF
C276 a_n1395_n194# VSUBS 0.24fF
C277 a_n1631_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6RUDQZ a_n594_n195# a_n1008_n140# a_n652_n140# a_652_n195#
+ a_772_n140# a_n60_n195# a_n474_n140# a_n416_n195# a_474_n195# a_594_n140# a_n296_n140#
+ a_n238_n195# a_60_n140# a_296_n195# a_416_n140# a_n118_n140# a_118_n195# a_238_n140#
+ a_n772_n195# a_n830_n140# a_830_n195# VSUBS
X0 a_772_n140# a_652_n195# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n195# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n195# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n195# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n195# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_830_n195# a_830_n195# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n1008_n140# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n195# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n195# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n195# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n195# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n60_n195# a_830_n195# 0.01fF
C1 a_n238_n195# a_118_n195# 0.03fF
C2 a_830_n195# a_n296_n140# 0.01fF
C3 a_n1008_n140# a_n830_n140# 0.06fF
C4 a_416_n140# a_238_n140# 0.06fF
C5 a_n772_n195# a_n60_n195# 0.01fF
C6 a_60_n140# a_n474_n140# 0.02fF
C7 a_n652_n140# a_830_n195# 0.01fF
C8 a_n118_n140# a_60_n140# 0.06fF
C9 a_n1008_n140# a_238_n140# 0.01fF
C10 a_416_n140# a_n296_n140# 0.01fF
C11 a_238_n140# a_n830_n140# 0.01fF
C12 a_n1008_n140# a_n60_n195# 0.01fF
C13 a_772_n140# a_n474_n140# 0.01fF
C14 a_416_n140# a_n652_n140# 0.01fF
C15 a_772_n140# a_n118_n140# 0.01fF
C16 a_n1008_n140# a_n296_n140# 0.01fF
C17 a_n594_n195# a_830_n195# 0.00fF
C18 a_652_n195# a_830_n195# 0.06fF
C19 a_594_n140# a_n474_n140# 0.01fF
C20 a_594_n140# a_n118_n140# 0.01fF
C21 a_n830_n140# a_n296_n140# 0.02fF
C22 a_n1008_n140# a_n652_n140# 0.03fF
C23 a_474_n195# a_830_n195# 0.02fF
C24 a_n772_n195# a_n594_n195# 0.10fF
C25 a_n830_n140# a_n652_n140# 0.06fF
C26 a_60_n140# a_830_n195# 0.01fF
C27 a_n772_n195# a_652_n195# 0.01fF
C28 a_238_n140# a_n296_n140# 0.02fF
C29 a_296_n195# a_830_n195# 0.01fF
C30 a_474_n195# a_n772_n195# 0.01fF
C31 a_n416_n195# a_830_n195# 0.00fF
C32 a_238_n140# a_n652_n140# 0.01fF
C33 a_772_n140# a_830_n195# 0.06fF
C34 a_416_n140# a_60_n140# 0.03fF
C35 a_n1008_n140# a_n594_n195# 0.02fF
C36 a_n1008_n140# a_652_n195# 0.00fF
C37 a_n772_n195# a_296_n195# 0.01fF
C38 a_594_n140# a_830_n195# 0.03fF
C39 a_n772_n195# a_n416_n195# 0.03fF
C40 a_118_n195# a_830_n195# 0.01fF
C41 a_474_n195# a_n1008_n140# 0.00fF
C42 a_n652_n140# a_n296_n140# 0.03fF
C43 a_n238_n195# a_830_n195# 0.01fF
C44 a_n1008_n140# a_60_n140# 0.01fF
C45 a_416_n140# a_772_n140# 0.03fF
C46 a_n118_n140# a_n474_n140# 0.03fF
C47 a_n830_n140# a_60_n140# 0.01fF
C48 a_n772_n195# a_118_n195# 0.01fF
C49 a_n1008_n140# a_296_n195# 0.00fF
C50 a_n772_n195# a_n238_n195# 0.02fF
C51 a_594_n140# a_416_n140# 0.06fF
C52 a_n594_n195# a_n60_n195# 0.02fF
C53 a_652_n195# a_n60_n195# 0.01fF
C54 a_n1008_n140# a_n416_n195# 0.01fF
C55 a_238_n140# a_60_n140# 0.06fF
C56 a_772_n140# a_n830_n140# 0.01fF
C57 a_474_n195# a_n60_n195# 0.02fF
C58 a_594_n140# a_n1008_n140# 0.01fF
C59 a_n1008_n140# a_118_n195# 0.01fF
C60 a_n1008_n140# a_n238_n195# 0.01fF
C61 a_594_n140# a_n830_n140# 0.01fF
C62 a_60_n140# a_n296_n140# 0.03fF
C63 a_296_n195# a_n60_n195# 0.03fF
C64 a_772_n140# a_238_n140# 0.02fF
C65 a_n474_n140# a_830_n195# 0.01fF
C66 a_n118_n140# a_830_n195# 0.01fF
C67 a_n60_n195# a_n416_n195# 0.03fF
C68 a_n652_n140# a_60_n140# 0.01fF
C69 a_594_n140# a_238_n140# 0.03fF
C70 a_772_n140# a_n296_n140# 0.01fF
C71 a_416_n140# a_n474_n140# 0.01fF
C72 a_n60_n195# a_118_n195# 0.10fF
C73 a_652_n195# a_n594_n195# 0.01fF
C74 a_n238_n195# a_n60_n195# 0.10fF
C75 a_416_n140# a_n118_n140# 0.02fF
C76 a_772_n140# a_n652_n140# 0.01fF
C77 a_594_n140# a_n296_n140# 0.01fF
C78 a_474_n195# a_n594_n195# 0.01fF
C79 a_474_n195# a_652_n195# 0.10fF
C80 a_n1008_n140# a_n474_n140# 0.02fF
C81 a_594_n140# a_n652_n140# 0.01fF
C82 a_n1008_n140# a_n118_n140# 0.01fF
C83 a_n830_n140# a_n474_n140# 0.03fF
C84 a_n118_n140# a_n830_n140# 0.01fF
C85 a_296_n195# a_n594_n195# 0.01fF
C86 a_652_n195# a_296_n195# 0.03fF
C87 a_n594_n195# a_n416_n195# 0.10fF
C88 a_652_n195# a_n416_n195# 0.01fF
C89 a_n772_n195# a_830_n195# 0.00fF
C90 a_474_n195# a_296_n195# 0.10fF
C91 a_238_n140# a_n474_n140# 0.01fF
C92 a_n118_n140# a_238_n140# 0.03fF
C93 a_416_n140# a_830_n195# 0.02fF
C94 a_474_n195# a_n416_n195# 0.01fF
C95 a_n594_n195# a_118_n195# 0.01fF
C96 a_772_n140# a_60_n140# 0.01fF
C97 a_n238_n195# a_n594_n195# 0.03fF
C98 a_652_n195# a_118_n195# 0.02fF
C99 a_652_n195# a_n238_n195# 0.01fF
C100 a_n474_n140# a_n296_n140# 0.06fF
C101 a_296_n195# a_n416_n195# 0.01fF
C102 a_594_n140# a_60_n140# 0.02fF
C103 a_n118_n140# a_n296_n140# 0.06fF
C104 a_474_n195# a_118_n195# 0.03fF
C105 a_474_n195# a_n238_n195# 0.01fF
C106 a_n652_n140# a_n474_n140# 0.06fF
C107 a_n118_n140# a_n652_n140# 0.02fF
C108 a_n772_n195# a_n1008_n140# 0.06fF
C109 a_296_n195# a_118_n195# 0.10fF
C110 a_n238_n195# a_296_n195# 0.02fF
C111 a_594_n140# a_772_n140# 0.06fF
C112 a_n1008_n140# a_416_n140# 0.01fF
C113 a_n416_n195# a_118_n195# 0.02fF
C114 a_n238_n195# a_n416_n195# 0.10fF
C115 a_238_n140# a_830_n195# 0.01fF
C116 a_416_n140# a_n830_n140# 0.01fF
C117 a_772_n140# VSUBS 0.01fF
C118 a_594_n140# VSUBS 0.01fF
C119 a_416_n140# VSUBS 0.02fF
C120 a_238_n140# VSUBS 0.02fF
C121 a_60_n140# VSUBS 0.02fF
C122 a_n118_n140# VSUBS 0.02fF
C123 a_n296_n140# VSUBS 0.02fF
C124 a_n474_n140# VSUBS 0.02fF
C125 a_n652_n140# VSUBS 0.02fF
C126 a_n830_n140# VSUBS 0.02fF
C127 a_830_n195# VSUBS 0.31fF
C128 a_652_n195# VSUBS 0.19fF
C129 a_474_n195# VSUBS 0.20fF
C130 a_296_n195# VSUBS 0.21fF
C131 a_118_n195# VSUBS 0.22fF
C132 a_n60_n195# VSUBS 0.23fF
C133 a_n238_n195# VSUBS 0.23fF
C134 a_n416_n195# VSUBS 0.24fF
C135 a_n594_n195# VSUBS 0.24fF
C136 a_n772_n195# VSUBS 0.24fF
C137 a_n1008_n140# VSUBS 0.36fF
.ends

.subckt sky130_fd_pr__nfet_01v8_SD55Q9 a_352_607# a_644_607# a_174_607# a_60_607#
+ a_232_553# a_n232_n389# a_466_607# a_n524_n389# a_524_553# a_n410_n887# a_n702_n887#
+ a_n994_n887# a_644_n389# a_352_n389# a_60_n389# a_524_55# a_n60_55# a_n352_55# a_n232_n887#
+ a_n524_n887# a_174_n389# a_n352_n445# a_466_n389# a_n60_n445# a_n644_n445# a_644_n887#
+ a_352_n887# a_n118_n389# a_60_n887# a_174_n887# a_n352_n943# a_466_n887# a_n118_n887#
+ a_n60_n943# a_n644_n943# a_232_n445# a_n118_109# a_n410_109# a_758_n887# a_524_n445#
+ a_n232_109# a_n702_109# a_n644_55# a_n524_109# a_352_109# a_232_55# a_n352_553#
+ a_644_109# a_174_109# a_60_109# a_n644_553# a_n60_553# a_466_109# a_n410_607# a_524_n943#
+ a_232_n943# a_n410_n389# a_n118_607# a_n702_n389# a_n232_607# a_n702_607# a_n524_607#
+ VSUBS
X0 a_60_n389# a_n60_n445# a_n118_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_644_n887# a_524_n943# a_466_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_644_607# a_524_553# a_466_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n524_607# a_n644_553# a_n702_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_352_n389# a_232_n445# a_174_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_644_n389# a_524_n445# a_466_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n232_n887# a_n352_n943# a_n410_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_644_109# a_524_55# a_466_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n524_n887# a_n644_n943# a_n702_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_352_607# a_232_553# a_174_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n524_109# a_n644_55# a_n702_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n232_607# a_n352_553# a_n410_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n232_n389# a_n352_n445# a_n410_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n524_n389# a_n644_n445# a_n702_n389# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_60_607# a_n60_553# a_n118_607# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_352_109# a_232_55# a_174_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n232_109# a_n352_55# a_n410_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_60_n887# a_n60_n943# a_n118_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_758_n887# a_758_n887# a_758_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_60_109# a_n60_55# a_n118_109# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_n994_n887# a_n994_n887# a_n994_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_352_n887# a_232_n943# a_174_n887# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_n702_n887# a_n232_n887# 0.04fF
C1 a_524_55# a_524_n445# 0.15fF
C2 a_758_n887# a_n232_n887# 0.04fF
C3 a_n232_n887# a_644_n887# 0.02fF
C4 a_n644_55# a_n644_n943# 0.03fF
C5 a_60_109# a_n524_109# 0.03fF
C6 a_n702_n887# a_466_n887# 0.02fF
C7 a_352_n389# a_352_109# 0.01fF
C8 a_60_109# a_758_n887# 0.05fF
C9 a_352_n887# a_n232_n887# 0.03fF
C10 a_758_n887# a_466_n887# 0.12fF
C11 a_n702_607# a_n702_109# 0.01fF
C12 a_466_n887# a_644_n887# 0.13fF
C13 a_n644_n445# a_n352_n445# 0.04fF
C14 a_644_109# a_174_109# 0.04fF
C15 a_n994_n887# a_n60_n943# 0.01fF
C16 a_352_n887# a_466_n887# 0.25fF
C17 a_466_109# a_644_109# 0.13fF
C18 a_524_n943# a_n644_n943# 0.01fF
C19 a_n994_n887# a_n410_109# 0.08fF
C20 a_n410_n389# a_n410_109# 0.01fF
C21 a_644_607# a_60_607# 0.03fF
C22 a_n644_55# a_n994_n887# 0.05fF
C23 a_n524_607# a_n410_607# 0.25fF
C24 a_n352_n445# a_524_n445# 0.01fF
C25 a_n232_n389# a_60_n389# 0.07fF
C26 a_60_n389# a_466_n389# 0.05fF
C27 a_644_n389# a_n994_n887# 0.02fF
C28 a_n410_n389# a_644_n389# 0.02fF
C29 a_n60_553# a_n60_55# 0.15fF
C30 a_n60_n445# a_n352_n445# 0.04fF
C31 a_n118_n389# a_60_n389# 0.13fF
C32 a_466_109# a_466_n389# 0.01fF
C33 a_524_n943# a_n994_n887# 0.01fF
C34 a_n232_607# a_174_607# 0.05fF
C35 a_n644_n943# a_232_n943# 0.01fF
C36 a_60_109# a_n702_109# 0.03fF
C37 a_758_n887# a_352_n389# 0.08fF
C38 a_n702_n887# a_n702_n389# 0.01fF
C39 a_352_607# a_644_607# 0.07fF
C40 a_644_109# a_644_607# 0.01fF
C41 a_758_n887# a_n702_n389# 0.02fF
C42 a_n118_607# a_n232_607# 0.25fF
C43 a_n352_55# a_n994_n887# 0.02fF
C44 a_n118_109# a_n118_n887# 0.00fF
C45 a_352_n887# a_352_n389# 0.01fF
C46 a_n994_n887# a_n232_607# 0.06fF
C47 a_758_n887# a_n60_553# 0.01fF
C48 a_n994_n887# a_352_109# 0.03fF
C49 a_60_n887# a_n118_n887# 0.13fF
C50 a_466_n887# a_n232_n887# 0.03fF
C51 a_n524_607# a_n524_n389# 0.00fF
C52 a_n524_n887# a_n702_n887# 0.13fF
C53 a_n524_n887# a_n524_109# 0.00fF
C54 a_n994_n887# a_232_n943# 0.01fF
C55 a_n524_n887# a_758_n887# 0.03fF
C56 a_n524_607# a_60_607# 0.03fF
C57 a_n524_n887# a_644_n887# 0.02fF
C58 a_524_55# a_524_553# 0.15fF
C59 a_n702_607# a_n702_n389# 0.00fF
C60 a_758_n887# a_n644_n943# 0.01fF
C61 a_n410_109# a_174_109# 0.03fF
C62 a_n232_109# a_644_109# 0.02fF
C63 a_n524_n887# a_352_n887# 0.02fF
C64 a_n60_55# a_n994_n887# 0.01fF
C65 a_466_109# a_n410_109# 0.02fF
C66 a_n410_607# a_466_607# 0.02fF
C67 a_n60_553# a_n644_553# 0.02fF
C68 a_60_n887# a_174_n887# 0.25fF
C69 a_n702_109# a_n702_n389# 0.01fF
C70 a_n352_553# a_n352_n445# 0.03fF
C71 a_60_n389# a_644_n389# 0.03fF
C72 a_n352_553# a_232_553# 0.02fF
C73 a_758_n887# a_174_607# 0.06fF
C74 a_n644_55# a_n644_n445# 0.15fF
C75 a_174_n389# a_352_n389# 0.13fF
C76 a_n524_607# a_352_607# 0.02fF
C77 a_758_n887# a_n118_607# 0.04fF
C78 a_174_n389# a_n702_n389# 0.02fF
C79 a_n702_n887# a_n994_n887# 0.33fF
C80 a_n994_n887# a_n524_109# 0.12fF
C81 a_n352_553# a_n352_n943# 0.01fF
C82 a_232_n943# a_232_n445# 0.15fF
C83 a_758_n887# a_n994_n887# 0.07fF
C84 a_758_n887# a_n410_n389# 0.03fF
C85 a_n232_109# a_n232_n389# 0.01fF
C86 a_n644_n943# a_n644_553# 0.01fF
C87 a_n994_n887# a_644_n887# 0.02fF
C88 a_n60_n445# a_n60_n943# 0.15fF
C89 a_352_n887# a_n994_n887# 0.03fF
C90 a_232_553# a_524_553# 0.04fF
C91 a_n702_607# a_174_607# 0.02fF
C92 a_174_n887# a_n118_n887# 0.07fF
C93 a_352_109# a_174_109# 0.13fF
C94 a_60_n887# a_60_607# 0.00fF
C95 a_466_109# a_352_109# 0.25fF
C96 a_n702_607# a_n118_607# 0.03fF
C97 a_466_607# a_60_607# 0.05fF
C98 a_n524_n887# a_n232_n887# 0.07fF
C99 a_644_n389# a_644_607# 0.00fF
C100 a_n994_n887# a_n644_553# 0.05fF
C101 a_n702_607# a_n994_n887# 0.33fF
C102 a_524_n943# a_524_n445# 0.15fF
C103 a_n118_109# a_644_109# 0.03fF
C104 a_758_n887# a_232_n445# 0.02fF
C105 a_n524_n887# a_466_n887# 0.02fF
C106 a_n410_n887# a_60_n887# 0.04fF
C107 a_n994_n887# a_232_55# 0.01fF
C108 a_174_n389# a_174_607# 0.00fF
C109 a_n702_109# a_n994_n887# 0.33fF
C110 a_n232_109# a_n410_109# 0.13fF
C111 a_466_607# a_352_607# 0.25fF
C112 a_n232_607# a_644_607# 0.02fF
C113 a_174_n389# a_n994_n887# 0.04fF
C114 a_n410_n389# a_174_n389# 0.03fF
C115 a_352_n389# a_n702_n389# 0.02fF
C116 a_758_n887# a_60_n389# 0.05fF
C117 a_n994_n887# a_n232_n887# 0.06fF
C118 a_n524_109# a_174_109# 0.03fF
C119 a_758_n887# a_174_109# 0.06fF
C120 a_466_109# a_n524_109# 0.02fF
C121 a_466_109# a_758_n887# 0.12fF
C122 a_60_109# a_n994_n887# 0.04fF
C123 a_n410_n887# a_n118_n887# 0.07fF
C124 a_466_n887# a_n994_n887# 0.03fF
C125 a_n410_607# a_60_607# 0.04fF
C126 a_n118_109# a_n118_n389# 0.01fF
C127 a_758_n887# a_n644_n445# 0.01fF
C128 a_232_55# a_232_n445# 0.15fF
C129 a_466_n389# a_466_607# 0.00fF
C130 a_n60_n445# a_n60_55# 0.15fF
C131 a_n232_109# a_n232_607# 0.01fF
C132 a_n410_n887# a_n410_607# 0.00fF
C133 a_n232_109# a_352_109# 0.03fF
C134 a_n410_n887# a_174_n887# 0.03fF
C135 a_758_n887# a_524_n445# 0.06fF
C136 a_n410_607# a_352_607# 0.03fF
C137 a_758_n887# a_644_607# 0.33fF
C138 a_n644_n445# a_n644_553# 0.03fF
C139 a_644_n887# a_644_607# 0.00fF
C140 a_n524_607# a_n232_607# 0.07fF
C141 a_n352_55# a_n352_553# 0.15fF
C142 a_n60_n445# a_758_n887# 0.01fF
C143 a_n702_109# a_174_109# 0.02fF
C144 a_n118_109# a_n410_109# 0.07fF
C145 a_60_n389# a_174_n389# 0.25fF
C146 a_466_109# a_n702_109# 0.02fF
C147 a_352_n389# a_n994_n887# 0.03fF
C148 a_n410_n389# a_352_n389# 0.03fF
C149 a_n994_n887# a_n702_n389# 0.33fF
C150 a_174_n389# a_174_109# 0.01fF
C151 a_n410_n389# a_n702_n389# 0.07fF
C152 a_n118_n389# a_n118_n887# 0.01fF
C153 a_524_n943# a_524_553# 0.01fF
C154 a_n60_553# a_n994_n887# 0.01fF
C155 a_60_109# a_60_n389# 0.01fF
C156 a_n702_607# a_644_607# 0.01fF
C157 a_n232_109# a_n524_109# 0.07fF
C158 a_60_109# a_174_109# 0.25fF
C159 a_n232_109# a_758_n887# 0.04fF
C160 a_60_109# a_466_109# 0.05fF
C161 a_466_109# a_466_n887# 0.00fF
C162 a_n524_n887# a_n994_n887# 0.12fF
C163 a_352_607# a_60_607# 0.07fF
C164 a_n994_n887# a_n644_n943# 0.05fF
C165 a_n524_607# a_n524_109# 0.01fF
C166 a_n118_109# a_352_109# 0.04fF
C167 a_n524_607# a_758_n887# 0.03fF
C168 a_n118_607# a_174_607# 0.07fF
C169 a_n352_n943# a_n352_n445# 0.15fF
C170 a_758_n887# a_n352_553# 0.01fF
C171 a_n994_n887# a_174_607# 0.04fF
C172 a_466_607# a_n232_607# 0.03fF
C173 a_n232_n389# a_n524_n389# 0.07fF
C174 a_466_n389# a_n524_n389# 0.02fF
C175 a_n118_607# a_n994_n887# 0.05fF
C176 a_n410_607# a_n410_109# 0.01fF
C177 a_60_n389# a_352_n389# 0.07fF
C178 a_60_n389# a_n702_n389# 0.03fF
C179 a_n118_n389# a_n524_n389# 0.05fF
C180 a_n410_n389# a_n994_n887# 0.08fF
C181 a_n232_109# a_n702_109# 0.04fF
C182 a_n702_607# a_n524_607# 0.13fF
C183 a_758_n887# a_524_553# 0.05fF
C184 a_n352_553# a_n644_553# 0.04fF
C185 a_n644_55# a_524_55# 0.01fF
C186 a_n118_109# a_n524_109# 0.05fF
C187 a_n232_109# a_n232_n887# 0.00fF
C188 a_n118_109# a_758_n887# 0.04fF
C189 a_n702_n887# a_60_n887# 0.03fF
C190 a_60_n887# a_758_n887# 0.05fF
C191 a_60_109# a_n232_109# 0.07fF
C192 a_60_n887# a_644_n887# 0.03fF
C193 a_n410_607# a_n232_607# 0.13fF
C194 a_n994_n887# a_232_n445# 0.01fF
C195 a_758_n887# a_466_607# 0.12fF
C196 a_524_553# a_n644_553# 0.01fF
C197 a_524_n943# a_524_55# 0.03fF
C198 a_60_n887# a_352_n887# 0.07fF
C199 a_n644_n445# a_n644_n943# 0.15fF
C200 a_n352_55# a_524_55# 0.01fF
C201 a_n232_n389# a_466_n389# 0.03fF
C202 a_174_607# a_174_109# 0.01fF
C203 a_644_n389# a_n524_n389# 0.02fF
C204 a_n410_n887# a_n410_109# 0.00fF
C205 a_n232_n389# a_n118_n389# 0.25fF
C206 a_60_n389# a_n994_n887# 0.04fF
C207 a_n60_n445# a_n60_553# 0.03fF
C208 a_n352_n943# a_n60_n943# 0.04fF
C209 a_n410_n389# a_60_n389# 0.04fF
C210 a_n118_n389# a_466_n389# 0.03fF
C211 a_n702_n887# a_n118_n887# 0.03fF
C212 a_n118_109# a_n702_109# 0.03fF
C213 a_n994_n887# a_174_109# 0.04fF
C214 a_644_109# a_n410_109# 0.02fF
C215 a_758_n887# a_n118_n887# 0.04fF
C216 a_n702_607# a_466_607# 0.02fF
C217 a_466_109# a_n994_n887# 0.03fF
C218 a_n118_n887# a_644_n887# 0.03fF
C219 a_n644_n445# a_n994_n887# 0.05fF
C220 a_352_n887# a_n118_n887# 0.04fF
C221 a_n232_607# a_60_607# 0.07fF
C222 a_n60_55# a_524_55# 0.02fF
C223 a_644_109# a_644_n389# 0.01fF
C224 a_758_n887# a_n410_607# 0.03fF
C225 a_174_607# a_644_607# 0.04fF
C226 a_n352_55# a_n352_n445# 0.15fF
C227 a_n702_n887# a_174_n887# 0.02fF
C228 a_60_109# a_n118_109# 0.13fF
C229 a_524_n943# a_n352_n943# 0.01fF
C230 a_60_n887# a_n232_n887# 0.07fF
C231 a_174_n887# a_758_n887# 0.06fF
C232 a_n118_607# a_644_607# 0.03fF
C233 a_174_n887# a_644_n887# 0.04fF
C234 a_n994_n887# a_524_n445# 0.01fF
C235 a_n994_n887# a_644_607# 0.02fF
C236 a_60_109# a_60_n887# 0.00fF
C237 a_n352_55# a_n352_n943# 0.03fF
C238 a_174_n887# a_352_n887# 0.13fF
C239 a_60_n887# a_466_n887# 0.05fF
C240 a_758_n887# a_524_55# 0.05fF
C241 a_352_607# a_n232_607# 0.03fF
C242 a_n60_n445# a_n994_n887# 0.01fF
C243 a_466_n887# a_466_607# 0.00fF
C244 a_232_553# a_232_n943# 0.01fF
C245 a_352_607# a_352_109# 0.01fF
C246 a_n644_n445# a_232_n445# 0.01fF
C247 a_n232_n389# a_644_n389# 0.02fF
C248 a_644_109# a_352_109# 0.07fF
C249 a_n352_553# a_n60_553# 0.04fF
C250 a_466_n389# a_644_n389# 0.13fF
C251 a_n702_607# a_n410_607# 0.07fF
C252 a_n524_n887# a_n524_607# 0.00fF
C253 a_n352_n943# a_232_n943# 0.02fF
C254 a_n524_n389# a_n524_109# 0.01fF
C255 a_n118_n389# a_644_n389# 0.03fF
C256 a_758_n887# a_n524_n389# 0.03fF
C257 a_n232_n887# a_n118_n887# 0.25fF
C258 a_758_n887# a_60_607# 0.05fF
C259 a_n232_n389# a_n232_607# 0.00fF
C260 a_232_n445# a_524_n445# 0.04fF
C261 a_466_109# a_174_109# 0.07fF
C262 a_n232_109# a_n994_n887# 0.06fF
C263 a_n60_553# a_524_553# 0.02fF
C264 a_466_n887# a_n118_n887# 0.03fF
C265 a_n524_607# a_174_607# 0.03fF
C266 a_n60_n445# a_232_n445# 0.04fF
C267 a_524_55# a_232_55# 0.04fF
C268 a_758_n887# a_n352_n445# 0.01fF
C269 a_n410_n887# a_n702_n887# 0.07fF
C270 a_758_n887# a_232_553# 0.02fF
C271 a_174_n887# a_174_n389# 0.01fF
C272 a_n410_n887# a_758_n887# 0.03fF
C273 a_n524_607# a_n118_607# 0.05fF
C274 a_n410_n887# a_644_n887# 0.02fF
C275 a_174_n887# a_n232_n887# 0.05fF
C276 a_644_109# a_n524_109# 0.02fF
C277 a_n524_607# a_n994_n887# 0.12fF
C278 a_524_n943# a_n60_n943# 0.02fF
C279 a_758_n887# a_644_109# 0.33fF
C280 a_758_n887# a_352_607# 0.08fF
C281 a_758_n887# a_n352_n943# 0.01fF
C282 a_n410_n887# a_352_n887# 0.03fF
C283 a_644_109# a_644_n887# 0.00fF
C284 a_n702_607# a_60_607# 0.03fF
C285 a_n352_553# a_n994_n887# 0.02fF
C286 a_174_n887# a_466_n887# 0.07fF
C287 a_352_n887# a_352_607# 0.00fF
C288 a_n524_n887# a_60_n887# 0.03fF
C289 a_n644_n445# a_524_n445# 0.01fF
C290 a_232_553# a_n644_553# 0.01fF
C291 a_174_n389# a_n524_n389# 0.03fF
C292 a_n352_55# a_n644_55# 0.04fF
C293 a_n60_n445# a_n644_n445# 0.02fF
C294 a_n410_109# a_352_109# 0.03fF
C295 a_758_n887# a_n232_n389# 0.04fF
C296 a_n60_n943# a_232_n943# 0.04fF
C297 a_232_553# a_232_55# 0.15fF
C298 a_758_n887# a_466_n389# 0.12fF
C299 a_n702_607# a_352_607# 0.02fF
C300 a_n994_n887# a_524_553# 0.01fF
C301 a_n118_109# a_n118_607# 0.01fF
C302 a_758_n887# a_n118_n389# 0.04fF
C303 a_n118_109# a_n994_n887# 0.05fF
C304 a_n702_109# a_644_109# 0.01fF
C305 a_n60_55# a_n60_n943# 0.03fF
C306 a_466_607# a_174_607# 0.07fF
C307 a_60_109# a_60_607# 0.01fF
C308 a_n232_109# a_174_109# 0.05fF
C309 a_n60_n445# a_524_n445# 0.02fF
C310 a_n232_109# a_466_109# 0.03fF
C311 a_n118_607# a_466_607# 0.03fF
C312 a_60_n887# a_n994_n887# 0.04fF
C313 a_n524_n887# a_n118_n887# 0.05fF
C314 a_n410_n887# a_n232_n887# 0.13fF
C315 a_n644_55# a_n60_55# 0.02fF
C316 a_n994_n887# a_466_607# 0.03fF
C317 a_524_n943# a_232_n943# 0.04fF
C318 a_n410_n887# a_466_n887# 0.02fF
C319 a_758_n887# a_n60_n943# 0.01fF
C320 a_n410_109# a_n524_109# 0.25fF
C321 a_60_109# a_644_109# 0.03fF
C322 a_758_n887# a_n410_109# 0.03fF
C323 a_n524_n887# a_174_n887# 0.03fF
C324 a_758_n887# a_n644_55# 0.01fF
C325 a_n232_n389# a_174_n389# 0.05fF
C326 a_n118_607# a_n118_n887# 0.00fF
C327 a_466_n389# a_174_n389# 0.07fF
C328 a_352_n389# a_n524_n389# 0.02fF
C329 a_n702_n389# a_n524_n389# 0.13fF
C330 a_n352_55# a_n60_55# 0.04fF
C331 a_n994_n887# a_n118_n887# 0.05fF
C332 a_n232_n389# a_n232_n887# 0.01fF
C333 a_758_n887# a_644_n389# 0.33fF
C334 a_n118_n389# a_174_n389# 0.07fF
C335 a_n410_607# a_174_607# 0.03fF
C336 a_644_n389# a_644_n887# 0.01fF
C337 a_n118_607# a_n410_607# 0.07fF
C338 a_524_n943# a_758_n887# 0.05fF
C339 a_n524_607# a_644_607# 0.02fF
C340 a_174_n887# a_174_607# 0.00fF
C341 a_466_n887# a_466_n389# 0.01fF
C342 a_n410_607# a_n994_n887# 0.08fF
C343 a_n410_n389# a_n410_607# 0.00fF
C344 a_n644_55# a_n644_553# 0.15fF
C345 a_n118_109# a_174_109# 0.07fF
C346 a_n352_55# a_758_n887# 0.01fF
C347 a_60_n887# a_60_n389# 0.01fF
C348 a_n524_n887# a_n524_n389# 0.01fF
C349 a_n118_109# a_466_109# 0.03fF
C350 a_758_n887# a_n232_607# 0.04fF
C351 a_174_n887# a_n994_n887# 0.04fF
C352 a_n524_109# a_352_109# 0.02fF
C353 a_352_n389# a_352_607# 0.00fF
C354 a_n702_109# a_n410_109# 0.07fF
C355 a_758_n887# a_352_109# 0.08fF
C356 a_n644_55# a_232_55# 0.01fF
C357 a_n60_553# a_232_553# 0.04fF
C358 a_n994_n887# a_524_55# 0.01fF
C359 a_758_n887# a_232_n943# 0.02fF
C360 a_466_109# a_466_607# 0.01fF
C361 a_352_n887# a_352_109# 0.00fF
C362 a_524_553# a_524_n445# 0.03fF
C363 a_n524_n887# a_n410_n887# 0.25fF
C364 a_174_607# a_60_607# 0.25fF
C365 a_758_n887# a_n60_55# 0.01fF
C366 a_n232_n389# a_352_n389# 0.03fF
C367 a_60_109# a_n410_109# 0.04fF
C368 a_n702_607# a_n232_607# 0.04fF
C369 a_644_n389# a_174_n389# 0.04fF
C370 a_466_n389# a_352_n389# 0.25fF
C371 a_n118_607# a_60_607# 0.13fF
C372 a_n994_n887# a_n524_n389# 0.12fF
C373 a_n232_n389# a_n702_n389# 0.04fF
C374 a_n410_n389# a_n524_n389# 0.25fF
C375 a_466_n389# a_n702_n389# 0.02fF
C376 a_n352_55# a_232_55# 0.02fF
C377 a_n644_n943# a_n352_n943# 0.04fF
C378 a_n994_n887# a_60_607# 0.04fF
C379 a_n118_n389# a_352_n389# 0.04fF
C380 a_n118_n389# a_n702_n389# 0.03fF
C381 a_466_607# a_644_607# 0.13fF
C382 a_n702_n887# a_758_n887# 0.02fF
C383 a_758_n887# a_n524_109# 0.03fF
C384 a_n702_109# a_352_109# 0.02fF
C385 a_n702_n887# a_644_n887# 0.01fF
C386 a_352_607# a_174_607# 0.13fF
C387 a_n994_n887# a_n352_n445# 0.02fF
C388 a_232_55# a_232_n943# 0.03fF
C389 a_758_n887# a_644_n887# 0.33fF
C390 a_n994_n887# a_232_553# 0.01fF
C391 a_n410_n887# a_n410_n389# 0.01fF
C392 a_n410_n887# a_n994_n887# 0.08fF
C393 a_n702_n887# a_352_n887# 0.02fF
C394 a_n118_607# a_352_607# 0.04fF
C395 a_758_n887# a_352_n887# 0.08fF
C396 a_n232_n887# a_n232_607# 0.00fF
C397 a_352_n887# a_644_n887# 0.07fF
C398 a_n994_n887# a_352_607# 0.03fF
C399 a_644_109# a_n994_n887# 0.02fF
C400 a_n994_n887# a_n352_n943# 0.02fF
C401 a_174_n887# a_174_109# 0.00fF
C402 a_n232_109# a_n118_109# 0.25fF
C403 a_n60_55# a_232_55# 0.04fF
C404 a_60_109# a_352_109# 0.07fF
C405 a_n702_n887# a_n702_607# 0.00fF
C406 a_n352_553# a_524_553# 0.01fF
C407 a_758_n887# a_n644_553# 0.01fF
C408 a_n702_607# a_758_n887# 0.02fF
C409 a_n60_553# a_n60_n943# 0.01fF
C410 a_n352_n445# a_232_n445# 0.02fF
C411 a_758_n887# a_232_55# 0.02fF
C412 a_232_553# a_232_n445# 0.03fF
C413 a_n702_n887# a_n702_109# 0.00fF
C414 a_n702_109# a_n524_109# 0.13fF
C415 a_60_n389# a_n524_n389# 0.03fF
C416 a_n232_n389# a_n994_n887# 0.06fF
C417 a_n410_n389# a_n232_n389# 0.13fF
C418 a_644_n389# a_352_n389# 0.07fF
C419 a_466_n389# a_n994_n887# 0.03fF
C420 a_758_n887# a_n702_109# 0.02fF
C421 a_n410_607# a_644_607# 0.02fF
C422 a_n410_n389# a_466_n389# 0.02fF
C423 a_n118_n389# a_n118_607# 0.00fF
C424 a_644_n389# a_n702_n389# 0.01fF
C425 a_60_n389# a_60_607# 0.00fF
C426 a_n524_607# a_466_607# 0.02fF
C427 a_n410_n389# a_n118_n389# 0.07fF
C428 a_n644_n943# a_n60_n943# 0.02fF
C429 a_n118_n389# a_n994_n887# 0.05fF
C430 a_758_n887# a_174_n389# 0.06fF
C431 a_644_n887# VSUBS 0.01fF
C432 a_466_n887# VSUBS 0.01fF
C433 a_352_n887# VSUBS 0.01fF
C434 a_174_n887# VSUBS 0.01fF
C435 a_60_n887# VSUBS 0.01fF
C436 a_n118_n887# VSUBS 0.01fF
C437 a_n232_n887# VSUBS 0.01fF
C438 a_n410_n887# VSUBS 0.01fF
C439 a_n524_n887# VSUBS 0.01fF
C440 a_n702_n887# VSUBS 0.01fF
C441 a_524_n943# VSUBS 0.17fF
C442 a_232_n943# VSUBS 0.19fF
C443 a_n60_n943# VSUBS 0.20fF
C444 a_n352_n943# VSUBS 0.21fF
C445 a_n644_n943# VSUBS 0.22fF
C446 a_644_n389# VSUBS 0.01fF
C447 a_466_n389# VSUBS 0.01fF
C448 a_352_n389# VSUBS 0.01fF
C449 a_174_n389# VSUBS 0.01fF
C450 a_60_n389# VSUBS 0.01fF
C451 a_n118_n389# VSUBS 0.01fF
C452 a_n232_n389# VSUBS 0.01fF
C453 a_n410_n389# VSUBS 0.01fF
C454 a_n524_n389# VSUBS 0.01fF
C455 a_n702_n389# VSUBS 0.01fF
C456 a_524_n445# VSUBS 0.16fF
C457 a_232_n445# VSUBS 0.17fF
C458 a_n60_n445# VSUBS 0.18fF
C459 a_n352_n445# VSUBS 0.19fF
C460 a_n644_n445# VSUBS 0.20fF
C461 a_644_109# VSUBS 0.01fF
C462 a_466_109# VSUBS 0.01fF
C463 a_352_109# VSUBS 0.01fF
C464 a_174_109# VSUBS 0.01fF
C465 a_60_109# VSUBS 0.01fF
C466 a_n118_109# VSUBS 0.01fF
C467 a_n232_109# VSUBS 0.01fF
C468 a_n410_109# VSUBS 0.01fF
C469 a_n524_109# VSUBS 0.01fF
C470 a_n702_109# VSUBS 0.01fF
C471 a_524_55# VSUBS 0.17fF
C472 a_232_55# VSUBS 0.18fF
C473 a_n60_55# VSUBS 0.19fF
C474 a_n352_55# VSUBS 0.20fF
C475 a_n644_55# VSUBS 0.21fF
C476 a_644_607# VSUBS 0.02fF
C477 a_466_607# VSUBS 0.02fF
C478 a_352_607# VSUBS 0.02fF
C479 a_174_607# VSUBS 0.02fF
C480 a_60_607# VSUBS 0.02fF
C481 a_n118_607# VSUBS 0.02fF
C482 a_n232_607# VSUBS 0.02fF
C483 a_n410_607# VSUBS 0.02fF
C484 a_n524_607# VSUBS 0.02fF
C485 a_n702_607# VSUBS 0.02fF
C486 a_758_n887# VSUBS 1.42fF
C487 a_524_553# VSUBS 0.20fF
C488 a_232_553# VSUBS 0.22fF
C489 a_n60_553# VSUBS 0.23fF
C490 a_n352_553# VSUBS 0.24fF
C491 a_n644_553# VSUBS 0.25fF
C492 a_n994_n887# VSUBS 1.66fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EZNTQN a_n830_109# a_n652_n887# a_n652_109# a_n772_55#
+ a_118_553# a_594_n389# a_n772_n445# a_60_607# a_772_n887# a_n474_109# a_772_109#
+ a_n296_109# a_n772_553# a_n296_n389# a_594_109# a_n594_55# a_n594_553# a_n474_n887#
+ a_118_n943# a_60_n389# a_n594_n445# a_n60_55# a_n830_607# a_n772_n943# a_416_n389#
+ a_n652_607# a_594_n887# a_652_n445# a_n416_55# a_n474_607# a_772_607# a_n296_607#
+ a_n60_n445# a_594_607# a_n296_n887# a_n118_n389# a_652_553# a_60_n887# a_n238_55#
+ a_474_553# a_n594_n943# a_238_n389# a_n416_n445# a_416_n887# a_474_n445# a_296_553#
+ a_652_n943# a_n830_n389# a_652_55# a_n118_n887# a_n60_n943# a_n118_109# a_n238_n445#
+ a_416_109# a_n416_553# a_296_n445# a_238_109# a_474_55# a_n238_553# a_238_n887#
+ a_n416_n943# a_n1110_n1061# a_474_n943# a_n652_n389# a_n830_n887# a_60_109# a_772_n389#
+ a_n60_553# a_296_55# a_n118_607# a_n238_n943# a_416_607# a_296_n943# a_n474_n389#
+ a_118_n445# a_118_55# a_238_607#
X0 a_n652_109# a_n772_55# a_n830_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_60_n389# a_n60_n445# a_n118_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_594_n389# a_474_n445# a_416_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1110_n1061# a_n1110_n1061# a_772_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=3.248e+12p pd=2.704e+07u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n830_n887# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n474_n887# a_n594_n943# a_n652_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_594_607# a_474_553# a_416_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_109# a_n416_55# a_n474_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_416_n887# a_296_n943# a_238_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n474_607# a_n594_553# a_n652_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n296_n887# a_n416_n943# a_n474_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1110_n1061# a_n1110_n1061# a_772_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1110_n1061# a_n1110_n1061# a_772_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_238_607# a_118_553# a_60_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_238_n887# a_118_n943# a_60_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n830_n389# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n474_n389# a_n594_n445# a_n652_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_n830_607# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n118_607# a_n238_553# a_n296_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_594_109# a_474_55# a_416_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_416_n389# a_296_n445# a_238_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_772_n887# a_652_n943# a_594_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n474_109# a_n594_55# a_n652_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n296_n389# a_n416_n445# a_n474_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1110_n1061# a_n1110_n1061# a_772_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_238_109# a_118_55# a_60_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X26 a_238_n389# a_118_n445# a_60_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_607# a_296_553# a_238_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n830_109# a_n1110_n1061# a_n1110_n1061# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n118_109# a_n238_55# a_n296_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n118_n887# a_n238_n943# a_n296_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_60_607# a_n60_553# a_n118_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_772_n389# a_652_n445# a_594_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_772_607# a_652_553# a_594_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_n652_n887# a_n772_n943# a_n830_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_594_n887# a_474_n943# a_416_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_n652_607# a_n772_553# a_n830_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_60_n887# a_n60_n943# a_n118_n887# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_416_109# a_296_55# a_238_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n118_n389# a_n238_n445# a_n296_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_60_109# a_n60_55# a_n118_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X41 a_n296_607# a_n416_553# a_n474_607# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X42 a_772_109# a_652_55# a_594_109# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_n652_n389# a_n772_n445# a_n830_n389# a_n1110_n1061# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n296_n389# a_n296_607# 0.00fF
C1 a_118_n445# a_652_n445# 0.02fF
C2 a_474_n445# a_n60_n445# 0.02fF
C3 a_n238_55# a_652_55# 0.01fF
C4 a_594_n887# a_n652_n887# 0.01fF
C5 a_n772_553# a_652_553# 0.01fF
C6 a_594_n389# a_n118_n389# 0.01fF
C7 a_n60_55# a_n60_n445# 0.15fF
C8 a_n772_553# a_n416_553# 0.03fF
C9 a_n296_607# a_n296_n887# 0.00fF
C10 a_n238_n943# a_296_n943# 0.02fF
C11 a_n474_n389# a_772_n389# 0.01fF
C12 a_416_n389# a_594_n389# 0.06fF
C13 a_n238_553# a_n60_553# 0.10fF
C14 a_n830_n389# a_n830_109# 0.00fF
C15 a_118_n445# a_118_553# 0.03fF
C16 a_n772_n943# a_n60_n943# 0.01fF
C17 a_296_n943# a_118_n943# 0.10fF
C18 a_n416_55# a_n60_55# 0.03fF
C19 a_238_607# a_60_607# 0.06fF
C20 a_n296_n389# a_n118_n389# 0.06fF
C21 a_n474_n887# a_n474_607# 0.00fF
C22 a_n60_553# a_296_553# 0.03fF
C23 a_n830_607# a_n296_607# 0.02fF
C24 a_772_109# a_772_n389# 0.00fF
C25 a_416_n389# a_n296_n389# 0.01fF
C26 a_652_n943# a_652_55# 0.03fF
C27 a_296_55# a_296_553# 0.15fF
C28 a_n474_n887# a_n830_n887# 0.03fF
C29 a_416_109# a_238_109# 0.06fF
C30 a_60_n389# a_n118_n389# 0.06fF
C31 a_n416_55# a_n416_553# 0.15fF
C32 a_n474_n389# a_n474_607# 0.00fF
C33 a_n652_109# a_n652_n887# 0.00fF
C34 a_60_n887# a_238_n887# 0.06fF
C35 a_n60_n943# a_n594_n943# 0.02fF
C36 a_416_n389# a_60_n389# 0.03fF
C37 a_60_109# a_n474_109# 0.02fF
C38 a_652_553# a_n416_553# 0.01fF
C39 a_n772_n943# a_652_n943# 0.01fF
C40 a_n118_109# a_60_109# 0.06fF
C41 a_n118_607# a_60_607# 0.06fF
C42 a_238_607# a_n830_607# 0.01fF
C43 a_n238_n445# a_n238_55# 0.15fF
C44 a_296_n445# a_n594_n445# 0.01fF
C45 a_772_n887# a_n652_n887# 0.01fF
C46 a_416_607# a_416_n887# 0.00fF
C47 a_n474_n887# a_n474_109# 0.00fF
C48 a_n652_n887# a_n296_n887# 0.03fF
C49 a_n238_n943# a_n60_n943# 0.10fF
C50 a_n238_n943# a_n238_55# 0.03fF
C51 a_416_109# a_n296_109# 0.01fF
C52 a_60_n887# a_60_109# 0.00fF
C53 a_238_n389# a_n652_n389# 0.01fF
C54 a_n60_n943# a_118_n943# 0.10fF
C55 a_n594_n943# a_652_n943# 0.01fF
C56 a_n474_n389# a_n474_109# 0.00fF
C57 a_n416_n943# a_n772_n943# 0.03fF
C58 a_772_607# a_60_607# 0.01fF
C59 a_n238_553# a_n772_553# 0.02fF
C60 a_652_n445# a_652_55# 0.15fF
C61 a_238_109# a_n830_109# 0.01fF
C62 a_118_55# a_118_n445# 0.15fF
C63 a_n416_n445# a_n60_n445# 0.03fF
C64 a_n416_n445# a_474_n445# 0.01fF
C65 a_n594_n943# a_n594_n445# 0.15fF
C66 a_n118_607# a_n830_607# 0.01fF
C67 a_n474_n887# a_60_n887# 0.02fF
C68 a_n772_553# a_296_553# 0.01fF
C69 a_n238_n445# a_n594_n445# 0.03fF
C70 a_772_109# a_n474_109# 0.01fF
C71 a_594_607# a_594_n887# 0.00fF
C72 a_772_607# a_772_n887# 0.00fF
C73 a_238_607# a_238_n887# 0.00fF
C74 a_416_109# a_n652_109# 0.01fF
C75 a_772_109# a_n118_109# 0.01fF
C76 a_296_n943# a_n60_n943# 0.03fF
C77 a_n238_n943# a_652_n943# 0.01fF
C78 a_n416_n445# a_n416_55# 0.15fF
C79 a_296_n445# a_652_n445# 0.03fF
C80 a_n474_n389# a_n652_n389# 0.06fF
C81 a_118_n943# a_652_n943# 0.02fF
C82 a_n416_n943# a_n594_n943# 0.10fF
C83 a_416_n887# a_n830_n887# 0.01fF
C84 a_n830_n389# a_594_n389# 0.01fF
C85 a_n772_55# a_652_55# 0.01fF
C86 a_772_607# a_n830_607# 0.01fF
C87 a_n416_n445# a_n416_553# 0.03fF
C88 a_416_607# a_n474_607# 0.01fF
C89 a_n594_n445# a_n772_n445# 0.10fF
C90 a_n652_n887# a_238_n887# 0.01fF
C91 a_474_55# a_652_55# 0.10fF
C92 a_594_109# a_n474_109# 0.01fF
C93 a_n238_553# a_652_553# 0.01fF
C94 a_238_n389# a_n118_n389# 0.03fF
C95 a_594_607# a_594_n389# 0.00fF
C96 a_594_109# a_n118_109# 0.01fF
C97 a_238_607# a_238_n389# 0.00fF
C98 a_n238_553# a_n416_553# 0.10fF
C99 a_n830_109# a_n296_109# 0.02fF
C100 a_n830_n389# a_n296_n389# 0.02fF
C101 a_652_553# a_296_553# 0.03fF
C102 a_n238_n943# a_n416_n943# 0.10fF
C103 a_118_n445# a_n60_n445# 0.10fF
C104 a_474_n445# a_118_n445# 0.03fF
C105 a_416_n389# a_238_n389# 0.06fF
C106 a_296_n943# a_652_n943# 0.03fF
C107 a_n772_n943# a_n772_55# 0.03fF
C108 a_296_553# a_n416_553# 0.01fF
C109 a_n594_553# a_n594_n445# 0.03fF
C110 a_594_607# a_60_607# 0.02fF
C111 a_n416_n943# a_118_n943# 0.02fF
C112 a_n238_n445# a_652_n445# 0.01fF
C113 a_n118_n887# a_594_n887# 0.01fF
C114 a_n830_n389# a_60_n389# 0.01fF
C115 a_296_55# a_652_55# 0.03fF
C116 a_n772_n943# a_474_n943# 0.01fF
C117 a_n830_109# a_n652_109# 0.06fF
C118 a_n474_n389# a_n118_n389# 0.03fF
C119 a_n830_n389# a_n830_607# 0.00fF
C120 a_416_n389# a_n474_n389# 0.01fF
C121 a_n416_n943# a_296_n943# 0.01fF
C122 a_652_n445# a_n772_n445# 0.01fF
C123 a_n474_n887# a_n652_n887# 0.06fF
C124 a_296_55# a_296_n445# 0.15fF
C125 a_416_607# a_n652_607# 0.01fF
C126 a_60_n887# a_416_n887# 0.03fF
C127 a_238_109# a_n296_109# 0.02fF
C128 a_594_607# a_n830_607# 0.01fF
C129 a_n594_553# a_474_553# 0.01fF
C130 a_474_n943# a_n594_n943# 0.01fF
C131 a_118_55# a_652_55# 0.02fF
C132 a_n830_607# a_n830_109# 0.00fF
C133 a_118_n943# a_118_553# 0.01fF
C134 a_n60_n943# a_652_n943# 0.01fF
C135 a_n772_55# a_n772_n445# 0.15fF
C136 a_238_109# a_n652_109# 0.01fF
C137 a_n594_55# a_652_55# 0.01fF
C138 a_772_n389# a_n652_n389# 0.01fF
C139 a_n118_n887# a_772_n887# 0.01fF
C140 a_n238_n943# a_474_n943# 0.01fF
C141 a_416_109# a_60_109# 0.03fF
C142 a_n474_607# a_n474_109# 0.00fF
C143 a_416_607# a_n296_607# 0.01fF
C144 a_594_n887# a_594_n389# 0.00fF
C145 a_n594_553# a_118_553# 0.01fF
C146 a_n118_n887# a_n296_n887# 0.06fF
C147 a_474_n943# a_118_n943# 0.03fF
C148 a_n238_553# a_296_553# 0.02fF
C149 a_n652_607# a_n474_607# 0.06fF
C150 a_n416_n943# a_n60_n943# 0.03fF
C151 a_n416_n445# a_118_n445# 0.02fF
C152 a_416_n389# a_416_n887# 0.00fF
C153 a_n772_n943# a_n772_553# 0.01fF
C154 a_594_n887# a_772_n887# 0.06fF
C155 a_772_607# a_772_109# 0.00fF
C156 a_296_n943# a_474_n943# 0.10fF
C157 a_n830_n389# a_238_n389# 0.01fF
C158 a_416_607# a_238_607# 0.06fF
C159 a_n60_55# a_652_55# 0.01fF
C160 a_594_n887# a_n296_n887# 0.01fF
C161 a_60_n887# a_n830_n887# 0.01fF
C162 a_n60_553# a_n594_553# 0.02fF
C163 a_n416_55# a_652_55# 0.01fF
C164 a_n652_109# a_n296_109# 0.03fF
C165 a_416_607# a_416_n389# 0.00fF
C166 a_296_n445# a_n60_n445# 0.03fF
C167 a_n296_n389# a_n296_109# 0.00fF
C168 a_296_n445# a_474_n445# 0.10fF
C169 a_n594_n943# a_n594_55# 0.03fF
C170 a_n652_n887# a_416_n887# 0.01fF
C171 a_772_n389# a_n118_n389# 0.01fF
C172 a_652_553# a_652_55# 0.15fF
C173 a_n474_607# a_n296_607# 0.06fF
C174 a_416_109# a_772_109# 0.03fF
C175 a_n118_109# a_n474_109# 0.03fF
C176 a_296_55# a_296_n943# 0.03fF
C177 a_n296_n389# a_594_n389# 0.01fF
C178 a_n416_n943# a_652_n943# 0.01fF
C179 a_416_n389# a_772_n389# 0.03fF
C180 a_n830_109# a_60_109# 0.01fF
C181 a_n296_n887# a_n296_109# 0.00fF
C182 a_118_55# a_118_n943# 0.03fF
C183 a_n118_n887# a_238_n887# 0.03fF
C184 a_n830_n389# a_n474_n389# 0.03fF
C185 a_416_607# a_n118_607# 0.02fF
C186 a_238_109# a_238_n887# 0.00fF
C187 a_60_n389# a_594_n389# 0.02fF
C188 a_594_109# a_416_109# 0.06fF
C189 a_238_607# a_n474_607# 0.01fF
C190 a_n238_n445# a_n60_n445# 0.10fF
C191 a_n652_607# a_n652_n389# 0.00fF
C192 a_n772_55# a_n238_55# 0.02fF
C193 a_n238_n445# a_474_n445# 0.01fF
C194 a_652_n943# a_652_n445# 0.15fF
C195 a_60_607# a_60_n389# 0.00fF
C196 a_474_55# a_n238_55# 0.01fF
C197 a_n296_n389# a_n296_n887# 0.00fF
C198 a_n772_553# a_n772_n445# 0.03fF
C199 a_n296_n389# a_60_n389# 0.03fF
C200 a_n594_n445# a_652_n445# 0.01fF
C201 a_474_n943# a_n60_n943# 0.02fF
C202 a_594_n887# a_238_n887# 0.03fF
C203 a_772_n887# a_n296_n887# 0.01fF
C204 a_n594_553# a_n594_55# 0.15fF
C205 a_416_607# a_772_607# 0.03fF
C206 a_60_607# a_n830_607# 0.01fF
C207 a_416_109# a_416_n887# 0.00fF
C208 a_238_109# a_60_109# 0.06fF
C209 a_n60_553# a_n60_n943# 0.01fF
C210 a_n652_607# a_n296_607# 0.03fF
C211 a_772_109# a_n830_109# 0.01fF
C212 a_n772_n445# a_n60_n445# 0.01fF
C213 a_238_109# a_238_n389# 0.00fF
C214 a_474_n445# a_n772_n445# 0.01fF
C215 a_n594_553# a_n772_553# 0.10fF
C216 a_n474_n887# a_n118_n887# 0.03fF
C217 a_n118_607# a_n474_607# 0.03fF
C218 a_n652_n887# a_n830_n887# 0.06fF
C219 a_296_55# a_n238_55# 0.02fF
C220 a_416_607# a_416_109# 0.00fF
C221 a_772_607# a_772_n389# 0.00fF
C222 a_594_109# a_594_607# 0.00fF
C223 a_n118_109# a_n118_n389# 0.00fF
C224 a_474_n943# a_652_n943# 0.10fF
C225 a_594_109# a_n830_109# 0.01fF
C226 a_238_607# a_n652_607# 0.01fF
C227 a_n416_n445# a_296_n445# 0.01fF
C228 a_n474_n887# a_594_n887# 0.01fF
C229 a_n118_n389# a_n652_n389# 0.02fF
C230 a_772_607# a_n474_607# 0.01fF
C231 a_60_109# a_n296_109# 0.03fF
C232 a_118_55# a_n238_55# 0.03fF
C233 a_n594_553# a_652_553# 0.01fF
C234 a_772_109# a_238_109# 0.02fF
C235 a_416_n389# a_n652_n389# 0.01fF
C236 a_772_n887# a_238_n887# 0.02fF
C237 a_474_553# a_118_553# 0.03fF
C238 a_416_607# a_594_607# 0.06fF
C239 a_n594_553# a_n416_553# 0.10fF
C240 a_296_n445# a_296_553# 0.03fF
C241 a_n416_n943# a_474_n943# 0.01fF
C242 a_238_n887# a_n296_n887# 0.02fF
C243 a_n830_n389# a_772_n389# 0.01fF
C244 a_n652_607# a_n652_n887# 0.00fF
C245 a_594_n389# a_238_n389# 0.03fF
C246 a_n118_607# a_n118_109# 0.00fF
C247 a_474_55# a_474_553# 0.15fF
C248 a_n238_55# a_n594_55# 0.03fF
C249 a_238_607# a_n296_607# 0.02fF
C250 a_n652_109# a_60_109# 0.01fF
C251 a_n118_607# a_n652_607# 0.02fF
C252 a_60_607# a_60_109# 0.00fF
C253 a_n652_n887# a_n652_n389# 0.00fF
C254 a_474_n943# a_474_553# 0.01fF
C255 a_n238_n445# a_n416_n445# 0.10fF
C256 a_60_n887# a_n652_n887# 0.01fF
C257 a_594_109# a_238_109# 0.03fF
C258 a_n296_n389# a_238_n389# 0.02fF
C259 a_296_n445# a_118_n445# 0.10fF
C260 a_n60_553# a_474_553# 0.02fF
C261 a_n238_553# a_n238_n445# 0.03fF
C262 a_n60_n943# a_n60_n445# 0.15fF
C263 a_60_n389# a_60_109# 0.00fF
C264 a_n474_n389# a_594_n389# 0.01fF
C265 a_772_109# a_n296_109# 0.01fF
C266 a_n118_n887# a_416_n887# 0.02fF
C267 a_60_n389# a_238_n389# 0.06fF
C268 a_n830_n389# a_n830_n887# 0.00fF
C269 a_772_607# a_n652_607# 0.01fF
C270 a_n474_n887# a_772_n887# 0.01fF
C271 a_594_109# a_594_n887# 0.00fF
C272 a_n416_n445# a_n772_n445# 0.03fF
C273 a_n60_n943# a_n60_55# 0.03fF
C274 a_594_607# a_n474_607# 0.01fF
C275 a_416_n389# a_n118_n389# 0.02fF
C276 a_416_109# a_n474_109# 0.01fF
C277 a_n118_607# a_n296_607# 0.06fF
C278 a_n238_553# a_n238_n943# 0.01fF
C279 a_n238_55# a_n60_55# 0.10fF
C280 a_n594_55# a_n594_n445# 0.15fF
C281 a_474_55# a_n772_55# 0.01fF
C282 a_n474_n887# a_n296_n887# 0.06fF
C283 a_n416_55# a_n238_55# 0.10fF
C284 a_n474_n389# a_n296_n389# 0.06fF
C285 a_416_109# a_n118_109# 0.02fF
C286 a_n60_553# a_118_553# 0.10fF
C287 a_772_109# a_n652_109# 0.01fF
C288 a_474_55# a_474_n943# 0.03fF
C289 a_594_109# a_n296_109# 0.01fF
C290 a_n238_n445# a_118_n445# 0.03fF
C291 a_594_n887# a_416_n887# 0.06fF
C292 a_n830_109# a_n830_n887# 0.00fF
C293 a_n474_n389# a_60_n389# 0.02fF
C294 a_772_109# a_772_n887# 0.00fF
C295 a_n118_607# a_n118_n389# 0.00fF
C296 a_n238_553# a_n594_553# 0.03fF
C297 a_296_55# a_n772_55# 0.01fF
C298 a_594_109# a_594_n389# 0.00fF
C299 a_772_607# a_n296_607# 0.01fF
C300 a_n594_n445# a_n60_n445# 0.02fF
C301 a_474_n445# a_n594_n445# 0.01fF
C302 a_n118_607# a_238_607# 0.03fF
C303 a_296_55# a_474_55# 0.10fF
C304 a_n594_553# a_296_553# 0.01fF
C305 a_594_109# a_n652_109# 0.01fF
C306 a_118_n445# a_n772_n445# 0.01fF
C307 a_296_n943# a_296_553# 0.01fF
C308 a_118_n445# a_118_n943# 0.15fF
C309 a_652_553# a_652_n943# 0.01fF
C310 a_238_n887# a_238_n389# 0.00fF
C311 a_n772_553# a_474_553# 0.01fF
C312 a_n830_n389# a_n652_n389# 0.06fF
C313 a_594_607# a_n652_607# 0.01fF
C314 a_118_55# a_118_553# 0.15fF
C315 a_n830_109# a_n474_109# 0.03fF
C316 a_n118_n887# a_n830_n887# 0.01fF
C317 a_n474_n887# a_238_n887# 0.01fF
C318 a_772_607# a_238_607# 0.02fF
C319 a_n118_109# a_n830_109# 0.01fF
C320 a_118_55# a_n772_55# 0.01fF
C321 a_474_55# a_118_55# 0.03fF
C322 a_n416_n943# a_n416_55# 0.03fF
C323 a_474_553# a_474_n445# 0.03fF
C324 a_772_n887# a_416_n887# 0.03fF
C325 a_652_n445# a_n60_n445# 0.01fF
C326 a_n772_55# a_n594_55# 0.10fF
C327 a_474_n445# a_652_n445# 0.10fF
C328 a_416_607# a_60_607# 0.03fF
C329 a_416_109# a_416_n389# 0.00fF
C330 a_n416_n943# a_n416_553# 0.01fF
C331 a_n772_553# a_118_553# 0.01fF
C332 a_474_55# a_n594_55# 0.01fF
C333 a_772_n389# a_594_n389# 0.06fF
C334 a_416_n887# a_n296_n887# 0.01fF
C335 a_594_607# a_n296_607# 0.01fF
C336 a_594_n887# a_n830_n887# 0.01fF
C337 a_474_553# a_652_553# 0.10fF
C338 a_n772_553# a_n772_55# 0.15fF
C339 a_296_55# a_118_55# 0.10fF
C340 a_n118_607# a_772_607# 0.01fF
C341 a_n238_553# a_n238_55# 0.15fF
C342 a_474_553# a_n416_553# 0.01fF
C343 a_n118_109# a_n118_n887# 0.00fF
C344 a_238_109# a_n474_109# 0.01fF
C345 a_n830_n389# a_n118_n389# 0.01fF
C346 a_772_n389# a_n296_n389# 0.01fF
C347 a_652_553# a_652_n445# 0.03fF
C348 a_n118_109# a_238_109# 0.03fF
C349 a_772_n389# a_772_n887# 0.00fF
C350 a_n830_n389# a_416_n389# 0.01fF
C351 a_n474_n389# a_238_n389# 0.01fF
C352 a_296_55# a_n594_55# 0.01fF
C353 a_474_55# a_474_n445# 0.15fF
C354 a_416_607# a_n830_607# 0.01fF
C355 a_n60_553# a_n772_553# 0.01fF
C356 a_772_n389# a_60_n389# 0.01fF
C357 a_n772_55# a_n60_55# 0.01fF
C358 a_594_607# a_238_607# 0.03fF
C359 a_n118_n887# a_60_n887# 0.06fF
C360 a_772_109# a_60_109# 0.01fF
C361 a_n416_55# a_n772_55# 0.03fF
C362 a_474_55# a_n60_55# 0.02fF
C363 a_n474_n389# a_n474_n887# 0.00fF
C364 a_n416_n445# a_n594_n445# 0.10fF
C365 a_474_n943# a_474_n445# 0.15fF
C366 a_60_607# a_n474_607# 0.02fF
C367 a_652_553# a_118_553# 0.02fF
C368 a_n772_n943# a_n594_n943# 0.10fF
C369 a_474_55# a_n416_55# 0.01fF
C370 a_n238_n445# a_296_n445# 0.02fF
C371 a_n416_553# a_118_553# 0.02fF
C372 a_n60_553# a_n60_n445# 0.03fF
C373 a_238_n887# a_416_n887# 0.06fF
C374 a_n474_109# a_n296_109# 0.06fF
C375 a_n60_553# a_n60_55# 0.15fF
C376 a_118_55# a_n594_55# 0.01fF
C377 a_772_n887# a_n830_n887# 0.01fF
C378 a_n416_n943# a_n416_n445# 0.15fF
C379 a_594_109# a_60_109# 0.02fF
C380 a_n238_n943# a_n772_n943# 0.02fF
C381 a_60_n887# a_594_n887# 0.02fF
C382 a_n118_109# a_n296_109# 0.06fF
C383 a_296_55# a_n60_55# 0.03fF
C384 a_n830_n887# a_n296_n887# 0.02fF
C385 a_n118_607# a_594_607# 0.01fF
C386 a_296_n445# a_n772_n445# 0.01fF
C387 a_296_55# a_n416_55# 0.01fF
C388 a_n60_553# a_652_553# 0.01fF
C389 a_n772_n943# a_118_n943# 0.01fF
C390 a_n772_n943# a_n772_n445# 0.15fF
C391 a_n830_607# a_n474_607# 0.03fF
C392 a_n60_553# a_n416_553# 0.03fF
C393 a_n118_n887# a_n118_n389# 0.00fF
C394 a_n652_109# a_n474_109# 0.06fF
C395 a_n830_607# a_n830_n887# 0.00fF
C396 a_118_n445# a_n594_n445# 0.01fF
C397 a_n416_n445# a_652_n445# 0.01fF
C398 a_n238_553# a_474_553# 0.01fF
C399 a_n118_109# a_n652_109# 0.02fF
C400 a_238_607# a_238_109# 0.00fF
C401 a_n238_n943# a_n594_n943# 0.03fF
C402 a_594_n389# a_n652_n389# 0.01fF
C403 a_296_n943# a_296_n445# 0.15fF
C404 a_n652_607# a_60_607# 0.01fF
C405 a_n652_607# a_n652_109# 0.00fF
C406 a_772_607# a_594_607# 0.06fF
C407 a_474_553# a_296_553# 0.10fF
C408 a_n772_n943# a_296_n943# 0.01fF
C409 a_118_55# a_n60_55# 0.10fF
C410 a_n238_n943# a_n238_n445# 0.15fF
C411 a_n416_55# a_118_55# 0.02fF
C412 a_118_n943# a_n594_n943# 0.01fF
C413 a_n474_n887# a_416_n887# 0.01fF
C414 a_n296_607# a_n296_109# 0.00fF
C415 a_n652_109# a_n652_n389# 0.00fF
C416 a_n238_n445# a_n772_n445# 0.02fF
C417 a_60_607# a_60_n887# 0.00fF
C418 a_n118_n887# a_n652_n887# 0.02fF
C419 a_594_109# a_772_109# 0.06fF
C420 a_n296_n389# a_n652_n389# 0.03fF
C421 a_n594_55# a_n60_55# 0.02fF
C422 a_n118_607# a_n118_n887# 0.00fF
C423 a_n416_55# a_n594_55# 0.10fF
C424 a_772_n389# a_238_n389# 0.02fF
C425 a_60_n887# a_772_n887# 0.01fF
C426 a_n238_553# a_118_553# 0.03fF
C427 a_n594_553# a_n594_n943# 0.01fF
C428 a_n238_n943# a_118_n943# 0.03fF
C429 a_238_n887# a_n830_n887# 0.01fF
C430 a_416_109# a_n830_109# 0.01fF
C431 a_296_n943# a_n594_n943# 0.01fF
C432 a_60_n389# a_n652_n389# 0.01fF
C433 a_60_607# a_n296_607# 0.03fF
C434 a_60_n887# a_n296_n887# 0.03fF
C435 a_296_553# a_118_553# 0.10fF
C436 a_n652_607# a_n830_607# 0.06fF
C437 a_60_n389# a_60_n887# 0.00fF
C438 a_772_n887# a_n1110_n1061# 0.10fF
C439 a_594_n887# a_n1110_n1061# 0.06fF
C440 a_416_n887# a_n1110_n1061# 0.05fF
C441 a_238_n887# a_n1110_n1061# 0.05fF
C442 a_60_n887# a_n1110_n1061# 0.04fF
C443 a_n118_n887# a_n1110_n1061# 0.04fF
C444 a_n296_n887# a_n1110_n1061# 0.05fF
C445 a_n474_n887# a_n1110_n1061# 0.05fF
C446 a_n652_n887# a_n1110_n1061# 0.06fF
C447 a_n830_n887# a_n1110_n1061# 0.10fF
C448 a_652_n943# a_n1110_n1061# 0.27fF
C449 a_474_n943# a_n1110_n1061# 0.24fF
C450 a_296_n943# a_n1110_n1061# 0.24fF
C451 a_118_n943# a_n1110_n1061# 0.24fF
C452 a_n60_n943# a_n1110_n1061# 0.25fF
C453 a_n238_n943# a_n1110_n1061# 0.26fF
C454 a_n416_n943# a_n1110_n1061# 0.26fF
C455 a_n594_n943# a_n1110_n1061# 0.27fF
C456 a_n772_n943# a_n1110_n1061# 0.32fF
C457 a_772_n389# a_n1110_n1061# 0.10fF
C458 a_594_n389# a_n1110_n1061# 0.06fF
C459 a_416_n389# a_n1110_n1061# 0.05fF
C460 a_238_n389# a_n1110_n1061# 0.04fF
C461 a_60_n389# a_n1110_n1061# 0.04fF
C462 a_n118_n389# a_n1110_n1061# 0.04fF
C463 a_n296_n389# a_n1110_n1061# 0.04fF
C464 a_n474_n389# a_n1110_n1061# 0.05fF
C465 a_n652_n389# a_n1110_n1061# 0.06fF
C466 a_n830_n389# a_n1110_n1061# 0.10fF
C467 a_652_n445# a_n1110_n1061# 0.22fF
C468 a_474_n445# a_n1110_n1061# 0.19fF
C469 a_296_n445# a_n1110_n1061# 0.19fF
C470 a_118_n445# a_n1110_n1061# 0.19fF
C471 a_n60_n445# a_n1110_n1061# 0.20fF
C472 a_n238_n445# a_n1110_n1061# 0.21fF
C473 a_n416_n445# a_n1110_n1061# 0.21fF
C474 a_n594_n445# a_n1110_n1061# 0.22fF
C475 a_n772_n445# a_n1110_n1061# 0.27fF
C476 a_772_109# a_n1110_n1061# 0.10fF
C477 a_594_109# a_n1110_n1061# 0.06fF
C478 a_416_109# a_n1110_n1061# 0.05fF
C479 a_238_109# a_n1110_n1061# 0.05fF
C480 a_60_109# a_n1110_n1061# 0.04fF
C481 a_n118_109# a_n1110_n1061# 0.04fF
C482 a_n296_109# a_n1110_n1061# 0.05fF
C483 a_n474_109# a_n1110_n1061# 0.05fF
C484 a_n652_109# a_n1110_n1061# 0.06fF
C485 a_n830_109# a_n1110_n1061# 0.10fF
C486 a_652_55# a_n1110_n1061# 0.23fF
C487 a_474_55# a_n1110_n1061# 0.20fF
C488 a_296_55# a_n1110_n1061# 0.20fF
C489 a_118_55# a_n1110_n1061# 0.21fF
C490 a_n60_55# a_n1110_n1061# 0.21fF
C491 a_n238_55# a_n1110_n1061# 0.22fF
C492 a_n416_55# a_n1110_n1061# 0.23fF
C493 a_n594_55# a_n1110_n1061# 0.24fF
C494 a_n772_55# a_n1110_n1061# 0.28fF
C495 a_772_607# a_n1110_n1061# 0.10fF
C496 a_594_607# a_n1110_n1061# 0.06fF
C497 a_416_607# a_n1110_n1061# 0.06fF
C498 a_238_607# a_n1110_n1061# 0.05fF
C499 a_60_607# a_n1110_n1061# 0.05fF
C500 a_n118_607# a_n1110_n1061# 0.05fF
C501 a_n296_607# a_n1110_n1061# 0.05fF
C502 a_n474_607# a_n1110_n1061# 0.06fF
C503 a_n652_607# a_n1110_n1061# 0.07fF
C504 a_n830_607# a_n1110_n1061# 0.10fF
C505 a_652_553# a_n1110_n1061# 0.30fF
C506 a_474_553# a_n1110_n1061# 0.27fF
C507 a_296_553# a_n1110_n1061# 0.27fF
C508 a_118_553# a_n1110_n1061# 0.27fF
C509 a_n60_553# a_n1110_n1061# 0.28fF
C510 a_n238_553# a_n1110_n1061# 0.29fF
C511 a_n416_553# a_n1110_n1061# 0.29fF
C512 a_n594_553# a_n1110_n1061# 0.30fF
C513 a_n772_553# a_n1110_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_JJWXCM a_n207_n140# a_29_n205# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n205# a_563_n205# a_n741_n140# a_n327_n205# a_n563_n140# a_385_n205#
+ w_n777_n241# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n327_n205# a_n385_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_563_n205# a_563_n205# a_505_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n29_n140# a_n149_n205# a_n207_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_505_n140# a_385_n205# a_327_n140# w_n777_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n385_n140# a_n741_n140# 0.03fF
C1 a_n207_n140# a_563_n205# 0.01fF
C2 a_n563_n140# a_n29_n140# 0.04fF
C3 a_563_n205# a_207_n205# 0.02fF
C4 a_n149_n205# a_n327_n205# 0.10fF
C5 a_n385_n140# w_n777_n241# 0.02fF
C6 a_149_n140# a_n741_n140# 0.01fF
C7 a_n327_n205# a_n505_n205# 0.10fF
C8 a_385_n205# a_n741_n140# 0.01fF
C9 a_563_n205# a_n327_n205# 0.01fF
C10 a_n385_n140# a_505_n140# 0.02fF
C11 a_149_n140# w_n777_n241# 0.02fF
C12 a_385_n205# w_n777_n241# 0.14fF
C13 a_327_n140# a_n29_n140# 0.06fF
C14 a_327_n140# a_n563_n140# 0.02fF
C15 a_149_n140# a_505_n140# 0.06fF
C16 a_n385_n140# a_563_n205# 0.01fF
C17 a_29_n205# a_207_n205# 0.10fF
C18 a_385_n205# a_n149_n205# 0.02fF
C19 a_n207_n140# a_n29_n140# 0.13fF
C20 a_n563_n140# a_n207_n140# 0.06fF
C21 a_149_n140# a_563_n205# 0.02fF
C22 a_n741_n140# w_n777_n241# 0.33fF
C23 a_385_n205# a_n505_n205# 0.01fF
C24 a_29_n205# a_n327_n205# 0.03fF
C25 a_385_n205# a_563_n205# 0.07fF
C26 a_n741_n140# a_505_n140# 0.01fF
C27 a_n149_n205# a_n741_n140# 0.01fF
C28 w_n777_n241# a_505_n140# 0.02fF
C29 a_n741_n140# a_n505_n205# 0.07fF
C30 a_n149_n205# w_n777_n241# 0.17fF
C31 a_327_n140# a_n207_n140# 0.04fF
C32 a_n741_n140# a_563_n205# 0.01fF
C33 w_n777_n241# a_n505_n205# 0.19fF
C34 a_n385_n140# a_n29_n140# 0.06fF
C35 a_n385_n140# a_n563_n140# 0.13fF
C36 w_n777_n241# a_563_n205# 0.28fF
C37 a_385_n205# a_29_n205# 0.03fF
C38 a_149_n140# a_n29_n140# 0.13fF
C39 a_149_n140# a_n563_n140# 0.03fF
C40 a_n149_n205# a_n505_n205# 0.03fF
C41 a_505_n140# a_563_n205# 0.06fF
C42 a_n149_n205# a_563_n205# 0.01fF
C43 a_563_n205# a_n505_n205# 0.01fF
C44 a_29_n205# a_n741_n140# 0.01fF
C45 a_327_n140# a_n385_n140# 0.03fF
C46 a_n327_n205# a_207_n205# 0.02fF
C47 a_29_n205# w_n777_n241# 0.16fF
C48 a_n741_n140# a_n29_n140# 0.01fF
C49 a_n563_n140# a_n741_n140# 0.06fF
C50 a_149_n140# a_327_n140# 0.13fF
C51 a_n385_n140# a_n207_n140# 0.13fF
C52 w_n777_n241# a_n29_n140# 0.02fF
C53 a_n563_n140# w_n777_n241# 0.02fF
C54 a_29_n205# a_n149_n205# 0.10fF
C55 a_149_n140# a_n207_n140# 0.06fF
C56 a_29_n205# a_n505_n205# 0.02fF
C57 a_505_n140# a_n29_n140# 0.04fF
C58 a_n563_n140# a_505_n140# 0.02fF
C59 a_29_n205# a_563_n205# 0.01fF
C60 a_385_n205# a_207_n205# 0.10fF
C61 a_327_n140# a_n741_n140# 0.01fF
C62 a_563_n205# a_n29_n140# 0.01fF
C63 a_n563_n140# a_563_n205# 0.01fF
C64 a_327_n140# w_n777_n241# 0.02fF
C65 a_385_n205# a_n327_n205# 0.01fF
C66 a_n741_n140# a_n207_n140# 0.02fF
C67 a_n741_n140# a_207_n205# 0.01fF
C68 a_327_n140# a_505_n140# 0.13fF
C69 a_149_n140# a_n385_n140# 0.04fF
C70 w_n777_n241# a_n207_n140# 0.02fF
C71 w_n777_n241# a_207_n205# 0.15fF
C72 a_n741_n140# a_n327_n205# 0.02fF
C73 a_n207_n140# a_505_n140# 0.03fF
C74 a_327_n140# a_563_n205# 0.03fF
C75 w_n777_n241# a_n327_n205# 0.18fF
C76 a_n149_n205# a_207_n205# 0.03fF
C77 a_207_n205# a_n505_n205# 0.01fF
C78 w_n777_n241# VSUBS 2.25fF
.ends

.subckt sky130_fd_pr__nfet_01v8_LJREPQ a_n149_n195# a_n207_n140# a_207_n195# a_n29_n140#
+ a_149_n140# a_29_n195# a_n385_n140# VSUBS
X0 a_n29_n140# a_n149_n195# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_207_n195# a_207_n195# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n195# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X3 a_n207_n140# a_n385_n140# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_29_n195# a_207_n195# 0.06fF
C1 a_n29_n140# a_n207_n140# 0.06fF
C2 a_n385_n140# a_n29_n140# 0.03fF
C3 a_207_n195# a_149_n140# 0.06fF
C4 a_29_n195# a_n385_n140# 0.02fF
C5 a_n149_n195# a_29_n195# 0.10fF
C6 a_207_n195# a_n207_n140# 0.02fF
C7 a_n207_n140# a_149_n140# 0.03fF
C8 a_n385_n140# a_207_n195# 0.03fF
C9 a_n149_n195# a_207_n195# 0.02fF
C10 a_n385_n140# a_149_n140# 0.02fF
C11 a_n29_n140# a_207_n195# 0.03fF
C12 a_n385_n140# a_n207_n140# 0.06fF
C13 a_n29_n140# a_149_n140# 0.06fF
C14 a_n149_n195# a_n385_n140# 0.06fF
C15 a_149_n140# VSUBS 0.01fF
C16 a_n29_n140# VSUBS 0.01fF
C17 a_n207_n140# VSUBS 0.02fF
C18 a_207_n195# VSUBS 0.31fF
C19 a_29_n195# VSUBS 0.19fF
C20 a_n149_n195# VSUBS 0.20fF
C21 a_n385_n140# VSUBS 0.33fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SAWXCM a_n207_n140# a_29_n204# a_327_n140# a_n29_n140#
+ a_149_n140# a_n505_n204# a_563_n204# a_n741_n140# a_n327_n204# a_385_n204# a_n563_n140#
+ a_n149_n204# w_n777_n240# a_n385_n140# a_207_n204# a_505_n140# VSUBS
X0 a_505_n140# a_385_n204# a_327_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n385_n140# a_n505_n204# a_n563_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_327_n140# a_207_n204# a_149_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_149_n140# a_29_n204# a_n29_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n204# a_n385_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_563_n204# a_563_n204# a_505_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n29_n140# a_n149_n204# a_n207_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_n563_n140# a_n741_n140# a_n741_n140# w_n777_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_385_n204# a_n505_n204# 0.01fF
C1 a_149_n140# a_n563_n140# 0.03fF
C2 a_563_n204# a_207_n204# 0.02fF
C3 a_327_n140# w_n777_n240# 0.02fF
C4 a_327_n140# a_505_n140# 0.13fF
C5 a_n29_n140# a_n741_n140# 0.01fF
C6 a_149_n140# a_563_n204# 0.02fF
C7 w_n777_n240# a_n505_n204# 0.19fF
C8 a_n207_n140# w_n777_n240# 0.02fF
C9 a_n207_n140# a_505_n140# 0.03fF
C10 a_327_n140# a_n385_n140# 0.03fF
C11 a_n741_n140# a_385_n204# 0.01fF
C12 a_n327_n204# a_n505_n204# 0.10fF
C13 a_n29_n140# w_n777_n240# 0.02fF
C14 a_n29_n140# a_505_n140# 0.04fF
C15 a_n149_n204# a_n505_n204# 0.03fF
C16 a_n207_n140# a_n385_n140# 0.13fF
C17 a_n741_n140# w_n777_n240# 0.33fF
C18 a_505_n140# a_n741_n140# 0.01fF
C19 a_327_n140# a_n563_n140# 0.02fF
C20 a_29_n204# a_n505_n204# 0.02fF
C21 a_n29_n140# a_n385_n140# 0.06fF
C22 a_327_n140# a_563_n204# 0.03fF
C23 w_n777_n240# a_385_n204# 0.14fF
C24 a_n741_n140# a_n385_n140# 0.03fF
C25 a_n327_n204# a_n741_n140# 0.02fF
C26 a_n207_n140# a_n563_n140# 0.06fF
C27 a_149_n140# a_327_n140# 0.13fF
C28 a_207_n204# a_n505_n204# 0.01fF
C29 a_563_n204# a_n505_n204# 0.01fF
C30 a_n149_n204# a_n741_n140# 0.01fF
C31 a_505_n140# w_n777_n240# 0.02fF
C32 a_n207_n140# a_563_n204# 0.01fF
C33 a_29_n204# a_n741_n140# 0.01fF
C34 a_n327_n204# a_385_n204# 0.01fF
C35 a_n29_n140# a_n563_n140# 0.04fF
C36 a_149_n140# a_n207_n140# 0.06fF
C37 a_n741_n140# a_n563_n140# 0.06fF
C38 a_n149_n204# a_385_n204# 0.02fF
C39 a_n29_n140# a_563_n204# 0.01fF
C40 w_n777_n240# a_n385_n140# 0.02fF
C41 a_505_n140# a_n385_n140# 0.02fF
C42 a_n327_n204# w_n777_n240# 0.18fF
C43 a_n741_n140# a_207_n204# 0.01fF
C44 a_563_n204# a_n741_n140# 0.01fF
C45 a_29_n204# a_385_n204# 0.03fF
C46 a_149_n140# a_n29_n140# 0.13fF
C47 a_n149_n204# w_n777_n240# 0.17fF
C48 a_149_n140# a_n741_n140# 0.01fF
C49 a_29_n204# w_n777_n240# 0.16fF
C50 a_385_n204# a_207_n204# 0.10fF
C51 a_563_n204# a_385_n204# 0.07fF
C52 w_n777_n240# a_n563_n140# 0.02fF
C53 a_505_n140# a_n563_n140# 0.02fF
C54 a_n149_n204# a_n327_n204# 0.10fF
C55 w_n777_n240# a_207_n204# 0.15fF
C56 a_563_n204# w_n777_n240# 0.28fF
C57 a_563_n204# a_505_n140# 0.06fF
C58 a_n207_n140# a_327_n140# 0.04fF
C59 a_n327_n204# a_29_n204# 0.03fF
C60 a_n385_n140# a_n563_n140# 0.13fF
C61 a_149_n140# w_n777_n240# 0.02fF
C62 a_149_n140# a_505_n140# 0.06fF
C63 a_n149_n204# a_29_n204# 0.10fF
C64 a_n29_n140# a_327_n140# 0.06fF
C65 a_563_n204# a_n385_n140# 0.01fF
C66 a_n327_n204# a_207_n204# 0.02fF
C67 a_n327_n204# a_563_n204# 0.01fF
C68 a_327_n140# a_n741_n140# 0.01fF
C69 a_149_n140# a_n385_n140# 0.04fF
C70 a_n149_n204# a_207_n204# 0.03fF
C71 a_n149_n204# a_563_n204# 0.01fF
C72 a_n741_n140# a_n505_n204# 0.07fF
C73 a_n207_n140# a_n29_n140# 0.13fF
C74 a_29_n204# a_207_n204# 0.10fF
C75 a_563_n204# a_29_n204# 0.01fF
C76 a_n207_n140# a_n741_n140# 0.02fF
C77 a_563_n204# a_n563_n140# 0.01fF
C78 w_n777_n240# VSUBS 2.24fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_28TRYY a_385_553# a_n1097_109# a_n149_55# a_919_n445#
+ a_29_55# a_n29_n389# a_n207_n887# a_1097_n943# a_n1555_n1061# a_n1097_n389# a_n327_n445#
+ a_149_n389# a_n207_109# a_385_n445# a_563_55# a_n505_n943# a_n1275_n887# a_327_n887#
+ a_505_109# a_563_n943# a_n505_553# a_n741_n389# a_327_109# a_n327_553# a_n1275_607#
+ a_n1217_55# a_861_n389# a_149_109# a_n149_553# a_n1097_607# a_385_55# a_n149_n445#
+ a_n29_109# a_919_n943# a_n29_n887# a_n327_n943# a_n1097_n887# a_149_n887# a_n207_607#
+ a_207_n445# a_385_n943# a_n563_n389# a_1097_553# a_n1039_55# a_1217_n389# a_207_55#
+ a_n1217_n445# a_505_607# a_n741_n887# a_327_607# a_n861_n445# a_683_n389# a_n861_55#
+ a_149_607# a_861_n887# a_n919_n389# a_207_553# a_n741_109# a_n919_109# a_n29_607#
+ a_n149_n943# a_1217_109# a_n563_109# a_919_55# a_n1217_553# a_n385_n389# a_1039_109#
+ a_1039_n389# a_861_109# a_n1039_n445# a_n385_109# a_207_n943# a_n861_553# a_n683_55#
+ a_n563_n887# a_n1039_553# a_29_n445# a_1217_n887# a_683_109# a_n683_n445# a_n1217_n943#
+ a_n683_553# a_29_553# a_505_n389# a_n861_n943# a_683_n887# a_741_n445# a_n505_55#
+ a_n919_n887# a_n741_607# a_n919_607# a_1217_607# a_n563_607# a_1097_55# a_1097_n445#
+ a_n207_n389# a_n385_n887# a_1039_607# a_1039_n887# a_861_607# a_n1039_n943# a_n385_607#
+ a_29_n943# a_n327_55# a_n1275_n389# a_683_607# a_n505_n445# a_327_n389# a_n683_n943#
+ a_919_553# a_741_553# a_563_n445# a_505_n887# a_563_553# a_741_n943# a_741_55# a_n1275_109#
X0 a_n919_607# a_n1039_553# a_n1097_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1039_607# a_919_553# a_861_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_109# a_29_55# a_n29_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n1097_n887# a_n1217_n943# a_n1275_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_683_n887# a_563_n943# a_505_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n207_n389# a_n327_n445# a_n385_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n207_607# a_n327_553# a_n385_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n1275_109# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=3.248e+12p ps=2.704e+07u w=1.4e+06u l=600000u
X8 a_683_109# a_563_55# a_505_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_1217_n389# a_1097_n445# a_1039_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1275_n389# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n563_109# a_n683_55# a_n741_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n1555_n1061# a_n1555_n1061# a_1217_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_n741_n389# a_n861_n445# a_n919_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n29_n887# a_n149_n943# a_n207_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n919_109# a_n1039_55# a_n1097_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_327_109# a_207_55# a_149_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1039_109# a_919_55# a_861_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1097_n389# a_n1217_n445# a_n1275_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_683_n389# a_563_n445# a_505_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_1039_n389# a_919_n445# a_861_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_505_607# a_385_553# a_327_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n207_109# a_n327_55# a_n385_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X23 a_n563_n887# a_n683_n943# a_n741_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X24 a_1217_607# a_1097_553# a_1039_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n919_n887# a_n1039_n943# a_n1097_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_505_n887# a_385_n943# a_327_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_861_607# a_741_553# a_683_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_n29_n389# a_n149_n445# a_n207_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n385_n887# a_n505_n943# a_n563_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n741_607# a_n861_553# a_n919_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_n1555_n1061# a_n1555_n1061# a_1217_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X32 a_n29_607# a_n149_553# a_n207_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_505_109# a_385_55# a_327_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_327_n887# a_207_n943# a_149_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X35 a_n563_n389# a_n683_n445# a_n741_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X36 a_149_n887# a_29_n943# a_n29_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_n1097_607# a_n1217_553# a_n1275_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X38 a_1217_109# a_1097_55# a_1039_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n919_n389# a_n1039_n445# a_n1097_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 a_505_n389# a_385_n445# a_327_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X41 a_n385_607# a_n505_553# a_n563_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X42 a_861_109# a_741_55# a_683_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_861_n887# a_741_n943# a_683_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X44 a_n385_n389# a_n505_n445# a_n563_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X45 a_n741_109# a_n861_55# a_n919_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X46 a_n1555_n1061# a_n1555_n1061# a_1217_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X47 a_n29_109# a_n149_55# a_n207_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X48 a_327_n389# a_207_n445# a_149_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X49 a_149_n389# a_29_n445# a_n29_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X50 a_149_607# a_29_553# a_n29_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X51 a_n1097_109# a_n1217_55# a_n1275_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X52 a_n207_n887# a_n327_n943# a_n385_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X53 a_n1275_607# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X54 a_683_607# a_563_553# a_505_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X55 a_n385_109# a_n505_55# a_n563_109# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X56 a_861_n389# a_741_n445# a_683_n389# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X57 a_1217_n887# a_1097_n943# a_1039_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X58 a_n1275_n887# a_n1555_n1061# a_n1555_n1061# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X59 a_n563_607# a_n683_553# a_n741_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X60 a_n1555_n1061# a_n1555_n1061# a_1217_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X61 a_n741_n887# a_n861_n943# a_n919_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X62 a_327_607# a_207_553# a_149_607# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X63 a_1039_n887# a_919_n943# a_861_n887# a_n1555_n1061# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_327_n389# a_n919_n389# 0.01fF
C1 a_207_553# a_n1039_553# 0.01fF
C2 a_1217_n389# a_1217_607# 0.00fF
C3 a_n385_607# a_149_607# 0.02fF
C4 a_n505_553# a_1097_553# 0.01fF
C5 a_1217_109# a_1217_n389# 0.00fF
C6 a_919_55# a_n683_55# 0.01fF
C7 a_n563_n887# a_505_n887# 0.01fF
C8 a_n29_607# a_n563_607# 0.02fF
C9 a_n207_607# a_n1275_607# 0.01fF
C10 a_919_55# a_919_n445# 0.15fF
C11 a_n385_109# a_505_109# 0.01fF
C12 a_207_n943# a_n1217_n943# 0.01fF
C13 a_563_553# a_1097_553# 0.02fF
C14 a_919_553# a_n505_553# 0.01fF
C15 a_149_607# a_505_607# 0.03fF
C16 a_n861_n943# a_n149_n943# 0.01fF
C17 a_29_n445# a_919_n445# 0.01fF
C18 a_1097_55# a_385_55# 0.01fF
C19 a_919_553# a_563_553# 0.03fF
C20 a_n563_109# a_n563_607# 0.00fF
C21 a_n1039_553# a_n1039_n445# 0.03fF
C22 a_n29_n887# a_149_n887# 0.06fF
C23 a_1097_55# a_1097_553# 0.15fF
C24 a_n741_n887# a_327_n887# 0.01fF
C25 a_n29_n389# a_n29_109# 0.00fF
C26 a_n861_n943# a_741_n943# 0.01fF
C27 a_741_553# a_741_n445# 0.03fF
C28 a_29_n445# a_385_n445# 0.03fF
C29 a_385_553# a_207_553# 0.10fF
C30 a_327_109# a_1039_109# 0.01fF
C31 a_1039_n389# a_1039_607# 0.00fF
C32 a_n327_553# a_n1217_553# 0.01fF
C33 a_n861_553# a_29_553# 0.01fF
C34 a_207_n445# a_n861_n445# 0.01fF
C35 a_n1039_n445# a_n683_n445# 0.03fF
C36 a_n207_n887# a_n741_n887# 0.02fF
C37 a_n29_n887# a_n919_n887# 0.01fF
C38 a_563_n445# a_563_n943# 0.15fF
C39 a_n29_n887# a_683_n887# 0.01fF
C40 a_919_n943# a_919_n445# 0.15fF
C41 a_n563_109# a_n207_109# 0.03fF
C42 a_919_55# a_741_55# 0.10fF
C43 a_327_n389# a_327_607# 0.00fF
C44 a_861_607# a_1039_607# 0.06fF
C45 a_n29_n389# a_861_n389# 0.01fF
C46 a_207_553# a_n149_553# 0.03fF
C47 a_n385_n887# a_n385_n389# 0.00fF
C48 a_n683_553# a_n1217_553# 0.02fF
C49 a_29_55# a_n1217_55# 0.01fF
C50 a_n563_n887# a_n563_n389# 0.00fF
C51 a_1097_n445# a_919_n445# 0.10fF
C52 a_n149_n943# a_n1217_n943# 0.01fF
C53 a_n1275_109# a_n1275_n389# 0.00fF
C54 a_n1275_n389# a_n741_n389# 0.02fF
C55 a_n149_n445# a_n683_n445# 0.02fF
C56 a_n505_n445# a_n505_55# 0.15fF
C57 a_861_n887# a_505_n887# 0.03fF
C58 a_29_55# a_n149_55# 0.10fF
C59 a_385_n445# a_1097_n445# 0.01fF
C60 a_n1097_109# a_n385_109# 0.01fF
C61 a_n1217_n445# a_n683_n445# 0.02fF
C62 a_327_n389# a_n741_n389# 0.01fF
C63 a_1039_607# a_1217_607# 0.06fF
C64 a_n861_n943# a_385_n943# 0.01fF
C65 a_1097_55# a_207_55# 0.01fF
C66 a_n385_n389# a_861_n389# 0.01fF
C67 a_563_n445# a_29_n445# 0.02fF
C68 a_n741_607# a_n1275_607# 0.02fF
C69 a_149_109# a_1039_109# 0.01fF
C70 a_n563_n887# a_149_n887# 0.01fF
C71 a_149_n389# a_n563_n389# 0.01fF
C72 a_327_n389# a_n1275_n389# 0.01fF
C73 a_207_553# a_n861_553# 0.01fF
C74 a_n505_553# a_563_553# 0.01fF
C75 a_n919_607# a_683_607# 0.01fF
C76 a_29_553# a_n1217_553# 0.01fF
C77 a_861_109# a_505_109# 0.03fF
C78 a_n683_n943# a_29_n943# 0.01fF
C79 a_207_n445# a_919_n445# 0.01fF
C80 a_1217_n389# a_n207_n389# 0.01fF
C81 a_n563_n887# a_n919_n887# 0.03fF
C82 a_n149_n445# a_n149_553# 0.03fF
C83 a_n563_n887# a_683_n887# 0.01fF
C84 a_149_607# a_1039_607# 0.01fF
C85 a_29_55# a_n1039_55# 0.01fF
C86 a_n505_55# a_n327_55# 0.10fF
C87 a_n1039_n943# a_n1039_n445# 0.15fF
C88 a_n207_607# a_n1097_607# 0.01fF
C89 a_207_n445# a_385_n445# 0.10fF
C90 a_563_n445# a_1097_n445# 0.02fF
C91 a_505_n389# a_505_607# 0.00fF
C92 a_1217_n389# a_683_n389# 0.02fF
C93 a_385_n943# a_n1217_n943# 0.01fF
C94 a_n29_n389# a_n29_607# 0.00fF
C95 a_327_607# a_n1275_607# 0.01fF
C96 a_n149_55# a_563_55# 0.01fF
C97 a_149_n389# a_149_n887# 0.00fF
C98 a_741_n943# a_741_55# 0.03fF
C99 a_505_n389# a_1217_n389# 0.01fF
C100 a_n563_n389# a_n919_n389# 0.03fF
C101 a_n29_n887# a_327_n887# 0.03fF
C102 a_n327_n445# a_n861_n445# 0.02fF
C103 a_1217_109# a_505_109# 0.01fF
C104 a_n207_607# a_861_607# 0.01fF
C105 a_n1097_n887# a_505_n887# 0.01fF
C106 a_29_n943# a_n1039_n943# 0.01fF
C107 a_n1097_109# a_n1097_607# 0.00fF
C108 a_n1275_109# a_n1275_607# 0.00fF
C109 a_385_553# a_385_55# 0.15fF
C110 a_n29_109# a_1039_109# 0.01fF
C111 a_385_n943# a_385_n445# 0.15fF
C112 a_29_55# a_n683_55# 0.01fF
C113 a_n207_n887# a_n29_n887# 0.06fF
C114 a_n861_n445# a_741_n445# 0.01fF
C115 a_385_553# a_1097_553# 0.01fF
C116 a_149_n389# a_1039_n389# 0.01fF
C117 a_861_n887# a_149_n887# 0.01fF
C118 a_n861_55# a_n327_55# 0.02fF
C119 a_207_553# a_n1217_553# 0.01fF
C120 a_n861_n943# a_n505_n943# 0.03fF
C121 a_563_n445# a_207_n445# 0.03fF
C122 a_385_553# a_919_553# 0.02fF
C123 a_n385_n887# a_n385_607# 0.00fF
C124 a_n1039_55# a_563_55# 0.01fF
C125 a_n149_553# a_1097_553# 0.01fF
C126 a_29_n445# a_29_553# 0.03fF
C127 a_n207_607# a_1217_607# 0.01fF
C128 a_n1275_n389# a_n1275_607# 0.00fF
C129 a_n919_607# a_n563_607# 0.03fF
C130 a_1039_n887# a_505_n887# 0.02fF
C131 a_n919_607# a_n29_607# 0.01fF
C132 a_861_n887# a_683_n887# 0.06fF
C133 a_n1275_109# a_n385_109# 0.01fF
C134 a_919_553# a_n149_553# 0.01fF
C135 a_n919_n887# a_n919_n389# 0.00fF
C136 a_861_109# a_861_n887# 0.00fF
C137 a_n741_607# a_n1097_607# 0.03fF
C138 a_683_607# a_n385_607# 0.01fF
C139 a_1217_n887# a_1217_n389# 0.00fF
C140 a_n385_n887# a_n741_n887# 0.03fF
C141 a_861_607# a_861_n887# 0.00fF
C142 a_29_55# a_741_55# 0.01fF
C143 a_n563_n887# a_327_n887# 0.01fF
C144 a_385_55# a_n505_55# 0.01fF
C145 a_n327_n445# a_919_n445# 0.01fF
C146 a_n505_553# a_n1039_553# 0.02fF
C147 a_n505_n943# a_n1217_n943# 0.01fF
C148 a_n207_607# a_149_607# 0.03fF
C149 a_683_109# a_n385_109# 0.01fF
C150 a_563_55# a_n683_55# 0.01fF
C151 a_683_607# a_505_607# 0.06fF
C152 a_29_n445# a_n505_n445# 0.02fF
C153 a_n563_n389# a_n741_n389# 0.06fF
C154 a_n1039_553# a_563_553# 0.01fF
C155 a_n563_n887# a_n207_n887# 0.03fF
C156 a_n327_n445# a_385_n445# 0.01fF
C157 a_n741_607# a_861_607# 0.01fF
C158 a_741_n445# a_919_n445# 0.10fF
C159 a_n1217_n445# a_n1217_553# 0.03fF
C160 a_n29_n389# a_n1097_n389# 0.01fF
C161 a_1217_n389# a_861_n389# 0.03fF
C162 a_149_n389# a_149_607# 0.00fF
C163 a_n919_109# a_505_109# 0.01fF
C164 a_741_n445# a_385_n445# 0.03fF
C165 a_327_607# a_n1097_607# 0.01fF
C166 a_n207_n887# a_n207_607# 0.00fF
C167 a_n741_n887# a_n741_109# 0.00fF
C168 a_n1097_n887# a_149_n887# 0.01fF
C169 a_207_553# a_207_n943# 0.01fF
C170 a_n563_n389# a_n1275_n389# 0.01fF
C171 a_327_109# a_505_109# 0.06fF
C172 a_385_553# a_n505_553# 0.01fF
C173 a_n149_55# a_n1217_55# 0.01fF
C174 a_n1097_607# a_n1097_n887# 0.00fF
C175 a_n683_n943# a_n327_n943# 0.03fF
C176 a_385_55# a_n861_55# 0.01fF
C177 a_919_55# a_n327_55# 0.01fF
C178 a_327_n389# a_n563_n389# 0.01fF
C179 a_n505_n445# a_1097_n445# 0.01fF
C180 a_n741_n887# a_n1275_n887# 0.02fF
C181 a_n919_n887# a_n1097_n887# 0.06fF
C182 a_207_55# a_n505_55# 0.01fF
C183 a_741_55# a_741_n445# 0.15fF
C184 a_n385_n389# a_n1097_n389# 0.01fF
C185 a_741_55# a_563_55# 0.10fF
C186 a_385_553# a_563_553# 0.10fF
C187 a_1039_109# a_n207_109# 0.01fF
C188 a_327_607# a_861_607# 0.02fF
C189 a_n505_553# a_n149_553# 0.03fF
C190 a_n327_n445# a_563_n445# 0.01fF
C191 a_563_n943# a_29_n943# 0.02fF
C192 a_n385_607# a_n563_607# 0.06fF
C193 a_n29_607# a_n385_607# 0.03fF
C194 a_n563_109# a_1039_109# 0.01fF
C195 a_29_n445# a_n1039_n445# 0.01fF
C196 a_861_n887# a_327_n887# 0.02fF
C197 a_1039_n887# a_149_n887# 0.01fF
C198 a_n29_n389# a_n385_n389# 0.03fF
C199 a_n149_553# a_563_553# 0.01fF
C200 a_563_n445# a_741_n445# 0.10fF
C201 a_563_n445# a_563_55# 0.15fF
C202 a_505_n389# a_505_109# 0.00fF
C203 a_n741_607# a_149_607# 0.01fF
C204 a_n207_607# a_n207_n389# 0.00fF
C205 a_n207_n887# a_861_n887# 0.01fF
C206 a_n563_607# a_505_607# 0.01fF
C207 a_n1217_55# a_n1039_55# 0.10fF
C208 a_327_607# a_1217_607# 0.01fF
C209 a_n29_607# a_505_607# 0.02fF
C210 a_1217_n887# a_n29_n887# 0.01fF
C211 a_29_n445# a_n149_n445# 0.10fF
C212 a_1039_n887# a_683_n887# 0.03fF
C213 a_n327_n445# a_n327_553# 0.03fF
C214 a_n327_n943# a_n1039_n943# 0.01fF
C215 a_29_n445# a_n1217_n445# 0.01fF
C216 a_741_553# a_741_55# 0.15fF
C217 a_683_109# a_683_n887# 0.00fF
C218 a_149_109# a_505_109# 0.03fF
C219 a_n1097_109# a_n919_109# 0.06fF
C220 a_n505_553# a_n505_55# 0.15fF
C221 a_29_n943# a_29_n445# 0.15fF
C222 a_207_n445# a_n505_n445# 0.01fF
C223 a_1039_n389# a_1039_n887# 0.00fF
C224 a_n385_n887# a_n29_n887# 0.03fF
C225 a_149_n389# a_n207_n389# 0.03fF
C226 a_207_55# a_n861_55# 0.01fF
C227 a_n149_55# a_n1039_55# 0.01fF
C228 a_683_109# a_861_109# 0.06fF
C229 a_683_607# a_1039_607# 0.03fF
C230 a_n1097_109# a_327_109# 0.01fF
C231 a_29_n943# a_207_n943# 0.10fF
C232 a_n29_n887# a_n29_109# 0.00fF
C233 a_n861_553# a_n505_553# 0.03fF
C234 a_327_n389# a_1039_n389# 0.01fF
C235 a_29_55# a_29_553# 0.15fF
C236 a_207_553# a_207_n445# 0.03fF
C237 a_149_n389# a_683_n389# 0.02fF
C238 a_n861_n943# a_n861_n445# 0.15fF
C239 a_n1217_55# a_n1217_n943# 0.03fF
C240 a_n861_553# a_563_553# 0.01fF
C241 a_29_n943# a_919_n943# 0.01fF
C242 a_327_607# a_149_607# 0.06fF
C243 a_1097_55# a_n505_55# 0.01fF
C244 a_n919_n389# a_n919_109# 0.00fF
C245 a_n1217_55# a_n683_55# 0.02fF
C246 a_n149_n445# a_1097_n445# 0.01fF
C247 a_327_607# a_327_n887# 0.00fF
C248 a_505_n389# a_149_n389# 0.03fF
C249 a_919_55# a_385_55# 0.02fF
C250 a_n919_n389# a_n207_n389# 0.01fF
C251 a_n149_55# a_n683_55# 0.02fF
C252 a_1217_109# a_683_109# 0.02fF
C253 a_741_553# a_n327_553# 0.01fF
C254 a_n1097_n887# a_327_n887# 0.01fF
C255 a_n149_n943# a_n149_n445# 0.15fF
C256 a_207_n445# a_n1039_n445# 0.01fF
C257 a_149_n389# a_149_109# 0.00fF
C258 a_n29_109# a_505_109# 0.02fF
C259 a_919_55# a_919_553# 0.15fF
C260 a_n149_n943# a_29_n943# 0.10fF
C261 a_n919_n389# a_683_n389# 0.01fF
C262 a_149_109# a_n1097_109# 0.01fF
C263 a_385_553# a_n1039_553# 0.01fF
C264 a_741_553# a_n683_553# 0.01fF
C265 a_n207_n887# a_n1097_n887# 0.01fF
C266 a_n29_n887# a_n1275_n887# 0.01fF
C267 a_n861_n943# a_n1217_n943# 0.03fF
C268 a_n563_n887# a_n385_n887# 0.06fF
C269 a_149_n887# a_505_n887# 0.03fF
C270 a_n1275_607# a_n1097_607# 0.06fF
C271 a_741_n943# a_29_n943# 0.01fF
C272 a_n505_553# a_n1217_553# 0.01fF
C273 a_505_n389# a_n919_n389# 0.01fF
C274 a_207_n445# a_n149_n445# 0.03fF
C275 a_n149_553# a_n1039_553# 0.01fF
C276 a_207_n445# a_n1217_n445# 0.01fF
C277 a_1039_n887# a_327_n887# 0.01fF
C278 a_n563_607# a_1039_607# 0.01fF
C279 a_n683_n943# a_n683_n445# 0.15fF
C280 a_n29_607# a_1039_607# 0.01fF
C281 a_n1039_55# a_n683_55# 0.03fF
C282 a_n919_n887# a_505_n887# 0.01fF
C283 a_505_n887# a_683_n887# 0.06fF
C284 a_n741_109# a_505_109# 0.01fF
C285 a_327_607# a_327_109# 0.00fF
C286 a_741_55# a_n149_55# 0.01fF
C287 a_207_55# a_919_55# 0.01fF
C288 a_919_553# a_919_n943# 0.01fF
C289 a_327_n389# a_327_n887# 0.00fF
C290 a_1097_n445# a_1097_553# 0.03fF
C291 a_n861_n445# a_385_n445# 0.01fF
C292 a_n207_n887# a_1039_n887# 0.01fF
C293 a_n327_n445# a_n505_n445# 0.10fF
C294 a_n29_n887# a_n29_607# 0.00fF
C295 a_29_55# a_n327_55# 0.03fF
C296 a_683_607# a_n207_607# 0.01fF
C297 a_n1039_553# a_n1039_n943# 0.01fF
C298 a_n1275_109# a_n919_109# 0.03fF
C299 a_563_n943# a_n327_n943# 0.01fF
C300 a_741_553# a_29_553# 0.01fF
C301 a_207_55# a_207_n943# 0.03fF
C302 a_n505_n445# a_741_n445# 0.01fF
C303 a_n1275_109# a_327_109# 0.01fF
C304 a_n385_n389# a_n385_607# 0.00fF
C305 a_29_n943# a_385_n943# 0.03fF
C306 a_385_553# a_n149_553# 0.02fF
C307 a_n1097_109# a_n29_109# 0.01fF
C308 a_563_n943# a_563_553# 0.01fF
C309 a_n505_n445# a_n505_n943# 0.15fF
C310 a_1217_n887# a_861_n887# 0.03fF
C311 a_n29_n389# a_1217_n389# 0.01fF
C312 a_861_109# a_n385_109# 0.01fF
C313 a_n741_n389# a_n207_n389# 0.02fF
C314 a_n861_553# a_n1039_553# 0.10fF
C315 a_n563_n887# a_n1275_n887# 0.01fF
C316 a_149_n389# a_861_n389# 0.01fF
C317 a_683_109# a_n919_109# 0.01fF
C318 a_n385_n887# a_861_n887# 0.01fF
C319 a_29_n943# a_1097_n943# 0.01fF
C320 a_n741_n389# a_683_n389# 0.01fF
C321 a_563_n445# a_n861_n445# 0.01fF
C322 a_29_n943# a_29_55# 0.03fF
C323 a_n327_n445# a_n327_55# 0.15fF
C324 a_327_109# a_683_109# 0.03fF
C325 a_n919_607# a_n385_607# 0.02fF
C326 a_n1275_n389# a_n207_n389# 0.01fF
C327 a_n327_n445# a_n1039_n445# 0.01fF
C328 a_n683_n943# a_n1039_n943# 0.03fF
C329 a_327_n389# a_327_109# 0.00fF
C330 a_n385_n389# a_1217_n389# 0.01fF
C331 a_505_n389# a_n741_n389# 0.01fF
C332 a_n1097_109# a_n741_109# 0.03fF
C333 a_n327_n943# a_207_n943# 0.02fF
C334 a_n563_n389# a_1039_n389# 0.01fF
C335 a_n327_55# a_563_55# 0.01fF
C336 a_385_n445# a_919_n445# 0.02fF
C337 a_327_n389# a_n207_n389# 0.02fF
C338 a_861_n887# a_861_n389# 0.00fF
C339 a_n563_n887# a_n563_607# 0.00fF
C340 a_n1275_607# a_149_607# 0.01fF
C341 a_1097_55# a_919_55# 0.10fF
C342 a_683_109# a_683_n389# 0.00fF
C343 a_n919_607# a_505_607# 0.01fF
C344 a_n207_109# a_505_109# 0.01fF
C345 a_385_55# a_385_n943# 0.03fF
C346 a_1217_109# a_n385_109# 0.01fF
C347 a_385_553# a_n861_553# 0.01fF
C348 a_207_553# a_741_553# 0.02fF
C349 a_149_109# a_n1275_109# 0.01fF
C350 a_n327_n943# a_919_n943# 0.01fF
C351 a_741_55# a_n683_55# 0.01fF
C352 a_n563_109# a_505_109# 0.01fF
C353 a_327_n389# a_683_n389# 0.03fF
C354 a_n327_n445# a_n149_n445# 0.10fF
C355 a_n741_607# a_683_607# 0.01fF
C356 a_n919_n887# a_149_n887# 0.01fF
C357 a_n327_n445# a_n1217_n445# 0.01fF
C358 a_n207_607# a_n563_607# 0.03fF
C359 a_149_n887# a_683_n887# 0.02fF
C360 a_327_n887# a_505_n887# 0.06fF
C361 a_n207_607# a_n29_607# 0.06fF
C362 a_n861_553# a_n149_553# 0.01fF
C363 a_207_55# a_207_n445# 0.15fF
C364 a_327_n389# a_505_n389# 0.06fF
C365 a_n563_n887# a_n563_109# 0.00fF
C366 a_n1039_553# a_n1217_553# 0.10fF
C367 a_n149_n445# a_741_n445# 0.01fF
C368 a_1097_n943# a_1097_553# 0.01fF
C369 a_29_55# a_385_55# 0.03fF
C370 a_n741_607# a_n741_109# 0.00fF
C371 a_n207_n887# a_505_n887# 0.01fF
C372 a_149_109# a_683_109# 0.02fF
C373 a_n919_n887# a_683_n887# 0.01fF
C374 a_n207_607# a_n207_109# 0.00fF
C375 a_n149_n943# a_n327_n943# 0.10fF
C376 a_29_n943# a_n505_n943# 0.02fF
C377 a_563_n445# a_919_n445# 0.03fF
C378 a_1097_55# a_1097_n445# 0.15fF
C379 a_n385_n887# a_n1097_n887# 0.01fF
C380 a_563_n445# a_385_n445# 0.10fF
C381 a_n29_n389# a_n29_n887# 0.00fF
C382 a_327_607# a_683_607# 0.03fF
C383 a_741_n943# a_n327_n943# 0.01fF
C384 a_861_607# a_861_109# 0.00fF
C385 a_n1097_109# a_n207_109# 0.01fF
C386 a_385_553# a_n1217_553# 0.01fF
C387 a_n1275_109# a_n29_109# 0.01fF
C388 a_1217_n887# a_1039_n887# 0.06fF
C389 a_n1097_109# a_n563_109# 0.02fF
C390 a_n683_553# a_n683_55# 0.15fF
C391 a_207_55# a_29_55# 0.10fF
C392 a_n385_n887# a_1039_n887# 0.01fF
C393 a_385_55# a_563_55# 0.10fF
C394 a_n149_553# a_n1217_553# 0.01fF
C395 a_n741_n389# a_861_n389# 0.01fF
C396 a_n741_607# a_n563_607# 0.06fF
C397 a_n385_607# a_505_607# 0.01fF
C398 a_n741_607# a_n29_607# 0.01fF
C399 a_n505_55# a_n861_55# 0.03fF
C400 a_n919_109# a_n385_109# 0.02fF
C401 a_n29_109# a_683_109# 0.01fF
C402 a_1217_109# a_861_109# 0.03fF
C403 a_327_109# a_n385_109# 0.01fF
C404 a_149_607# a_149_n887# 0.00fF
C405 a_n327_n943# a_385_n943# 0.01fF
C406 a_n1275_109# a_n741_109# 0.02fF
C407 a_861_607# a_1217_607# 0.03fF
C408 a_n861_553# a_n861_55# 0.15fF
C409 a_n741_n389# a_n741_109# 0.00fF
C410 a_n683_n943# a_563_n943# 0.01fF
C411 a_149_n887# a_327_n887# 0.06fF
C412 a_683_607# a_683_109# 0.00fF
C413 a_n1097_607# a_149_607# 0.01fF
C414 a_n1275_n887# a_n1097_n887# 0.06fF
C415 a_505_n389# a_505_n887# 0.00fF
C416 a_n505_n445# a_n861_n445# 0.03fF
C417 a_29_n445# a_n683_n445# 0.01fF
C418 a_n1217_55# a_n327_55# 0.01fF
C419 a_n327_n943# a_1097_n943# 0.01fF
C420 a_327_n389# a_861_n389# 0.02fF
C421 a_n1275_109# a_n1275_n887# 0.00fF
C422 a_n207_n887# a_149_n887# 0.03fF
C423 a_n919_n887# a_327_n887# 0.01fF
C424 a_327_n887# a_683_n887# 0.03fF
C425 a_683_109# a_n741_109# 0.01fF
C426 a_n149_55# a_n327_55# 0.10fF
C427 a_741_553# a_1097_553# 0.03fF
C428 a_327_607# a_n563_607# 0.01fF
C429 a_327_607# a_n29_607# 0.03fF
C430 a_n861_553# a_n1217_553# 0.03fF
C431 a_1217_109# a_1217_607# 0.00fF
C432 a_n563_n389# a_n207_n389# 0.03fF
C433 a_861_607# a_149_607# 0.01fF
C434 a_207_55# a_563_55# 0.03fF
C435 a_n207_n887# a_n919_n887# 0.01fF
C436 a_741_553# a_919_553# 0.10fF
C437 a_n207_n887# a_683_n887# 0.01fF
C438 a_149_n389# a_n1097_n389# 0.01fF
C439 a_1097_55# a_1097_n943# 0.03fF
C440 a_563_n943# a_n1039_n943# 0.01fF
C441 a_n683_n943# a_207_n943# 0.01fF
C442 a_n1275_n389# a_n1275_n887# 0.00fF
C443 a_n1217_55# a_n1217_n445# 0.15fF
C444 a_n563_n389# a_683_n389# 0.01fF
C445 a_149_109# a_n385_109# 0.02fF
C446 a_1097_55# a_29_55# 0.01fF
C447 a_n1097_109# a_n1097_n389# 0.00fF
C448 a_n29_n389# a_149_n389# 0.06fF
C449 a_1039_109# a_1039_607# 0.00fF
C450 a_n149_n445# a_n149_55# 0.15fF
C451 a_n861_n445# a_n1039_n445# 0.10fF
C452 a_n683_n943# a_919_n943# 0.01fF
C453 a_149_607# a_1217_607# 0.01fF
C454 a_n327_n445# a_n327_n943# 0.15fF
C455 a_505_n389# a_n563_n389# 0.01fF
C456 a_1217_n887# a_505_n887# 0.01fF
C457 a_n1039_55# a_n327_55# 0.01fF
C458 a_n919_n887# a_n919_109# 0.00fF
C459 a_n683_553# a_n327_553# 0.03fF
C460 a_n505_n445# a_919_n445# 0.01fF
C461 a_n1275_109# a_n207_109# 0.01fF
C462 a_n1039_55# a_n1039_n445# 0.15fF
C463 a_919_55# a_n505_55# 0.01fF
C464 a_n385_n887# a_505_n887# 0.01fF
C465 a_n1275_109# a_n563_109# 0.01fF
C466 a_n385_607# a_1039_607# 0.01fF
C467 a_n1097_n389# a_n919_n389# 0.06fF
C468 a_n505_553# a_n505_n943# 0.01fF
C469 a_n861_n445# a_n149_n445# 0.01fF
C470 a_n505_n445# a_385_n445# 0.01fF
C471 a_149_n389# a_n385_n389# 0.02fF
C472 a_n505_n943# a_n327_n943# 0.10fF
C473 a_207_n943# a_n1039_n943# 0.01fF
C474 a_563_553# a_563_55# 0.15fF
C475 a_n861_n445# a_n1217_n445# 0.03fF
C476 a_327_109# a_861_109# 0.02fF
C477 a_n919_607# a_n207_607# 0.01fF
C478 a_207_n445# a_n683_n445# 0.01fF
C479 a_n29_n389# a_n919_n389# 0.01fF
C480 a_n861_n943# a_29_n943# 0.01fF
C481 a_n683_n943# a_n149_n943# 0.02fF
C482 a_1039_n389# a_n207_n389# 0.01fF
C483 a_683_109# a_n207_109# 0.01fF
C484 a_385_55# a_n1217_55# 0.01fF
C485 a_1039_607# a_505_607# 0.02fF
C486 a_683_n389# a_683_n887# 0.00fF
C487 a_n385_n887# a_n385_109# 0.00fF
C488 a_n563_109# a_683_109# 0.01fF
C489 a_1097_55# a_563_55# 0.02fF
C490 a_n327_55# a_n683_55# 0.03fF
C491 a_n149_n943# a_n149_553# 0.01fF
C492 a_n29_109# a_n385_109# 0.03fF
C493 a_n683_n943# a_741_n943# 0.01fF
C494 a_1039_n389# a_683_n389# 0.03fF
C495 a_385_55# a_n149_55# 0.02fF
C496 a_741_553# a_n505_553# 0.01fF
C497 a_149_109# a_149_n887# 0.00fF
C498 a_n327_553# a_29_553# 0.03fF
C499 a_1039_109# a_505_109# 0.02fF
C500 a_n29_n887# a_n741_n887# 0.01fF
C501 a_n385_n389# a_n919_n389# 0.02fF
C502 a_505_n389# a_1039_n389# 0.02fF
C503 a_741_553# a_563_553# 0.10fF
C504 a_n1275_607# a_n1275_n887# 0.00fF
C505 a_n207_n887# a_327_n887# 0.02fF
C506 a_563_n445# a_n505_n445# 0.01fF
C507 a_327_109# a_1217_109# 0.01fF
C508 a_n683_553# a_29_553# 0.01fF
C509 a_n1217_n445# a_n1217_n943# 0.15fF
C510 a_385_n445# a_n1039_n445# 0.01fF
C511 a_29_n943# a_n1217_n943# 0.01fF
C512 a_n149_n943# a_n1039_n943# 0.01fF
C513 a_n385_109# a_n741_109# 0.03fF
C514 a_149_109# a_861_109# 0.01fF
C515 a_n1097_n389# a_n1097_n887# 0.00fF
C516 a_n149_n445# a_919_n445# 0.01fF
C517 a_385_553# a_385_n943# 0.01fF
C518 a_207_55# a_n1217_55# 0.01fF
C519 a_n919_607# a_n919_n389# 0.00fF
C520 a_n683_n943# a_385_n943# 0.01fF
C521 a_741_55# a_n327_55# 0.01fF
C522 a_1217_n887# a_149_n887# 0.01fF
C523 a_385_55# a_n1039_55# 0.01fF
C524 a_n563_n389# a_861_n389# 0.01fF
C525 a_n1097_n389# a_n741_n389# 0.03fF
C526 a_n149_n445# a_385_n445# 0.02fF
C527 a_n741_607# a_n919_607# 0.06fF
C528 a_n1275_607# a_n563_607# 0.01fF
C529 a_505_109# a_505_607# 0.00fF
C530 a_n29_607# a_n1275_607# 0.01fF
C531 a_n1217_n445# a_385_n445# 0.01fF
C532 a_207_55# a_n149_55# 0.03fF
C533 a_n385_n887# a_149_n887# 0.02fF
C534 a_327_109# a_327_n887# 0.00fF
C535 a_n29_n389# a_n741_n389# 0.01fF
C536 a_1217_n887# a_683_n887# 0.02fF
C537 a_207_553# a_n327_553# 0.02fF
C538 a_n207_607# a_n385_607# 0.06fF
C539 a_563_n445# a_n1039_n445# 0.01fF
C540 a_149_109# a_1217_109# 0.01fF
C541 a_n1275_n389# a_n1097_n389# 0.06fF
C542 a_n385_n887# a_n919_n887# 0.02fF
C543 a_n563_n887# a_n741_n887# 0.06fF
C544 a_n385_n887# a_683_n887# 0.01fF
C545 a_n207_n887# a_n207_n389# 0.00fF
C546 a_n327_n445# a_n683_n445# 0.03fF
C547 a_327_n389# a_n1097_n389# 0.01fF
C548 a_207_553# a_n683_553# 0.01fF
C549 a_385_55# a_n683_55# 0.01fF
C550 a_385_n943# a_n1039_n943# 0.01fF
C551 a_n207_607# a_505_607# 0.01fF
C552 a_n29_n389# a_n1275_n389# 0.01fF
C553 a_n29_109# a_861_109# 0.01fF
C554 a_n327_553# a_n327_55# 0.15fF
C555 a_563_n943# a_207_n943# 0.03fF
C556 a_n385_n389# a_n741_n389# 0.03fF
C557 a_327_607# a_n919_607# 0.01fF
C558 a_327_n389# a_n29_n389# 0.03fF
C559 a_563_n445# a_n149_n445# 0.01fF
C560 a_741_n445# a_n683_n445# 0.01fF
C561 a_683_607# a_683_n887# 0.00fF
C562 a_207_55# a_n1039_55# 0.01fF
C563 a_149_109# a_149_607# 0.00fF
C564 a_327_109# a_n919_109# 0.01fF
C565 a_n385_109# a_n207_109# 0.06fF
C566 a_385_55# a_385_n445# 0.15fF
C567 a_1217_n887# a_1217_607# 0.00fF
C568 a_1039_n389# a_861_n389# 0.06fF
C569 a_861_109# a_861_n389# 0.00fF
C570 a_563_n943# a_919_n943# 0.03fF
C571 a_919_553# a_919_n445# 0.03fF
C572 a_n563_109# a_n385_109# 0.06fF
C573 a_1217_n887# a_1217_109# 0.00fF
C574 a_683_607# a_861_607# 0.06fF
C575 a_29_55# a_n505_55# 0.02fF
C576 a_n1275_n887# a_149_n887# 0.01fF
C577 a_n563_n389# a_n563_607# 0.00fF
C578 a_n385_n389# a_n1275_n389# 0.01fF
C579 a_861_607# a_861_n389# 0.00fF
C580 a_149_n389# a_1217_n389# 0.01fF
C581 a_861_109# a_n741_109# 0.01fF
C582 a_327_n389# a_n385_n389# 0.01fF
C583 a_1097_55# a_n149_55# 0.01fF
C584 a_n861_n943# a_n327_n943# 0.02fF
C585 a_385_55# a_741_55# 0.03fF
C586 a_207_553# a_29_553# 0.10fF
C587 a_n683_n943# a_n505_n943# 0.10fF
C588 a_1217_109# a_n29_109# 0.01fF
C589 a_919_55# a_919_n943# 0.03fF
C590 a_n919_n887# a_n1275_n887# 0.03fF
C591 a_207_55# a_n683_55# 0.01fF
C592 a_n741_607# a_n385_607# 0.03fF
C593 a_n741_n887# a_861_n887# 0.01fF
C594 a_563_n943# a_n149_n943# 0.01fF
C595 a_n207_n389# a_683_n389# 0.01fF
C596 a_683_607# a_1217_607# 0.02fF
C597 a_n563_n389# a_n563_109# 0.00fF
C598 a_1217_n887# a_327_n887# 0.01fF
C599 a_207_n943# a_919_n943# 0.01fF
C600 a_29_n445# a_1097_n445# 0.01fF
C601 a_563_n943# a_741_n943# 0.10fF
C602 a_385_553# a_741_553# 0.03fF
C603 a_505_n389# a_n207_n389# 0.01fF
C604 a_n741_607# a_505_607# 0.01fF
C605 a_149_109# a_n919_109# 0.01fF
C606 a_n1097_607# a_n563_607# 0.02fF
C607 a_n741_607# a_n741_n887# 0.00fF
C608 a_n29_607# a_n1097_607# 0.01fF
C609 a_29_55# a_n861_55# 0.01fF
C610 a_n385_n887# a_327_n887# 0.01fF
C611 a_1217_n887# a_n207_n887# 0.01fF
C612 a_149_109# a_327_109# 0.06fF
C613 a_n505_55# a_563_55# 0.01fF
C614 a_n327_n943# a_n1217_n943# 0.01fF
C615 a_n505_n943# a_n1039_n943# 0.02fF
C616 a_505_n389# a_683_n389# 0.06fF
C617 a_741_553# a_n149_553# 0.01fF
C618 a_683_607# a_149_607# 0.02fF
C619 a_n505_n943# a_n505_55# 0.03fF
C620 a_327_607# a_n385_607# 0.01fF
C621 a_n563_n887# a_n29_n887# 0.02fF
C622 a_n207_607# a_1039_607# 0.01fF
C623 a_n385_n887# a_n207_n887# 0.06fF
C624 a_207_55# a_741_55# 0.02fF
C625 a_n149_n943# a_207_n943# 0.03fF
C626 a_n327_553# a_1097_553# 0.01fF
C627 a_861_607# a_n563_607# 0.01fF
C628 a_861_607# a_n29_607# 0.01fF
C629 a_29_n943# a_29_553# 0.01fF
C630 a_919_553# a_n327_553# 0.01fF
C631 a_861_109# a_n207_109# 0.01fF
C632 a_563_n943# a_385_n943# 0.10fF
C633 a_741_n943# a_207_n943# 0.02fF
C634 a_327_607# a_505_607# 0.06fF
C635 a_1039_109# a_1039_n887# 0.00fF
C636 a_207_n445# a_29_n445# 0.10fF
C637 a_n149_n943# a_919_n943# 0.01fF
C638 a_n505_n445# a_n1039_n445# 0.02fF
C639 a_n563_109# a_861_109# 0.01fF
C640 a_683_109# a_1039_109# 0.03fF
C641 a_207_n445# a_207_n943# 0.15fF
C642 a_919_553# a_n683_553# 0.01fF
C643 a_n861_55# a_563_55# 0.01fF
C644 a_563_n943# a_1097_n943# 0.02fF
C645 a_n741_n887# a_n1097_n887# 0.03fF
C646 a_741_n943# a_919_n943# 0.10fF
C647 a_n29_607# a_1217_607# 0.01fF
C648 a_n29_109# a_n919_109# 0.01fF
C649 a_741_553# a_n861_553# 0.01fF
C650 a_n563_n389# a_n1097_n389# 0.02fF
C651 a_n1275_n887# a_327_n887# 0.01fF
C652 a_n505_n445# a_n149_n445# 0.03fF
C653 a_n919_607# a_n1275_607# 0.03fF
C654 a_327_109# a_n29_109# 0.03fF
C655 a_n741_n887# a_n741_n389# 0.00fF
C656 a_n505_n445# a_n1217_n445# 0.01fF
C657 a_n29_n389# a_n563_n389# 0.02fF
C658 a_n385_n389# a_n385_109# 0.00fF
C659 a_1217_109# a_n207_109# 0.01fF
C660 a_207_n445# a_1097_n445# 0.01fF
C661 a_n207_n887# a_n1275_n887# 0.01fF
C662 a_207_n943# a_385_n943# 0.10fF
C663 a_n29_n887# a_861_n887# 0.01fF
C664 a_29_55# a_919_55# 0.01fF
C665 a_1097_553# a_29_553# 0.01fF
C666 a_741_n943# a_n149_n943# 0.01fF
C667 a_n207_n389# a_861_n389# 0.01fF
C668 a_n1039_55# a_n1039_553# 0.15fF
C669 a_n919_109# a_n741_109# 0.06fF
C670 a_149_607# a_n563_607# 0.01fF
C671 a_n29_607# a_149_607# 0.06fF
C672 a_n861_n445# a_n683_n445# 0.10fF
C673 a_1097_55# a_741_55# 0.03fF
C674 a_563_n445# a_563_553# 0.03fF
C675 a_29_55# a_29_n445# 0.15fF
C676 a_385_n943# a_919_n943# 0.02fF
C677 a_207_n943# a_1097_n943# 0.01fF
C678 a_919_553# a_29_553# 0.01fF
C679 a_327_109# a_n741_109# 0.01fF
C680 a_683_607# a_683_n389# 0.00fF
C681 a_n1097_n389# a_n1097_607# 0.00fF
C682 a_683_n389# a_861_n389# 0.06fF
C683 a_n385_n389# a_n563_n389# 0.06fF
C684 a_n149_55# a_n149_553# 0.15fF
C685 a_n327_553# a_n505_553# 0.10fF
C686 a_n1097_109# a_505_109# 0.01fF
C687 a_327_n389# a_1217_n389# 0.01fF
C688 a_n327_553# a_n327_n943# 0.01fF
C689 a_919_n943# a_1097_n943# 0.10fF
C690 a_n149_n445# a_n1039_n445# 0.01fF
C691 a_563_n943# a_563_55# 0.03fF
C692 a_149_109# a_n29_109# 0.06fF
C693 a_505_n389# a_861_n389# 0.03fF
C694 a_n861_n943# a_n683_n943# 0.10fF
C695 a_n1217_n445# a_n1039_n445# 0.10fF
C696 a_n327_553# a_563_553# 0.01fF
C697 a_563_n943# a_n505_n943# 0.01fF
C698 a_n505_55# a_n1217_55# 0.01fF
C699 a_n683_553# a_n505_553# 0.10fF
C700 a_1097_n445# a_1097_n943# 0.15fF
C701 a_327_607# a_1039_607# 0.01fF
C702 a_n149_n943# a_385_n943# 0.02fF
C703 a_n207_n887# a_n207_109# 0.00fF
C704 a_n29_n389# a_1039_n389# 0.01fF
C705 a_n327_n445# a_29_n445# 0.03fF
C706 a_n683_553# a_563_553# 0.01fF
C707 a_n505_55# a_n149_55# 0.03fF
C708 a_919_55# a_563_55# 0.03fF
C709 a_n149_n445# a_n1217_n445# 0.01fF
C710 a_207_553# a_1097_553# 0.01fF
C711 a_n683_n445# a_n683_55# 0.15fF
C712 a_741_n943# a_385_n943# 0.03fF
C713 a_n563_n887# a_861_n887# 0.01fF
C714 a_n149_n943# a_1097_n943# 0.01fF
C715 a_1217_n887# a_n385_n887# 0.01fF
C716 a_149_109# a_n741_109# 0.01fF
C717 a_n1275_607# a_n385_607# 0.01fF
C718 a_29_n445# a_741_n445# 0.01fF
C719 a_919_n445# a_n683_n445# 0.01fF
C720 a_207_553# a_919_553# 0.01fF
C721 a_n29_n887# a_n1097_n887# 0.01fF
C722 a_1039_109# a_n385_109# 0.01fF
C723 a_741_n943# a_1097_n943# 0.03fF
C724 a_n683_n943# a_n1217_n943# 0.02fF
C725 a_n861_n943# a_n1039_n943# 0.10fF
C726 a_n919_109# a_n207_109# 0.01fF
C727 a_385_55# a_n327_55# 0.01fF
C728 a_n385_n389# a_1039_n389# 0.01fF
C729 a_n505_n943# a_207_n943# 0.01fF
C730 a_385_n445# a_n683_n445# 0.01fF
C731 a_n563_109# a_n919_109# 0.03fF
C732 a_n683_n943# a_n683_55# 0.03fF
C733 a_n861_55# a_n1217_55# 0.03fF
C734 a_327_109# a_n207_109# 0.02fF
C735 a_n919_607# a_n1097_607# 0.06fF
C736 a_n327_n445# a_1097_n445# 0.01fF
C737 a_n505_553# a_29_553# 0.02fF
C738 a_n1039_55# a_n1039_n943# 0.03fF
C739 a_1039_n887# a_1039_607# 0.00fF
C740 a_n207_n389# a_n207_109# 0.00fF
C741 a_n861_553# a_n861_n445# 0.03fF
C742 a_327_109# a_n563_109# 0.01fF
C743 a_n505_55# a_n1039_55# 0.02fF
C744 a_n919_607# a_n919_n887# 0.00fF
C745 a_n861_n943# a_n861_553# 0.01fF
C746 a_505_607# a_505_n887# 0.00fF
C747 a_n505_n943# a_919_n943# 0.01fF
C748 a_n385_607# a_n385_109# 0.00fF
C749 a_n741_607# a_n207_607# 0.02fF
C750 a_n741_n887# a_505_n887# 0.01fF
C751 a_n149_55# a_n861_55# 0.01fF
C752 a_563_553# a_29_553# 0.02fF
C753 a_741_n445# a_1097_n445# 0.03fF
C754 a_385_553# a_385_n445# 0.03fF
C755 a_n29_n887# a_1039_n887# 0.01fF
C756 a_207_553# a_207_55# 0.15fF
C757 a_149_n389# a_n919_n389# 0.01fF
C758 a_n1217_55# a_n1217_553# 0.15fF
C759 a_n1217_n943# a_n1039_n943# 0.10fF
C760 a_385_n943# a_1097_n943# 0.01fF
C761 a_n29_109# a_n741_109# 0.01fF
C762 a_n861_n445# a_n861_55# 0.15fF
C763 a_563_n445# a_n683_n445# 0.01fF
C764 a_n505_n445# a_n505_553# 0.03fF
C765 a_n861_n943# a_n861_55# 0.03fF
C766 a_n149_n943# a_n505_n943# 0.03fF
C767 a_207_55# a_n327_55# 0.02fF
C768 a_n327_n445# a_207_n445# 0.02fF
C769 a_n505_55# a_n683_55# 0.10fF
C770 a_n385_n887# a_n1275_n887# 0.01fF
C771 a_n563_n887# a_n1097_n887# 0.02fF
C772 a_741_n943# a_741_n445# 0.15fF
C773 a_149_109# a_n207_109# 0.03fF
C774 a_n327_553# a_n1039_553# 0.01fF
C775 a_327_607# a_n207_607# 0.02fF
C776 a_n861_55# a_n1039_55# 0.10fF
C777 a_741_n943# a_n505_n943# 0.01fF
C778 a_149_109# a_n563_109# 0.01fF
C779 a_207_553# a_n505_553# 0.01fF
C780 a_207_n445# a_741_n445# 0.02fF
C781 a_n683_553# a_n1039_553# 0.03fF
C782 a_683_109# a_505_109# 0.06fF
C783 a_207_553# a_563_553# 0.03fF
C784 a_1039_n389# a_1039_109# 0.00fF
C785 a_861_109# a_1039_109# 0.06fF
C786 a_n563_n887# a_1039_n887# 0.01fF
C787 a_n683_553# a_n683_n445# 0.03fF
C788 a_n385_607# a_n1097_607# 0.01fF
C789 a_n327_n943# a_n327_55# 0.03fF
C790 a_741_n943# a_741_553# 0.01fF
C791 a_n919_607# a_149_607# 0.01fF
C792 a_n1097_n389# a_n207_n389# 0.01fF
C793 a_385_553# a_n327_553# 0.01fF
C794 a_741_55# a_n505_55# 0.01fF
C795 a_n29_607# a_n29_109# 0.00fF
C796 a_n861_55# a_n683_55# 0.10fF
C797 a_n1097_109# a_n1097_n887# 0.00fF
C798 a_919_55# a_n149_55# 0.01fF
C799 a_n741_n887# a_149_n887# 0.01fF
C800 a_149_n389# a_n741_n389# 0.01fF
C801 a_n505_n943# a_385_n943# 0.01fF
C802 a_n29_n389# a_n207_n389# 0.06fF
C803 a_919_553# a_1097_553# 0.10fF
C804 a_n861_n943# a_563_n943# 0.01fF
C805 a_683_607# a_n563_607# 0.01fF
C806 a_n1097_607# a_505_607# 0.01fF
C807 a_683_607# a_n29_607# 0.01fF
C808 a_n1097_109# a_n1275_109# 0.06fF
C809 a_n327_553# a_n149_553# 0.10fF
C810 a_385_553# a_n683_553# 0.01fF
C811 a_n683_n943# a_n683_553# 0.01fF
C812 a_n29_109# a_n207_109# 0.06fF
C813 a_861_607# a_n385_607# 0.01fF
C814 a_n1039_553# a_29_553# 0.01fF
C815 a_n1217_n943# a_n1217_553# 0.01fF
C816 a_1097_55# a_n327_55# 0.01fF
C817 a_n29_n887# a_505_n887# 0.02fF
C818 a_n919_n887# a_n741_n887# 0.06fF
C819 a_n563_109# a_n29_109# 0.02fF
C820 a_n505_n943# a_1097_n943# 0.01fF
C821 a_n29_n389# a_683_n389# 0.01fF
C822 a_29_55# a_563_55# 0.02fF
C823 a_n741_n887# a_683_n887# 0.01fF
C824 a_505_n389# a_n1097_n389# 0.01fF
C825 a_1217_109# a_1039_109# 0.06fF
C826 a_n683_553# a_n149_553# 0.02fF
C827 a_327_607# a_n741_607# 0.01fF
C828 a_149_n389# a_n1275_n389# 0.01fF
C829 a_29_n943# a_n327_n943# 0.03fF
C830 a_207_55# a_385_55# 0.10fF
C831 a_505_n389# a_n29_n389# 0.02fF
C832 a_327_n389# a_149_n389# 0.06fF
C833 a_861_607# a_505_607# 0.03fF
C834 a_n385_n389# a_n207_n389# 0.06fF
C835 a_29_n445# a_n861_n445# 0.01fF
C836 a_741_55# a_n861_55# 0.01fF
C837 a_n741_n389# a_n919_n389# 0.06fF
C838 a_n385_607# a_1217_607# 0.01fF
C839 a_1039_n389# a_1217_n389# 0.06fF
C840 a_n741_109# a_n207_109# 0.02fF
C841 a_n919_607# a_n919_109# 0.00fF
C842 a_n861_n943# a_207_n943# 0.01fF
C843 a_n385_n389# a_683_n389# 0.01fF
C844 a_n563_109# a_n741_109# 0.06fF
C845 a_861_n887# a_1039_n887# 0.06fF
C846 a_n741_607# a_n741_n389# 0.00fF
C847 a_385_553# a_29_553# 0.03fF
C848 a_n861_553# a_n327_553# 0.02fF
C849 a_n327_n445# a_741_n445# 0.01fF
C850 a_505_607# a_1217_607# 0.01fF
C851 a_505_109# a_505_n887# 0.00fF
C852 a_n1275_n389# a_n919_n389# 0.03fF
C853 a_505_n389# a_n385_n389# 0.01fF
C854 a_n149_n943# a_n149_55# 0.03fF
C855 a_n861_553# a_n683_553# 0.10fF
C856 a_n149_553# a_29_553# 0.10fF
C857 a_n505_n445# a_n683_n445# 0.10fF
C858 a_1217_n887# a_n1555_n1061# 0.10fF
C859 a_1039_n887# a_n1555_n1061# 0.05fF
C860 a_861_n887# a_n1555_n1061# 0.04fF
C861 a_683_n887# a_n1555_n1061# 0.03fF
C862 a_505_n887# a_n1555_n1061# 0.03fF
C863 a_327_n887# a_n1555_n1061# 0.03fF
C864 a_149_n887# a_n1555_n1061# 0.03fF
C865 a_n29_n887# a_n1555_n1061# 0.03fF
C866 a_n207_n887# a_n1555_n1061# 0.03fF
C867 a_n385_n887# a_n1555_n1061# 0.03fF
C868 a_n563_n887# a_n1555_n1061# 0.03fF
C869 a_n741_n887# a_n1555_n1061# 0.03fF
C870 a_n919_n887# a_n1555_n1061# 0.04fF
C871 a_n1097_n887# a_n1555_n1061# 0.05fF
C872 a_n1275_n887# a_n1555_n1061# 0.10fF
C873 a_1097_n943# a_n1555_n1061# 0.27fF
C874 a_919_n943# a_n1555_n1061# 0.23fF
C875 a_741_n943# a_n1555_n1061# 0.23fF
C876 a_563_n943# a_n1555_n1061# 0.24fF
C877 a_385_n943# a_n1555_n1061# 0.24fF
C878 a_207_n943# a_n1555_n1061# 0.25fF
C879 a_29_n943# a_n1555_n1061# 0.26fF
C880 a_n149_n943# a_n1555_n1061# 0.26fF
C881 a_n327_n943# a_n1555_n1061# 0.26fF
C882 a_n505_n943# a_n1555_n1061# 0.26fF
C883 a_n683_n943# a_n1555_n1061# 0.26fF
C884 a_n861_n943# a_n1555_n1061# 0.26fF
C885 a_n1039_n943# a_n1555_n1061# 0.27fF
C886 a_n1217_n943# a_n1555_n1061# 0.32fF
C887 a_1217_n389# a_n1555_n1061# 0.10fF
C888 a_1039_n389# a_n1555_n1061# 0.05fF
C889 a_861_n389# a_n1555_n1061# 0.04fF
C890 a_683_n389# a_n1555_n1061# 0.03fF
C891 a_505_n389# a_n1555_n1061# 0.03fF
C892 a_327_n389# a_n1555_n1061# 0.02fF
C893 a_149_n389# a_n1555_n1061# 0.03fF
C894 a_n29_n389# a_n1555_n1061# 0.03fF
C895 a_n207_n389# a_n1555_n1061# 0.03fF
C896 a_n385_n389# a_n1555_n1061# 0.02fF
C897 a_n563_n389# a_n1555_n1061# 0.03fF
C898 a_n741_n389# a_n1555_n1061# 0.03fF
C899 a_n919_n389# a_n1555_n1061# 0.04fF
C900 a_n1097_n389# a_n1555_n1061# 0.05fF
C901 a_n1275_n389# a_n1555_n1061# 0.10fF
C902 a_1097_n445# a_n1555_n1061# 0.22fF
C903 a_919_n445# a_n1555_n1061# 0.18fF
C904 a_741_n445# a_n1555_n1061# 0.18fF
C905 a_563_n445# a_n1555_n1061# 0.19fF
C906 a_385_n445# a_n1555_n1061# 0.19fF
C907 a_207_n445# a_n1555_n1061# 0.20fF
C908 a_29_n445# a_n1555_n1061# 0.21fF
C909 a_n149_n445# a_n1555_n1061# 0.21fF
C910 a_n327_n445# a_n1555_n1061# 0.21fF
C911 a_n505_n445# a_n1555_n1061# 0.21fF
C912 a_n683_n445# a_n1555_n1061# 0.21fF
C913 a_n861_n445# a_n1555_n1061# 0.21fF
C914 a_n1039_n445# a_n1555_n1061# 0.22fF
C915 a_n1217_n445# a_n1555_n1061# 0.27fF
C916 a_1217_109# a_n1555_n1061# 0.10fF
C917 a_1039_109# a_n1555_n1061# 0.05fF
C918 a_861_109# a_n1555_n1061# 0.04fF
C919 a_683_109# a_n1555_n1061# 0.03fF
C920 a_505_109# a_n1555_n1061# 0.03fF
C921 a_327_109# a_n1555_n1061# 0.03fF
C922 a_149_109# a_n1555_n1061# 0.03fF
C923 a_n29_109# a_n1555_n1061# 0.03fF
C924 a_n207_109# a_n1555_n1061# 0.03fF
C925 a_n385_109# a_n1555_n1061# 0.03fF
C926 a_n563_109# a_n1555_n1061# 0.03fF
C927 a_n741_109# a_n1555_n1061# 0.03fF
C928 a_n919_109# a_n1555_n1061# 0.04fF
C929 a_n1097_109# a_n1555_n1061# 0.06fF
C930 a_n1275_109# a_n1555_n1061# 0.10fF
C931 a_1097_55# a_n1555_n1061# 0.23fF
C932 a_919_55# a_n1555_n1061# 0.20fF
C933 a_741_55# a_n1555_n1061# 0.20fF
C934 a_563_55# a_n1555_n1061# 0.20fF
C935 a_385_55# a_n1555_n1061# 0.21fF
C936 a_207_55# a_n1555_n1061# 0.21fF
C937 a_29_55# a_n1555_n1061# 0.22fF
C938 a_n149_55# a_n1555_n1061# 0.22fF
C939 a_n327_55# a_n1555_n1061# 0.22fF
C940 a_n505_55# a_n1555_n1061# 0.22fF
C941 a_n683_55# a_n1555_n1061# 0.22fF
C942 a_n861_55# a_n1555_n1061# 0.23fF
C943 a_n1039_55# a_n1555_n1061# 0.23fF
C944 a_n1217_55# a_n1555_n1061# 0.28fF
C945 a_1217_607# a_n1555_n1061# 0.10fF
C946 a_1039_607# a_n1555_n1061# 0.06fF
C947 a_861_607# a_n1555_n1061# 0.05fF
C948 a_683_607# a_n1555_n1061# 0.04fF
C949 a_505_607# a_n1555_n1061# 0.03fF
C950 a_327_607# a_n1555_n1061# 0.03fF
C951 a_149_607# a_n1555_n1061# 0.03fF
C952 a_n29_607# a_n1555_n1061# 0.04fF
C953 a_n207_607# a_n1555_n1061# 0.03fF
C954 a_n385_607# a_n1555_n1061# 0.03fF
C955 a_n563_607# a_n1555_n1061# 0.03fF
C956 a_n741_607# a_n1555_n1061# 0.04fF
C957 a_n919_607# a_n1555_n1061# 0.05fF
C958 a_n1097_607# a_n1555_n1061# 0.06fF
C959 a_n1275_607# a_n1555_n1061# 0.10fF
C960 a_1097_553# a_n1555_n1061# 0.30fF
C961 a_919_553# a_n1555_n1061# 0.26fF
C962 a_741_553# a_n1555_n1061# 0.26fF
C963 a_563_553# a_n1555_n1061# 0.27fF
C964 a_385_553# a_n1555_n1061# 0.27fF
C965 a_207_553# a_n1555_n1061# 0.28fF
C966 a_29_553# a_n1555_n1061# 0.29fF
C967 a_n149_553# a_n1555_n1061# 0.29fF
C968 a_n327_553# a_n1555_n1061# 0.29fF
C969 a_n505_553# a_n1555_n1061# 0.29fF
C970 a_n683_553# a_n1555_n1061# 0.29fF
C971 a_n861_553# a_n1555_n1061# 0.29fF
C972 a_n1039_553# a_n1555_n1061# 0.30fF
C973 a_n1217_553# a_n1555_n1061# 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EL6FQZ a_n1008_n140# a_1306_n140# a_n652_n140# a_652_n194#
+ a_n1662_n194# a_772_n140# a_n1720_n140# a_n60_n194# a_2076_n194# a_1008_n194# a_2196_n140#
+ a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194# a_594_n140# a_n1542_n140#
+ a_1720_n194# a_1840_n140# a_n238_n194# a_n296_n140# a_n1898_n140# a_296_n194# a_2018_n140#
+ a_60_n140# a_n1306_n194# a_n1364_n140# a_1542_n194# a_416_n140# a_n950_n194# a_n2432_n140#
+ a_1662_n140# a_1898_n194# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194# a_238_n140#
+ a_n1186_n140# a_n2254_n140# a_1364_n194# a_n772_n194# a_1484_n140# a_n830_n140#
+ a_830_n194# a_n1840_n194# a_950_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2254_n194# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2254_n140# a_n2432_n140# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_594_n140# a_2196_n140# 0.01fF
C1 a_n1484_n194# a_n2196_n194# 0.01fF
C2 a_n652_n140# a_n1542_n140# 0.01fF
C3 a_n416_n194# a_n1306_n194# 0.01fF
C4 a_n238_n194# a_830_n194# 0.01fF
C5 a_n594_n194# a_n2196_n194# 0.01fF
C6 a_296_n194# a_n1128_n194# 0.01fF
C7 a_238_n140# a_950_n140# 0.01fF
C8 a_1542_n194# a_2076_n194# 0.02fF
C9 a_416_n140# a_n296_n140# 0.01fF
C10 a_474_n194# a_118_n194# 0.03fF
C11 a_n416_n194# a_1008_n194# 0.01fF
C12 a_416_n140# a_1128_n140# 0.01fF
C13 a_n772_n194# a_830_n194# 0.01fF
C14 a_474_n194# a_n594_n194# 0.01fF
C15 a_n1364_n140# a_n2076_n140# 0.01fF
C16 a_60_n140# a_1662_n140# 0.01fF
C17 a_n474_n140# a_n830_n140# 0.03fF
C18 a_1542_n194# a_2254_n194# 0.01fF
C19 a_594_n140# a_772_n140# 0.06fF
C20 a_1364_n194# a_652_n194# 0.01fF
C21 a_1542_n194# a_n60_n194# 0.01fF
C22 a_n772_n194# a_n2018_n194# 0.01fF
C23 a_n1306_n194# a_n238_n194# 0.01fF
C24 a_118_n194# a_1720_n194# 0.01fF
C25 a_118_n194# a_830_n194# 0.01fF
C26 a_652_n194# a_1186_n194# 0.02fF
C27 a_n238_n194# a_1008_n194# 0.01fF
C28 a_n2432_n140# a_n2196_n194# 0.06fF
C29 a_n1306_n194# a_n772_n194# 0.02fF
C30 a_1484_n140# a_1662_n140# 0.06fF
C31 a_60_n140# a_n652_n140# 0.01fF
C32 a_n594_n194# a_830_n194# 0.01fF
C33 a_416_n140# a_1306_n140# 0.01fF
C34 a_n1186_n140# a_n2076_n140# 0.01fF
C35 a_n1484_n194# a_n2018_n194# 0.02fF
C36 a_416_n140# a_n830_n140# 0.01fF
C37 a_416_n140# a_n474_n140# 0.01fF
C38 a_n594_n194# a_n2018_n194# 0.01fF
C39 a_n1898_n140# a_n1542_n140# 0.03fF
C40 a_118_n194# a_n1306_n194# 0.01fF
C41 a_n1484_n194# a_n1306_n194# 0.10fF
C42 a_2018_n140# a_1840_n140# 0.06fF
C43 a_652_n194# a_2076_n194# 0.01fF
C44 a_118_n194# a_1008_n194# 0.01fF
C45 a_n1840_n194# a_n416_n194# 0.01fF
C46 a_n594_n194# a_n1306_n194# 0.01fF
C47 a_1662_n140# a_950_n140# 0.01fF
C48 a_n594_n194# a_1008_n194# 0.01fF
C49 a_2254_n194# a_652_n194# 0.00fF
C50 a_n2254_n140# a_n1542_n140# 0.01fF
C51 a_n1128_n194# a_n2196_n194# 0.01fF
C52 a_n60_n194# a_652_n194# 0.01fF
C53 a_2018_n140# a_2254_n194# 0.03fF
C54 a_238_n140# a_1662_n140# 0.01fF
C55 a_n1008_n140# a_n2076_n140# 0.01fF
C56 a_1484_n140# a_2196_n140# 0.01fF
C57 a_n2432_n140# a_n2018_n194# 0.02fF
C58 a_n1840_n194# a_n238_n194# 0.01fF
C59 a_n652_n140# a_950_n140# 0.01fF
C60 a_474_n194# a_296_n194# 0.10fF
C61 a_474_n194# a_n1128_n194# 0.01fF
C62 a_60_n140# a_772_n140# 0.01fF
C63 a_594_n140# a_n118_n140# 0.01fF
C64 a_n1306_n194# a_n2432_n140# 0.01fF
C65 a_n1840_n194# a_n772_n194# 0.01fF
C66 a_n416_n194# a_1186_n194# 0.01fF
C67 a_238_n140# a_n652_n140# 0.01fF
C68 a_n1898_n140# a_n2432_n140# 0.02fF
C69 a_1484_n140# a_772_n140# 0.01fF
C70 a_1720_n194# a_296_n194# 0.01fF
C71 a_1128_n140# a_2018_n140# 0.01fF
C72 a_296_n194# a_830_n194# 0.02fF
C73 a_950_n140# a_2196_n140# 0.01fF
C74 a_n1720_n140# a_n652_n140# 0.01fF
C75 a_n238_n194# a_1364_n194# 0.01fF
C76 a_652_n194# a_n950_n194# 0.01fF
C77 a_n1484_n194# a_n1840_n194# 0.03fF
C78 a_n238_n194# a_1186_n194# 0.01fF
C79 a_296_n194# a_1898_n194# 0.01fF
C80 a_n1840_n194# a_n594_n194# 0.01fF
C81 a_n2254_n140# a_n2432_n140# 0.06fF
C82 a_n118_n140# a_n1542_n140# 0.01fF
C83 a_n1128_n194# a_n2018_n194# 0.01fF
C84 a_n1364_n140# a_n1542_n140# 0.06fF
C85 a_594_n140# a_1840_n140# 0.01fF
C86 a_n1306_n194# a_296_n194# 0.01fF
C87 a_n1306_n194# a_n1128_n194# 0.10fF
C88 a_1306_n140# a_2018_n140# 0.01fF
C89 a_772_n140# a_950_n140# 0.06fF
C90 a_n2076_n140# a_n830_n140# 0.01fF
C91 a_118_n194# a_1364_n194# 0.01fF
C92 a_296_n194# a_1008_n194# 0.01fF
C93 a_n416_n194# a_n60_n194# 0.03fF
C94 a_n474_n140# a_n2076_n140# 0.01fF
C95 a_n1662_n194# a_n416_n194# 0.01fF
C96 a_118_n194# a_1186_n194# 0.01fF
C97 a_238_n140# a_772_n140# 0.02fF
C98 a_n1840_n194# a_n2432_n140# 0.01fF
C99 a_n1186_n140# a_n1542_n140# 0.03fF
C100 a_60_n140# a_n118_n140# 0.06fF
C101 a_594_n140# a_n1008_n140# 0.01fF
C102 a_n1720_n140# a_n1898_n140# 0.06fF
C103 a_60_n140# a_n1364_n140# 0.01fF
C104 a_n60_n194# a_n238_n194# 0.10fF
C105 a_n1662_n194# a_n238_n194# 0.01fF
C106 a_n60_n194# a_n772_n194# 0.01fF
C107 a_416_n140# a_2018_n140# 0.01fF
C108 a_n1364_n140# a_n2432_n140# 0.01fF
C109 a_n1662_n194# a_n772_n194# 0.01fF
C110 a_1484_n140# a_n118_n140# 0.01fF
C111 a_n416_n194# a_n950_n194# 0.02fF
C112 a_594_n140# a_n296_n140# 0.01fF
C113 a_594_n140# a_1128_n140# 0.02fF
C114 a_1662_n140# a_2196_n140# 0.02fF
C115 a_n2254_n140# a_n1720_n140# 0.02fF
C116 a_474_n194# a_1720_n194# 0.01fF
C117 a_n1008_n140# a_n1542_n140# 0.02fF
C118 a_118_n194# a_n60_n194# 0.10fF
C119 a_n1186_n140# a_60_n140# 0.01fF
C120 a_n1484_n194# a_n60_n194# 0.01fF
C121 a_n1840_n194# a_n1128_n194# 0.01fF
C122 a_474_n194# a_830_n194# 0.03fF
C123 a_n1484_n194# a_n1662_n194# 0.10fF
C124 a_n2018_n194# a_n2196_n194# 0.10fF
C125 a_n238_n194# a_n950_n194# 0.01fF
C126 a_n594_n194# a_n60_n194# 0.02fF
C127 a_n1662_n194# a_n594_n194# 0.01fF
C128 a_n1186_n140# a_n2432_n140# 0.01fF
C129 a_474_n194# a_1898_n194# 0.01fF
C130 a_n118_n140# a_950_n140# 0.01fF
C131 a_n1306_n194# a_n2196_n194# 0.01fF
C132 a_n296_n140# a_n1542_n140# 0.01fF
C133 a_n772_n194# a_n950_n194# 0.10fF
C134 a_772_n140# a_1662_n140# 0.01fF
C135 a_1306_n140# a_594_n140# 0.01fF
C136 a_1542_n194# a_652_n194# 0.01fF
C137 a_1720_n194# a_830_n194# 0.01fF
C138 a_1484_n140# a_1840_n140# 0.03fF
C139 a_238_n140# a_n118_n140# 0.03fF
C140 a_296_n194# a_1364_n194# 0.01fF
C141 a_594_n140# a_n830_n140# 0.01fF
C142 a_594_n140# a_n474_n140# 0.01fF
C143 a_238_n140# a_n1364_n140# 0.01fF
C144 a_1720_n194# a_1898_n194# 0.10fF
C145 a_474_n194# a_1008_n194# 0.02fF
C146 a_60_n140# a_n1008_n140# 0.01fF
C147 a_296_n194# a_1186_n194# 0.01fF
C148 a_772_n140# a_n652_n140# 0.01fF
C149 a_118_n194# a_n950_n194# 0.01fF
C150 a_n1898_n140# a_n652_n140# 0.01fF
C151 a_830_n194# a_1898_n194# 0.01fF
C152 a_n1484_n194# a_n950_n194# 0.02fF
C153 a_n1720_n140# a_n118_n140# 0.01fF
C154 a_n1662_n194# a_n2432_n140# 0.01fF
C155 a_1484_n140# a_2254_n194# 0.01fF
C156 a_n594_n194# a_n950_n194# 0.03fF
C157 a_n1008_n140# a_n2432_n140# 0.01fF
C158 a_n1364_n140# a_n1720_n140# 0.03fF
C159 a_60_n140# a_n296_n140# 0.03fF
C160 a_1720_n194# a_1008_n194# 0.01fF
C161 a_1840_n140# a_950_n140# 0.01fF
C162 a_60_n140# a_1128_n140# 0.01fF
C163 a_1008_n194# a_830_n194# 0.10fF
C164 a_416_n140# a_594_n140# 0.06fF
C165 a_n830_n140# a_n1542_n140# 0.01fF
C166 a_n2254_n140# a_n652_n140# 0.01fF
C167 a_n1186_n140# a_238_n140# 0.01fF
C168 a_n474_n140# a_n1542_n140# 0.01fF
C169 a_772_n140# a_2196_n140# 0.01fF
C170 a_n1306_n194# a_n2018_n194# 0.01fF
C171 a_238_n140# a_1840_n140# 0.01fF
C172 a_1008_n194# a_1898_n194# 0.01fF
C173 a_1484_n140# a_1128_n140# 0.03fF
C174 a_2254_n194# a_950_n140# 0.01fF
C175 a_n1840_n194# a_n2196_n194# 0.03fF
C176 a_n1186_n140# a_n1720_n140# 0.02fF
C177 a_n2432_n140# a_n950_n194# 0.00fF
C178 a_n60_n194# a_296_n194# 0.03fF
C179 a_n60_n194# a_n1128_n194# 0.01fF
C180 a_n1662_n194# a_n1128_n194# 0.02fF
C181 a_1306_n140# a_60_n140# 0.01fF
C182 a_60_n140# a_n830_n140# 0.01fF
C183 a_238_n140# a_n1008_n140# 0.01fF
C184 a_60_n140# a_n474_n140# 0.02fF
C185 a_n296_n140# a_950_n140# 0.01fF
C186 a_1306_n140# a_1484_n140# 0.06fF
C187 a_1128_n140# a_950_n140# 0.06fF
C188 a_n830_n140# a_n2432_n140# 0.01fF
C189 a_n118_n140# a_n652_n140# 0.02fF
C190 a_n1008_n140# a_n1720_n140# 0.01fF
C191 a_n2254_n140# a_n1898_n140# 0.03fF
C192 a_n1364_n140# a_n652_n140# 0.01fF
C193 a_238_n140# a_n296_n140# 0.02fF
C194 a_474_n194# a_1364_n194# 0.01fF
C195 a_238_n140# a_1128_n140# 0.01fF
C196 a_296_n194# a_n950_n194# 0.01fF
C197 a_n950_n194# a_n1128_n194# 0.10fF
C198 a_474_n194# a_1186_n194# 0.01fF
C199 a_416_n140# a_60_n140# 0.03fF
C200 a_n1840_n194# a_n2018_n194# 0.10fF
C201 a_n1720_n140# a_n296_n140# 0.01fF
C202 a_1662_n140# a_1840_n140# 0.06fF
C203 a_1720_n194# a_1364_n194# 0.03fF
C204 a_1306_n140# a_950_n140# 0.03fF
C205 a_n1840_n194# a_n1306_n194# 0.02fF
C206 a_1364_n194# a_830_n194# 0.02fF
C207 a_1542_n194# a_118_n194# 0.01fF
C208 a_n416_n194# a_652_n194# 0.01fF
C209 a_1720_n194# a_1186_n194# 0.02fF
C210 a_n1186_n140# a_n652_n140# 0.02fF
C211 a_416_n140# a_1484_n140# 0.01fF
C212 a_1306_n140# a_238_n140# 0.01fF
C213 a_830_n194# a_1186_n194# 0.03fF
C214 a_n474_n140# a_950_n140# 0.01fF
C215 a_1364_n194# a_1898_n194# 0.02fF
C216 a_1662_n140# a_2254_n194# 0.01fF
C217 a_474_n194# a_2076_n194# 0.01fF
C218 a_238_n140# a_n830_n140# 0.01fF
C219 a_1898_n194# a_1186_n194# 0.01fF
C220 a_594_n140# a_2018_n140# 0.01fF
C221 a_n1662_n194# a_n2196_n194# 0.02fF
C222 a_238_n140# a_n474_n140# 0.01fF
C223 a_772_n140# a_n118_n140# 0.01fF
C224 a_n238_n194# a_652_n194# 0.01fF
C225 a_n1364_n140# a_n1898_n140# 0.02fF
C226 a_474_n194# a_n60_n194# 0.02fF
C227 a_1008_n194# a_1364_n194# 0.03fF
C228 a_1720_n194# a_2076_n194# 0.03fF
C229 a_n1720_n140# a_n830_n140# 0.01fF
C230 a_n772_n194# a_652_n194# 0.01fF
C231 a_n474_n140# a_n1720_n140# 0.01fF
C232 a_416_n140# a_950_n140# 0.02fF
C233 a_830_n194# a_2076_n194# 0.01fF
C234 a_1840_n140# a_2196_n140# 0.03fF
C235 a_n1008_n140# a_n652_n140# 0.03fF
C236 a_1008_n194# a_1186_n194# 0.10fF
C237 a_1128_n140# a_1662_n140# 0.02fF
C238 a_n2076_n140# a_n1542_n140# 0.02fF
C239 a_2076_n194# a_1898_n194# 0.10fF
C240 a_1720_n194# a_2254_n194# 0.01fF
C241 a_416_n140# a_238_n140# 0.06fF
C242 a_n1364_n140# a_n2254_n140# 0.01fF
C243 a_2254_n194# a_830_n194# 0.00fF
C244 a_n60_n194# a_830_n194# 0.01fF
C245 a_118_n194# a_652_n194# 0.02fF
C246 a_n950_n194# a_n2196_n194# 0.01fF
C247 a_2254_n194# a_2196_n140# 0.06fF
C248 a_n652_n140# a_n296_n140# 0.03fF
C249 a_n1186_n140# a_n1898_n140# 0.01fF
C250 a_2254_n194# a_1898_n194# 0.02fF
C251 a_n594_n194# a_652_n194# 0.01fF
C252 a_772_n140# a_1840_n140# 0.01fF
C253 a_474_n194# a_n950_n194# 0.01fF
C254 a_1008_n194# a_2076_n194# 0.01fF
C255 a_n1662_n194# a_n2018_n194# 0.03fF
C256 a_1306_n140# a_1662_n140# 0.03fF
C257 a_n60_n194# a_n1306_n194# 0.01fF
C258 a_n1186_n140# a_n2254_n140# 0.01fF
C259 a_n1662_n194# a_n1306_n194# 0.03fF
C260 a_2254_n194# a_1008_n194# 0.00fF
C261 a_772_n140# a_2254_n194# 0.01fF
C262 a_1542_n194# a_296_n194# 0.01fF
C263 a_n60_n194# a_1008_n194# 0.01fF
C264 a_1128_n140# a_2196_n140# 0.01fF
C265 a_n1008_n140# a_n1898_n140# 0.01fF
C266 a_n416_n194# a_n238_n194# 0.10fF
C267 a_n2076_n140# a_n2432_n140# 0.03fF
C268 a_n1364_n140# a_n118_n140# 0.01fF
C269 a_n652_n140# a_n830_n140# 0.06fF
C270 a_n416_n194# a_n772_n194# 0.03fF
C271 a_n474_n140# a_n652_n140# 0.06fF
C272 a_1484_n140# a_2018_n140# 0.02fF
C273 a_n950_n194# a_n2018_n194# 0.01fF
C274 a_n1898_n140# a_n296_n140# 0.01fF
C275 a_772_n140# a_n296_n140# 0.01fF
C276 a_416_n140# a_1662_n140# 0.01fF
C277 a_1128_n140# a_772_n140# 0.03fF
C278 a_n2254_n140# a_n1008_n140# 0.01fF
C279 a_n1306_n194# a_n950_n194# 0.03fF
C280 a_1306_n140# a_2196_n140# 0.01fF
C281 a_n416_n194# a_118_n194# 0.02fF
C282 a_1364_n194# a_1186_n194# 0.10fF
C283 a_n1484_n194# a_n416_n194# 0.01fF
C284 a_n238_n194# a_n772_n194# 0.02fF
C285 a_n416_n194# a_n594_n194# 0.10fF
C286 a_n1186_n140# a_n118_n140# 0.01fF
C287 a_416_n140# a_n652_n140# 0.01fF
C288 a_n1186_n140# a_n1364_n140# 0.06fF
C289 a_2018_n140# a_950_n140# 0.01fF
C290 a_296_n194# a_652_n194# 0.03fF
C291 a_n1662_n194# a_n1840_n194# 0.10fF
C292 a_1306_n140# a_772_n140# 0.02fF
C293 a_118_n194# a_n238_n194# 0.03fF
C294 a_n1484_n194# a_n238_n194# 0.01fF
C295 a_1364_n194# a_2076_n194# 0.01fF
C296 a_n1898_n140# a_n830_n140# 0.01fF
C297 a_772_n140# a_n830_n140# 0.01fF
C298 a_n594_n194# a_n238_n194# 0.03fF
C299 a_118_n194# a_n772_n194# 0.01fF
C300 a_n474_n140# a_772_n140# 0.01fF
C301 a_n474_n140# a_n1898_n140# 0.01fF
C302 a_n1484_n194# a_n772_n194# 0.01fF
C303 a_2076_n194# a_1186_n194# 0.01fF
C304 a_n1720_n140# a_n2076_n140# 0.03fF
C305 a_60_n140# a_594_n140# 0.02fF
C306 a_n594_n194# a_n772_n194# 0.10fF
C307 a_2254_n194# a_1364_n194# 0.01fF
C308 a_n1008_n140# a_n118_n140# 0.01fF
C309 a_n60_n194# a_1364_n194# 0.01fF
C310 a_n1364_n140# a_n1008_n140# 0.03fF
C311 a_474_n194# a_1542_n194# 0.01fF
C312 a_2254_n194# a_1186_n194# 0.01fF
C313 a_n60_n194# a_1186_n194# 0.01fF
C314 a_n2254_n140# a_n830_n140# 0.01fF
C315 a_n1840_n194# a_n950_n194# 0.01fF
C316 a_n1484_n194# a_118_n194# 0.01fF
C317 a_1484_n140# a_594_n140# 0.01fF
C318 a_n594_n194# a_118_n194# 0.01fF
C319 a_n118_n140# a_n296_n140# 0.06fF
C320 a_n1484_n194# a_n594_n194# 0.01fF
C321 a_416_n140# a_772_n140# 0.03fF
C322 a_1128_n140# a_n118_n140# 0.01fF
C323 a_n1364_n140# a_n296_n140# 0.01fF
C324 a_1542_n194# a_1720_n194# 0.10fF
C325 a_n772_n194# a_n2432_n140# 0.00fF
C326 a_60_n140# a_n1542_n140# 0.01fF
C327 a_1542_n194# a_830_n194# 0.01fF
C328 a_2254_n194# a_1840_n140# 0.02fF
C329 a_n1186_n140# a_n1008_n140# 0.06fF
C330 a_2254_n194# a_2076_n194# 0.06fF
C331 a_n416_n194# a_296_n194# 0.01fF
C332 a_n416_n194# a_n1128_n194# 0.01fF
C333 a_1542_n194# a_1898_n194# 0.03fF
C334 a_n2432_n140# a_n1542_n140# 0.01fF
C335 a_2018_n140# a_1662_n140# 0.03fF
C336 a_594_n140# a_950_n140# 0.03fF
C337 a_1306_n140# a_n118_n140# 0.01fF
C338 a_n1484_n194# a_n2432_n140# 0.01fF
C339 a_n1186_n140# a_n296_n140# 0.01fF
C340 a_n1662_n194# a_n60_n194# 0.01fF
C341 a_n2076_n140# a_n652_n140# 0.01fF
C342 a_n118_n140# a_n830_n140# 0.01fF
C343 a_238_n140# a_594_n140# 0.03fF
C344 a_474_n194# a_652_n194# 0.10fF
C345 a_1128_n140# a_1840_n140# 0.01fF
C346 a_1542_n194# a_1008_n194# 0.02fF
C347 a_296_n194# a_n238_n194# 0.02fF
C348 a_n474_n140# a_n118_n140# 0.03fF
C349 a_n238_n194# a_n1128_n194# 0.01fF
C350 a_n1364_n140# a_n830_n140# 0.02fF
C351 a_n1364_n140# a_n474_n140# 0.01fF
C352 a_296_n194# a_n772_n194# 0.01fF
C353 a_n772_n194# a_n1128_n194# 0.03fF
C354 a_1720_n194# a_652_n194# 0.01fF
C355 a_1128_n140# a_2254_n194# 0.01fF
C356 a_60_n140# a_1484_n140# 0.01fF
C357 a_830_n194# a_652_n194# 0.10fF
C358 a_n1008_n140# a_n296_n140# 0.01fF
C359 a_416_n140# a_n118_n140# 0.02fF
C360 a_118_n194# a_296_n194# 0.10fF
C361 a_1306_n140# a_1840_n140# 0.02fF
C362 a_118_n194# a_n1128_n194# 0.01fF
C363 a_n60_n194# a_n950_n194# 0.01fF
C364 a_2018_n140# a_2196_n140# 0.06fF
C365 a_652_n194# a_1898_n194# 0.01fF
C366 a_n1662_n194# a_n950_n194# 0.01fF
C367 a_n1484_n194# a_n1128_n194# 0.03fF
C368 a_n1186_n140# a_n830_n140# 0.03fF
C369 a_n594_n194# a_296_n194# 0.01fF
C370 a_n1186_n140# a_n474_n140# 0.01fF
C371 a_n594_n194# a_n1128_n194# 0.02fF
C372 a_n1720_n140# a_n1542_n140# 0.06fF
C373 a_1128_n140# a_n296_n140# 0.01fF
C374 a_1306_n140# a_2254_n194# 0.01fF
C375 a_n1898_n140# a_n2076_n140# 0.06fF
C376 a_1008_n194# a_652_n194# 0.03fF
C377 a_60_n140# a_950_n140# 0.01fF
C378 a_772_n140# a_2018_n140# 0.01fF
C379 a_594_n140# a_1662_n140# 0.01fF
C380 a_474_n194# a_n416_n194# 0.01fF
C381 a_416_n140# a_n1186_n140# 0.01fF
C382 a_60_n140# a_238_n140# 0.06fF
C383 a_n1008_n140# a_n830_n140# 0.06fF
C384 a_416_n140# a_1840_n140# 0.01fF
C385 a_n474_n140# a_n1008_n140# 0.02fF
C386 a_n2432_n140# a_n1128_n194# 0.00fF
C387 a_1484_n140# a_950_n140# 0.02fF
C388 a_n2254_n140# a_n2076_n140# 0.06fF
C389 a_1306_n140# a_n296_n140# 0.01fF
C390 a_594_n140# a_n652_n140# 0.01fF
C391 a_1306_n140# a_1128_n140# 0.06fF
C392 a_1542_n194# a_1364_n194# 0.10fF
C393 a_238_n140# a_1484_n140# 0.01fF
C394 a_n772_n194# a_n2196_n194# 0.01fF
C395 a_n296_n140# a_n830_n140# 0.02fF
C396 a_474_n194# a_n238_n194# 0.01fF
C397 a_n416_n194# a_830_n194# 0.01fF
C398 a_1542_n194# a_1186_n194# 0.03fF
C399 a_n474_n140# a_n296_n140# 0.06fF
C400 a_1128_n140# a_n474_n140# 0.01fF
C401 a_n1720_n140# a_n2432_n140# 0.01fF
C402 a_474_n194# a_n772_n194# 0.01fF
C403 a_416_n140# a_n1008_n140# 0.01fF
C404 a_n416_n194# a_n2018_n194# 0.01fF
C405 a_2196_n140# VSUBS 0.01fF
C406 a_2018_n140# VSUBS 0.01fF
C407 a_1840_n140# VSUBS 0.02fF
C408 a_1662_n140# VSUBS 0.02fF
C409 a_1484_n140# VSUBS 0.02fF
C410 a_1306_n140# VSUBS 0.02fF
C411 a_1128_n140# VSUBS 0.02fF
C412 a_950_n140# VSUBS 0.02fF
C413 a_772_n140# VSUBS 0.02fF
C414 a_594_n140# VSUBS 0.02fF
C415 a_416_n140# VSUBS 0.02fF
C416 a_238_n140# VSUBS 0.02fF
C417 a_60_n140# VSUBS 0.02fF
C418 a_n118_n140# VSUBS 0.02fF
C419 a_n296_n140# VSUBS 0.02fF
C420 a_n474_n140# VSUBS 0.02fF
C421 a_n652_n140# VSUBS 0.02fF
C422 a_n830_n140# VSUBS 0.02fF
C423 a_n1008_n140# VSUBS 0.02fF
C424 a_n1186_n140# VSUBS 0.02fF
C425 a_n1364_n140# VSUBS 0.02fF
C426 a_n1542_n140# VSUBS 0.02fF
C427 a_n1720_n140# VSUBS 0.02fF
C428 a_n1898_n140# VSUBS 0.02fF
C429 a_n2076_n140# VSUBS 0.02fF
C430 a_n2254_n140# VSUBS 0.02fF
C431 a_2254_n194# VSUBS 0.31fF
C432 a_2076_n194# VSUBS 0.19fF
C433 a_1898_n194# VSUBS 0.20fF
C434 a_1720_n194# VSUBS 0.21fF
C435 a_1542_n194# VSUBS 0.22fF
C436 a_1364_n194# VSUBS 0.23fF
C437 a_1186_n194# VSUBS 0.23fF
C438 a_1008_n194# VSUBS 0.24fF
C439 a_830_n194# VSUBS 0.24fF
C440 a_652_n194# VSUBS 0.24fF
C441 a_474_n194# VSUBS 0.24fF
C442 a_296_n194# VSUBS 0.24fF
C443 a_118_n194# VSUBS 0.24fF
C444 a_n60_n194# VSUBS 0.24fF
C445 a_n238_n194# VSUBS 0.24fF
C446 a_n416_n194# VSUBS 0.24fF
C447 a_n594_n194# VSUBS 0.24fF
C448 a_n772_n194# VSUBS 0.24fF
C449 a_n950_n194# VSUBS 0.24fF
C450 a_n1128_n194# VSUBS 0.24fF
C451 a_n1306_n194# VSUBS 0.24fF
C452 a_n1484_n194# VSUBS 0.24fF
C453 a_n1662_n194# VSUBS 0.24fF
C454 a_n1840_n194# VSUBS 0.24fF
C455 a_n2018_n194# VSUBS 0.24fF
C456 a_n2196_n194# VSUBS 0.24fF
C457 a_n2432_n140# VSUBS 0.36fF
.ends

.subckt bias_circuit bias_c bias_e i_bias VDD m1_1243_5997# m1_3443_5997# bias_a m1_7347_1428#
+ m1_7639_1420# m1_7169_923# m1_7461_921# m1_7347_423# m1_7639_427# bias_b VSS m1_3551_3596#
+ m1_5643_5997# bias_d
Xsky130_fd_pr__nfet_01v8_6RUDQZ_0 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_1 bias_a VSS VSS bias_a VSS bias_a li_3433_399# bias_a
+ bias_a li_3433_399# VSS bias_a VSS bias_a VSS li_3433_399# bias_a li_3433_399# bias_a
+ li_3433_399# VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_2 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_6RUDQZ_3 bias_d VSS li_3433_399# bias_d li_3433_399# bias_d
+ bias_a bias_d bias_d bias_a li_3433_399# bias_d li_3433_399# bias_d li_3433_399#
+ bias_a bias_d bias_a bias_d bias_a VSS VSS sky130_fd_pr__nfet_01v8_6RUDQZ
Xsky130_fd_pr__nfet_01v8_SD55Q9_0 m1_7347_1428# m1_7639_1420# bias_e m1_7055_1417#
+ bias_e m1_6763_422# bias_e m1_6471_422# bias_e VSS VSS VSS m1_7639_427# m1_7347_423#
+ m1_7055_433# bias_e bias_e bias_e m1_6763_422# m1_6471_422# m1_7169_923# bias_e
+ m1_7461_921# bias_e bias_e m1_7639_427# m1_7347_423# m1_6877_922# m1_7055_433# VSS
+ bias_e VSS VSS bias_e bias_e bias_e m1_6877_922# m1_6585_923# VSS bias_e m1_6763_1422#
+ m1_6293_922# bias_e m1_6471_1426# m1_7347_1428# bias_e bias_e m1_7639_1420# m1_7169_923#
+ m1_7055_1417# bias_e bias_e m1_7461_921# bias_e bias_e bias_e m1_6585_923# bias_e
+ m1_6293_922# m1_6763_1422# bias_e m1_6471_1426# VSS sky130_fd_pr__nfet_01v8_SD55Q9
Xsky130_fd_pr__nfet_01v8_EZNTQN_0 bias_c VSS VSS i_bias i_bias i_bias i_bias VSS VSS
+ bias_c VSS VSS i_bias VSS bias_c i_bias i_bias i_bias i_bias VSS i_bias i_bias bias_c
+ i_bias VSS VSS i_bias i_bias i_bias bias_c VSS VSS i_bias bias_c VSS i_bias i_bias
+ VSS i_bias i_bias i_bias i_bias i_bias VSS i_bias i_bias i_bias i_bias i_bias i_bias
+ i_bias bias_c i_bias VSS i_bias i_bias bias_c i_bias i_bias i_bias i_bias VSS i_bias
+ VSS i_bias VSS VSS i_bias i_bias bias_c i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ sky130_fd_pr__nfet_01v8_EZNTQN
Xsky130_fd_pr__pfet_01v8_JJWXCM_0 bias_b bias_c m1_1243_5997# m1_1243_5997# bias_b
+ bias_c VDD VDD bias_c bias_b bias_c VDD bias_c m1_1243_5997# bias_c bias_b VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_1 m1_3551_3596# bias_c m1_3443_5997# m1_3443_5997#
+ m1_3551_3596# bias_c VDD VDD bias_c m1_3551_3596# bias_c VDD bias_c m1_3443_5997#
+ bias_c m1_3551_3596# VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__pfet_01v8_JJWXCM_2 bias_e bias_c m1_5643_5997# m1_5643_5997# bias_e
+ bias_c VDD VDD bias_c bias_e bias_c VDD bias_c m1_5643_5997# bias_c bias_e VSS sky130_fd_pr__pfet_01v8_JJWXCM
Xsky130_fd_pr__nfet_01v8_LJREPQ_0 m1_3551_3596# bias_d VSS bias_a bias_d m1_3551_3596#
+ VSS VSS sky130_fd_pr__nfet_01v8_LJREPQ
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_0 m1_1243_5997# bias_b VDD VDD m1_1243_5997# bias_b
+ VDD VDD bias_b bias_b m1_1243_5997# bias_b VDD VDD bias_b m1_1243_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_1 m1_3443_5997# bias_b VDD VDD m1_3443_5997# bias_b
+ VDD VDD bias_b bias_b m1_3443_5997# bias_b VDD VDD bias_b m1_3443_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__pfet_01v8_lvt_SAWXCM_2 m1_5643_5997# bias_b VDD VDD m1_5643_5997# bias_b
+ VDD VDD bias_b bias_b m1_5643_5997# bias_b VDD VDD bias_b m1_5643_5997# VSS sky130_fd_pr__pfet_01v8_lvt_SAWXCM
Xsky130_fd_pr__nfet_01v8_lvt_28TRYY_0 bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b VSS bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_c bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_c bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_b bias_c bias_b bias_b bias_b
+ bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_c
+ bias_c bias_b bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b bias_c
+ bias_b bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_b bias_b bias_b bias_c bias_c bias_c bias_b bias_b bias_c bias_b
+ bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b bias_b bias_b bias_b bias_b
+ bias_b bias_b sky130_fd_pr__nfet_01v8_lvt_28TRYY
Xsky130_fd_pr__nfet_01v8_EL6FQZ_0 bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d VSS m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
Xsky130_fd_pr__nfet_01v8_EL6FQZ_1 bias_d m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596#
+ bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d
+ m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596#
+ bias_d m1_3551_3596# bias_d m1_3551_3596# VSS m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d m1_3551_3596# m1_3551_3596# m1_3551_3596# m1_3551_3596#
+ m1_3551_3596# m1_3551_3596# bias_d VSS m1_3551_3596# VSS sky130_fd_pr__nfet_01v8_EL6FQZ
C0 m1_6471_1426# bias_d 0.01fF
C1 m1_7055_1417# m1_7055_433# -0.00fF
C2 li_3433_399# m1_6471_1426# 0.01fF
C3 li_3433_399# bias_d 5.36fF
C4 VDD m1_3443_5997# 0.84fF
C5 m1_6471_422# bias_a 0.01fF
C6 bias_b m1_5643_5997# 0.63fF
C7 m1_6763_422# m1_6471_422# 0.03fF
C8 bias_e m1_6471_422# 0.25fF
C9 m1_6471_1426# m1_7347_1428# 0.01fF
C10 m1_3443_5997# bias_c 0.44fF
C11 bias_d m1_7347_1428# 0.00fF
C12 bias_b bias_d 0.26fF
C13 m1_7055_433# m1_7347_423# 0.03fF
C14 VDD m1_1243_5997# 1.50fF
C15 m1_3551_3596# m1_5643_5997# 0.08fF
C16 bias_e m1_3443_5997# 0.02fF
C17 bias_a m1_7055_433# 0.01fF
C18 m1_3551_3596# bias_d 18.83fF
C19 m1_6763_422# m1_7055_433# 0.03fF
C20 m1_1243_5997# bias_c 0.52fF
C21 bias_e m1_7055_433# 0.26fF
C22 m1_3551_3596# li_3433_399# 0.03fF
C23 m1_7055_1417# bias_a 0.00fF
C24 m1_7055_1417# m1_6763_1422# 0.03fF
C25 m1_7639_427# m1_6471_422# 0.01fF
C26 VDD bias_c 4.90fF
C27 bias_e m1_7055_1417# 0.33fF
C28 m1_7055_1417# m1_7639_1420# 0.01fF
C29 bias_b m1_3551_3596# 0.71fF
C30 bias_e VDD 0.26fF
C31 m1_6585_923# bias_a 0.00fF
C32 m1_6471_422# m1_6471_1426# -0.00fF
C33 li_3433_399# m1_6471_422# 0.01fF
C34 bias_a m1_7347_423# 0.01fF
C35 bias_e m1_6585_923# 0.22fF
C36 bias_a bias_c 0.02fF
C37 m1_6763_422# m1_7347_423# 0.01fF
C38 bias_e m1_7347_423# 0.26fF
C39 m1_3443_5997# m1_5643_5997# 0.11fF
C40 m1_7639_427# m1_7055_433# 0.01fF
C41 i_bias bias_c 5.62fF
C42 bias_e bias_c 0.65fF
C43 m1_6585_923# m1_7169_923# 0.01fF
C44 bias_a m1_6763_1422# 0.00fF
C45 m1_3443_5997# bias_d 0.03fF
C46 i_bias bias_a 0.02fF
C47 m1_6763_422# bias_a 0.01fF
C48 bias_e bias_a 0.24fF
C49 bias_a m1_7639_1420# 0.00fF
C50 m1_6763_422# m1_6763_1422# -0.00fF
C51 bias_e m1_6763_1422# 0.33fF
C52 m1_6763_1422# m1_7639_1420# 0.01fF
C53 m1_6293_922# m1_6585_923# 0.03fF
C54 bias_e m1_6763_422# 0.26fF
C55 bias_e m1_7639_1420# 0.18fF
C56 bias_a m1_7169_923# 0.00fF
C57 m1_7055_1417# m1_6471_1426# 0.01fF
C58 m1_6585_923# m1_6877_922# 0.03fF
C59 m1_7055_1417# bias_d 0.00fF
C60 bias_e m1_7169_923# 0.22fF
C61 VDD m1_5643_5997# 1.16fF
C62 bias_b m1_3443_5997# 0.65fF
C63 m1_6293_922# bias_a 0.01fF
C64 m1_7639_427# m1_7347_423# 0.03fF
C65 bias_e m1_6293_922# 0.18fF
C66 VDD bias_d 0.07fF
C67 m1_6877_922# bias_a 0.00fF
C68 m1_5643_5997# bias_c 0.44fF
C69 m1_6585_923# bias_d 0.00fF
C70 m1_7639_427# bias_a 0.01fF
C71 m1_7055_1417# m1_7347_1428# 0.03fF
C72 li_3433_399# m1_6585_923# 0.01fF
C73 bias_e m1_6877_922# 0.22fF
C74 m1_6293_922# m1_7169_923# 0.01fF
C75 m1_3551_3596# m1_3443_5997# 0.98fF
C76 m1_6585_923# m1_7461_921# 0.01fF
C77 m1_6763_422# m1_7639_427# 0.01fF
C78 bias_e m1_7639_427# 0.18fF
C79 m1_7639_427# m1_7639_1420# -0.00fF
C80 bias_b m1_1243_5997# 0.77fF
C81 bias_c bias_d 0.90fF
C82 bias_e m1_5643_5997# 0.71fF
C83 m1_6877_922# m1_7169_923# 0.03fF
C84 bias_a m1_6471_1426# 0.01fF
C85 bias_b VDD 8.29fF
C86 bias_a bias_d 7.33fF
C87 m1_6471_1426# m1_6763_1422# 0.03fF
C88 li_3433_399# bias_a 7.53fF
C89 m1_6763_1422# bias_d 0.00fF
C90 bias_e m1_6471_1426# 0.34fF
C91 i_bias bias_d 0.00fF
C92 bias_a m1_7461_921# 0.00fF
C93 m1_6471_1426# m1_7639_1420# 0.01fF
C94 bias_e bias_d 0.26fF
C95 li_3433_399# i_bias 0.03fF
C96 bias_d m1_7639_1420# 0.00fF
C97 m1_6293_922# m1_6877_922# 0.01fF
C98 bias_e li_3433_399# 0.02fF
C99 m1_7347_423# m1_7347_1428# -0.00fF
C100 m1_3551_3596# m1_1243_5997# 0.03fF
C101 bias_e m1_7461_921# 0.21fF
C102 bias_b bias_c 22.44fF
C103 m1_3551_3596# VDD 0.64fF
C104 m1_6471_422# m1_7055_433# 0.01fF
C105 bias_a m1_7347_1428# 0.00fF
C106 m1_7169_923# m1_7461_921# 0.03fF
C107 m1_6763_1422# m1_7347_1428# 0.01fF
C108 bias_b i_bias 0.60fF
C109 bias_e m1_7347_1428# 0.32fF
C110 m1_6293_922# bias_d 0.00fF
C111 m1_7347_1428# m1_7639_1420# 0.03fF
C112 bias_e bias_b 0.07fF
C113 m1_6293_922# li_3433_399# 0.02fF
C114 m1_6293_922# m1_7461_921# 0.01fF
C115 m1_3551_3596# bias_c 2.13fF
C116 m1_3551_3596# bias_a 0.26fF
C117 m1_6877_922# m1_7461_921# 0.01fF
C118 bias_e m1_3551_3596# 0.76fF
C119 m1_5643_5997# bias_d 0.03fF
C120 m1_6471_422# m1_7347_423# 0.01fF
C121 m1_1243_5997# m1_3443_5997# 0.07fF
C122 m1_3551_3596# VSS -340.53fF
C123 bias_b VSS -284.38fF
C124 m1_5643_5997# VSS 38.06fF
C125 m1_3443_5997# VSS 35.86fF
C126 m1_1243_5997# VSS 25.05fF
C127 VDD VSS 131.74fF
C128 i_bias VSS -59.70fF
C129 bias_c VSS -50.79fF
C130 m1_7639_427# VSS 0.32fF
C131 m1_7347_423# VSS 0.27fF
C132 m1_7461_921# VSS 0.22fF
C133 m1_7169_923# VSS 0.20fF
C134 m1_7055_433# VSS 0.28fF
C135 m1_6763_422# VSS 0.35fF
C136 m1_6471_422# VSS 0.38fF
C137 m1_7639_1420# VSS 0.31fF
C138 m1_7347_1428# VSS 0.20fF
C139 m1_6877_922# VSS 0.21fF
C140 m1_6585_923# VSS 0.29fF
C141 m1_6293_922# VSS 0.32fF
C142 m1_7055_1417# VSS 0.20fF
C143 m1_6763_1422# VSS 0.29fF
C144 m1_6471_1426# VSS 0.30fF
C145 bias_e VSS 7.90fF
C146 bias_d VSS -76.91fF
C147 li_3433_399# VSS 5.57fF
C148 bias_a VSS -48.09fF
.ends

.subckt sky130_fd_pr__pfet_01v8_YVTMSC a_n207_n140# a_29_n205# a_327_n140# a_n683_n205#
+ a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140# a_n505_n205# a_n741_n140# a_563_n205#
+ a_861_n140# a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_683_n140# w_n1133_n241#
+ a_n919_n140# a_n149_n205# a_n385_n140# a_207_n205# a_505_n140# a_n861_n205# VSUBS
X0 a_n385_n140# a_n505_n205# a_n563_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_327_n140# a_207_n205# a_149_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_149_n140# a_29_n205# a_n29_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_861_n140# a_741_n205# a_683_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n207_n140# a_n327_n205# a_n385_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_n741_n140# a_n861_n205# a_n919_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_683_n140# a_563_n205# a_505_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_919_n205# a_919_n205# a_861_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_n29_n140# a_n149_n205# a_n207_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n563_n140# a_n683_n205# a_n741_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_n919_n140# a_n1097_n140# a_n1097_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_505_n140# a_385_n205# a_327_n140# w_n1133_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n563_n140# a_n29_n140# 0.02fF
C1 a_327_n140# a_n1097_n140# 0.01fF
C2 a_385_n205# a_29_n205# 0.03fF
C3 a_327_n140# a_n207_n140# 0.02fF
C4 a_207_n205# a_n1097_n140# 0.00fF
C5 a_n683_n205# a_n149_n205# 0.02fF
C6 a_861_n140# a_n207_n140# 0.01fF
C7 a_n563_n140# a_n741_n140# 0.06fF
C8 a_327_n140# a_n385_n140# 0.01fF
C9 a_563_n205# w_n1133_n241# 0.15fF
C10 a_563_n205# a_n861_n205# 0.01fF
C11 a_861_n140# a_n385_n140# 0.01fF
C12 a_n327_n205# a_n149_n205# 0.10fF
C13 a_327_n140# a_919_n205# 0.01fF
C14 a_n1097_n140# a_n505_n205# 0.01fF
C15 a_385_n205# a_n149_n205# 0.02fF
C16 a_919_n205# a_207_n205# 0.01fF
C17 w_n1133_n241# a_n919_n140# 0.02fF
C18 a_919_n205# a_861_n140# 0.06fF
C19 a_n1097_n140# a_29_n205# 0.01fF
C20 a_327_n140# a_683_n140# 0.03fF
C21 a_741_n205# a_207_n205# 0.02fF
C22 a_861_n140# a_683_n140# 0.06fF
C23 a_919_n205# a_n505_n205# 0.00fF
C24 a_n563_n140# a_505_n140# 0.01fF
C25 a_149_n140# a_n919_n140# 0.01fF
C26 a_563_n205# a_n683_n205# 0.01fF
C27 a_n29_n140# a_n919_n140# 0.01fF
C28 a_919_n205# a_29_n205# 0.01fF
C29 a_n1097_n140# a_n149_n205# 0.01fF
C30 a_563_n205# a_n327_n205# 0.01fF
C31 a_741_n205# a_n505_n205# 0.01fF
C32 a_n563_n140# a_n1097_n140# 0.02fF
C33 a_n563_n140# a_n207_n140# 0.03fF
C34 a_n741_n140# a_n919_n140# 0.06fF
C35 a_n861_n205# w_n1133_n241# 0.20fF
C36 a_563_n205# a_385_n205# 0.10fF
C37 a_n563_n140# a_n385_n140# 0.06fF
C38 a_741_n205# a_29_n205# 0.01fF
C39 a_149_n140# w_n1133_n241# 0.02fF
C40 a_327_n140# a_861_n140# 0.02fF
C41 a_919_n205# a_n149_n205# 0.01fF
C42 a_n563_n140# a_919_n205# 0.01fF
C43 w_n1133_n241# a_n29_n140# 0.02fF
C44 a_741_n205# a_n149_n205# 0.01fF
C45 a_n563_n140# a_683_n140# 0.01fF
C46 a_n683_n205# w_n1133_n241# 0.20fF
C47 a_n861_n205# a_n683_n205# 0.10fF
C48 a_n741_n140# w_n1133_n241# 0.02fF
C49 a_505_n140# a_n919_n140# 0.01fF
C50 a_563_n205# a_n1097_n140# 0.00fF
C51 a_207_n205# a_n505_n205# 0.01fF
C52 a_149_n140# a_n29_n140# 0.06fF
C53 a_n327_n205# w_n1133_n241# 0.19fF
C54 a_n327_n205# a_n861_n205# 0.02fF
C55 a_207_n205# a_29_n205# 0.10fF
C56 a_149_n140# a_n741_n140# 0.01fF
C57 a_385_n205# w_n1133_n241# 0.16fF
C58 a_n1097_n140# a_n919_n140# 0.06fF
C59 a_385_n205# a_n861_n205# 0.01fF
C60 a_n207_n140# a_n919_n140# 0.01fF
C61 a_n741_n140# a_n29_n140# 0.01fF
C62 a_563_n205# a_919_n205# 0.02fF
C63 a_n385_n140# a_n919_n140# 0.02fF
C64 a_n505_n205# a_29_n205# 0.02fF
C65 w_n1133_n241# a_505_n140# 0.02fF
C66 a_327_n140# a_n563_n140# 0.01fF
C67 a_207_n205# a_n149_n205# 0.03fF
C68 a_741_n205# a_563_n205# 0.10fF
C69 a_n327_n205# a_n683_n205# 0.03fF
C70 a_n563_n140# a_861_n140# 0.01fF
C71 a_385_n205# a_n683_n205# 0.01fF
C72 w_n1133_n241# a_n1097_n140# 0.33fF
C73 a_n861_n205# a_n1097_n140# 0.07fF
C74 a_n919_n140# a_683_n140# 0.01fF
C75 w_n1133_n241# a_n207_n140# 0.02fF
C76 a_149_n140# a_505_n140# 0.03fF
C77 a_n505_n205# a_n149_n205# 0.03fF
C78 a_n385_n140# w_n1133_n241# 0.02fF
C79 a_505_n140# a_n29_n140# 0.02fF
C80 a_385_n205# a_n327_n205# 0.01fF
C81 a_149_n140# a_n1097_n140# 0.01fF
C82 a_n741_n140# a_505_n140# 0.01fF
C83 a_149_n140# a_n207_n140# 0.03fF
C84 a_n149_n205# a_29_n205# 0.10fF
C85 a_919_n205# w_n1133_n241# 0.28fF
C86 a_n1097_n140# a_n29_n140# 0.01fF
C87 a_n207_n140# a_n29_n140# 0.06fF
C88 a_149_n140# a_n385_n140# 0.02fF
C89 a_563_n205# a_207_n205# 0.03fF
C90 a_n385_n140# a_n29_n140# 0.03fF
C91 a_n683_n205# a_n1097_n140# 0.02fF
C92 a_n741_n140# a_n1097_n140# 0.03fF
C93 a_n741_n140# a_n207_n140# 0.02fF
C94 w_n1133_n241# a_683_n140# 0.01fF
C95 a_741_n205# w_n1133_n241# 0.14fF
C96 a_741_n205# a_n861_n205# 0.01fF
C97 a_149_n140# a_919_n205# 0.01fF
C98 a_327_n140# a_n919_n140# 0.01fF
C99 a_n741_n140# a_n385_n140# 0.03fF
C100 a_n327_n205# a_n1097_n140# 0.01fF
C101 a_919_n205# a_n29_n140# 0.01fF
C102 a_563_n205# a_n505_n205# 0.01fF
C103 a_385_n205# a_n1097_n140# 0.00fF
C104 a_149_n140# a_683_n140# 0.02fF
C105 a_919_n205# a_n683_n205# 0.00fF
C106 a_n29_n140# a_683_n140# 0.01fF
C107 a_563_n205# a_29_n205# 0.02fF
C108 a_919_n205# a_n327_n205# 0.00fF
C109 a_n741_n140# a_683_n140# 0.01fF
C110 a_741_n205# a_n683_n205# 0.01fF
C111 a_n1097_n140# a_505_n140# 0.01fF
C112 a_505_n140# a_n207_n140# 0.01fF
C113 a_919_n205# a_385_n205# 0.01fF
C114 a_327_n140# w_n1133_n241# 0.02fF
C115 a_207_n205# w_n1133_n241# 0.17fF
C116 a_n861_n205# a_207_n205# 0.01fF
C117 a_n385_n140# a_505_n140# 0.01fF
C118 a_741_n205# a_n327_n205# 0.01fF
C119 a_861_n140# w_n1133_n241# 0.01fF
C120 a_563_n205# a_n149_n205# 0.01fF
C121 a_n1097_n140# a_n207_n140# 0.01fF
C122 a_741_n205# a_385_n205# 0.03fF
C123 a_327_n140# a_149_n140# 0.06fF
C124 a_919_n205# a_505_n140# 0.02fF
C125 a_n385_n140# a_n1097_n140# 0.01fF
C126 a_n385_n140# a_n207_n140# 0.06fF
C127 w_n1133_n241# a_n505_n205# 0.20fF
C128 a_n861_n205# a_n505_n205# 0.03fF
C129 a_327_n140# a_n29_n140# 0.03fF
C130 a_149_n140# a_861_n140# 0.01fF
C131 a_n563_n140# a_n919_n140# 0.03fF
C132 a_861_n140# a_n29_n140# 0.01fF
C133 a_505_n140# a_683_n140# 0.06fF
C134 a_327_n140# a_n741_n140# 0.01fF
C135 w_n1133_n241# a_29_n205# 0.18fF
C136 a_919_n205# a_n207_n140# 0.01fF
C137 a_n861_n205# a_29_n205# 0.01fF
C138 a_n683_n205# a_207_n205# 0.01fF
C139 a_861_n140# a_n741_n140# 0.01fF
C140 a_919_n205# a_n385_n140# 0.01fF
C141 a_n327_n205# a_207_n205# 0.02fF
C142 a_n207_n140# a_683_n140# 0.01fF
C143 a_385_n205# a_207_n205# 0.10fF
C144 a_n385_n140# a_683_n140# 0.01fF
C145 a_n683_n205# a_n505_n205# 0.10fF
C146 w_n1133_n241# a_n149_n205# 0.19fF
C147 a_n861_n205# a_n149_n205# 0.01fF
C148 a_n563_n140# w_n1133_n241# 0.02fF
C149 a_n327_n205# a_n505_n205# 0.10fF
C150 a_n683_n205# a_29_n205# 0.01fF
C151 a_919_n205# a_683_n140# 0.03fF
C152 a_741_n205# a_919_n205# 0.07fF
C153 a_327_n140# a_505_n140# 0.06fF
C154 a_385_n205# a_n505_n205# 0.01fF
C155 a_861_n140# a_505_n140# 0.03fF
C156 a_n563_n140# a_149_n140# 0.01fF
C157 a_n327_n205# a_29_n205# 0.03fF
C158 w_n1133_n241# VSUBS 3.28fF
.ends

.subckt ota_v2_without_cmfb in bias_c bias_e op on i_bias VDD VSS bias_circuit_0/m1_3551_3596#
+ cmc li_14138_570# bias_circuit_0/bias_d li_11121_570# li_11122_5650# li_8434_570#
+ bias_b li_8436_5651# bias_circuit_0/m1_1243_5997# bias_circuit_0/m1_3443_5997# bias_a
+ ip bias_circuit_0/m1_5643_5997#
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_0 VDD bias_b bias_b li_8436_5651# bias_b VDD bias_b
+ li_8436_5651# VDD li_8436_5651# VDD bias_b li_8436_5651# bias_b VDD VDD bias_b bias_b
+ VDD bias_b li_8436_5651# VDD bias_b li_8436_5651# li_8436_5651# bias_b VDD bias_b
+ VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_8 bias_circuit_0/bias_d li_8434_570# bias_circuit_0/bias_d
+ on VSS bias_circuit_0/bias_d on li_8434_570# on bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on bias_circuit_0/bias_d li_8434_570# VSS li_8434_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on li_8434_570# bias_circuit_0/bias_d on on bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_1 VDD bias_b bias_b li_11122_5650# bias_b VDD
+ bias_b li_11122_5650# VDD li_11122_5650# VDD bias_b li_11122_5650# bias_b VDD VDD
+ bias_b bias_b VDD bias_b li_11122_5650# VDD bias_b li_11122_5650# li_11122_5650#
+ bias_b VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_AKSJZW_9 bias_circuit_0/bias_d li_11121_570# bias_circuit_0/bias_d
+ op VSS bias_circuit_0/bias_d op li_11121_570# op bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op bias_circuit_0/bias_d li_11121_570# VSS li_11121_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op li_11121_570# bias_circuit_0/bias_d op op bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_2 VDD bias_b bias_b li_8436_5651# bias_b VDD bias_b
+ li_8436_5651# VDD li_8436_5651# VDD bias_b li_8436_5651# bias_b VDD VDD bias_b bias_b
+ VDD bias_b li_8436_5651# VDD bias_b li_8436_5651# li_8436_5651# bias_b VDD bias_b
+ VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__pfet_01v8_lvt_YVTR7C_3 VDD bias_b bias_b li_11122_5650# bias_b VDD
+ bias_b li_11122_5650# VDD li_11122_5650# VDD bias_b li_11122_5650# bias_b VDD VDD
+ bias_b bias_b VDD bias_b li_11122_5650# VDD bias_b li_11122_5650# li_11122_5650#
+ bias_b VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_YVTR7C
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_0 VSS li_8436_5651# li_14138_570# ip li_8436_5651#
+ li_8436_5651# ip li_14138_570# li_8436_5651# li_14138_570# li_14138_570# li_8436_5651#
+ li_8436_5651# ip ip li_14138_570# ip li_14138_570# ip VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_lvt_K7HVMB_1 VSS li_11122_5650# li_14138_570# in li_11122_5650#
+ li_11122_5650# in li_14138_570# li_11122_5650# li_14138_570# li_14138_570# li_11122_5650#
+ li_11122_5650# in in li_14138_570# in li_14138_570# in VSS VSS sky130_fd_pr__nfet_01v8_lvt_K7HVMB
Xsky130_fd_pr__nfet_01v8_AKSJZW_10 bias_circuit_0/bias_d li_11121_570# bias_circuit_0/bias_d
+ op VSS bias_circuit_0/bias_d op li_11121_570# op bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op bias_circuit_0/bias_d li_11121_570# VSS li_11121_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op li_11121_570# bias_circuit_0/bias_d op op bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_0 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_AKSJZW_11 bias_circuit_0/bias_d li_11121_570# bias_circuit_0/bias_d
+ op VSS bias_circuit_0/bias_d op li_11121_570# op bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op bias_circuit_0/bias_d li_11121_570# VSS li_11121_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d op li_11121_570# bias_circuit_0/bias_d op op bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_11121_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_S6RQQZ_1 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_2 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_3 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_4 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_5 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_6 cmc VSS cmc VSS cmc li_14138_570# VSS cmc li_14138_570#
+ cmc VSS li_14138_570# cmc cmc cmc li_14138_570# li_14138_570# cmc VSS cmc cmc VSS
+ cmc VSS li_14138_570# VSS cmc VSS cmc li_14138_570# li_14138_570# cmc cmc VSS li_14138_570#
+ VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_7 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_8 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_9 bias_a VSS bias_a VSS bias_a li_14138_570# VSS bias_a
+ li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570# li_14138_570#
+ bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS bias_a li_14138_570#
+ li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_10 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xsky130_fd_pr__nfet_01v8_S6RQQZ_11 bias_a VSS bias_a VSS bias_a li_14138_570# VSS
+ bias_a li_14138_570# bias_a VSS li_14138_570# bias_a bias_a bias_a li_14138_570#
+ li_14138_570# bias_a VSS bias_a bias_a VSS bias_a VSS li_14138_570# VSS bias_a VSS
+ bias_a li_14138_570# li_14138_570# bias_a bias_a VSS li_14138_570# VSS sky130_fd_pr__nfet_01v8_S6RQQZ
Xbias_circuit_0 bias_c bias_e i_bias VDD bias_circuit_0/m1_1243_5997# bias_circuit_0/m1_3443_5997#
+ bias_a bias_circuit_0/m1_7347_1428# bias_circuit_0/m1_7639_1420# bias_circuit_0/m1_7169_923#
+ bias_circuit_0/m1_7461_921# bias_circuit_0/m1_7347_423# bias_circuit_0/m1_7639_427#
+ bias_b VSS bias_circuit_0/m1_3551_3596# bias_circuit_0/m1_5643_5997# bias_circuit_0/bias_d
+ bias_circuit
Xsky130_fd_pr__pfet_01v8_YVTMSC_0 on bias_c li_8436_5651# bias_c bias_c li_8436_5651#
+ on VDD bias_c li_8436_5651# bias_c on VDD bias_c on bias_c li_8436_5651# VDD on
+ bias_c li_8436_5651# bias_c on bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_1 on bias_c li_8436_5651# bias_c bias_c li_8436_5651#
+ on VDD bias_c li_8436_5651# bias_c on VDD bias_c on bias_c li_8436_5651# VDD on
+ bias_c li_8436_5651# bias_c on bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_0 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__pfet_01v8_YVTMSC_2 op bias_c li_11122_5650# bias_c bias_c li_11122_5650#
+ op VDD bias_c li_11122_5650# bias_c op VDD bias_c op bias_c li_11122_5650# VDD op
+ bias_c li_11122_5650# bias_c op bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__pfet_01v8_YVTMSC_3 op bias_c li_11122_5650# bias_c bias_c li_11122_5650#
+ op VDD bias_c li_11122_5650# bias_c op VDD bias_c op bias_c li_11122_5650# VDD op
+ bias_c li_11122_5650# bias_c op bias_c VSS sky130_fd_pr__pfet_01v8_YVTMSC
Xsky130_fd_pr__nfet_01v8_AKSJZW_2 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_1 bias_a VSS bias_a li_8434_570# VSS bias_a li_8434_570#
+ VSS li_8434_570# bias_a bias_a bias_a li_8434_570# bias_a VSS VSS VSS bias_a bias_a
+ li_8434_570# VSS bias_a li_8434_570# li_8434_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_3 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_4 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_5 bias_a VSS bias_a li_11121_570# VSS bias_a li_11121_570#
+ VSS li_11121_570# bias_a bias_a bias_a li_11121_570# bias_a VSS VSS VSS bias_a bias_a
+ li_11121_570# VSS bias_a li_11121_570# li_11121_570# bias_a bias_a VSS VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_6 bias_circuit_0/bias_d li_8434_570# bias_circuit_0/bias_d
+ on VSS bias_circuit_0/bias_d on li_8434_570# on bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on bias_circuit_0/bias_d li_8434_570# VSS li_8434_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on li_8434_570# bias_circuit_0/bias_d on on bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
Xsky130_fd_pr__nfet_01v8_AKSJZW_7 bias_circuit_0/bias_d li_8434_570# bias_circuit_0/bias_d
+ on VSS bias_circuit_0/bias_d on li_8434_570# on bias_circuit_0/bias_d bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on bias_circuit_0/bias_d li_8434_570# VSS li_8434_570# bias_circuit_0/bias_d
+ bias_circuit_0/bias_d on li_8434_570# bias_circuit_0/bias_d on on bias_circuit_0/bias_d
+ bias_circuit_0/bias_d li_8434_570# VSS sky130_fd_pr__nfet_01v8_AKSJZW
C0 bias_c VDD 6.22fF
C1 li_11122_5650# VDD 3.68fF
C2 cmc li_11122_5650# 0.13fF
C3 m1_17097_3928# li_14138_570# 0.00fF
C4 bias_b VDD 12.49fF
C5 on li_8434_570# 4.15fF
C6 on bias_e 0.01fF
C7 ip in 0.03fF
C8 bias_a bias_circuit_0/m1_7639_427# 0.01fF
C9 li_8434_570# bias_c 0.12fF
C10 li_11121_570# li_14138_570# 0.23fF
C11 ip m1_17393_3568# 0.00fF
C12 on li_11121_570# 0.17fF
C13 li_8436_5651# VDD 4.67fF
C14 bias_a bias_circuit_0/bias_d 2.87fF
C15 bias_a bias_circuit_0/m1_7639_1420# 0.00fF
C16 li_11121_570# bias_c 0.12fF
C17 li_11121_570# li_11122_5650# 0.16fF
C18 op bias_circuit_0/bias_d 9.36fF
C19 ip li_14138_570# 1.47fF
C20 li_8434_570# li_8436_5651# 0.16fF
C21 li_8434_570# bias_circuit_0/m1_7461_921# 0.01fF
C22 m1_18877_3928# cmc 0.01fF
C23 ip li_11122_5650# 0.01fF
C24 bias_a li_14138_570# 27.43fF
C25 op li_14138_570# 0.08fF
C26 on bias_a 0.48fF
C27 on op 0.59fF
C28 li_8434_570# VDD 0.03fF
C29 op bias_c 4.25fF
C30 op li_11122_5650# 2.52fF
C31 op bias_b 0.27fF
C32 ip li_8436_5651# 1.22fF
C33 li_11121_570# VDD 0.02fF
C34 ip m1_15613_3568# 0.01fF
C35 li_8434_570# bias_e 0.00fF
C36 bias_circuit_0/bias_d bias_circuit_0/m1_7639_1420# 0.00fF
C37 bias_a li_8436_5651# 0.14fF
C38 op li_8436_5651# 0.12fF
C39 bias_a m1_15613_3568# 0.01fF
C40 li_8434_570# li_11121_570# 0.52fF
C41 in m1_17393_3568# 0.01fF
C42 li_14138_570# bias_circuit_0/bias_d 0.02fF
C43 li_14138_570# in 1.51fF
C44 bias_a cmc 0.78fF
C45 bias_circuit_0/m1_3551_3596# bias_circuit_0/bias_d 0.03fF
C46 on bias_circuit_0/bias_d 10.13fF
C47 m1_17097_3928# ip 0.01fF
C48 on bias_circuit_0/m1_7639_1420# 0.00fF
C49 op VDD 0.65fF
C50 li_14138_570# m1_17393_3568# 0.01fF
C51 bias_c bias_circuit_0/bias_d 2.13fF
C52 li_11122_5650# bias_circuit_0/bias_d 0.28fF
C53 li_11122_5650# in 1.14fF
C54 bias_b bias_circuit_0/bias_d 0.02fF
C55 li_8434_570# bias_a 10.56fF
C56 li_11122_5650# m1_17393_3568# 0.00fF
C57 bias_a bias_e 0.00fF
C58 li_8434_570# op 0.17fF
C59 li_11121_570# bias_a 10.56fF
C60 on bias_circuit_0/m1_3551_3596# 0.00fF
C61 li_11121_570# op 4.14fF
C62 bias_circuit_0/bias_d li_8436_5651# 0.66fF
C63 in li_8436_5651# 0.01fF
C64 li_14138_570# li_11122_5650# 0.78fF
C65 bias_circuit_0/m1_3551_3596# bias_c 0.00fF
C66 on bias_c 4.65fF
C67 on li_11122_5650# 0.12fF
C68 on bias_b 0.27fF
C69 bias_circuit_0/m1_5643_5997# VDD -0.00fF
C70 bias_c li_11122_5650# 3.17fF
C71 bias_a ip 0.31fF
C72 bias_c bias_b 1.94fF
C73 bias_b li_11122_5650# 4.93fF
C74 m1_18877_3928# in 0.01fF
C75 li_14138_570# li_8436_5651# 0.80fF
C76 bias_circuit_0/bias_d VDD 3.37fF
C77 cmc in 0.31fF
C78 on li_8436_5651# 2.52fF
C79 li_8434_570# bias_circuit_0/m1_7639_427# 0.01fF
C80 li_14138_570# m1_15613_3568# 0.01fF
C81 op bias_a 0.52fF
C82 bias_c li_8436_5651# 4.18fF
C83 li_11122_5650# li_8436_5651# 1.47fF
C84 li_8434_570# bias_circuit_0/bias_d 6.56fF
C85 li_8434_570# bias_circuit_0/m1_7639_1420# 0.01fF
C86 m1_17097_3928# in 0.00fF
C87 bias_b li_8436_5651# 4.46fF
C88 m1_18877_3928# li_14138_570# 0.00fF
C89 cmc li_14138_570# 26.78fF
C90 bias_circuit_0/m1_3551_3596# VDD 0.15fF
C91 on VDD 0.63fF
C92 li_11121_570# bias_circuit_0/bias_d 6.30fF
C93 m1_17393_3568# VSS 0.09fF $ **FLOATING
C94 m1_15613_3568# VSS 0.12fF $ **FLOATING
C95 m1_18877_3928# VSS 0.10fF $ **FLOATING
C96 m1_17097_3928# VSS 0.06fF $ **FLOATING
C97 on VSS 5.53fF
C98 li_11121_570# VSS 10.99fF
C99 li_11122_5650# VSS -33.02fF
C100 li_8434_570# VSS 10.90fF
C101 bias_a VSS -274.59fF
C102 li_8436_5651# VSS 3.30fF
C103 bias_circuit_0/m1_3551_3596# VSS -342.21fF
C104 bias_b VSS -360.90fF
C105 bias_circuit_0/m1_5643_5997# VSS 38.05fF
C106 bias_circuit_0/m1_3443_5997# VSS 35.85fF
C107 bias_circuit_0/m1_1243_5997# VSS 25.03fF
C108 VDD VSS 288.24fF
C109 i_bias VSS -60.68fF
C110 bias_c VSS -128.43fF
C111 bias_circuit_0/m1_7639_427# VSS 0.13fF
C112 bias_circuit_0/m1_7347_423# VSS 0.13fF
C113 bias_circuit_0/m1_7461_921# VSS 0.14fF
C114 bias_circuit_0/m1_7169_923# VSS 0.14fF
C115 bias_circuit_0/m1_7055_433# VSS 0.14fF
C116 bias_circuit_0/m1_6763_422# VSS 0.20fF
C117 bias_circuit_0/m1_6471_422# VSS 0.20fF
C118 bias_circuit_0/m1_7639_1420# VSS 0.13fF
C119 bias_circuit_0/m1_7347_1428# VSS 0.14fF
C120 bias_circuit_0/m1_6877_922# VSS 0.14fF
C121 bias_circuit_0/m1_6585_923# VSS 0.22fF
C122 bias_circuit_0/m1_6293_922# VSS 0.16fF
C123 bias_circuit_0/m1_7055_1417# VSS 0.14fF
C124 bias_circuit_0/m1_6763_1422# VSS 0.22fF
C125 bias_circuit_0/m1_6471_1426# VSS 0.22fF
C126 bias_e VSS 3.22fF
C127 bias_circuit_0/bias_d VSS -237.66fF
C128 bias_circuit_0/li_3433_399# VSS 4.65fF
C129 li_14138_570# VSS 26.06fF
C130 cmc VSS -107.67fF
C131 op VSS 5.29fF
C132 in VSS -27.57fF
C133 ip VSS -26.06fF
.ends

.subckt pmos_tgate a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136# a_64_n136# a_160_n136#
+ a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136# a_n512_n234# a_256_n136#
+ VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_64_n136# a_160_n136# 0.33fF
C1 a_n320_n136# a_256_n136# 0.03fF
C2 a_n32_n136# a_448_n136# 0.04fF
C3 a_448_n136# a_n128_n136# 0.03fF
C4 a_n508_n136# w_n646_n356# 0.13fF
C5 a_n32_n136# a_352_n136# 0.05fF
C6 a_n224_n136# a_256_n136# 0.04fF
C7 a_352_n136# a_n128_n136# 0.04fF
C8 a_n32_n136# a_n416_n136# 0.05fF
C9 a_n416_n136# a_n128_n136# 0.07fF
C10 a_n512_n234# a_256_n136# 0.03fF
C11 a_n508_n136# a_448_n136# 0.02fF
C12 a_n32_n136# a_160_n136# 0.12fF
C13 a_n508_n136# a_352_n136# 0.02fF
C14 a_160_n136# a_n128_n136# 0.07fF
C15 a_n416_n136# a_n508_n136# 0.33fF
C16 a_64_n136# a_256_n136# 0.12fF
C17 a_n224_n136# a_n320_n136# 0.33fF
C18 a_n320_n136# a_n512_n234# 0.03fF
C19 a_n508_n136# a_160_n136# 0.03fF
C20 a_n224_n136# a_n512_n234# 0.03fF
C21 w_n646_n356# a_448_n136# 0.13fF
C22 a_352_n136# w_n646_n356# 0.08fF
C23 a_n416_n136# w_n646_n356# 0.08fF
C24 a_64_n136# a_n320_n136# 0.05fF
C25 a_n32_n136# a_256_n136# 0.07fF
C26 a_256_n136# a_n128_n136# 0.05fF
C27 a_n224_n136# a_64_n136# 0.07fF
C28 a_352_n136# a_448_n136# 0.33fF
C29 a_64_n136# a_n512_n234# 0.03fF
C30 a_n416_n136# a_448_n136# 0.02fF
C31 a_160_n136# w_n646_n356# 0.06fF
C32 a_n416_n136# a_352_n136# 0.02fF
C33 a_n508_n136# a_256_n136# 0.02fF
C34 a_160_n136# a_448_n136# 0.07fF
C35 a_n32_n136# a_n320_n136# 0.07fF
C36 a_n320_n136# a_n128_n136# 0.12fF
C37 a_160_n136# a_352_n136# 0.12fF
C38 a_n416_n136# a_160_n136# 0.03fF
C39 a_n224_n136# a_n32_n136# 0.12fF
C40 a_n224_n136# a_n128_n136# 0.33fF
C41 a_n32_n136# a_n512_n234# 0.03fF
C42 a_n512_n234# a_n128_n136# 0.03fF
C43 w_n646_n356# a_256_n136# 0.06fF
C44 a_n320_n136# a_n508_n136# 0.12fF
C45 a_n224_n136# a_n508_n136# 0.07fF
C46 a_n512_n234# a_n508_n136# 0.03fF
C47 a_n32_n136# a_64_n136# 0.33fF
C48 a_64_n136# a_n128_n136# 0.12fF
C49 a_256_n136# a_448_n136# 0.12fF
C50 a_352_n136# a_256_n136# 0.33fF
C51 a_n416_n136# a_256_n136# 0.03fF
C52 a_n320_n136# w_n646_n356# 0.06fF
C53 a_64_n136# a_n508_n136# 0.03fF
C54 a_n224_n136# w_n646_n356# 0.06fF
C55 a_n512_n234# w_n646_n356# 1.47fF
C56 a_160_n136# a_256_n136# 0.33fF
C57 a_n320_n136# a_448_n136# 0.02fF
C58 a_n32_n136# a_n128_n136# 0.33fF
C59 a_n320_n136# a_352_n136# 0.03fF
C60 a_n320_n136# a_n416_n136# 0.33fF
C61 a_n224_n136# a_448_n136# 0.03fF
C62 a_n512_n234# a_448_n136# 0.03fF
C63 a_n224_n136# a_352_n136# 0.03fF
C64 a_64_n136# w_n646_n356# 0.05fF
C65 a_n224_n136# a_n416_n136# 0.12fF
C66 a_n512_n234# a_352_n136# 0.03fF
C67 a_n32_n136# a_n508_n136# 0.04fF
C68 a_n416_n136# a_n512_n234# 0.03fF
C69 a_n508_n136# a_n128_n136# 0.05fF
C70 a_n320_n136# a_160_n136# 0.04fF
C71 a_n224_n136# a_160_n136# 0.05fF
C72 a_64_n136# a_448_n136# 0.05fF
C73 a_n512_n234# a_160_n136# 0.03fF
C74 a_64_n136# a_352_n136# 0.07fF
C75 a_64_n136# a_n416_n136# 0.04fF
C76 a_n32_n136# w_n646_n356# 0.05fF
C77 w_n646_n356# a_n128_n136# 0.05fF
C78 w_n646_n356# VSUBS 2.52fF
.ends

.subckt nmos_tgate a_256_n52# a_n32_n52# a_n224_n52# a_448_n52# a_n416_n52# a_160_n52#
+ a_n610_n226# a_n128_n52# a_352_n52# a_n320_n52# a_n508_n52# a_n512_n149# a_64_n52#
X0 a_n32_n52# a_n512_n149# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n149# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n149# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n149# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n149# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n149# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n149# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n149# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n149# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n149# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_256_n52# a_n416_n52# 0.01fF
C1 a_64_n52# a_n32_n52# 0.13fF
C2 a_n320_n52# a_n508_n52# 0.05fF
C3 a_160_n52# a_448_n52# 0.03fF
C4 a_n32_n52# a_n224_n52# 0.05fF
C5 a_448_n52# a_n512_n149# 0.03fF
C6 a_n320_n52# a_n416_n52# 0.13fF
C7 a_256_n52# a_n128_n52# 0.02fF
C8 a_64_n52# a_448_n52# 0.02fF
C9 a_256_n52# a_160_n52# 0.13fF
C10 a_n320_n52# a_n128_n52# 0.05fF
C11 a_448_n52# a_n224_n52# 0.01fF
C12 a_256_n52# a_n512_n149# 0.03fF
C13 a_n32_n52# a_448_n52# 0.02fF
C14 a_n508_n52# a_352_n52# 0.01fF
C15 a_256_n52# a_64_n52# 0.05fF
C16 a_n416_n52# a_352_n52# 0.01fF
C17 a_n320_n52# a_160_n52# 0.02fF
C18 a_n320_n52# a_n512_n149# 0.03fF
C19 a_256_n52# a_n224_n52# 0.02fF
C20 a_n320_n52# a_64_n52# 0.02fF
C21 a_256_n52# a_n32_n52# 0.03fF
C22 a_n128_n52# a_352_n52# 0.02fF
C23 a_n320_n52# a_n224_n52# 0.13fF
C24 a_n320_n52# a_n32_n52# 0.03fF
C25 a_160_n52# a_352_n52# 0.05fF
C26 a_256_n52# a_448_n52# 0.05fF
C27 a_352_n52# a_n512_n149# 0.03fF
C28 a_64_n52# a_352_n52# 0.03fF
C29 a_n320_n52# a_448_n52# 0.01fF
C30 a_352_n52# a_n224_n52# 0.01fF
C31 a_n32_n52# a_352_n52# 0.02fF
C32 a_256_n52# a_n320_n52# 0.01fF
C33 a_n508_n52# a_n416_n52# 0.13fF
C34 a_448_n52# a_352_n52# 0.13fF
C35 a_n508_n52# a_n128_n52# 0.02fF
C36 a_n128_n52# a_n416_n52# 0.03fF
C37 a_256_n52# a_352_n52# 0.13fF
C38 a_n508_n52# a_160_n52# 0.01fF
C39 a_n508_n52# a_n512_n149# 0.03fF
C40 a_160_n52# a_n416_n52# 0.01fF
C41 a_n416_n52# a_n512_n149# 0.03fF
C42 a_n508_n52# a_64_n52# 0.01fF
C43 a_n320_n52# a_352_n52# 0.01fF
C44 a_64_n52# a_n416_n52# 0.02fF
C45 a_n508_n52# a_n224_n52# 0.03fF
C46 a_n128_n52# a_160_n52# 0.03fF
C47 a_n128_n52# a_n512_n149# 0.03fF
C48 a_n508_n52# a_n32_n52# 0.02fF
C49 a_n416_n52# a_n224_n52# 0.05fF
C50 a_n32_n52# a_n416_n52# 0.02fF
C51 a_64_n52# a_n128_n52# 0.05fF
C52 a_160_n52# a_n512_n149# 0.03fF
C53 a_n128_n52# a_n224_n52# 0.13fF
C54 a_n508_n52# a_448_n52# 0.01fF
C55 a_64_n52# a_160_n52# 0.13fF
C56 a_n32_n52# a_n128_n52# 0.13fF
C57 a_64_n52# a_n512_n149# 0.03fF
C58 a_n416_n52# a_448_n52# 0.01fF
C59 a_160_n52# a_n224_n52# 0.02fF
C60 a_n224_n52# a_n512_n149# 0.03fF
C61 a_n32_n52# a_160_n52# 0.05fF
C62 a_n32_n52# a_n512_n149# 0.03fF
C63 a_256_n52# a_n508_n52# 0.01fF
C64 a_n128_n52# a_448_n52# 0.01fF
C65 a_64_n52# a_n224_n52# 0.03fF
C66 a_448_n52# a_n610_n226# 0.07fF
C67 a_352_n52# a_n610_n226# 0.05fF
C68 a_256_n52# a_n610_n226# 0.04fF
C69 a_160_n52# a_n610_n226# 0.04fF
C70 a_64_n52# a_n610_n226# 0.04fF
C71 a_n32_n52# a_n610_n226# 0.04fF
C72 a_n128_n52# a_n610_n226# 0.04fF
C73 a_n224_n52# a_n610_n226# 0.04fF
C74 a_n320_n52# a_n610_n226# 0.04fF
C75 a_n416_n52# a_n610_n226# 0.05fF
C76 a_n508_n52# a_n610_n226# 0.07fF
C77 a_n512_n149# a_n610_n226# 1.83fF
.ends

.subckt transmission_gate en en_b VDD in out VSS
Xpmos_tgate_0 in in out in out in out VDD in out out en_b out VSS pmos_tgate
Xnmos_tgate_0 out in in out in in VSS out in out out en out nmos_tgate
C0 in en_b 0.15fF
C1 VDD out 0.29fF
C2 out en 0.01fF
C3 VDD en 0.12fF
C4 in out 0.77fF
C5 VDD in 0.70fF
C6 in en 0.13fF
C7 out en_b 0.01fF
C8 VDD en_b -0.11fF
C9 en_b en 0.07fF
C10 en VSS 1.70fF
C11 out VSS 0.57fF
C12 in VSS 1.13fF
C13 en_b VSS 0.09fF
C14 VDD VSS 3.16fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 m3_n630_n580# c1_n530_n480# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb cm op cmc p2_b p2 on unit_cap_mim_m3m4_30/m3_n630_n580# transmission_gate_4/out
+ transmission_gate_8/in bias_a p1 VDD transmission_gate_3/out transmission_gate_7/in
+ VSS p1_b
Xtransmission_gate_10 p1 p1_b VDD transmission_gate_3/out on VSS transmission_gate
Xtransmission_gate_11 p1 p1_b VDD transmission_gate_4/out op VSS transmission_gate
Xtransmission_gate_0 p1 p1_b VDD cm transmission_gate_7/in VSS transmission_gate
Xtransmission_gate_1 p1 p1_b VDD cm transmission_gate_6/in VSS transmission_gate
Xtransmission_gate_2 p1 p1_b VDD bias_a transmission_gate_8/in VSS transmission_gate
Xtransmission_gate_3 p2 p2_b VDD cm transmission_gate_3/out VSS transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 p2_b VDD cm transmission_gate_4/out VSS transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 p2_b VDD bias_a transmission_gate_9/in VSS transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 p2_b VDD transmission_gate_6/in op VSS transmission_gate
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 p2_b VDD transmission_gate_7/in on VSS transmission_gate
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 p2_b VDD transmission_gate_8/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 p1_b VDD transmission_gate_9/in cmc VSS transmission_gate
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 p1_b unit_cap_mim_m3m4_18/m3_n630_n580# 0.06fF
C1 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C2 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_23/c1_n530_n480# -0.19fF
C3 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.12fF
C4 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580# 0.17fF
C5 p2 on 0.24fF
C6 transmission_gate_3/out transmission_gate_9/in 1.40fF
C7 transmission_gate_4/out p1_b 0.55fF
C8 p1 VDD 1.10fF
C9 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_7/in -0.56fF
C10 cmc unit_cap_mim_m3m4_27/m3_n630_n580# 0.10fF
C11 p1 unit_cap_mim_m3m4_22/m3_n630_n580# 0.06fF
C12 p1_b transmission_gate_7/in 0.40fF
C13 cmc transmission_gate_9/in 6.62fF
C14 p1_b p2_b 2.92fF
C15 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_27/m3_n630_n580# 0.12fF
C16 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_26/c1_n530_n480# -0.35fF
C17 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_34/m3_n630_n580# 0.17fF
C18 cmc transmission_gate_3/out 0.97fF
C19 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.17fF
C20 unit_cap_mim_m3m4_24/m3_n630_n580# p1 0.08fF
C21 op on 2.00fF
C22 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C23 unit_cap_mim_m3m4_25/c1_n530_n480# p2 0.04fF
C24 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580# -0.29fF
C25 VDD transmission_gate_9/in -0.11fF
C26 p1 p2 2.82fF
C27 transmission_gate_6/in on 0.40fF
C28 bias_a cm 1.15fF
C29 unit_cap_mim_m3m4_31/c1_n530_n480# op 0.05fF
C30 op unit_cap_mim_m3m4_29/m3_n630_n580# 0.39fF
C31 VDD transmission_gate_3/out -0.05fF
C32 transmission_gate_8/in cm 0.03fF
C33 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C34 p1 unit_cap_mim_m3m4_17/m3_n630_n580# 0.08fF
C35 unit_cap_mim_m3m4_20/m3_n630_n580# p1_b 0.05fF
C36 unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_9/in -0.80fF
C37 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_34/m3_n630_n580# 0.17fF
C38 unit_cap_mim_m3m4_26/m3_n630_n580# cmc 0.10fF
C39 unit_cap_mim_m3m4_23/c1_n530_n480# transmission_gate_3/out -0.24fF
C40 transmission_gate_6/in unit_cap_mim_m3m4_29/m3_n630_n580# -0.80fF
C41 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480# -0.20fF
C42 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580# -0.18fF
C43 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580# -0.20fF
C44 unit_cap_mim_m3m4_24/m3_n630_n580# transmission_gate_9/in 0.17fF
C45 cmc VDD 1.23fF
C46 p1 unit_cap_mim_m3m4_29/c1_n530_n480# 0.11fF
C47 transmission_gate_4/out unit_cap_mim_m3m4_31/m3_n630_n580# 0.32fF
C48 p1 op 0.52fF
C49 unit_cap_mim_m3m4_26/c1_n530_n480# p2 0.04fF
C50 transmission_gate_4/out cm 0.07fF
C51 p2 transmission_gate_9/in 0.14fF
C52 unit_cap_mim_m3m4_20/c1_n530_n480# transmission_gate_7/in -0.18fF
C53 cmc unit_cap_mim_m3m4_22/m3_n630_n580# 0.71fF
C54 p1 unit_cap_mim_m3m4_21/m3_n630_n580# 0.06fF
C55 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580# -0.32fF
C56 unit_cap_mim_m3m4_23/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580# 0.12fF
C57 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C58 p2 transmission_gate_3/out 0.15fF
C59 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_27/m3_n630_n580# 0.12fF
C60 transmission_gate_6/in p1 0.38fF
C61 cmc unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C62 transmission_gate_7/in cm 0.10fF
C63 unit_cap_mim_m3m4_17/m3_n630_n580# transmission_gate_3/out -0.23fF
C64 p2_b cm 1.01fF
C65 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_34/c1_n530_n480# -0.14fF
C66 unit_cap_mim_m3m4_28/c1_n530_n480# p2 0.04fF
C67 p1 unit_cap_mim_m3m4_16/m3_n630_n580# 0.08fF
C68 p1_b unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C69 cmc p2 0.25fF
C70 op unit_cap_mim_m3m4_27/m3_n630_n580# 0.48fF
C71 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_28/c1_n530_n480# -0.33fF
C72 p1 unit_cap_mim_m3m4_30/m3_n630_n580# 0.06fF
C73 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C74 op transmission_gate_9/in 0.67fF
C75 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_20/c1_n530_n480# -0.19fF
C76 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580# -0.13fF
C77 cmc unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C78 transmission_gate_8/in unit_cap_mim_m3m4_35/m3_n630_n580# -0.15fF
C79 op transmission_gate_3/out 0.56fF
C80 transmission_gate_8/in on 0.88fF
C81 transmission_gate_6/in unit_cap_mim_m3m4_27/m3_n630_n580# 0.13fF
C82 transmission_gate_6/in transmission_gate_9/in 0.09fF
C83 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C84 unit_cap_mim_m3m4_25/m3_n630_n580# transmission_gate_9/in 0.38fF
C85 VDD p2 4.16fF
C86 unit_cap_mim_m3m4_28/c1_n530_n480# op 0.17fF
C87 transmission_gate_6/in transmission_gate_3/out 0.76fF
C88 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C89 p1_b cm 1.15fF
C90 unit_cap_mim_m3m4_16/m3_n630_n580# transmission_gate_9/in 0.17fF
C91 cmc op 4.24fF
C92 transmission_gate_6/in unit_cap_mim_m3m4_28/c1_n530_n480# 0.05fF
C93 cmc unit_cap_mim_m3m4_21/m3_n630_n580# 0.69fF
C94 transmission_gate_4/out on 3.24fF
C95 unit_cap_mim_m3m4_24/m3_n630_n580# p2 0.05fF
C96 transmission_gate_6/in cmc 1.15fF
C97 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C98 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C99 p1 bias_a 0.81fF
C100 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C101 unit_cap_mim_m3m4_31/c1_n530_n480# transmission_gate_4/out 0.05fF
C102 op VDD 0.89fF
C103 transmission_gate_7/in on 3.12fF
C104 p1 transmission_gate_8/in 0.39fF
C105 p2_b on 0.34fF
C106 unit_cap_mim_m3m4_21/c1_n530_n480# on 0.06fF
C107 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C108 p1 unit_cap_mim_m3m4_27/c1_n530_n480# 0.11fF
C109 op unit_cap_mim_m3m4_23/c1_n530_n480# 0.13fF
C110 p1 unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C111 transmission_gate_6/in VDD 0.03fF
C112 op unit_cap_mim_m3m4_30/c1_n530_n480# 0.18fF
C113 unit_cap_mim_m3m4_17/m3_n630_n580# p2 0.04fF
C114 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.17fF
C115 transmission_gate_4/out unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C116 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580# -0.21fF
C117 p1 transmission_gate_4/out 0.80fF
C118 unit_cap_mim_m3m4_29/c1_n530_n480# p2 0.04fF
C119 bias_a transmission_gate_9/in 0.02fF
C120 unit_cap_mim_m3m4_20/m3_n630_n580# on 0.61fF
C121 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C122 op p2 0.16fF
C123 transmission_gate_8/in transmission_gate_9/in 3.35fF
C124 bias_a transmission_gate_3/out 0.07fF
C125 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580# -0.37fF
C126 p1_b unit_cap_mim_m3m4_35/m3_n630_n580# 0.01fF
C127 transmission_gate_7/in unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C128 p1_b on 0.45fF
C129 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C130 transmission_gate_8/in transmission_gate_3/out 0.24fF
C131 p1 transmission_gate_7/in 0.39fF
C132 transmission_gate_8/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C133 p1 p2_b 2.16fF
C134 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580# -0.12fF
C135 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.10fF
C136 transmission_gate_6/in p2 0.61fF
C137 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.10fF
C138 unit_cap_mim_m3m4_28/m3_n630_n580# op 0.66fF
C139 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C140 p1_b unit_cap_mim_m3m4_29/m3_n630_n580# 0.05fF
C141 unit_cap_mim_m3m4_23/m3_n630_n580# p1_b 0.05fF
C142 unit_cap_mim_m3m4_28/m3_n630_n580# transmission_gate_6/in -0.13fF
C143 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C144 unit_cap_mim_m3m4_16/m3_n630_n580# p2 0.05fF
C145 cmc transmission_gate_8/in 8.44fF
C146 op unit_cap_mim_m3m4_29/c1_n530_n480# 0.03fF
C147 transmission_gate_4/out transmission_gate_9/in 3.02fF
C148 transmission_gate_4/out transmission_gate_3/out 0.37fF
C149 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.17fF
C150 cmc unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C151 transmission_gate_6/in unit_cap_mim_m3m4_29/c1_n530_n480# -0.37fF
C152 unit_cap_mim_m3m4_20/m3_n630_n580# p1 0.06fF
C153 p1_b unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C154 transmission_gate_7/in transmission_gate_9/in 0.02fF
C155 bias_a VDD 0.99fF
C156 transmission_gate_6/in op 0.60fF
C157 p2_b transmission_gate_9/in 0.01fF
C158 transmission_gate_7/in transmission_gate_3/out 0.29fF
C159 transmission_gate_8/in VDD -0.07fF
C160 p1 p1_b 8.88fF
C161 transmission_gate_7/in unit_cap_mim_m3m4_19/m3_n630_n580# -0.28fF
C162 p2_b transmission_gate_3/out 0.10fF
C163 cmc transmission_gate_4/out 0.10fF
C164 unit_cap_mim_m3m4_28/c1_n530_n480# transmission_gate_7/in 0.06fF
C165 unit_cap_mim_m3m4_20/c1_n530_n480# on 0.15fF
C166 op unit_cap_mim_m3m4_30/m3_n630_n580# 0.56fF
C167 cmc transmission_gate_7/in 0.07fF
C168 cmc p2_b 0.12fF
C169 unit_cap_mim_m3m4_21/c1_n530_n480# cmc 0.13fF
C170 transmission_gate_4/out VDD -0.06fF
C171 unit_cap_mim_m3m4_18/c1_n530_n480# on 0.06fF
C172 bias_a p2 0.60fF
C173 unit_cap_mim_m3m4_26/c1_n530_n480# p1_b 0.06fF
C174 transmission_gate_4/out unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C175 p1_b transmission_gate_9/in 0.59fF
C176 transmission_gate_8/in p2 0.63fF
C177 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_24/c1_n530_n480# 0.06fF
C178 transmission_gate_4/out unit_cap_mim_m3m4_30/c1_n530_n480# -0.37fF
C179 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_16/c1_n530_n480# -0.21fF
C180 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# -0.25fF
C181 op unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C182 p1_b transmission_gate_3/out 0.59fF
C183 VDD transmission_gate_7/in -0.16fF
C184 p1_b unit_cap_mim_m3m4_19/m3_n630_n580# 0.06fF
C185 unit_cap_mim_m3m4_27/c1_n530_n480# p2 0.04fF
C186 p1 unit_cap_mim_m3m4_24/c1_n530_n480# 0.11fF
C187 p2_b VDD 1.67fF
C188 unit_cap_mim_m3m4_28/m3_n630_n580# transmission_gate_8/in 0.10fF
C189 unit_cap_mim_m3m4_28/c1_n530_n480# p1_b 0.06fF
C190 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C191 cmc p1_b 0.53fF
C192 transmission_gate_4/out p2 0.15fF
C193 unit_cap_mim_m3m4_22/c1_n530_n480# transmission_gate_9/in -0.37fF
C194 op transmission_gate_8/in 0.86fF
C195 p1 cm 1.50fF
C196 unit_cap_mim_m3m4_21/m3_n630_n580# transmission_gate_8/in -1.15fF
C197 transmission_gate_6/in bias_a 0.07fF
C198 op unit_cap_mim_m3m4_27/c1_n530_n480# 0.01fF
C199 transmission_gate_7/in p2 0.60fF
C200 transmission_gate_6/in transmission_gate_8/in -0.31fF
C201 p2_b p2 6.58fF
C202 p1_b VDD 1.01fF
C203 transmission_gate_6/in unit_cap_mim_m3m4_27/c1_n530_n480# -0.13fF
C204 cmc unit_cap_mim_m3m4_22/c1_n530_n480# 0.13fF
C205 transmission_gate_6/in unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C206 transmission_gate_8/in unit_cap_mim_m3m4_34/m3_n630_n580# 0.57fF
C207 p1_b unit_cap_mim_m3m4_22/m3_n630_n580# 0.05fF
C208 transmission_gate_4/out op 1.08fF
C209 unit_cap_mim_m3m4_24/m3_n630_n580# p1_b 0.06fF
C210 unit_cap_mim_m3m4_31/m3_n630_n580# transmission_gate_9/in 0.12fF
C211 transmission_gate_6/in transmission_gate_4/out 0.46fF
C212 transmission_gate_9/in cm 0.04fF
C213 op transmission_gate_7/in 2.63fF
C214 transmission_gate_3/out cm 0.17fF
C215 unit_cap_mim_m3m4_23/m3_n630_n580# on 0.47fF
C216 op p2_b 0.40fF
C217 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C218 p1_b p2 5.94fF
C219 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480# -0.19fF
C220 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580# -0.19fF
C221 transmission_gate_4/out unit_cap_mim_m3m4_16/m3_n630_n580# -0.28fF
C222 transmission_gate_6/in transmission_gate_7/in 0.45fF
C223 transmission_gate_6/in p2_b 0.42fF
C224 transmission_gate_4/out unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C225 p1_b unit_cap_mim_m3m4_17/m3_n630_n580# 0.06fF
C226 transmission_gate_4/out unit_cap_mim_m3m4_30/m3_n630_n580# -0.80fF
C227 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C228 p1 unit_cap_mim_m3m4_35/m3_n630_n580# 0.07fF
C229 p1 on 0.49fF
C230 unit_cap_mim_m3m4_29/c1_n530_n480# p1_b 0.06fF
C231 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_24/c1_n530_n480# -0.30fF
C232 bias_a transmission_gate_8/in 0.04fF
C233 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_17/c1_n530_n480# -0.20fF
C234 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.17fF
C235 op p1_b 0.28fF
C236 p1 unit_cap_mim_m3m4_29/m3_n630_n580# 0.06fF
C237 VDD cm 1.83fF
C238 unit_cap_mim_m3m4_23/m3_n630_n580# p1 0.06fF
C239 p1_b unit_cap_mim_m3m4_21/m3_n630_n580# 0.05fF
C240 unit_cap_mim_m3m4_24/c1_n530_n480# p2 0.04fF
C241 transmission_gate_6/in p1_b 0.41fF
C242 unit_cap_mim_m3m4_32/c1_n530_n480# on 0.06fF
C243 op unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C244 unit_cap_mim_m3m4_26/c1_n530_n480# on 0.06fF
C245 cmc unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C246 on transmission_gate_9/in 1.05fF
C247 p1 unit_cap_mim_m3m4_25/c1_n530_n480# 0.11fF
C248 transmission_gate_4/out bias_a 0.10fF
C249 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_32/m3_n630_n580# 0.12fF
C250 p1_b unit_cap_mim_m3m4_16/m3_n630_n580# 0.06fF
C251 unit_cap_mim_m3m4_19/c1_n530_n480# transmission_gate_7/in 0.06fF
C252 op unit_cap_mim_m3m4_22/c1_n530_n480# 0.07fF
C253 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C254 transmission_gate_3/out on 0.40fF
C255 transmission_gate_4/out transmission_gate_8/in 0.26fF
C256 p1_b unit_cap_mim_m3m4_30/m3_n630_n580# 0.01fF
C257 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C258 bias_a transmission_gate_7/in 0.11fF
C259 p2 cm 1.33fF
C260 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_9/in 0.17fF
C261 p2_b bias_a 0.48fF
C262 transmission_gate_8/in transmission_gate_7/in 0.81fF
C263 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_3/out -0.30fF
C264 p2_b transmission_gate_8/in 0.40fF
C265 unit_cap_mim_m3m4_21/c1_n530_n480# transmission_gate_8/in -0.41fF
C266 cmc on 1.91fF
C267 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C268 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_20/c1_n530_n480# 0.06fF
C269 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C270 p1 unit_cap_mim_m3m4_26/c1_n530_n480# 0.11fF
C271 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C272 p1 transmission_gate_9/in 0.70fF
C273 transmission_gate_4/out transmission_gate_7/in 0.61fF
C274 VDD on 0.88fF
C275 op unit_cap_mim_m3m4_31/m3_n630_n580# 0.03fF
C276 p1 transmission_gate_3/out 0.72fF
C277 p1 unit_cap_mim_m3m4_19/m3_n630_n580# 0.08fF
C278 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C279 transmission_gate_4/out p2_b 0.05fF
C280 unit_cap_mim_m3m4_20/m3_n630_n580# transmission_gate_8/in 0.17fF
C281 unit_cap_mim_m3m4_23/c1_n530_n480# on 0.19fF
C282 p1_b bias_a 0.52fF
C283 p1 unit_cap_mim_m3m4_28/c1_n530_n480# 0.11fF
C284 transmission_gate_6/in cm 0.17fF
C285 p1_b transmission_gate_8/in 0.17fF
C286 p2_b transmission_gate_7/in 0.41fF
C287 p1_b unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C288 p1 cmc 0.49fF
C289 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C290 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.39fF
C291 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C292 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.51fF
C293 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C294 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.74fF
C295 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C296 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.51fF
C297 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.51fF
C298 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.82fF
C299 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.60fF
C300 cmc VSS -31.94fF
C301 transmission_gate_9/in VSS 3.96fF
C302 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.61fF
C303 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.61fF
C304 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C305 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C306 p2 VSS 148.24fF
C307 p2_b VSS 41.62fF
C308 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.84fF
C309 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C310 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.39fF
C311 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C312 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.04fF
C313 transmission_gate_4/out VSS -3.74fF
C314 transmission_gate_3/out VSS 2.28fF
C315 p1 VSS 111.99fF
C316 transmission_gate_8/in VSS 2.29fF
C317 bias_a VSS 11.61fF
C318 transmission_gate_6/in VSS -13.31fF
C319 transmission_gate_7/in VSS 9.28fF
C320 cm VSS 13.12fF
C321 op VSS -1.36fF
C322 p1_b VSS 173.74fF
C323 VDD VSS 71.01fF
C324 on VSS -23.21fF
.ends

.subckt ota_w_test_v2 ip in p1 p1_b p2 p2_b op on i_bias cm bias_a bias_b bias_c bias_d
+ cmc VDD VSS
Xota_v2_without_cmfb_0 in bias_c cm op on i_bias VDD VSS ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596#
+ cmc ota_v2_without_cmfb_0/li_14138_570# bias_d ota_v2_without_cmfb_0/li_11121_570#
+ ota_v2_without_cmfb_0/li_11122_5650# ota_v2_without_cmfb_0/li_8434_570# bias_b ota_v2_without_cmfb_0/li_8436_5651#
+ ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997#
+ bias_a ip ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# ota_v2_without_cmfb
Xsc_cmfb_0 cm op cmc p2_b p2 on sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_4/out
+ sc_cmfb_0/transmission_gate_8/in bias_a p1 VDD sc_cmfb_0/transmission_gate_3/out
+ sc_cmfb_0/transmission_gate_7/in VSS p1_b sc_cmfb
C0 ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VDD 0.00fF
C1 p1_b p1 0.00fF
C2 bias_c cm 2.51fF
C3 ota_v2_without_cmfb_0/li_14138_570# ota_v2_without_cmfb_0/li_8436_5651# 0.00fF
C4 ip op 0.01fF
C5 op p1 0.01fF
C6 ota_v2_without_cmfb_0/li_11121_570# bias_d -0.00fF
C7 ota_v2_without_cmfb_0/li_8436_5651# on 0.26fF
C8 cmc op 0.38fF
C9 bias_a cm 3.21fF
C10 cm VDD -0.07fF
C11 ota_v2_without_cmfb_0/li_8434_570# on 0.98fF
C12 ota_v2_without_cmfb_0/li_14138_570# op 0.00fF
C13 cm bias_d 4.04fF
C14 p1_b on 0.02fF
C15 op on 3.07fF
C16 sc_cmfb_0/transmission_gate_4/out VDD 0.04fF
C17 ota_v2_without_cmfb_0/li_14138_570# in -0.00fF
C18 ip ota_v2_without_cmfb_0/li_14138_570# -0.00fF
C19 p1 sc_cmfb_0/transmission_gate_8/in 0.00fF
C20 bias_c ota_v2_without_cmfb_0/li_8436_5651# 0.00fF
C21 cmc p1 -0.00fF
C22 VDD sc_cmfb_0/transmission_gate_7/in 0.01fF
C23 cm ota_v2_without_cmfb_0/li_11121_570# 0.38fF
C24 cmc sc_cmfb_0/transmission_gate_8/in -0.03fF
C25 p1 on 0.01fF
C26 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.02fF
C27 cmc ota_v2_without_cmfb_0/li_14138_570# 0.03fF
C28 ota_v2_without_cmfb_0/li_8436_5651# ota_v2_without_cmfb_0/li_11122_5650# -0.01fF
C29 ota_v2_without_cmfb_0/li_8436_5651# VDD -0.11fF
C30 bias_c op 1.79fF
C31 cmc on 0.30fF
C32 ota_v2_without_cmfb_0/li_14138_570# on 0.54fF
C33 bias_c i_bias 0.00fF
C34 ota_v2_without_cmfb_0/li_8434_570# bias_a -0.00fF
C35 ota_v2_without_cmfb_0/li_8434_570# bias_d -0.00fF
C36 p1_b VDD -0.01fF
C37 bias_a p1_b 0.00fF
C38 op ota_v2_without_cmfb_0/li_11122_5650# 0.94fF
C39 op VDD 0.52fF
C40 ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VDD 0.00fF
C41 op bias_d -0.00fF
C42 bias_c bias_b 0.26fF
C43 bias_a p1 0.00fF
C44 bias_c on 0.00fF
C45 op ota_v2_without_cmfb_0/li_11121_570# -0.00fF
C46 VDD ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# 0.00fF
C47 VDD sc_cmfb_0/transmission_gate_8/in 0.02fF
C48 bias_a sc_cmfb_0/transmission_gate_8/in 0.00fF
C49 ota_v2_without_cmfb_0/li_8434_570# cm 0.37fF
C50 cmc VDD -0.06fF
C51 ota_v2_without_cmfb_0/li_14138_570# bias_a -0.04fF
C52 p1_b cm 0.01fF
C53 bias_b ota_v2_without_cmfb_0/li_11122_5650# -0.00fF
C54 bias_a bias_b 0.15fF
C55 bias_b VDD 0.16fF
C56 ota_v2_without_cmfb_0/li_11122_5650# on 0.43fF
C57 op cm 1.40fF
C58 VDD on 2.12fF
C59 bias_a on 0.27fF
C60 cmc p2 0.01fF
C61 on bias_d 12.62fF
C62 sc_cmfb_0/transmission_gate_4/out p1_b 0.00fF
C63 p2_b p1 0.00fF
C64 bias_c ota_v2_without_cmfb_0/li_11122_5650# 0.00fF
C65 ota_v2_without_cmfb_0/li_11121_570# on 1.99fF
C66 bias_c bias_a 2.52fF
C67 sc_cmfb_0/transmission_gate_3/out p1 -0.00fF
C68 cmc cm -2.78fF
C69 sc_cmfb_0/transmission_gate_4/out p1 0.05fF
C70 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# cm 0.23fF
C71 ota_v2_without_cmfb_0/li_14138_570# cm 1.28fF
C72 ota_v2_without_cmfb_0/li_8436_5651# op 0.62fF
C73 bias_b cm 3.45fF
C74 cm on 3.38fF
C75 ota_v2_without_cmfb_0/li_11122_5650# VDD 0.21fF
C76 bias_a VDD 0.02fF
C77 op p1_b 0.01fF
C78 bias_a bias_d -0.00fF
C79 sc_cmfb_0/transmission_gate_3/out on 0.01fF
C80 ip ota_v2_without_cmfb_0/li_8436_5651# -0.00fF
C81 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C82 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C83 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C84 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C85 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C86 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C87 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C88 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C89 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C90 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.37fF
C91 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C92 sc_cmfb_0/transmission_gate_9/in VSS 2.57fF
C93 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C94 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C95 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C96 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C97 p2 VSS 147.98fF
C98 p2_b VSS 40.26fF
C99 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C100 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C101 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C102 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C103 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.86fF
C104 sc_cmfb_0/transmission_gate_4/out VSS -4.88fF
C105 sc_cmfb_0/transmission_gate_3/out VSS 1.20fF
C106 p1 VSS 111.49fF
C107 sc_cmfb_0/transmission_gate_8/in VSS 1.02fF
C108 sc_cmfb_0/transmission_gate_6/in VSS -14.71fF
C109 sc_cmfb_0/transmission_gate_7/in VSS 7.86fF
C110 cm VSS 33.63fF
C111 op VSS 8.47fF
C112 p1_b VSS 173.22fF
C113 on VSS -28.09fF
C114 ota_v2_without_cmfb_0/m1_17393_3568# VSS 0.03fF $ **FLOATING
C115 ota_v2_without_cmfb_0/m1_15613_3568# VSS 0.05fF $ **FLOATING
C116 ota_v2_without_cmfb_0/m1_18877_3928# VSS 0.05fF $ **FLOATING
C117 ota_v2_without_cmfb_0/m1_17097_3928# VSS 0.04fF $ **FLOATING
C118 ota_v2_without_cmfb_0/li_11121_570# VSS 9.30fF
C119 ota_v2_without_cmfb_0/li_11122_5650# VSS -33.11fF
C120 ota_v2_without_cmfb_0/li_8434_570# VSS 9.00fF
C121 bias_a VSS -301.05fF
C122 ota_v2_without_cmfb_0/li_8436_5651# VSS 3.26fF
C123 ota_v2_without_cmfb_0/bias_circuit_0/m1_3551_3596# VSS -342.20fF
C124 bias_b VSS -361.59fF
C125 ota_v2_without_cmfb_0/bias_circuit_0/m1_5643_5997# VSS 38.05fF
C126 ota_v2_without_cmfb_0/bias_circuit_0/m1_3443_5997# VSS 35.85fF
C127 ota_v2_without_cmfb_0/bias_circuit_0/m1_1243_5997# VSS 25.03fF
C128 VDD VSS 358.95fF
C129 i_bias VSS -61.82fF
C130 bias_c VSS -130.38fF
C131 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_427# VSS 0.11fF
C132 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_423# VSS 0.11fF
C133 ota_v2_without_cmfb_0/bias_circuit_0/m1_7461_921# VSS 0.12fF
C134 ota_v2_without_cmfb_0/bias_circuit_0/m1_7169_923# VSS 0.13fF
C135 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_433# VSS 0.14fF
C136 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_422# VSS 0.20fF
C137 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_422# VSS 0.20fF
C138 ota_v2_without_cmfb_0/bias_circuit_0/m1_7639_1420# VSS 0.12fF
C139 ota_v2_without_cmfb_0/bias_circuit_0/m1_7347_1428# VSS 0.13fF
C140 ota_v2_without_cmfb_0/bias_circuit_0/m1_6877_922# VSS 0.14fF
C141 ota_v2_without_cmfb_0/bias_circuit_0/m1_6585_923# VSS 0.22fF
C142 ota_v2_without_cmfb_0/bias_circuit_0/m1_6293_922# VSS 0.16fF
C143 ota_v2_without_cmfb_0/bias_circuit_0/m1_7055_1417# VSS 0.14fF
C144 ota_v2_without_cmfb_0/bias_circuit_0/m1_6763_1422# VSS 0.22fF
C145 ota_v2_without_cmfb_0/bias_circuit_0/m1_6471_1426# VSS 0.22fF
C146 bias_d VSS -231.85fF
C147 ota_v2_without_cmfb_0/bias_circuit_0/li_3433_399# VSS 4.65fF
C148 ota_v2_without_cmfb_0/li_14138_570# VSS 17.77fF
C149 cmc VSS -141.66fF
C150 in VSS -28.55fF
C151 ip VSS -27.04fF
.ends

