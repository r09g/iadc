magic
tech sky130A
magscale 1 2
timestamp 1654766757
<< pwell >>
rect 388066 484631 388240 485269
rect 388002 463587 388176 464225
rect 251604 454544 251778 455182
rect 388034 442623 388208 443261
rect 251590 433523 251764 434161
rect 385510 422705 386148 422879
rect 386152 421261 386790 421435
<< viali >>
rect 387972 485193 388088 485249
rect 388006 484815 388098 484863
rect 387908 464149 388024 464205
rect 387942 463771 388034 463819
rect 251510 455106 251626 455162
rect 251544 454728 251636 454776
rect 387940 443185 388056 443241
rect 387974 442807 388066 442855
rect 251496 434085 251612 434141
rect 251530 433707 251622 433755
rect 385694 422847 385742 422939
rect 386072 422857 386128 422973
rect 386336 421403 386384 421495
rect 386714 421413 386770 421529
<< metal1 >>
rect 266353 537651 266415 537727
rect 387960 485249 388100 485255
rect 387960 485193 387972 485249
rect 388088 485193 388100 485249
rect 387960 485187 388100 485193
rect 387994 484811 388006 484869
rect 388098 484811 388110 484869
rect 387994 484809 388110 484811
rect 387896 464205 388036 464211
rect 387896 464149 387908 464205
rect 388024 464149 388036 464205
rect 387896 464143 388036 464149
rect 387930 463767 387942 463825
rect 388034 463767 388046 463825
rect 387930 463765 388046 463767
rect 251498 455162 251638 455168
rect 251498 455106 251510 455162
rect 251626 455106 251638 455162
rect 251498 455100 251638 455106
rect 251532 454724 251544 454782
rect 251636 454724 251648 454782
rect 251532 454722 251648 454724
rect 387928 443241 388068 443247
rect 387928 443185 387940 443241
rect 388056 443185 388068 443241
rect 387928 443179 388068 443185
rect 387962 442803 387974 442861
rect 388066 442803 388078 442861
rect 387962 442801 388078 442803
rect 251484 434141 251624 434147
rect 251484 434085 251496 434141
rect 251612 434085 251624 434141
rect 251484 434079 251624 434085
rect 251518 433703 251530 433761
rect 251622 433703 251634 433761
rect 251518 433701 251634 433703
rect 386066 422973 386134 422985
rect 385688 422939 385748 422951
rect 385688 422847 385690 422939
rect 385688 422835 385748 422847
rect 386066 422857 386072 422973
rect 386128 422857 386134 422973
rect 386066 422845 386134 422857
rect 386708 421529 386776 421541
rect 386330 421495 386390 421507
rect 386330 421403 386332 421495
rect 386330 421391 386390 421403
rect 386708 421413 386714 421529
rect 386770 421413 386776 421529
rect 386708 421401 386776 421413
<< via1 >>
rect 387972 485193 388088 485249
rect 388006 484863 388098 484869
rect 388006 484815 388098 484863
rect 388006 484811 388098 484815
rect 387908 464149 388024 464205
rect 387942 463819 388034 463825
rect 387942 463771 388034 463819
rect 387942 463767 388034 463771
rect 251510 455106 251626 455162
rect 251544 454776 251636 454782
rect 251544 454728 251636 454776
rect 251544 454724 251636 454728
rect 387940 443185 388056 443241
rect 387974 442855 388066 442861
rect 387974 442807 388066 442855
rect 387974 442803 388066 442807
rect 251496 434085 251612 434141
rect 251530 433755 251622 433761
rect 251530 433707 251622 433755
rect 251530 433703 251622 433707
rect 385690 422847 385694 422939
rect 385694 422847 385742 422939
rect 385742 422847 385748 422939
rect 386072 422857 386128 422973
rect 386332 421403 386336 421495
rect 386336 421403 386384 421495
rect 386384 421403 386390 421495
rect 386714 421413 386770 421529
<< metal2 >>
rect 266346 537652 266426 537724
rect 387972 485249 388088 485259
rect 387972 485183 388088 485193
rect 388006 484869 388098 484879
rect 388006 484801 388098 484811
rect 387908 464205 388024 464215
rect 387908 464139 388024 464149
rect 387942 463825 388034 463835
rect 387942 463757 388034 463767
rect 251510 455162 251626 455172
rect 251510 455096 251626 455106
rect 251544 454782 251636 454792
rect 251544 454714 251636 454724
rect 387940 443241 388056 443251
rect 387940 443175 388056 443185
rect 387974 442861 388066 442871
rect 387974 442793 388066 442803
rect 251496 434141 251612 434151
rect 251496 434075 251612 434085
rect 251530 433761 251622 433771
rect 251530 433693 251622 433703
rect 385680 422847 385690 422939
rect 385748 422847 385758 422939
rect 386062 422857 386072 422973
rect 386128 422857 386138 422973
rect 386322 421403 386332 421495
rect 386390 421403 386400 421495
rect 386704 421413 386714 421529
rect 386770 421413 386780 421529
<< via2 >>
rect 387972 485193 388088 485249
rect 388006 484811 388098 484869
rect 387908 464149 388024 464205
rect 387942 463767 388034 463825
rect 251510 455106 251626 455162
rect 251544 454724 251636 454782
rect 387940 443185 388056 443241
rect 387974 442803 388066 442861
rect 251496 434085 251612 434141
rect 251530 433703 251622 433761
rect 385690 422847 385748 422939
rect 386072 422857 386128 422973
rect 386332 421403 386390 421495
rect 386714 421413 386770 421529
<< metal3 >>
rect 15950 695660 21404 702751
rect 49800 695660 55254 695667
rect 15950 690206 55254 695660
rect 631 679916 41399 685370
rect 5444 648766 8456 648790
rect 878 643702 8456 648766
rect 13544 643702 13550 648790
rect 878 643700 6018 643702
rect 5444 638740 8464 638756
rect 878 633684 8464 638740
rect 13536 633684 13542 638756
rect 878 633674 6018 633684
rect 35945 617473 41399 679916
rect 49800 657879 55254 690206
rect 68171 673059 73394 702561
rect 119883 690210 125294 702715
rect 413264 690703 418526 702969
rect 119883 684799 260421 690210
rect 68171 667836 228031 673059
rect 49800 652425 203886 657879
rect 198432 646074 203886 652425
rect 222808 646074 228031 667836
rect 255010 646074 260421 684799
rect 285551 685441 418526 690703
rect 285551 646074 290813 685441
rect 465325 675451 470438 703028
rect 566483 693344 571777 703703
rect 308764 670338 470438 675451
rect 501812 688050 571777 693344
rect 308764 646074 313877 670338
rect 501812 655883 507106 688050
rect 571615 677583 583026 683351
rect 571615 665741 577383 677583
rect 342135 650589 507106 655883
rect 530234 659973 577383 665741
rect 342135 646074 347429 650589
rect 199583 623979 200583 646074
rect 224429 628120 225429 646074
rect 257917 640543 258917 646074
rect 238444 639543 258917 640543
rect 224429 627120 232372 628120
rect 199583 622979 217927 623979
rect 35945 615155 171274 617473
rect 35945 614155 210936 615155
rect 35945 612019 171274 614155
rect 209936 586305 210936 614155
rect 216927 586305 217927 622979
rect 231372 585884 232372 627120
rect 238444 587064 239444 639543
rect 287625 633521 288625 646074
rect 248446 632521 288625 633521
rect 248446 585722 249446 632521
rect 311030 628480 312030 646074
rect 259321 627480 312030 628480
rect 259321 585708 260321 627480
rect 344338 622358 345338 646074
rect 267631 621358 345338 622358
rect 267631 586608 268631 621358
rect 530234 618203 536002 659973
rect 570885 639606 570891 644708
rect 575993 644698 580085 644708
rect 575993 639606 583426 644698
rect 579000 639592 583426 639606
rect 579460 634688 583886 634762
rect 570940 629652 570946 634688
rect 575982 629656 583886 634688
rect 575982 629652 580085 629656
rect 356783 616237 536002 618203
rect 276971 615237 536002 616237
rect 276971 586610 277971 615237
rect 356783 612435 536002 615237
rect 286427 602572 481850 603572
rect 286427 584356 287427 602572
rect 288427 596104 482535 597104
rect 288427 586102 289427 596104
rect 290427 589091 479261 590091
rect 290427 585609 291427 589091
rect 336951 531611 366548 532611
rect 365548 522039 366548 531611
rect 365548 522021 368182 522039
rect 365548 521498 373220 522021
rect 365548 521438 374294 521498
rect 365548 521039 373220 521438
rect 367304 521021 373220 521039
rect 387975 507774 388242 507834
rect 387975 505419 388035 507774
rect 339054 504348 354532 505348
rect 337722 502341 352509 503341
rect 339853 500351 350532 501351
rect 336990 498341 348513 499341
rect 338721 496359 346532 497359
rect 340233 494344 344532 495344
rect 336760 492341 342546 493341
rect 341546 491341 342546 492341
rect 251027 455266 252027 458057
rect 251510 455167 251626 455266
rect 251500 455162 251636 455167
rect 251500 455106 251510 455162
rect 251626 455106 251636 455162
rect 251500 455101 251636 455106
rect 251534 454782 251646 454788
rect 251534 454724 251544 454782
rect 251636 454724 251646 454782
rect 251534 454464 251646 454724
rect 251027 434298 252027 454464
rect 339532 452388 340532 491341
rect 341532 490870 342546 491341
rect 341532 452388 342532 490870
rect 343532 452388 344532 494344
rect 345532 452388 346532 496359
rect 347513 491341 348513 498341
rect 347513 490897 348532 491341
rect 347532 452388 348532 490897
rect 349532 452388 350532 500351
rect 351509 491341 352509 502341
rect 351509 490298 352532 491341
rect 351532 452388 352532 490298
rect 353532 452388 354532 504348
rect 387498 485374 388498 505419
rect 387972 485254 388088 485374
rect 387962 485249 388098 485254
rect 387962 485193 387972 485249
rect 388088 485193 388098 485249
rect 387962 485188 388098 485193
rect 387996 484869 388108 484875
rect 387996 484811 388006 484869
rect 388098 484811 388108 484869
rect 387996 484534 388108 484811
rect 387498 464330 388498 484534
rect 387908 464210 388024 464330
rect 387898 464205 388034 464210
rect 387898 464149 387908 464205
rect 388024 464149 388034 464205
rect 387898 464144 388034 464149
rect 387932 463825 388044 463831
rect 387932 463767 387942 463825
rect 388034 463767 388044 463825
rect 387932 463476 388044 463767
rect 387498 443364 388498 463476
rect 387940 443246 388056 443364
rect 387930 443241 388066 443246
rect 387930 443185 387940 443241
rect 388056 443185 388066 443241
rect 387930 443180 388066 443185
rect 387964 442861 388076 442867
rect 387964 442803 387974 442861
rect 388066 442803 388076 442861
rect 387964 442534 388076 442803
rect 251496 434146 251612 434298
rect 251486 434141 251622 434146
rect 251486 434085 251496 434141
rect 251612 434085 251622 434141
rect 251486 434080 251622 434085
rect 251520 433761 251632 433767
rect 251520 433703 251530 433761
rect 251622 433703 251632 433761
rect 251520 433440 251632 433703
rect 251027 422028 252027 433440
rect 386067 422973 386133 422983
rect 385429 422939 385754 422949
rect 385429 422847 385690 422939
rect 385748 422847 385754 422939
rect 386067 422857 386072 422973
rect 386128 422857 386235 422973
rect 386067 422847 386133 422857
rect 385429 422837 385754 422847
rect 387498 422029 388498 442534
rect 251022 421030 251028 422028
rect 252026 421030 252032 422028
rect 386300 421372 386310 421531
rect 386409 421372 386419 421531
rect 386688 421402 386698 421554
rect 386788 421402 386798 421554
rect 251027 421029 252027 421030
rect 387492 421029 387498 422029
rect 388498 421029 388504 422029
rect 570568 191344 570574 196304
rect 575534 196302 580085 196304
rect 575534 191344 583140 196302
rect 579028 191326 583140 191344
rect 570481 181266 570487 186384
rect 575605 186382 580085 186384
rect 575605 185276 583718 186382
rect 575605 181270 583716 185276
rect 575605 181266 580085 181270
rect 1063 172756 13139 177874
rect 18257 172756 18263 177874
rect 881 162758 13447 167876
rect 18565 162758 18571 167876
<< via3 >>
rect 8456 643702 13544 648790
rect 8464 633684 13536 638756
rect 570891 639606 575993 644708
rect 570946 629652 575982 634688
rect 251028 421030 252026 422028
rect 386310 421495 386409 421531
rect 386310 421403 386332 421495
rect 386332 421403 386390 421495
rect 386390 421403 386409 421495
rect 386310 421372 386409 421403
rect 386698 421529 386788 421554
rect 386698 421413 386714 421529
rect 386714 421413 386770 421529
rect 386770 421413 386788 421529
rect 386698 421402 386788 421413
rect 387498 421029 388498 422029
rect 570574 191344 575534 196304
rect 570487 181266 575605 186384
rect 13139 172756 18257 177874
rect 13447 162758 18565 167876
<< metal4 >>
rect 131094 648766 136182 649988
rect 131094 643726 131292 648766
rect 131094 638732 136182 643726
rect 131094 633708 131116 638732
rect 136140 633708 136182 638732
rect 118401 580355 123519 614385
rect 131094 584249 136182 633708
rect 437148 605510 442248 629615
rect 378880 584090 379500 584289
rect 437148 584151 442236 605510
rect 396704 584094 397324 584150
rect 118401 577849 118427 580355
rect 123347 577849 123519 580355
rect 118401 467405 123519 577849
rect 118401 177850 123519 465142
rect 131094 463309 136182 581889
rect 377640 533154 378260 578117
rect 378880 533845 379500 582075
rect 396704 533938 397324 582079
rect 397944 580082 398564 580216
rect 437148 578620 442236 581974
rect 449741 580130 454859 612043
rect 397944 533213 398564 578067
rect 437148 530365 442248 578620
rect 442222 529695 442248 530365
rect 437148 513420 442248 529695
rect 449741 531582 454859 578012
rect 449741 530912 449785 531582
rect 437148 512750 437176 513420
rect 377640 467305 378260 509841
rect 377640 465251 378260 465299
rect 136108 461046 136182 463309
rect 378880 463303 379500 509113
rect 396704 463291 397324 509321
rect 397944 467304 398564 508905
rect 437148 463390 442248 512750
rect 449741 512189 454859 530912
rect 449741 511519 449744 512189
rect 454845 511519 454859 512189
rect 449741 467435 454859 511519
rect 449741 465172 449747 467435
rect 131094 201256 136182 461046
rect 387497 422029 388499 422030
rect 251027 422028 386010 422029
rect 251027 421030 251028 422028
rect 252026 421539 386010 422028
rect 386697 421554 386789 421555
rect 386960 421554 387498 422029
rect 252026 421531 386423 421539
rect 252026 421372 386310 421531
rect 386409 421372 386423 421531
rect 386692 421402 386698 421554
rect 386788 421402 387498 421554
rect 386697 421401 386789 421402
rect 252026 421366 386423 421372
rect 252026 421030 386010 421366
rect 251027 421029 386010 421030
rect 386960 421029 387498 421402
rect 388498 421029 388499 422029
rect 387497 421028 388499 421029
rect 437148 195286 442248 461127
rect 449741 196280 454859 465172
rect 454508 191368 454859 196280
rect 449741 186360 454859 191368
rect 575533 196304 575535 196305
rect 575534 191344 575535 196304
rect 575533 191343 575535 191344
rect 454587 181290 454859 186360
rect 123471 172780 123519 177850
rect 118401 167852 123519 172780
rect 123337 162782 123519 167852
rect 449741 177850 454859 181290
rect 449741 172780 449949 177850
rect 449741 167852 454859 172780
rect 449741 163009 449811 167852
rect 118401 160075 123519 162782
<< via4 >>
rect 8455 648790 13545 648791
rect 8455 643702 8456 648790
rect 8456 643702 13544 648790
rect 13544 643702 13545 648790
rect 8455 643701 13545 643702
rect 131292 643726 136332 648766
rect 8463 638756 13537 638757
rect 8463 633684 8464 638756
rect 8464 633684 13536 638756
rect 13536 633684 13537 638756
rect 8463 633683 13537 633684
rect 131116 633708 136140 638732
rect 437096 629615 442307 648816
rect 570890 644708 575994 644709
rect 570890 639606 570891 644708
rect 570891 639606 575993 644708
rect 575993 639606 575994 644708
rect 570890 639605 575994 639606
rect 570945 634688 575983 634689
rect 570945 629652 570946 634688
rect 570946 629652 575982 634688
rect 575982 629652 575983 634688
rect 570945 629651 575983 629652
rect 131057 581889 136194 584249
rect 378865 582075 379542 584090
rect 396657 582079 397334 584094
rect 118427 577849 123347 580355
rect 118375 465142 123527 467405
rect 13138 177874 18258 177875
rect 13138 172756 13139 177874
rect 13139 172756 18257 177874
rect 18257 172756 18258 177874
rect 13138 172755 18258 172756
rect 377518 578117 378369 580063
rect 437110 581974 442245 584151
rect 397931 578067 398608 580082
rect 449720 578012 454860 580130
rect 437121 529695 442222 530365
rect 449785 530912 454886 531582
rect 437176 512750 442277 513420
rect 377585 465299 378302 467305
rect 130956 461046 136108 463309
rect 378855 461297 379572 463303
rect 397927 465298 398644 467304
rect 449744 511519 454845 512189
rect 449747 465172 454899 467435
rect 396654 461285 397371 463291
rect 437131 461127 442283 463390
rect 449596 191368 454508 196280
rect 570573 196304 575533 196305
rect 570573 191344 570574 196304
rect 570574 191344 575533 196304
rect 570573 191343 575533 191344
rect 449517 181290 454587 186360
rect 118401 172780 123471 177850
rect 13446 167876 18566 167877
rect 13446 162758 13447 167876
rect 13447 162758 18565 167876
rect 18565 162758 18566 167876
rect 118267 162782 123337 167852
rect 570486 186384 575606 186385
rect 570486 181266 570487 186384
rect 570487 181266 575605 186384
rect 575605 181266 575606 186384
rect 570486 181265 575606 181266
rect 449949 172780 455019 177850
rect 449811 162782 454881 167852
rect 13446 162757 18566 162758
<< metal5 >>
rect 437072 648816 442331 648840
rect 8431 648791 13569 648815
rect 8431 643701 8455 648791
rect 13545 648790 13569 648791
rect 437072 648790 437096 648816
rect 13545 648766 437096 648790
rect 13545 643726 131292 648766
rect 136332 643726 437096 648766
rect 13545 643702 437096 643726
rect 13545 643701 13569 643702
rect 8431 643677 13569 643701
rect 8439 638757 13561 638781
rect 8439 633683 8463 638757
rect 13537 638756 13561 638757
rect 437072 638756 437096 643702
rect 13537 638732 437096 638756
rect 13537 633708 131116 638732
rect 136140 633708 437096 638732
rect 13537 633684 437096 633708
rect 13537 633683 13561 633684
rect 8439 633659 13561 633683
rect 437072 629615 437096 633684
rect 442307 644708 442331 648816
rect 570866 644709 576018 644733
rect 570866 644708 570890 644709
rect 442307 639606 570890 644708
rect 442307 634688 442331 639606
rect 570866 639605 570890 639606
rect 575994 639605 576018 644709
rect 570866 639581 576018 639605
rect 570921 634689 576007 634713
rect 570921 634688 570945 634689
rect 442307 629652 570945 634688
rect 442307 629615 442331 629652
rect 570921 629651 570945 629652
rect 575983 629651 576007 634689
rect 570921 629627 576007 629651
rect 437072 629591 442331 629615
rect 131033 584249 136218 584273
rect 131033 581889 131057 584249
rect 136194 584076 136218 584249
rect 437086 584151 442269 584175
rect 378841 584090 379566 584114
rect 378841 584076 378865 584090
rect 136194 582076 181001 584076
rect 338096 582076 378865 584076
rect 136194 581889 136218 582076
rect 378841 582075 378865 582076
rect 379542 584076 379566 584090
rect 396633 584094 397358 584118
rect 396633 584076 396657 584094
rect 379542 582079 396657 584076
rect 397334 584076 397358 584094
rect 437086 584076 437110 584151
rect 397334 582079 437110 584076
rect 379542 582076 437110 582079
rect 379542 582075 379566 582076
rect 378841 582051 379566 582075
rect 396633 582055 397358 582076
rect 437086 581974 437110 582076
rect 442245 581974 442269 584151
rect 437086 581950 442269 581974
rect 131033 581865 136218 581889
rect 118403 580355 123371 580379
rect 118403 577849 118427 580355
rect 123347 580076 123371 580355
rect 449696 580130 454884 580154
rect 377494 580076 378393 580087
rect 397907 580082 398632 580106
rect 397907 580076 397931 580082
rect 123347 578076 180266 580076
rect 337001 580063 397931 580076
rect 337001 578117 377518 580063
rect 378369 578117 397931 580063
rect 337001 578076 397931 578117
rect 123347 577849 123371 578076
rect 397907 578067 397931 578076
rect 398608 580076 398632 580082
rect 449696 580076 449720 580130
rect 398608 578076 449720 580076
rect 398608 578067 398632 578076
rect 397907 578043 398632 578067
rect 449696 578012 449720 578076
rect 454860 580076 454884 580130
rect 454860 578076 454920 580076
rect 454860 578012 454884 578076
rect 449696 577988 454884 578012
rect 118403 577825 123371 577849
rect 449761 531582 454910 531606
rect 449761 531562 449785 531582
rect 400694 530942 449785 531562
rect 449761 530912 449785 530942
rect 454886 530912 454910 531582
rect 449761 530888 454910 530912
rect 437097 530365 442246 530389
rect 437097 530322 437121 530365
rect 401112 529702 437121 530322
rect 437097 529695 437121 529702
rect 442222 529695 442246 530365
rect 437097 529671 442246 529695
rect 437152 513420 442301 513444
rect 437152 513382 437176 513420
rect 400486 512762 437176 513382
rect 437152 512750 437176 512762
rect 442277 512750 442301 513420
rect 437152 512726 442301 512750
rect 449720 512189 454869 512213
rect 449720 512142 449744 512189
rect 401112 511522 449744 512142
rect 449720 511519 449744 511522
rect 454845 511519 454869 512189
rect 449720 511495 454869 511519
rect 449723 467435 454923 467459
rect 118351 467405 123551 467429
rect 118351 467294 118375 467405
rect 118243 465294 118375 467294
rect 118351 465142 118375 465294
rect 123527 467294 123551 467405
rect 377561 467305 378326 467329
rect 377561 467294 377585 467305
rect 123527 465299 377585 467294
rect 378302 467294 378326 467305
rect 397903 467304 398668 467328
rect 397903 467294 397927 467304
rect 378302 465299 397927 467294
rect 123527 465298 397927 465299
rect 398644 467294 398668 467304
rect 449723 467294 449747 467435
rect 398644 465298 449747 467294
rect 123527 465294 449747 465298
rect 123527 465142 123551 465294
rect 377561 465275 378326 465294
rect 397903 465274 398668 465294
rect 449723 465172 449747 465294
rect 454899 465172 454923 467435
rect 449723 465148 454923 465172
rect 118351 465118 123551 465142
rect 437107 463390 442307 463414
rect 130932 463309 136132 463333
rect 130932 463294 130956 463309
rect 130507 461294 130956 463294
rect 130932 461046 130956 461294
rect 136108 463294 136132 463309
rect 378831 463303 379596 463327
rect 378831 463294 378855 463303
rect 136108 461294 201876 463294
rect 318684 461297 378855 463294
rect 379572 463294 379596 463303
rect 396630 463294 397395 463315
rect 437107 463294 437131 463390
rect 379572 463291 437131 463294
rect 379572 461297 396654 463291
rect 318684 461294 396654 461297
rect 136108 461046 136132 461294
rect 378831 461273 379596 461294
rect 396630 461285 396654 461294
rect 397371 461294 437131 463291
rect 397371 461285 397395 461294
rect 396630 461261 397395 461285
rect 437107 461127 437131 461294
rect 442283 463294 442307 463390
rect 442283 461294 442558 463294
rect 442283 461127 442307 461294
rect 437107 461103 442307 461127
rect 130932 461022 136132 461046
rect 570549 196305 575557 196329
rect 570549 196304 570573 196305
rect 449572 196280 570573 196304
rect 449572 191368 449596 196280
rect 454508 191368 570573 196280
rect 449572 191344 570573 191368
rect 570549 191343 570573 191344
rect 575533 191343 575557 196305
rect 570549 191319 575557 191343
rect 570462 186385 575630 186409
rect 570462 186384 570486 186385
rect 449493 186360 570486 186384
rect 449493 181290 449517 186360
rect 454587 181290 570486 186360
rect 449493 181266 570486 181290
rect 570462 181265 570486 181266
rect 575606 181265 575630 186385
rect 570462 181241 575630 181265
rect 13114 177875 18282 177899
rect 13114 172755 13138 177875
rect 18258 177874 18282 177875
rect 18258 177850 455043 177874
rect 18258 172780 118401 177850
rect 123471 172780 449949 177850
rect 455019 172780 455043 177850
rect 18258 172756 455043 172780
rect 18258 172755 18282 172756
rect 13114 172731 18282 172755
rect 13422 167877 18590 167901
rect 13422 162757 13446 167877
rect 18566 167876 18590 167877
rect 18566 167852 454905 167876
rect 18566 162782 118267 167852
rect 123337 162782 449811 167852
rect 454881 162782 454905 167852
rect 18566 162758 454905 162782
rect 18566 162757 18590 162758
rect 13422 162733 18590 162757
use analog_top  analog_top_0
timestamp 1654755406
transform 1 0 173563 0 1 497679
box 4703 -40917 166970 91353
use digital_top  digital_top_0
timestamp 1654755406
transform 1 0 373703 0 1 507665
box 0 0 28796 27744
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 0 -1 251799 1 0 454633
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_1
timestamp 1650294714
transform 0 -1 388261 1 0 484720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_2
timestamp 1650294714
transform 0 -1 251785 1 0 433612
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_3
timestamp 1650294714
transform 0 -1 388197 1 0 463676
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_4
timestamp 1650294714
transform 0 -1 388229 1 0 442712
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_5
timestamp 1650294714
transform 1 0 385599 0 1 422684
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_6
timestamp 1650294714
transform 1 0 386241 0 1 421240
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1654752884
transform 0 -1 251799 1 0 454541
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1654752884
transform 0 -1 388261 1 0 484628
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1654752884
transform 0 -1 251785 1 0 433520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1654752884
transform 0 -1 388197 1 0 463584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1654752884
transform 0 -1 388229 1 0 442620
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1654752884
transform 1 0 385507 0 1 422684
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1654752884
transform 1 0 386149 0 1 421240
box -38 -48 130 592
<< labels >>
flabel metal5 19178 643940 30500 648236 1 FreeSans 32000 0 0 0 VDD
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
