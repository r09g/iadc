magic
tech sky130A
magscale 1 2
timestamp 1653911004
<< metal1 >>
rect -2068 8268 -2022 8360
rect 6932 8182 6978 8360
rect -3494 7647 -2106 7681
rect -3494 -1319 -3419 7647
rect -1032 7631 -1022 7695
rect -958 7631 -948 7695
rect -485 7681 2411 7697
rect -723 7647 2411 7681
rect -485 7633 2411 7647
rect 6681 7633 6691 7697
rect 6755 7681 6765 7697
rect 6755 7647 6899 7681
rect 8265 7647 9310 7681
rect 6755 7633 6765 7647
rect -2068 7160 -2022 7246
rect -2068 6382 -2022 6560
rect 1618 6412 1628 6476
rect 1692 6412 1702 6476
rect -2886 5847 -2090 5881
rect -2886 481 -2811 5847
rect -1038 5831 -1028 5895
rect -964 5831 -954 5895
rect -487 5881 -477 5893
rect -739 5847 -477 5881
rect -487 5829 -477 5847
rect -413 5829 -403 5893
rect -2068 5360 -2022 5532
rect -2068 4582 -2022 4760
rect -2428 4047 -2100 4081
rect -2428 2281 -2353 4047
rect -1034 4031 -1024 4095
rect -960 4031 -950 4095
rect -444 4081 -434 4094
rect -719 4047 -434 4081
rect -444 4030 -434 4047
rect -370 4030 -360 4094
rect 1628 3846 1692 6412
rect 2347 4563 2411 7633
rect 6932 7160 6978 7332
rect 6932 6382 6978 6560
rect 6694 5831 6704 5895
rect 6768 5881 6778 5895
rect 6768 5847 6894 5881
rect 8281 5847 8799 5881
rect 6768 5831 6778 5847
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 3157 5084 3221 5494
rect 6932 5360 6978 5532
rect 3147 5020 3157 5084
rect 3221 5020 3231 5084
rect 3831 4928 6166 4932
rect 3758 4864 3768 4928
rect 3832 4868 6166 4928
rect 6230 4868 6240 4932
rect 3832 4864 3842 4868
rect 6932 4582 6978 4760
rect 2347 4499 3106 4563
rect 3170 4499 3180 4563
rect 4874 4326 5207 4390
rect 5271 4326 5281 4390
rect 3298 4148 3308 4212
rect 3372 4148 3382 4212
rect 3308 4085 3372 4148
rect 1628 3782 1866 3846
rect -2068 3560 -2022 3732
rect 323 3419 333 3483
rect 397 3419 1631 3483
rect 1695 3419 1705 3483
rect 1802 3154 1866 3782
rect 323 3090 333 3154
rect 397 3090 1866 3154
rect -2068 2782 -2022 2960
rect -2428 2247 -2106 2281
rect -1037 2231 -1027 2295
rect -963 2231 -953 2295
rect -444 2281 -434 2291
rect -719 2247 -434 2281
rect -444 2227 -434 2247
rect -370 2227 -360 2291
rect 3308 2223 3371 4085
rect 4874 3642 4938 4326
rect 6749 4031 6759 4095
rect 6823 4081 6833 4095
rect 8724 4081 8799 5847
rect 6823 4047 6894 4081
rect 8271 4047 8799 4081
rect 6823 4031 6833 4047
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 6932 3560 6978 3732
rect 6932 2782 6978 2960
rect 6754 2233 6764 2297
rect 6828 2281 6838 2297
rect 8724 2281 8799 4047
rect 6828 2247 6894 2281
rect 8275 2247 8799 2281
rect 6828 2233 6838 2247
rect 3298 2159 3308 2223
rect 3372 2159 3382 2223
rect -2068 1760 -2022 1932
rect 6932 1760 6978 1932
rect -364 1576 2330 1640
rect 2394 1576 2404 1640
rect -2068 982 -2022 1160
rect -2886 447 -2106 481
rect -1030 433 -1020 497
rect -956 433 -946 497
rect -364 481 -300 1576
rect 3592 1462 3602 1526
rect 3666 1462 6152 1526
rect 6216 1462 6226 1526
rect 160 1277 170 1341
rect 234 1277 4326 1341
rect 4390 1277 4400 1341
rect 6932 982 6978 1160
rect -729 447 -300 481
rect -364 446 -300 447
rect 6690 429 6700 493
rect 6764 481 6774 493
rect 8724 481 8799 2247
rect 6764 447 6895 481
rect 8277 447 8799 481
rect 6764 429 6774 447
rect -2068 -40 -2022 132
rect 6932 -40 6978 132
rect -2068 -818 -2022 -640
rect 6932 -818 6978 -640
rect -3494 -1353 -2106 -1319
rect -1029 -1368 -1019 -1304
rect -955 -1368 -945 -1304
rect -512 -1319 -502 -1301
rect -720 -1353 -502 -1319
rect -512 -1365 -502 -1353
rect -438 -1365 -428 -1301
rect 6708 -1363 6718 -1299
rect 6782 -1319 6792 -1299
rect 9235 -1319 9310 7647
rect 6782 -1353 6894 -1319
rect 8271 -1353 9310 -1319
rect 6782 -1363 6792 -1353
rect -2068 -1840 -2022 -1668
rect 6932 -1840 6978 -1668
<< via1 >>
rect -1022 7631 -958 7695
rect 6691 7633 6755 7697
rect 1628 6412 1692 6476
rect -1028 5831 -964 5895
rect -477 5829 -413 5893
rect -1024 4031 -960 4095
rect -434 4030 -370 4094
rect 6704 5831 6768 5895
rect 3157 5494 3221 5558
rect 3157 5020 3221 5084
rect 3768 4864 3832 4928
rect 6166 4868 6230 4932
rect 3106 4499 3170 4563
rect 5207 4326 5271 4390
rect 3308 4148 3372 4212
rect 333 3419 397 3483
rect 1631 3419 1695 3483
rect 333 3090 397 3154
rect -1027 2231 -963 2295
rect -434 2227 -370 2291
rect 6759 4031 6823 4095
rect 4874 3578 4938 3642
rect 6764 2233 6828 2297
rect 3308 2159 3372 2223
rect 2330 1576 2394 1640
rect -1020 433 -956 497
rect 3602 1462 3666 1526
rect 6152 1462 6216 1526
rect 170 1277 234 1341
rect 4326 1277 4390 1341
rect 6700 429 6764 493
rect -1019 -1368 -955 -1304
rect -502 -1365 -438 -1301
rect 6718 -1363 6782 -1299
<< metal2 >>
rect -2651 8198 -2587 8208
rect 8848 8198 8912 8208
rect -2587 8134 -1907 8186
rect 8303 8134 8848 8186
rect -2651 8124 -2587 8134
rect 8848 8124 8912 8134
rect -1022 7855 2060 7919
rect -1022 7695 -958 7855
rect -1022 7621 -958 7631
rect -2398 7390 -2334 7400
rect -2334 7326 -1922 7378
rect -2398 7316 -2334 7326
rect 1996 6756 2060 7855
rect 6691 7697 6755 7707
rect 6691 7623 6755 7633
rect 8595 7391 8659 7401
rect 8279 7327 8595 7379
rect 8595 7317 8659 7327
rect 1996 6682 2060 6692
rect 1628 6476 1692 6486
rect -2651 6398 -2587 6408
rect 1628 6402 1692 6412
rect 8848 6398 8912 6408
rect -2587 6334 -1907 6386
rect 8280 6334 8848 6386
rect -2651 6324 -2587 6334
rect 8848 6324 8912 6334
rect -1028 5895 -964 5905
rect -1028 5726 -964 5831
rect -477 5893 -413 5903
rect -477 5819 -413 5829
rect 6704 5895 6768 5905
rect 6704 5821 6768 5831
rect 3410 5781 3474 5791
rect -1028 5662 -133 5726
rect -2398 5590 -2334 5600
rect -2334 5526 -1906 5578
rect -2398 5516 -2334 5526
rect -197 5170 -133 5662
rect -197 5096 -133 5106
rect 1282 5612 1346 5622
rect -2651 4598 -2587 4608
rect -2587 4534 -1915 4586
rect -2651 4524 -2587 4534
rect 1282 4219 1346 5548
rect 1630 5613 1694 5623
rect 1428 4219 1492 4229
rect -434 4155 1428 4219
rect -1024 4095 -960 4105
rect -1024 3923 -960 4031
rect -434 4094 -370 4155
rect 1428 4145 1492 4155
rect -434 4020 -370 4030
rect -1024 3859 -369 3923
rect -2398 3790 -2334 3800
rect -2334 3726 -1918 3778
rect -2398 3716 -2334 3726
rect -433 3327 -369 3859
rect 1630 3843 1694 5549
rect 3157 5558 3221 5568
rect 3157 5484 3221 5494
rect 3410 5169 3474 5717
rect 8595 5591 8659 5601
rect 8280 5527 8595 5579
rect 8595 5517 8659 5527
rect 3410 5095 3474 5105
rect 4658 5106 4722 5116
rect 5418 5106 5482 5116
rect 3157 5084 3221 5094
rect 4722 5042 5418 5106
rect 4658 5032 4722 5042
rect 5418 5032 5482 5042
rect 3157 5010 3221 5020
rect 3768 4928 3832 4938
rect 3768 4854 3832 4864
rect 4084 4928 4148 4938
rect 5706 4928 5770 4938
rect 4148 4864 5706 4928
rect 4084 4854 4148 4864
rect 5706 4854 5770 4864
rect 6166 4932 6230 4942
rect 6166 4858 6230 4868
rect 8848 4598 8912 4608
rect 3106 4563 3170 4573
rect 8279 4534 8848 4586
rect 8848 4524 8912 4534
rect 3106 4489 3170 4499
rect 5207 4390 5271 4400
rect 5207 4316 5271 4326
rect 3308 4212 3372 4222
rect 3308 4138 3372 4148
rect 6759 4095 6823 4105
rect 5952 4031 6759 4095
rect 4876 3980 4940 3990
rect 5206 3980 5270 3990
rect 4940 3916 5206 3980
rect 4876 3906 4940 3916
rect 5206 3906 5270 3916
rect 3306 3862 3370 3872
rect 1630 3779 1866 3843
rect 333 3483 397 3493
rect 333 3409 397 3419
rect 765 3483 829 3493
rect 1408 3483 1472 3493
rect 829 3419 1408 3483
rect 765 3409 829 3419
rect 1408 3409 1472 3419
rect 1631 3483 1695 3493
rect 1631 3409 1695 3419
rect 333 3327 397 3337
rect -433 3307 333 3327
rect -434 3263 333 3307
rect 397 3263 402 3327
rect -2651 2798 -2587 2808
rect -2587 2734 -1936 2786
rect -2651 2724 -2587 2734
rect -434 2536 -370 3263
rect 333 3253 397 3263
rect 333 3154 397 3164
rect 333 3080 397 3090
rect 764 3153 828 3163
rect 1802 3153 1866 3779
rect 828 3089 1866 3153
rect 764 3079 828 3089
rect 3306 2623 3370 3798
rect 4874 3642 4938 3652
rect 4874 3568 4938 3578
rect 4510 3462 4574 3472
rect 5952 3462 6016 4031
rect 6759 4021 6823 4031
rect 8595 3791 8659 3801
rect 8291 3727 8595 3779
rect 8595 3717 8659 3727
rect 4574 3398 6016 3462
rect 4510 3388 4574 3398
rect 4508 3151 4572 3161
rect 4572 3087 6011 3151
rect 4508 3077 4572 3087
rect 3306 2549 3370 2559
rect -1027 2472 -370 2536
rect -1027 2295 -963 2472
rect -1027 2221 -963 2231
rect -434 2291 -370 2301
rect 5947 2297 6011 3087
rect 8848 2798 8912 2808
rect 8277 2734 8848 2786
rect 8848 2724 8912 2734
rect 6764 2297 6828 2307
rect 5947 2233 6764 2297
rect -2398 1990 -2334 2000
rect -2334 1926 -1921 1978
rect -2398 1916 -2334 1926
rect -434 1674 -370 2227
rect 3308 2223 3372 2233
rect 6764 2223 6828 2233
rect 3308 2149 3372 2159
rect 8595 1991 8659 2001
rect 8292 1927 8595 1979
rect 8595 1917 8659 1927
rect 4437 1704 4501 1714
rect 5426 1704 5490 1714
rect 540 1674 604 1684
rect 1830 1674 1894 1684
rect -434 1610 540 1674
rect 604 1610 1830 1674
rect 540 1600 604 1610
rect 1830 1600 1894 1610
rect 2330 1640 2394 1650
rect 4501 1640 5426 1704
rect 4437 1630 4501 1640
rect 5426 1630 5490 1640
rect 2330 1566 2394 1576
rect 3602 1526 3666 1536
rect 3602 1452 3666 1462
rect 3894 1522 3958 1532
rect 5736 1522 5800 1532
rect 3958 1458 5736 1522
rect 3894 1448 3958 1458
rect 5736 1448 5800 1458
rect 6152 1526 6216 1536
rect 6152 1452 6216 1462
rect 170 1341 234 1351
rect 170 1267 234 1277
rect 930 1341 994 1351
rect 3943 1341 4007 1351
rect 994 1277 3943 1341
rect 930 1267 994 1277
rect 3943 1267 4007 1277
rect 4326 1341 4390 1351
rect 4326 1267 4390 1277
rect -2651 998 -2587 1008
rect 8848 998 8912 1008
rect -2587 934 -1916 986
rect 8292 934 8848 986
rect -2651 924 -2587 934
rect 8848 924 8912 934
rect -1020 497 -956 507
rect -1020 348 -956 433
rect 6700 493 6764 503
rect 6700 419 6764 429
rect 1423 349 1487 359
rect -1020 285 1423 348
rect -1020 284 1487 285
rect 1423 275 1487 284
rect -2398 190 -2334 200
rect 8595 191 8659 201
rect -2334 126 -1925 178
rect 8279 127 8595 179
rect -2398 116 -2334 126
rect 8595 117 8659 127
rect 160 -218 224 -208
rect -2651 -802 -2587 -792
rect -2587 -866 -1906 -814
rect -2651 -876 -2587 -866
rect -364 -1074 -300 -1064
rect -1019 -1138 -364 -1074
rect -1019 -1304 -955 -1138
rect -364 -1148 -300 -1138
rect -1019 -1378 -955 -1368
rect -502 -1301 -438 -1291
rect 160 -1301 224 -282
rect 8848 -802 8912 -792
rect 8279 -866 8848 -814
rect 8848 -876 8912 -866
rect -438 -1365 224 -1301
rect 6718 -1299 6782 -1289
rect -502 -1375 -438 -1365
rect 6718 -1373 6782 -1363
rect -2398 -1610 -2334 -1600
rect 8595 -1609 8659 -1599
rect -2334 -1674 -1913 -1622
rect 8300 -1673 8595 -1621
rect -2398 -1684 -2334 -1674
rect 8595 -1683 8659 -1673
<< via2 >>
rect -2651 8134 -2587 8198
rect 8848 8134 8912 8198
rect -2398 7326 -2334 7390
rect 6691 7633 6755 7697
rect 8595 7327 8659 7391
rect 1996 6692 2060 6756
rect 1628 6412 1692 6476
rect -2651 6334 -2587 6398
rect 8848 6334 8912 6398
rect -477 5829 -413 5893
rect 6704 5831 6768 5895
rect -2398 5526 -2334 5590
rect 3410 5717 3474 5781
rect -197 5106 -133 5170
rect 1282 5548 1346 5612
rect -2651 4534 -2587 4598
rect 1630 5549 1694 5613
rect 1428 4155 1492 4219
rect -2398 3726 -2334 3790
rect 3157 5494 3221 5558
rect 8595 5527 8659 5591
rect 3410 5105 3474 5169
rect 3157 5020 3221 5084
rect 4658 5042 4722 5106
rect 5418 5042 5482 5106
rect 3768 4864 3832 4928
rect 4084 4864 4148 4928
rect 5706 4864 5770 4928
rect 6166 4868 6230 4932
rect 3106 4499 3170 4563
rect 8848 4534 8912 4598
rect 5207 4326 5271 4390
rect 3308 4148 3372 4212
rect 4876 3916 4940 3980
rect 5206 3916 5270 3980
rect 333 3419 397 3483
rect 765 3419 829 3483
rect 1408 3419 1472 3483
rect 1631 3419 1695 3483
rect 333 3263 397 3327
rect -2651 2734 -2587 2798
rect 333 3090 397 3154
rect 764 3089 828 3153
rect 3306 3798 3370 3862
rect 4874 3578 4938 3642
rect 8595 3727 8659 3791
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3306 2559 3370 2623
rect 8848 2734 8912 2798
rect -2398 1926 -2334 1990
rect 3308 2159 3372 2223
rect 8595 1927 8659 1991
rect 540 1610 604 1674
rect 1830 1610 1894 1674
rect 2330 1576 2394 1640
rect 4437 1640 4501 1704
rect 5426 1640 5490 1704
rect 3602 1462 3666 1526
rect 3894 1458 3958 1522
rect 5736 1458 5800 1522
rect 6152 1462 6216 1526
rect 170 1277 234 1341
rect 930 1277 994 1341
rect 3943 1277 4007 1341
rect 4326 1277 4390 1341
rect -2651 934 -2587 998
rect 8848 934 8912 998
rect 6700 429 6764 493
rect 1423 285 1487 349
rect -2398 126 -2334 190
rect 8595 127 8659 191
rect 160 -282 224 -218
rect -2651 -866 -2587 -802
rect -364 -1138 -300 -1074
rect 8848 -866 8912 -802
rect 6718 -1363 6782 -1299
rect -2398 -1674 -2334 -1610
rect 8595 -1673 8659 -1609
<< metal3 >>
rect -2651 8203 -2587 8208
rect 8848 8203 8912 8208
rect -2661 8198 -2577 8203
rect -2661 8134 -2651 8198
rect -2587 8134 -2577 8198
rect -2661 8129 -2577 8134
rect 8838 8198 8922 8203
rect 8838 8134 8848 8198
rect 8912 8134 8922 8198
rect 8838 8129 8922 8134
rect -2651 6403 -2587 8129
rect 6681 7697 6765 7702
rect 6681 7633 6691 7697
rect 6755 7633 6765 7697
rect 6681 7628 6765 7633
rect -2398 7395 -2334 7400
rect -2408 7390 -2324 7395
rect -2408 7326 -2398 7390
rect -2334 7326 -2324 7390
rect -2408 7321 -2324 7326
rect -2661 6398 -2577 6403
rect -2661 6334 -2651 6398
rect -2587 6334 -2577 6398
rect -2661 6329 -2577 6334
rect -2651 4603 -2587 6329
rect -2398 5595 -2334 7321
rect 1975 6756 2080 6780
rect 6691 6779 6755 7628
rect 8595 7396 8659 7401
rect 8585 7391 8669 7396
rect 8585 7327 8595 7391
rect 8659 7327 8669 7391
rect 8585 7322 8669 7327
rect 1975 6692 1996 6756
rect 2060 6692 2080 6756
rect 1975 6669 2080 6692
rect 6191 6715 6755 6779
rect 6191 6515 6255 6715
rect 1618 6476 1702 6481
rect 1618 6412 1628 6476
rect 1692 6412 1896 6476
rect 1618 6407 1702 6412
rect 3157 6133 3698 6197
rect -497 5893 -391 5915
rect -497 5829 -477 5893
rect -413 5829 -391 5893
rect -497 5808 -391 5829
rect 1272 5612 1356 5617
rect -2408 5590 -2324 5595
rect -2408 5526 -2398 5590
rect -2334 5526 -2324 5590
rect -2408 5521 -2324 5526
rect -2661 4598 -2577 4603
rect -2661 4534 -2651 4598
rect -2587 4534 -2577 4598
rect -2661 4529 -2577 4534
rect -2651 4524 -2587 4529
rect -2398 3795 -2334 5521
rect 544 5311 608 5551
rect 1110 5548 1282 5612
rect 1346 5548 1356 5612
rect 1272 5543 1356 5548
rect 1616 5613 1708 5646
rect 1616 5549 1630 5613
rect 1694 5549 1708 5613
rect 3157 5563 3221 6133
rect 6686 5895 6784 5914
rect 6686 5831 6704 5895
rect 6768 5831 6784 5895
rect 6686 5814 6784 5831
rect 3400 5781 3484 5810
rect 3400 5717 3410 5781
rect 3474 5717 3484 5781
rect 3400 5693 3484 5717
rect 8595 5596 8659 7322
rect 8848 6403 8912 8129
rect 8838 6398 8922 6403
rect 8838 6334 8848 6398
rect 8912 6334 8922 6398
rect 8838 6329 8922 6334
rect 8585 5591 8669 5596
rect 1616 5524 1708 5549
rect 3147 5558 3231 5563
rect 3147 5494 3157 5558
rect 3221 5494 3231 5558
rect 8585 5527 8595 5591
rect 8659 5527 8669 5591
rect 8585 5522 8669 5527
rect 3147 5489 3231 5494
rect 544 5247 5105 5311
rect -238 5170 -98 5201
rect -238 5106 -197 5170
rect -133 5106 -98 5170
rect -238 5072 -98 5106
rect 3379 5169 3508 5177
rect 3379 5105 3410 5169
rect 3474 5105 3508 5169
rect 3379 5097 3508 5105
rect 4648 5106 4732 5111
rect 3147 5084 3231 5089
rect 754 5020 3157 5084
rect 3221 5020 3231 5084
rect 4648 5042 4658 5106
rect 4722 5042 4732 5106
rect 4648 5037 4732 5042
rect 754 4663 818 5020
rect 3147 5015 3231 5020
rect 3758 4928 3842 4933
rect 1241 4864 3768 4928
rect 3832 4864 3842 4928
rect -2408 3790 -2324 3795
rect -2408 3726 -2398 3790
rect -2334 3726 -2324 3790
rect -2408 3721 -2324 3726
rect 333 3488 397 3761
rect 323 3483 407 3488
rect 323 3419 333 3483
rect 397 3419 407 3483
rect 323 3414 407 3419
rect 743 3483 849 3501
rect 743 3419 765 3483
rect 829 3419 849 3483
rect 333 3332 397 3414
rect 743 3404 849 3419
rect 323 3327 407 3332
rect 323 3263 333 3327
rect 397 3263 407 3327
rect 323 3258 407 3263
rect 333 3159 397 3258
rect 323 3154 407 3159
rect 323 3090 333 3154
rect 397 3090 407 3154
rect 323 3085 407 3090
rect 745 3158 837 3183
rect 745 3153 838 3158
rect 745 3089 764 3153
rect 828 3089 838 3153
rect 333 2812 397 3085
rect 745 3084 838 3089
rect 745 3061 837 3084
rect -2651 2803 -2587 2808
rect -2661 2798 -2577 2803
rect -2661 2734 -2651 2798
rect -2587 2734 -2577 2798
rect -2661 2729 -2577 2734
rect -2651 1003 -2587 2729
rect -2398 1995 -2334 2000
rect -2408 1990 -2324 1995
rect -2408 1926 -2398 1990
rect -2334 1926 -2324 1990
rect -2408 1921 -2324 1926
rect -2661 998 -2577 1003
rect -2661 934 -2651 998
rect -2587 934 -2577 998
rect -2661 929 -2577 934
rect -2651 -797 -2587 929
rect -2398 195 -2334 1921
rect 170 1346 234 1946
rect 530 1674 614 1679
rect 530 1610 540 1674
rect 604 1610 614 1674
rect 530 1605 614 1610
rect 160 1341 244 1346
rect 160 1277 170 1341
rect 234 1277 244 1341
rect 160 1272 244 1277
rect 540 1112 604 1605
rect 910 1341 1011 1357
rect 910 1277 930 1341
rect 994 1277 1011 1341
rect 910 1259 1011 1277
rect 1241 354 1305 4864
rect 3758 4859 3842 4864
rect 4061 4928 4171 4944
rect 4061 4864 4084 4928
rect 4148 4864 4171 4928
rect 4061 4850 4171 4864
rect 4658 4712 4722 5037
rect 3081 4563 3190 4586
rect 3081 4499 3106 4563
rect 3170 4499 3190 4563
rect 3081 4479 3190 4499
rect 1418 4219 1502 4224
rect 1418 4155 1428 4219
rect 1492 4155 1842 4219
rect 3298 4212 3382 4217
rect 1418 4150 1502 4155
rect 3298 4148 3308 4212
rect 3372 4148 3698 4212
rect 3298 4143 3382 4148
rect 4862 3980 4953 4019
rect 4862 3916 4876 3980
rect 4940 3916 4953 3980
rect 3283 3862 3389 3885
rect 4862 3879 4953 3916
rect 3283 3798 3306 3862
rect 3370 3798 3389 3862
rect 3283 3778 3389 3798
rect 1397 3483 1484 3517
rect 1397 3419 1408 3483
rect 1472 3419 1484 3483
rect 1397 3388 1484 3419
rect 1621 3483 1705 3488
rect 1621 3419 1631 3483
rect 1695 3419 1705 3483
rect 1621 3414 1705 3419
rect 2348 3432 2412 3740
rect 4864 3642 4948 3647
rect 4864 3578 4874 3642
rect 4938 3578 4948 3642
rect 4864 3573 4948 3578
rect 4479 3462 4604 3492
rect 999 290 1305 354
rect 1405 349 1503 380
rect 1405 285 1423 349
rect 1487 285 1503 349
rect 1631 365 1695 3414
rect 2348 3368 3912 3432
rect 4479 3398 4510 3462
rect 4574 3398 4604 3462
rect 4479 3371 4604 3398
rect 3848 2819 3912 3368
rect 4486 3151 4590 3171
rect 4486 3087 4508 3151
rect 4572 3087 4590 3151
rect 4486 3071 4590 3087
rect 3284 2623 3390 2645
rect 3284 2559 3306 2623
rect 3370 2559 3390 2623
rect 3284 2538 3390 2559
rect 3298 2223 3382 2228
rect 2887 2159 3308 2223
rect 3372 2159 3382 2223
rect 3298 2154 3382 2159
rect 1830 1679 1894 1868
rect 4437 1709 4501 1893
rect 4427 1704 4511 1709
rect 1820 1674 1904 1679
rect 1820 1610 1830 1674
rect 1894 1610 1904 1674
rect 1820 1605 1904 1610
rect 2307 1640 2415 1666
rect 2307 1576 2330 1640
rect 2394 1576 2415 1640
rect 4427 1640 4437 1704
rect 4501 1640 4511 1704
rect 4427 1635 4511 1640
rect 2307 1553 2415 1576
rect 3592 1526 3676 1531
rect 3083 1462 3602 1526
rect 3666 1462 3676 1526
rect 1631 301 1897 365
rect 3083 363 3147 1462
rect 3592 1457 3676 1462
rect 3873 1522 3978 1546
rect 3873 1458 3894 1522
rect 3958 1458 3978 1522
rect 3873 1437 3978 1458
rect 3923 1341 4024 1360
rect 3923 1277 3943 1341
rect 4007 1277 4024 1341
rect 3923 1262 4024 1277
rect 4316 1341 4400 1346
rect 4316 1277 4326 1341
rect 4390 1277 4400 1341
rect 4316 1272 4400 1277
rect 4326 1060 4390 1272
rect 4874 448 4938 3573
rect 5041 616 5105 5247
rect 5418 5111 5482 5460
rect 5408 5106 5492 5111
rect 5408 5042 5418 5106
rect 5482 5042 5492 5106
rect 5408 5037 5492 5042
rect 5683 4928 5793 4943
rect 6166 4937 6230 5491
rect 5683 4864 5706 4928
rect 5770 4864 5793 4928
rect 5683 4849 5793 4864
rect 6156 4932 6240 4937
rect 6156 4868 6166 4932
rect 6230 4868 6240 4932
rect 6156 4863 6240 4868
rect 5197 4390 5281 4395
rect 5197 4326 5207 4390
rect 5271 4326 5495 4390
rect 5197 4321 5281 4326
rect 5193 3980 5284 4018
rect 5193 3916 5206 3980
rect 5270 3916 5284 3980
rect 5193 3878 5284 3916
rect 8595 3796 8659 5522
rect 8848 4603 8912 6329
rect 8838 4598 8922 4603
rect 8838 4534 8848 4598
rect 8912 4534 8922 4598
rect 8838 4529 8922 4534
rect 8585 3791 8669 3796
rect 8585 3727 8595 3791
rect 8659 3727 8669 3791
rect 8585 3722 8669 3727
rect 8595 3717 8659 3722
rect 8848 2803 8912 2808
rect 8838 2798 8922 2803
rect 8838 2734 8848 2798
rect 8912 2734 8922 2798
rect 8838 2729 8922 2734
rect 8595 1996 8659 2001
rect 8585 1991 8669 1996
rect 8585 1927 8595 1991
rect 8659 1927 8669 1991
rect 8585 1922 8669 1927
rect 5416 1704 5500 1709
rect 5416 1640 5426 1704
rect 5490 1640 5500 1704
rect 5416 1635 5500 1640
rect 5426 1079 5490 1635
rect 5715 1522 5820 1544
rect 6152 1531 6216 1903
rect 5715 1458 5736 1522
rect 5800 1458 5820 1522
rect 5715 1435 5820 1458
rect 6142 1526 6226 1531
rect 6142 1462 6152 1526
rect 6216 1462 6226 1526
rect 6142 1457 6226 1462
rect 5041 552 5566 616
rect 6683 493 6785 514
rect 4610 384 4941 448
rect 6683 429 6700 493
rect 6764 429 6785 493
rect 6683 411 6785 429
rect 2812 299 3147 363
rect 1405 260 1503 285
rect 8595 196 8659 1922
rect 8848 1003 8912 2729
rect 8838 998 8922 1003
rect 8838 934 8848 998
rect 8912 934 8922 998
rect 8838 929 8922 934
rect -2408 190 -2324 195
rect -2408 126 -2398 190
rect -2334 126 -2324 190
rect -2408 121 -2324 126
rect 8585 191 8669 196
rect 8585 127 8595 191
rect 8659 127 8669 191
rect 8585 122 8669 127
rect -2661 -802 -2577 -797
rect -2661 -866 -2651 -802
rect -2587 -866 -2577 -802
rect -2661 -871 -2577 -866
rect -2651 -876 -2587 -871
rect -2398 -1605 -2334 121
rect 139 -218 245 -195
rect 139 -282 160 -218
rect 224 -282 245 -218
rect 139 -299 245 -282
rect 6179 -442 6243 116
rect 6179 -506 6782 -442
rect -378 -1074 -280 -1056
rect -378 -1138 -364 -1074
rect -300 -1138 -280 -1074
rect -378 -1159 -280 -1138
rect 6718 -1294 6782 -506
rect 6708 -1299 6792 -1294
rect 6708 -1363 6718 -1299
rect 6782 -1363 6792 -1299
rect 6708 -1368 6792 -1363
rect 6718 -1372 6782 -1368
rect 8595 -1604 8659 122
rect 8848 -797 8912 929
rect 8838 -802 8922 -797
rect 8838 -866 8848 -802
rect 8912 -866 8922 -802
rect 8838 -871 8922 -866
rect -2408 -1610 -2324 -1605
rect -2408 -1674 -2398 -1610
rect -2334 -1674 -2324 -1610
rect -2408 -1679 -2324 -1674
rect 8585 -1609 8669 -1604
rect 8585 -1673 8595 -1609
rect 8659 -1673 8669 -1609
rect 8585 -1678 8669 -1673
rect -2398 -1684 -2334 -1679
rect 8595 -1683 8659 -1678
<< via3 >>
rect 1996 6692 2060 6756
rect -477 5829 -413 5893
rect 1630 5549 1694 5613
rect 6704 5831 6768 5895
rect 3410 5717 3474 5781
rect -197 5106 -133 5170
rect 3410 5105 3474 5169
rect 765 3419 829 3483
rect 764 3089 828 3153
rect 930 1277 994 1341
rect 4084 4864 4148 4928
rect 3106 4499 3170 4563
rect 4876 3916 4940 3980
rect 3306 3798 3370 3862
rect 1408 3419 1472 3483
rect 1423 285 1487 349
rect 4510 3398 4574 3462
rect 4508 3087 4572 3151
rect 3306 2559 3370 2623
rect 2330 1576 2394 1640
rect 3894 1458 3958 1522
rect 3943 1277 4007 1341
rect 5706 4864 5770 4928
rect 5206 3916 5270 3980
rect 5736 1458 5800 1522
rect 6700 429 6764 493
rect 160 -282 224 -218
rect -364 -1138 -300 -1074
<< metal4 >>
rect 1995 6756 2061 6757
rect 1995 6692 1996 6756
rect 2060 6692 2061 6756
rect 1995 6691 2061 6692
rect 1996 6377 2060 6691
rect 6703 5895 6769 5896
rect -478 5893 -412 5894
rect -478 5829 -477 5893
rect -413 5829 155 5893
rect 6322 5831 6704 5895
rect 6768 5831 6769 5895
rect 6703 5830 6769 5831
rect -478 5828 -412 5829
rect 3409 5781 3475 5782
rect 3409 5717 3410 5781
rect 3474 5717 3744 5781
rect 3409 5716 3475 5717
rect 1629 5613 1695 5614
rect 544 5311 608 5551
rect 1629 5549 1630 5613
rect 1694 5549 1949 5613
rect 1629 5548 1695 5549
rect 544 5247 5105 5311
rect -198 5170 -132 5171
rect -198 5106 -197 5170
rect -133 5169 -132 5170
rect 3409 5169 3475 5170
rect -133 5106 3410 5169
rect -198 5105 3410 5106
rect 3474 5105 3475 5169
rect 320 4612 384 5105
rect 3409 5104 3475 5105
rect 4083 4928 4149 4929
rect 1242 4864 4084 4928
rect 4148 4864 4150 4928
rect 765 3484 829 3761
rect 764 3483 830 3484
rect 764 3419 765 3483
rect 829 3419 830 3483
rect 764 3418 830 3419
rect 763 3153 829 3154
rect 763 3089 764 3153
rect 828 3089 829 3153
rect 763 3088 829 3089
rect 764 2811 828 3088
rect -364 1985 213 2049
rect -364 -1073 -300 1985
rect 930 1342 994 1946
rect 929 1341 995 1342
rect 929 1277 930 1341
rect 994 1277 995 1341
rect 929 1276 995 1277
rect 1242 859 1306 4864
rect 4083 4863 4149 4864
rect 3105 4563 3171 4564
rect 2808 4499 3106 4563
rect 3170 4499 3171 4563
rect 3105 4498 3171 4499
rect 4875 3980 4941 3981
rect 4875 3916 4876 3980
rect 4940 3916 4941 3980
rect 4875 3915 4941 3916
rect 3305 3862 3371 3863
rect 3305 3798 3306 3862
rect 3370 3798 3746 3862
rect 3305 3797 3371 3798
rect 1407 3483 1473 3484
rect 1407 3419 1408 3483
rect 1472 3419 1473 3483
rect 1407 3418 1473 3419
rect 2348 3432 2412 3740
rect 4510 3463 4574 3790
rect 4509 3462 4575 3463
rect 998 795 1306 859
rect 1408 813 1472 3418
rect 2348 3368 3912 3432
rect 4509 3398 4510 3462
rect 4574 3398 4575 3462
rect 4509 3397 4575 3398
rect 3848 2820 3912 3368
rect 4507 3151 4573 3152
rect 4507 3087 4508 3151
rect 4572 3087 4573 3151
rect 4507 3086 4573 3087
rect 4508 2788 4572 3086
rect 3305 2623 3371 2624
rect 2816 2559 3306 2623
rect 3370 2559 3371 2623
rect 3305 2558 3371 2559
rect 2330 1641 2394 1961
rect 2329 1640 2395 1641
rect 2329 1576 2330 1640
rect 2394 1576 2395 1640
rect 2329 1575 2395 1576
rect 3893 1522 3959 1523
rect 3083 1458 3894 1522
rect 3958 1458 3959 1522
rect 1408 749 1954 813
rect 3083 812 3147 1458
rect 3893 1457 3959 1458
rect 3943 1342 4007 1345
rect 3942 1341 4008 1342
rect 3942 1277 3943 1341
rect 4007 1277 4008 1341
rect 3942 1276 4008 1277
rect 3943 1007 4007 1276
rect 4876 844 4940 3915
rect 2812 748 3147 812
rect 4609 780 4940 844
rect 5041 616 5105 5247
rect 5706 4929 5770 5552
rect 5705 4928 5771 4929
rect 5705 4864 5706 4928
rect 5770 4864 5771 4928
rect 5705 4863 5771 4864
rect 5205 3980 5271 3981
rect 5205 3916 5206 3980
rect 5270 3916 5546 3980
rect 5205 3915 5271 3916
rect 5736 1523 5800 1953
rect 5735 1522 5801 1523
rect 5735 1458 5736 1522
rect 5800 1458 5801 1522
rect 5735 1457 5801 1458
rect 5041 552 5566 616
rect 6699 493 6765 494
rect 6384 429 6700 493
rect 6764 429 6766 493
rect 6699 428 6765 429
rect 1422 349 1488 350
rect 1420 285 1423 349
rect 1487 285 1953 349
rect 1422 284 1488 285
rect 160 -217 224 179
rect 159 -218 225 -217
rect 159 -282 160 -218
rect 224 -282 225 -218
rect 159 -283 225 -282
rect -365 -1074 -299 -1073
rect -365 -1138 -364 -1074
rect -300 -1138 -299 -1074
rect -365 -1139 -299 -1138
use transmission_gate  transmission_gate_0 ~/ee372/incremental_delta_sigma_adc/design/analog_modulator/layout/transmission_gate
timestamp 1653911004
transform -1 0 8143 0 1 51
box -216 -51 1283 1063
use transmission_gate  transmission_gate_1
timestamp 1653911004
transform -1 0 8143 0 1 1851
box -216 -51 1283 1063
use transmission_gate  transmission_gate_2
timestamp 1653911004
transform -1 0 8143 0 1 -1749
box -216 -51 1283 1063
use transmission_gate  transmission_gate_3
timestamp 1653911004
transform -1 0 8143 0 1 3651
box -216 -51 1283 1063
use transmission_gate  transmission_gate_4
timestamp 1653911004
transform -1 0 8143 0 1 5451
box -216 -51 1283 1063
use transmission_gate  transmission_gate_5
timestamp 1653911004
transform -1 0 8143 0 1 7251
box -216 -51 1283 1063
use transmission_gate  transmission_gate_6
timestamp 1653911004
transform -1 0 -857 0 1 7251
box -216 -51 1283 1063
use transmission_gate  transmission_gate_7
timestamp 1653911004
transform -1 0 -857 0 1 5451
box -216 -51 1283 1063
use transmission_gate  transmission_gate_8
timestamp 1653911004
transform -1 0 -857 0 1 3651
box -216 -51 1283 1063
use transmission_gate  transmission_gate_9
timestamp 1653911004
transform -1 0 -857 0 1 1851
box -216 -51 1283 1063
use transmission_gate  transmission_gate_10
timestamp 1653911004
transform -1 0 -857 0 1 51
box -216 -51 1283 1063
use transmission_gate  transmission_gate_11
timestamp 1653911004
transform -1 0 -857 0 1 -1749
box -216 -51 1283 1063
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_0
timestamp 1653911004
transform 1 0 630 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_1
timestamp 1653911004
transform 1 0 2430 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_2
timestamp 1653911004
transform 1 0 4230 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_3
timestamp 1653911004
transform 1 0 6030 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_4
timestamp 1653911004
transform 1 0 6030 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_5
timestamp 1653911004
transform 1 0 4230 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_6
timestamp 1653911004
transform 1 0 2430 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_7
timestamp 1653911004
transform 1 0 630 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_8
timestamp 1653911004
transform 1 0 6030 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_9
timestamp 1653911004
transform 1 0 4230 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_10
timestamp 1653911004
transform 1 0 2430 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_11
timestamp 1653911004
transform 1 0 630 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_12
timestamp 1653911004
transform 1 0 6030 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_13
timestamp 1653911004
transform 1 0 4230 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_14
timestamp 1653911004
transform 1 0 2430 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_15
timestamp 1653911004
transform 1 0 630 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_16
timestamp 1653911004
transform 1 0 7830 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_17
timestamp 1653911004
transform 1 0 7830 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_18
timestamp 1653911004
transform 1 0 7830 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_19
timestamp 1653911004
transform 1 0 7830 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_20
timestamp 1653911004
transform 1 0 -1170 0 1 5980
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_21
timestamp 1653911004
transform 1 0 -1170 0 1 4180
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_22
timestamp 1653911004
transform 1 0 -1170 0 1 2380
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_23
timestamp 1653911004
transform 1 0 -1170 0 1 580
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_24
timestamp 1653911004
transform 1 0 7830 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_25
timestamp 1653911004
transform 1 0 6030 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_26
timestamp 1653911004
transform 1 0 4230 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_27
timestamp 1653911004
transform 1 0 2430 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_28
timestamp 1653911004
transform 1 0 630 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_29
timestamp 1653911004
transform 1 0 -1170 0 1 7780
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_30
timestamp 1653911004
transform 1 0 -1170 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_31
timestamp 1653911004
transform 1 0 630 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_32
timestamp 1653911004
transform 1 0 2430 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_33
timestamp 1653911004
transform 1 0 4230 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_34
timestamp 1653911004
transform 1 0 6030 0 1 -1220
box -630 -580 528 580
use unit_cap_mim_m3m4  unit_cap_mim_m3m4_35
timestamp 1653911004
transform 1 0 7830 0 1 -1220
box -630 -580 528 580
<< labels >>
flabel metal3 -2642 8019 -2642 8019 1 FreeSans 400 0 0 0 p2_b
flabel metal3 -2389 7236 -2389 7236 1 FreeSans 400 0 0 0 p2
flabel metal3 -2639 2626 -2639 2626 1 FreeSans 400 0 0 0 p1_b
flabel metal3 -2389 1840 -2389 1840 1 FreeSans 400 0 0 0 p1
flabel metal3 8645 -1537 8645 -1537 1 FreeSans 400 0 0 0 p1
flabel metal3 8898 -670 8898 -670 1 FreeSans 400 0 0 0 p1_b
flabel metal3 8648 7246 8648 7246 1 FreeSans 400 0 0 0 p2
flabel metal3 8904 8016 8904 8016 1 FreeSans 400 0 0 0 p2_b
flabel metal1 -3484 3369 -3484 3369 1 FreeSans 400 0 0 0 op
flabel metal1 -2872 3368 -2872 3368 1 FreeSans 400 0 0 0 on
flabel metal1 -2412 3371 -2412 3371 1 FreeSans 400 0 0 0 cmc
flabel metal1 8790 3295 8790 3295 1 FreeSans 400 0 0 0 cm
flabel metal1 9292 3298 9292 3298 1 FreeSans 400 0 0 0 bias_a
flabel metal1 -2046 8350 -2046 8350 1 FreeSans 400 0 0 0 VDD
flabel metal1 -2045 7178 -2045 7178 1 FreeSans 400 0 0 0 VSS
flabel metal1 -2043 6543 -2043 6543 1 FreeSans 400 0 0 0 VDD
flabel metal1 -2045 5370 -2045 5370 1 FreeSans 400 0 0 0 VSS
flabel metal1 -2043 4743 -2043 4743 1 FreeSans 400 0 0 0 VDD
flabel metal1 -2047 3574 -2047 3574 1 FreeSans 400 0 0 0 VSS
flabel metal1 -2047 2942 -2047 2942 1 FreeSans 400 0 0 0 VDD
flabel metal1 -2045 1776 -2045 1776 1 FreeSans 400 0 0 0 VSS
flabel metal1 -2043 1146 -2043 1146 1 FreeSans 400 0 0 0 VDD
flabel metal1 -2047 -27 -2047 -27 1 FreeSans 400 0 0 0 VSS
flabel metal1 -2045 -659 -2045 -659 1 FreeSans 400 0 0 0 VDD
flabel metal1 -2045 -1822 -2045 -1822 1 FreeSans 400 0 0 0 VSS
flabel metal1 6957 -1822 6957 -1822 1 FreeSans 400 0 0 0 VSS
flabel metal1 6954 -659 6954 -659 1 FreeSans 400 0 0 0 VDD
flabel metal1 6957 -26 6957 -26 1 FreeSans 400 0 0 0 VSS
flabel metal1 6952 1141 6952 1141 1 FreeSans 400 0 0 0 VDD
flabel metal1 6952 1776 6952 1776 1 FreeSans 400 0 0 0 VSS
flabel metal1 6954 2944 6954 2944 1 FreeSans 400 0 0 0 VDD
flabel metal1 6954 3579 6954 3579 1 FreeSans 400 0 0 0 VSS
flabel metal1 6957 4740 6957 4740 1 FreeSans 400 0 0 0 VDD
flabel metal1 6954 5375 6954 5375 1 FreeSans 400 0 0 0 VSS
flabel metal1 6952 6547 6952 6547 1 FreeSans 400 0 0 0 VDD
flabel metal1 6954 7180 6954 7180 1 FreeSans 400 0 0 0 VSS
flabel metal1 6954 8345 6954 8345 1 FreeSans 400 0 0 0 VDD
<< end >>
