* NGSPICE file created from sc_cmfb_flat.ext - technology: sky130A


* Top level circuit sc_cmfb_flat

.end

