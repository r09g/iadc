magic
tech sky130A
magscale 1 2
timestamp 1654572275
<< nmos >>
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
<< ndiff >>
rect -1453 128 -1395 140
rect -1453 -128 -1441 128
rect -1407 -128 -1395 128
rect -1453 -140 -1395 -128
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
rect 1395 128 1453 140
rect 1395 -128 1407 128
rect 1441 -128 1453 128
rect 1395 -140 1453 -128
<< ndiffc >>
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
<< poly >>
rect -1373 212 -1297 228
rect -1373 194 -1357 212
rect -1395 178 -1357 194
rect -1313 194 -1297 212
rect -1195 212 -1119 228
rect -1195 194 -1179 212
rect -1313 178 -1275 194
rect -1395 140 -1275 178
rect -1217 178 -1179 194
rect -1135 194 -1119 212
rect -1017 212 -941 228
rect -1017 194 -1001 212
rect -1135 178 -1097 194
rect -1217 140 -1097 178
rect -1039 178 -1001 194
rect -957 194 -941 212
rect -839 212 -763 228
rect -839 194 -823 212
rect -957 178 -919 194
rect -1039 140 -919 178
rect -861 178 -823 194
rect -779 194 -763 212
rect -661 212 -585 228
rect -661 194 -645 212
rect -779 178 -741 194
rect -861 140 -741 178
rect -683 178 -645 194
rect -601 194 -585 212
rect -483 212 -407 228
rect -483 194 -467 212
rect -601 178 -563 194
rect -683 140 -563 178
rect -505 178 -467 194
rect -423 194 -407 212
rect -305 212 -229 228
rect -305 194 -289 212
rect -423 178 -385 194
rect -505 140 -385 178
rect -327 178 -289 194
rect -245 194 -229 212
rect -127 212 -51 228
rect -127 194 -111 212
rect -245 178 -207 194
rect -327 140 -207 178
rect -149 178 -111 194
rect -67 194 -51 212
rect 51 212 127 228
rect 51 194 67 212
rect -67 178 -29 194
rect -149 140 -29 178
rect 29 178 67 194
rect 111 194 127 212
rect 229 212 305 228
rect 229 194 245 212
rect 111 178 149 194
rect 29 140 149 178
rect 207 178 245 194
rect 289 194 305 212
rect 407 212 483 228
rect 407 194 423 212
rect 289 178 327 194
rect 207 140 327 178
rect 385 178 423 194
rect 467 194 483 212
rect 585 212 661 228
rect 585 194 601 212
rect 467 178 505 194
rect 385 140 505 178
rect 563 178 601 194
rect 645 194 661 212
rect 763 212 839 228
rect 763 194 779 212
rect 645 178 683 194
rect 563 140 683 178
rect 741 178 779 194
rect 823 194 839 212
rect 941 212 1017 228
rect 941 194 957 212
rect 823 178 861 194
rect 741 140 861 178
rect 919 178 957 194
rect 1001 194 1017 212
rect 1119 212 1195 228
rect 1119 194 1135 212
rect 1001 178 1039 194
rect 919 140 1039 178
rect 1097 178 1135 194
rect 1179 194 1195 212
rect 1297 212 1373 228
rect 1297 194 1313 212
rect 1179 178 1217 194
rect 1097 140 1217 178
rect 1275 178 1313 194
rect 1357 194 1373 212
rect 1357 178 1395 194
rect 1275 140 1395 178
rect -1395 -178 -1275 -140
rect -1395 -194 -1357 -178
rect -1373 -212 -1357 -194
rect -1313 -194 -1275 -178
rect -1217 -178 -1097 -140
rect -1217 -194 -1179 -178
rect -1313 -212 -1297 -194
rect -1373 -228 -1297 -212
rect -1195 -212 -1179 -194
rect -1135 -194 -1097 -178
rect -1039 -178 -919 -140
rect -1039 -194 -1001 -178
rect -1135 -212 -1119 -194
rect -1195 -228 -1119 -212
rect -1017 -212 -1001 -194
rect -957 -194 -919 -178
rect -861 -178 -741 -140
rect -861 -194 -823 -178
rect -957 -212 -941 -194
rect -1017 -228 -941 -212
rect -839 -212 -823 -194
rect -779 -194 -741 -178
rect -683 -178 -563 -140
rect -683 -194 -645 -178
rect -779 -212 -763 -194
rect -839 -228 -763 -212
rect -661 -212 -645 -194
rect -601 -194 -563 -178
rect -505 -178 -385 -140
rect -505 -194 -467 -178
rect -601 -212 -585 -194
rect -661 -228 -585 -212
rect -483 -212 -467 -194
rect -423 -194 -385 -178
rect -327 -178 -207 -140
rect -327 -194 -289 -178
rect -423 -212 -407 -194
rect -483 -228 -407 -212
rect -305 -212 -289 -194
rect -245 -194 -207 -178
rect -149 -178 -29 -140
rect -149 -194 -111 -178
rect -245 -212 -229 -194
rect -305 -228 -229 -212
rect -127 -212 -111 -194
rect -67 -194 -29 -178
rect 29 -178 149 -140
rect 29 -194 67 -178
rect -67 -212 -51 -194
rect -127 -228 -51 -212
rect 51 -212 67 -194
rect 111 -194 149 -178
rect 207 -178 327 -140
rect 207 -194 245 -178
rect 111 -212 127 -194
rect 51 -228 127 -212
rect 229 -212 245 -194
rect 289 -194 327 -178
rect 385 -178 505 -140
rect 385 -194 423 -178
rect 289 -212 305 -194
rect 229 -228 305 -212
rect 407 -212 423 -194
rect 467 -194 505 -178
rect 563 -178 683 -140
rect 563 -194 601 -178
rect 467 -212 483 -194
rect 407 -228 483 -212
rect 585 -212 601 -194
rect 645 -194 683 -178
rect 741 -178 861 -140
rect 741 -194 779 -178
rect 645 -212 661 -194
rect 585 -228 661 -212
rect 763 -212 779 -194
rect 823 -194 861 -178
rect 919 -178 1039 -140
rect 919 -194 957 -178
rect 823 -212 839 -194
rect 763 -228 839 -212
rect 941 -212 957 -194
rect 1001 -194 1039 -178
rect 1097 -178 1217 -140
rect 1097 -194 1135 -178
rect 1001 -212 1017 -194
rect 941 -228 1017 -212
rect 1119 -212 1135 -194
rect 1179 -194 1217 -178
rect 1275 -178 1395 -140
rect 1275 -194 1313 -178
rect 1179 -212 1195 -194
rect 1119 -228 1195 -212
rect 1297 -212 1313 -194
rect 1357 -194 1395 -178
rect 1357 -212 1373 -194
rect 1297 -228 1373 -212
<< polycont >>
rect -1357 178 -1313 212
rect -1179 178 -1135 212
rect -1001 178 -957 212
rect -823 178 -779 212
rect -645 178 -601 212
rect -467 178 -423 212
rect -289 178 -245 212
rect -111 178 -67 212
rect 67 178 111 212
rect 245 178 289 212
rect 423 178 467 212
rect 601 178 645 212
rect 779 178 823 212
rect 957 178 1001 212
rect 1135 178 1179 212
rect 1313 178 1357 212
rect -1357 -212 -1313 -178
rect -1179 -212 -1135 -178
rect -1001 -212 -957 -178
rect -823 -212 -779 -178
rect -645 -212 -601 -178
rect -467 -212 -423 -178
rect -289 -212 -245 -178
rect -111 -212 -67 -178
rect 67 -212 111 -178
rect 245 -212 289 -178
rect 423 -212 467 -178
rect 601 -212 645 -178
rect 779 -212 823 -178
rect 957 -212 1001 -178
rect 1135 -212 1179 -178
rect 1313 -212 1357 -178
<< locali >>
rect -1373 178 -1357 212
rect -1313 178 -1297 212
rect -1195 178 -1179 212
rect -1135 178 -1119 212
rect -1017 178 -1001 212
rect -957 178 -941 212
rect -839 178 -823 212
rect -779 178 -763 212
rect -661 178 -645 212
rect -601 178 -585 212
rect -483 178 -467 212
rect -423 178 -407 212
rect -305 178 -289 212
rect -245 178 -229 212
rect -127 178 -111 212
rect -67 178 -51 212
rect 51 178 67 212
rect 111 178 127 212
rect 229 178 245 212
rect 289 178 305 212
rect 407 178 423 212
rect 467 178 483 212
rect 585 178 601 212
rect 645 178 661 212
rect 763 178 779 212
rect 823 178 839 212
rect 941 178 957 212
rect 1001 178 1017 212
rect 1119 178 1135 212
rect 1179 178 1195 212
rect 1297 178 1313 212
rect 1357 178 1373 212
rect -1441 128 -1407 144
rect -1441 -144 -1407 -128
rect -1263 128 -1229 144
rect -1263 -144 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 144
rect 1229 -144 1263 -128
rect 1407 128 1441 144
rect 1407 -144 1441 -128
rect -1373 -212 -1357 -178
rect -1313 -212 -1297 -178
rect -1195 -212 -1179 -178
rect -1135 -212 -1119 -178
rect -1017 -212 -1001 -178
rect -957 -212 -941 -178
rect -839 -212 -823 -178
rect -779 -212 -763 -178
rect -661 -212 -645 -178
rect -601 -212 -585 -178
rect -483 -212 -467 -178
rect -423 -212 -407 -178
rect -305 -212 -289 -178
rect -245 -212 -229 -178
rect -127 -212 -111 -178
rect -67 -212 -51 -178
rect 51 -212 67 -178
rect 111 -212 127 -178
rect 229 -212 245 -178
rect 289 -212 305 -178
rect 407 -212 423 -178
rect 467 -212 483 -178
rect 585 -212 601 -178
rect 645 -212 661 -178
rect 763 -212 779 -178
rect 823 -212 839 -178
rect 941 -212 957 -178
rect 1001 -212 1017 -178
rect 1119 -212 1135 -178
rect 1179 -212 1195 -178
rect 1297 -212 1313 -178
rect 1357 -212 1373 -178
<< viali >>
rect -1357 178 -1313 212
rect -1179 178 -1135 212
rect -1001 178 -957 212
rect -823 178 -779 212
rect -645 178 -601 212
rect -467 178 -423 212
rect -289 178 -245 212
rect -111 178 -67 212
rect 67 178 111 212
rect 245 178 289 212
rect 423 178 467 212
rect 601 178 645 212
rect 779 178 823 212
rect 957 178 1001 212
rect 1135 178 1179 212
rect 1313 178 1357 212
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
rect -1357 -212 -1313 -178
rect -1179 -212 -1135 -178
rect -1001 -212 -957 -178
rect -823 -212 -779 -178
rect -645 -212 -601 -178
rect -467 -212 -423 -178
rect -289 -212 -245 -178
rect -111 -212 -67 -178
rect 67 -212 111 -178
rect 245 -212 289 -178
rect 423 -212 467 -178
rect 601 -212 645 -178
rect 779 -212 823 -178
rect 957 -212 1001 -178
rect 1135 -212 1179 -178
rect 1313 -212 1357 -178
<< metal1 >>
rect -1373 212 -1297 228
rect -1373 178 -1357 212
rect -1313 178 -1297 212
rect -1373 172 -1297 178
rect -1195 212 -1119 228
rect -1195 178 -1179 212
rect -1135 178 -1119 212
rect -1195 172 -1119 178
rect -1017 212 -941 228
rect -1017 178 -1001 212
rect -957 178 -941 212
rect -1017 172 -941 178
rect -839 212 -763 228
rect -839 178 -823 212
rect -779 178 -763 212
rect -839 172 -763 178
rect -661 212 -585 228
rect -661 178 -645 212
rect -601 178 -585 212
rect -661 172 -585 178
rect -483 212 -407 228
rect -483 178 -467 212
rect -423 178 -407 212
rect -483 172 -407 178
rect -305 212 -229 228
rect -305 178 -289 212
rect -245 178 -229 212
rect -305 172 -229 178
rect -127 212 -51 228
rect -127 178 -111 212
rect -67 178 -51 212
rect -127 172 -51 178
rect 51 212 127 228
rect 51 178 67 212
rect 111 178 127 212
rect 51 172 127 178
rect 229 212 305 228
rect 229 178 245 212
rect 289 178 305 212
rect 229 172 305 178
rect 407 212 483 228
rect 407 178 423 212
rect 467 178 483 212
rect 407 172 483 178
rect 585 212 661 228
rect 585 178 601 212
rect 645 178 661 212
rect 585 172 661 178
rect 763 212 839 228
rect 763 178 779 212
rect 823 178 839 212
rect 763 172 839 178
rect 941 212 1017 228
rect 941 178 957 212
rect 1001 178 1017 212
rect 941 172 1017 178
rect 1119 212 1195 228
rect 1119 178 1135 212
rect 1179 178 1195 212
rect 1119 172 1195 178
rect 1297 212 1373 228
rect 1297 178 1313 212
rect 1357 178 1373 212
rect 1297 172 1373 178
rect -1447 128 -1401 140
rect -1447 -128 -1441 128
rect -1407 -128 -1401 128
rect -1447 -140 -1401 -128
rect -1269 128 -1223 140
rect -1269 -128 -1263 128
rect -1229 -128 -1223 128
rect -1269 -140 -1223 -128
rect -1091 128 -1045 140
rect -1091 -128 -1085 128
rect -1051 -128 -1045 128
rect -1091 -140 -1045 -128
rect -913 128 -867 140
rect -913 -128 -907 128
rect -873 -128 -867 128
rect -913 -140 -867 -128
rect -735 128 -689 140
rect -735 -128 -729 128
rect -695 -128 -689 128
rect -735 -140 -689 -128
rect -557 128 -511 140
rect -557 -128 -551 128
rect -517 -128 -511 128
rect -557 -140 -511 -128
rect -379 128 -333 140
rect -379 -128 -373 128
rect -339 -128 -333 128
rect -379 -140 -333 -128
rect -201 128 -155 140
rect -201 -128 -195 128
rect -161 -128 -155 128
rect -201 -140 -155 -128
rect -23 128 23 140
rect -23 -128 -17 128
rect 17 -128 23 128
rect -23 -140 23 -128
rect 155 128 201 140
rect 155 -128 161 128
rect 195 -128 201 128
rect 155 -140 201 -128
rect 333 128 379 140
rect 333 -128 339 128
rect 373 -128 379 128
rect 333 -140 379 -128
rect 511 128 557 140
rect 511 -128 517 128
rect 551 -128 557 128
rect 511 -140 557 -128
rect 689 128 735 140
rect 689 -128 695 128
rect 729 -128 735 128
rect 689 -140 735 -128
rect 867 128 913 140
rect 867 -128 873 128
rect 907 -128 913 128
rect 867 -140 913 -128
rect 1045 128 1091 140
rect 1045 -128 1051 128
rect 1085 -128 1091 128
rect 1045 -140 1091 -128
rect 1223 128 1269 140
rect 1223 -128 1229 128
rect 1263 -128 1269 128
rect 1223 -140 1269 -128
rect 1401 128 1447 140
rect 1401 -128 1407 128
rect 1441 -128 1447 128
rect 1401 -140 1447 -128
rect -1373 -178 -1297 -172
rect -1373 -212 -1357 -178
rect -1313 -212 -1297 -178
rect -1373 -228 -1297 -212
rect -1195 -178 -1119 -172
rect -1195 -212 -1179 -178
rect -1135 -212 -1119 -178
rect -1195 -228 -1119 -212
rect -1017 -178 -941 -172
rect -1017 -212 -1001 -178
rect -957 -212 -941 -178
rect -1017 -228 -941 -212
rect -839 -178 -763 -172
rect -839 -212 -823 -178
rect -779 -212 -763 -178
rect -839 -228 -763 -212
rect -661 -178 -585 -172
rect -661 -212 -645 -178
rect -601 -212 -585 -178
rect -661 -228 -585 -212
rect -483 -178 -407 -172
rect -483 -212 -467 -178
rect -423 -212 -407 -178
rect -483 -228 -407 -212
rect -305 -178 -229 -172
rect -305 -212 -289 -178
rect -245 -212 -229 -178
rect -305 -228 -229 -212
rect -127 -178 -51 -172
rect -127 -212 -111 -178
rect -67 -212 -51 -178
rect -127 -228 -51 -212
rect 51 -178 127 -172
rect 51 -212 67 -178
rect 111 -212 127 -178
rect 51 -228 127 -212
rect 229 -178 305 -172
rect 229 -212 245 -178
rect 289 -212 305 -178
rect 229 -228 305 -212
rect 407 -178 483 -172
rect 407 -212 423 -178
rect 467 -212 483 -178
rect 407 -228 483 -212
rect 585 -178 661 -172
rect 585 -212 601 -178
rect 645 -212 661 -178
rect 585 -228 661 -212
rect 763 -178 839 -172
rect 763 -212 779 -178
rect 823 -212 839 -178
rect 763 -228 839 -212
rect 941 -178 1017 -172
rect 941 -212 957 -178
rect 1001 -212 1017 -178
rect 941 -228 1017 -212
rect 1119 -178 1195 -172
rect 1119 -212 1135 -178
rect 1179 -212 1195 -178
rect 1119 -228 1195 -212
rect 1297 -178 1373 -172
rect 1297 -212 1313 -178
rect 1357 -212 1373 -178
rect 1297 -228 1373 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 16 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
