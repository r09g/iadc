magic
tech sky130A
timestamp 1654720150
<< nmos >>
rect -1187 -70 -1127 70
rect -1098 -70 -1038 70
rect -1009 -70 -949 70
rect -920 -70 -860 70
rect -831 -70 -771 70
rect -742 -70 -682 70
rect -653 -70 -593 70
rect -564 -70 -504 70
rect -475 -70 -415 70
rect -386 -70 -326 70
rect -297 -70 -237 70
rect -208 -70 -148 70
rect -119 -70 -59 70
rect -30 -70 30 70
rect 59 -70 119 70
rect 148 -70 208 70
rect 237 -70 297 70
rect 326 -70 386 70
rect 415 -70 475 70
rect 504 -70 564 70
rect 593 -70 653 70
rect 682 -70 742 70
rect 771 -70 831 70
rect 860 -70 920 70
rect 949 -70 1009 70
rect 1038 -70 1098 70
rect 1127 -70 1187 70
<< ndiff >>
rect -1216 64 -1187 70
rect -1216 -64 -1210 64
rect -1193 -64 -1187 64
rect -1216 -70 -1187 -64
rect -1127 64 -1098 70
rect -1127 -64 -1121 64
rect -1104 -64 -1098 64
rect -1127 -70 -1098 -64
rect -1038 64 -1009 70
rect -1038 -64 -1032 64
rect -1015 -64 -1009 64
rect -1038 -70 -1009 -64
rect -949 64 -920 70
rect -949 -64 -943 64
rect -926 -64 -920 64
rect -949 -70 -920 -64
rect -860 64 -831 70
rect -860 -64 -854 64
rect -837 -64 -831 64
rect -860 -70 -831 -64
rect -771 64 -742 70
rect -771 -64 -765 64
rect -748 -64 -742 64
rect -771 -70 -742 -64
rect -682 64 -653 70
rect -682 -64 -676 64
rect -659 -64 -653 64
rect -682 -70 -653 -64
rect -593 64 -564 70
rect -593 -64 -587 64
rect -570 -64 -564 64
rect -593 -70 -564 -64
rect -504 64 -475 70
rect -504 -64 -498 64
rect -481 -64 -475 64
rect -504 -70 -475 -64
rect -415 64 -386 70
rect -415 -64 -409 64
rect -392 -64 -386 64
rect -415 -70 -386 -64
rect -326 64 -297 70
rect -326 -64 -320 64
rect -303 -64 -297 64
rect -326 -70 -297 -64
rect -237 64 -208 70
rect -237 -64 -231 64
rect -214 -64 -208 64
rect -237 -70 -208 -64
rect -148 64 -119 70
rect -148 -64 -142 64
rect -125 -64 -119 64
rect -148 -70 -119 -64
rect -59 64 -30 70
rect -59 -64 -53 64
rect -36 -64 -30 64
rect -59 -70 -30 -64
rect 30 64 59 70
rect 30 -64 36 64
rect 53 -64 59 64
rect 30 -70 59 -64
rect 119 64 148 70
rect 119 -64 125 64
rect 142 -64 148 64
rect 119 -70 148 -64
rect 208 64 237 70
rect 208 -64 214 64
rect 231 -64 237 64
rect 208 -70 237 -64
rect 297 64 326 70
rect 297 -64 303 64
rect 320 -64 326 64
rect 297 -70 326 -64
rect 386 64 415 70
rect 386 -64 392 64
rect 409 -64 415 64
rect 386 -70 415 -64
rect 475 64 504 70
rect 475 -64 481 64
rect 498 -64 504 64
rect 475 -70 504 -64
rect 564 64 593 70
rect 564 -64 570 64
rect 587 -64 593 64
rect 564 -70 593 -64
rect 653 64 682 70
rect 653 -64 659 64
rect 676 -64 682 64
rect 653 -70 682 -64
rect 742 64 771 70
rect 742 -64 748 64
rect 765 -64 771 64
rect 742 -70 771 -64
rect 831 64 860 70
rect 831 -64 837 64
rect 854 -64 860 64
rect 831 -70 860 -64
rect 920 64 949 70
rect 920 -64 926 64
rect 943 -64 949 64
rect 920 -70 949 -64
rect 1009 64 1038 70
rect 1009 -64 1015 64
rect 1032 -64 1038 64
rect 1009 -70 1038 -64
rect 1098 64 1127 70
rect 1098 -64 1104 64
rect 1121 -64 1127 64
rect 1098 -70 1127 -64
rect 1187 64 1216 70
rect 1187 -64 1193 64
rect 1210 -64 1216 64
rect 1187 -70 1216 -64
<< ndiffc >>
rect -1210 -64 -1193 64
rect -1121 -64 -1104 64
rect -1032 -64 -1015 64
rect -943 -64 -926 64
rect -854 -64 -837 64
rect -765 -64 -748 64
rect -676 -64 -659 64
rect -587 -64 -570 64
rect -498 -64 -481 64
rect -409 -64 -392 64
rect -320 -64 -303 64
rect -231 -64 -214 64
rect -142 -64 -125 64
rect -53 -64 -36 64
rect 36 -64 53 64
rect 125 -64 142 64
rect 214 -64 231 64
rect 303 -64 320 64
rect 392 -64 409 64
rect 481 -64 498 64
rect 570 -64 587 64
rect 659 -64 676 64
rect 748 -64 765 64
rect 837 -64 854 64
rect 926 -64 943 64
rect 1015 -64 1032 64
rect 1104 -64 1121 64
rect 1193 -64 1210 64
<< poly >>
rect -1178 106 -1136 114
rect -1178 97 -1170 106
rect -1187 89 -1170 97
rect -1144 97 -1136 106
rect -1089 106 -1047 114
rect -1089 97 -1081 106
rect -1144 89 -1127 97
rect -1187 70 -1127 89
rect -1098 89 -1081 97
rect -1055 97 -1047 106
rect -1000 106 -958 114
rect -1000 97 -992 106
rect -1055 89 -1038 97
rect -1098 70 -1038 89
rect -1009 89 -992 97
rect -966 97 -958 106
rect -911 106 -869 114
rect -911 97 -903 106
rect -966 89 -949 97
rect -1009 70 -949 89
rect -920 89 -903 97
rect -877 97 -869 106
rect -822 106 -780 114
rect -822 97 -814 106
rect -877 89 -860 97
rect -920 70 -860 89
rect -831 89 -814 97
rect -788 97 -780 106
rect -733 106 -691 114
rect -733 97 -725 106
rect -788 89 -771 97
rect -831 70 -771 89
rect -742 89 -725 97
rect -699 97 -691 106
rect -644 106 -602 114
rect -644 97 -636 106
rect -699 89 -682 97
rect -742 70 -682 89
rect -653 89 -636 97
rect -610 97 -602 106
rect -555 106 -513 114
rect -555 97 -547 106
rect -610 89 -593 97
rect -653 70 -593 89
rect -564 89 -547 97
rect -521 97 -513 106
rect -466 106 -424 114
rect -466 97 -458 106
rect -521 89 -504 97
rect -564 70 -504 89
rect -475 89 -458 97
rect -432 97 -424 106
rect -377 106 -335 114
rect -377 97 -369 106
rect -432 89 -415 97
rect -475 70 -415 89
rect -386 89 -369 97
rect -343 97 -335 106
rect -288 106 -246 114
rect -288 97 -280 106
rect -343 89 -326 97
rect -386 70 -326 89
rect -297 89 -280 97
rect -254 97 -246 106
rect -199 106 -157 114
rect -199 97 -191 106
rect -254 89 -237 97
rect -297 70 -237 89
rect -208 89 -191 97
rect -165 97 -157 106
rect -110 106 -68 114
rect -110 97 -102 106
rect -165 89 -148 97
rect -208 70 -148 89
rect -119 89 -102 97
rect -76 97 -68 106
rect -21 106 21 114
rect -21 97 -13 106
rect -76 89 -59 97
rect -119 70 -59 89
rect -30 89 -13 97
rect 13 97 21 106
rect 68 106 110 114
rect 68 97 76 106
rect 13 89 30 97
rect -30 70 30 89
rect 59 89 76 97
rect 102 97 110 106
rect 157 106 199 114
rect 157 97 165 106
rect 102 89 119 97
rect 59 70 119 89
rect 148 89 165 97
rect 191 97 199 106
rect 246 106 288 114
rect 246 97 254 106
rect 191 89 208 97
rect 148 70 208 89
rect 237 89 254 97
rect 280 97 288 106
rect 335 106 377 114
rect 335 97 343 106
rect 280 89 297 97
rect 237 70 297 89
rect 326 89 343 97
rect 369 97 377 106
rect 424 106 466 114
rect 424 97 432 106
rect 369 89 386 97
rect 326 70 386 89
rect 415 89 432 97
rect 458 97 466 106
rect 513 106 555 114
rect 513 97 521 106
rect 458 89 475 97
rect 415 70 475 89
rect 504 89 521 97
rect 547 97 555 106
rect 602 106 644 114
rect 602 97 610 106
rect 547 89 564 97
rect 504 70 564 89
rect 593 89 610 97
rect 636 97 644 106
rect 691 106 733 114
rect 691 97 699 106
rect 636 89 653 97
rect 593 70 653 89
rect 682 89 699 97
rect 725 97 733 106
rect 780 106 822 114
rect 780 97 788 106
rect 725 89 742 97
rect 682 70 742 89
rect 771 89 788 97
rect 814 97 822 106
rect 869 106 911 114
rect 869 97 877 106
rect 814 89 831 97
rect 771 70 831 89
rect 860 89 877 97
rect 903 97 911 106
rect 958 106 1000 114
rect 958 97 966 106
rect 903 89 920 97
rect 860 70 920 89
rect 949 89 966 97
rect 992 97 1000 106
rect 1047 106 1089 114
rect 1047 97 1055 106
rect 992 89 1009 97
rect 949 70 1009 89
rect 1038 89 1055 97
rect 1081 97 1089 106
rect 1136 106 1178 114
rect 1136 97 1144 106
rect 1081 89 1098 97
rect 1038 70 1098 89
rect 1127 89 1144 97
rect 1170 97 1178 106
rect 1170 89 1187 97
rect 1127 70 1187 89
rect -1187 -89 -1127 -70
rect -1187 -97 -1170 -89
rect -1178 -106 -1170 -97
rect -1144 -97 -1127 -89
rect -1098 -89 -1038 -70
rect -1098 -97 -1081 -89
rect -1144 -106 -1136 -97
rect -1178 -114 -1136 -106
rect -1089 -106 -1081 -97
rect -1055 -97 -1038 -89
rect -1009 -89 -949 -70
rect -1009 -97 -992 -89
rect -1055 -106 -1047 -97
rect -1089 -114 -1047 -106
rect -1000 -106 -992 -97
rect -966 -97 -949 -89
rect -920 -89 -860 -70
rect -920 -97 -903 -89
rect -966 -106 -958 -97
rect -1000 -114 -958 -106
rect -911 -106 -903 -97
rect -877 -97 -860 -89
rect -831 -89 -771 -70
rect -831 -97 -814 -89
rect -877 -106 -869 -97
rect -911 -114 -869 -106
rect -822 -106 -814 -97
rect -788 -97 -771 -89
rect -742 -89 -682 -70
rect -742 -97 -725 -89
rect -788 -106 -780 -97
rect -822 -114 -780 -106
rect -733 -106 -725 -97
rect -699 -97 -682 -89
rect -653 -89 -593 -70
rect -653 -97 -636 -89
rect -699 -106 -691 -97
rect -733 -114 -691 -106
rect -644 -106 -636 -97
rect -610 -97 -593 -89
rect -564 -89 -504 -70
rect -564 -97 -547 -89
rect -610 -106 -602 -97
rect -644 -114 -602 -106
rect -555 -106 -547 -97
rect -521 -97 -504 -89
rect -475 -89 -415 -70
rect -475 -97 -458 -89
rect -521 -106 -513 -97
rect -555 -114 -513 -106
rect -466 -106 -458 -97
rect -432 -97 -415 -89
rect -386 -89 -326 -70
rect -386 -97 -369 -89
rect -432 -106 -424 -97
rect -466 -114 -424 -106
rect -377 -106 -369 -97
rect -343 -97 -326 -89
rect -297 -89 -237 -70
rect -297 -97 -280 -89
rect -343 -106 -335 -97
rect -377 -114 -335 -106
rect -288 -106 -280 -97
rect -254 -97 -237 -89
rect -208 -89 -148 -70
rect -208 -97 -191 -89
rect -254 -106 -246 -97
rect -288 -114 -246 -106
rect -199 -106 -191 -97
rect -165 -97 -148 -89
rect -119 -89 -59 -70
rect -119 -97 -102 -89
rect -165 -106 -157 -97
rect -199 -114 -157 -106
rect -110 -106 -102 -97
rect -76 -97 -59 -89
rect -30 -89 30 -70
rect -30 -97 -13 -89
rect -76 -106 -68 -97
rect -110 -114 -68 -106
rect -21 -106 -13 -97
rect 13 -97 30 -89
rect 59 -89 119 -70
rect 59 -97 76 -89
rect 13 -106 21 -97
rect -21 -114 21 -106
rect 68 -106 76 -97
rect 102 -97 119 -89
rect 148 -89 208 -70
rect 148 -97 165 -89
rect 102 -106 110 -97
rect 68 -114 110 -106
rect 157 -106 165 -97
rect 191 -97 208 -89
rect 237 -89 297 -70
rect 237 -97 254 -89
rect 191 -106 199 -97
rect 157 -114 199 -106
rect 246 -106 254 -97
rect 280 -97 297 -89
rect 326 -89 386 -70
rect 326 -97 343 -89
rect 280 -106 288 -97
rect 246 -114 288 -106
rect 335 -106 343 -97
rect 369 -97 386 -89
rect 415 -89 475 -70
rect 415 -97 432 -89
rect 369 -106 377 -97
rect 335 -114 377 -106
rect 424 -106 432 -97
rect 458 -97 475 -89
rect 504 -89 564 -70
rect 504 -97 521 -89
rect 458 -106 466 -97
rect 424 -114 466 -106
rect 513 -106 521 -97
rect 547 -97 564 -89
rect 593 -89 653 -70
rect 593 -97 610 -89
rect 547 -106 555 -97
rect 513 -114 555 -106
rect 602 -106 610 -97
rect 636 -97 653 -89
rect 682 -89 742 -70
rect 682 -97 699 -89
rect 636 -106 644 -97
rect 602 -114 644 -106
rect 691 -106 699 -97
rect 725 -97 742 -89
rect 771 -89 831 -70
rect 771 -97 788 -89
rect 725 -106 733 -97
rect 691 -114 733 -106
rect 780 -106 788 -97
rect 814 -97 831 -89
rect 860 -89 920 -70
rect 860 -97 877 -89
rect 814 -106 822 -97
rect 780 -114 822 -106
rect 869 -106 877 -97
rect 903 -97 920 -89
rect 949 -89 1009 -70
rect 949 -97 966 -89
rect 903 -106 911 -97
rect 869 -114 911 -106
rect 958 -106 966 -97
rect 992 -97 1009 -89
rect 1038 -89 1098 -70
rect 1038 -97 1055 -89
rect 992 -106 1000 -97
rect 958 -114 1000 -106
rect 1047 -106 1055 -97
rect 1081 -97 1098 -89
rect 1127 -89 1187 -70
rect 1127 -97 1144 -89
rect 1081 -106 1089 -97
rect 1047 -114 1089 -106
rect 1136 -106 1144 -97
rect 1170 -97 1187 -89
rect 1170 -106 1178 -97
rect 1136 -114 1178 -106
<< polycont >>
rect -1170 89 -1144 106
rect -1081 89 -1055 106
rect -992 89 -966 106
rect -903 89 -877 106
rect -814 89 -788 106
rect -725 89 -699 106
rect -636 89 -610 106
rect -547 89 -521 106
rect -458 89 -432 106
rect -369 89 -343 106
rect -280 89 -254 106
rect -191 89 -165 106
rect -102 89 -76 106
rect -13 89 13 106
rect 76 89 102 106
rect 165 89 191 106
rect 254 89 280 106
rect 343 89 369 106
rect 432 89 458 106
rect 521 89 547 106
rect 610 89 636 106
rect 699 89 725 106
rect 788 89 814 106
rect 877 89 903 106
rect 966 89 992 106
rect 1055 89 1081 106
rect 1144 89 1170 106
rect -1170 -106 -1144 -89
rect -1081 -106 -1055 -89
rect -992 -106 -966 -89
rect -903 -106 -877 -89
rect -814 -106 -788 -89
rect -725 -106 -699 -89
rect -636 -106 -610 -89
rect -547 -106 -521 -89
rect -458 -106 -432 -89
rect -369 -106 -343 -89
rect -280 -106 -254 -89
rect -191 -106 -165 -89
rect -102 -106 -76 -89
rect -13 -106 13 -89
rect 76 -106 102 -89
rect 165 -106 191 -89
rect 254 -106 280 -89
rect 343 -106 369 -89
rect 432 -106 458 -89
rect 521 -106 547 -89
rect 610 -106 636 -89
rect 699 -106 725 -89
rect 788 -106 814 -89
rect 877 -106 903 -89
rect 966 -106 992 -89
rect 1055 -106 1081 -89
rect 1144 -106 1170 -89
<< locali >>
rect -1210 89 -1170 106
rect -1144 89 -1136 106
rect -1089 89 -1081 106
rect -1055 89 -1047 106
rect -1000 89 -992 106
rect -966 89 -958 106
rect -911 89 -903 106
rect -877 89 -869 106
rect -822 89 -814 106
rect -788 89 -780 106
rect -733 89 -725 106
rect -699 89 -691 106
rect -644 89 -636 106
rect -610 89 -602 106
rect -555 89 -547 106
rect -521 89 -513 106
rect -466 89 -458 106
rect -432 89 -424 106
rect -377 89 -369 106
rect -343 89 -335 106
rect -288 89 -280 106
rect -254 89 -246 106
rect -199 89 -191 106
rect -165 89 -157 106
rect -110 89 -102 106
rect -76 89 -68 106
rect -21 89 -13 106
rect 13 89 21 106
rect 68 89 76 106
rect 102 89 110 106
rect 157 89 165 106
rect 191 89 199 106
rect 246 89 254 106
rect 280 89 288 106
rect 335 89 343 106
rect 369 89 377 106
rect 424 89 432 106
rect 458 89 466 106
rect 513 89 521 106
rect 547 89 555 106
rect 602 89 610 106
rect 636 89 644 106
rect 691 89 699 106
rect 725 89 733 106
rect 780 89 788 106
rect 814 89 822 106
rect 869 89 877 106
rect 903 89 911 106
rect 958 89 966 106
rect 992 89 1000 106
rect 1047 89 1055 106
rect 1081 89 1089 106
rect 1136 89 1144 106
rect 1170 89 1210 106
rect -1210 64 -1193 89
rect -1210 -89 -1193 -64
rect -1121 64 -1104 72
rect -1121 -72 -1104 -64
rect -1032 64 -1015 72
rect -1032 -72 -1015 -64
rect -943 64 -926 72
rect -943 -72 -926 -64
rect -854 64 -837 72
rect -854 -72 -837 -64
rect -765 64 -748 72
rect -765 -72 -748 -64
rect -676 64 -659 72
rect -676 -72 -659 -64
rect -587 64 -570 72
rect -587 -72 -570 -64
rect -498 64 -481 72
rect -498 -72 -481 -64
rect -409 64 -392 72
rect -409 -72 -392 -64
rect -320 64 -303 72
rect -320 -72 -303 -64
rect -231 64 -214 72
rect -231 -72 -214 -64
rect -142 64 -125 72
rect -142 -72 -125 -64
rect -53 64 -36 72
rect -53 -72 -36 -64
rect 36 64 53 72
rect 36 -72 53 -64
rect 125 64 142 72
rect 125 -72 142 -64
rect 214 64 231 72
rect 214 -72 231 -64
rect 303 64 320 72
rect 303 -72 320 -64
rect 392 64 409 72
rect 392 -72 409 -64
rect 481 64 498 72
rect 481 -72 498 -64
rect 570 64 587 72
rect 570 -72 587 -64
rect 659 64 676 72
rect 659 -72 676 -64
rect 748 64 765 72
rect 748 -72 765 -64
rect 837 64 854 72
rect 837 -72 854 -64
rect 926 64 943 72
rect 926 -72 943 -64
rect 1015 64 1032 72
rect 1015 -72 1032 -64
rect 1104 64 1121 72
rect 1104 -72 1121 -64
rect 1193 64 1210 89
rect 1193 -89 1210 -64
rect -1210 -106 -1170 -89
rect -1144 -106 -1136 -89
rect -1089 -106 -1081 -89
rect -1055 -106 -1047 -89
rect -1000 -106 -992 -89
rect -966 -106 -958 -89
rect -911 -106 -903 -89
rect -877 -106 -869 -89
rect -822 -106 -814 -89
rect -788 -106 -780 -89
rect -733 -106 -725 -89
rect -699 -106 -691 -89
rect -644 -106 -636 -89
rect -610 -106 -602 -89
rect -555 -106 -547 -89
rect -521 -106 -513 -89
rect -466 -106 -458 -89
rect -432 -106 -424 -89
rect -377 -106 -369 -89
rect -343 -106 -335 -89
rect -288 -106 -280 -89
rect -254 -106 -246 -89
rect -199 -106 -191 -89
rect -165 -106 -157 -89
rect -110 -106 -102 -89
rect -76 -106 -68 -89
rect -21 -106 -13 -89
rect 13 -106 21 -89
rect 68 -106 76 -89
rect 102 -106 110 -89
rect 157 -106 165 -89
rect 191 -106 199 -89
rect 246 -106 254 -89
rect 280 -106 288 -89
rect 335 -106 343 -89
rect 369 -106 377 -89
rect 424 -106 432 -89
rect 458 -106 466 -89
rect 513 -106 521 -89
rect 547 -106 555 -89
rect 602 -106 610 -89
rect 636 -106 644 -89
rect 691 -106 699 -89
rect 725 -106 733 -89
rect 780 -106 788 -89
rect 814 -106 822 -89
rect 869 -106 877 -89
rect 903 -106 911 -89
rect 958 -106 966 -89
rect 992 -106 1000 -89
rect 1047 -106 1055 -89
rect 1081 -106 1089 -89
rect 1136 -106 1144 -89
rect 1170 -106 1210 -89
<< viali >>
rect -1081 89 -1055 106
rect -992 89 -966 106
rect -903 89 -877 106
rect -814 89 -788 106
rect -725 89 -699 106
rect -636 89 -610 106
rect -547 89 -521 106
rect -458 89 -432 106
rect -369 89 -343 106
rect -280 89 -254 106
rect -191 89 -165 106
rect -102 89 -76 106
rect -13 89 13 106
rect 76 89 102 106
rect 165 89 191 106
rect 254 89 280 106
rect 343 89 369 106
rect 432 89 458 106
rect 521 89 547 106
rect 610 89 636 106
rect 699 89 725 106
rect 788 89 814 106
rect 877 89 903 106
rect 966 89 992 106
rect 1055 89 1081 106
rect -1081 -106 -1055 -89
rect -992 -106 -966 -89
rect -903 -106 -877 -89
rect -814 -106 -788 -89
rect -725 -106 -699 -89
rect -636 -106 -610 -89
rect -547 -106 -521 -89
rect -458 -106 -432 -89
rect -369 -106 -343 -89
rect -280 -106 -254 -89
rect -191 -106 -165 -89
rect -102 -106 -76 -89
rect -13 -106 13 -89
rect 76 -106 102 -89
rect 165 -106 191 -89
rect 254 -106 280 -89
rect 343 -106 369 -89
rect 432 -106 458 -89
rect 521 -106 547 -89
rect 610 -106 636 -89
rect 699 -106 725 -89
rect 788 -106 814 -89
rect 877 -106 903 -89
rect 966 -106 992 -89
rect 1055 -106 1081 -89
<< metal1 >>
rect -1087 106 -1049 109
rect -1087 89 -1081 106
rect -1055 89 -1049 106
rect -1087 86 -1049 89
rect -998 106 -960 109
rect -998 89 -992 106
rect -966 89 -960 106
rect -998 86 -960 89
rect -909 106 -871 109
rect -909 89 -903 106
rect -877 89 -871 106
rect -909 86 -871 89
rect -820 106 -782 109
rect -820 89 -814 106
rect -788 89 -782 106
rect -820 86 -782 89
rect -731 106 -693 109
rect -731 89 -725 106
rect -699 89 -693 106
rect -731 86 -693 89
rect -642 106 -604 109
rect -642 89 -636 106
rect -610 89 -604 106
rect -642 86 -604 89
rect -553 106 -515 109
rect -553 89 -547 106
rect -521 89 -515 106
rect -553 86 -515 89
rect -464 106 -426 109
rect -464 89 -458 106
rect -432 89 -426 106
rect -464 86 -426 89
rect -375 106 -337 109
rect -375 89 -369 106
rect -343 89 -337 106
rect -375 86 -337 89
rect -286 106 -248 109
rect -286 89 -280 106
rect -254 89 -248 106
rect -286 86 -248 89
rect -197 106 -159 109
rect -197 89 -191 106
rect -165 89 -159 106
rect -197 86 -159 89
rect -108 106 -70 109
rect -108 89 -102 106
rect -76 89 -70 106
rect -108 86 -70 89
rect -19 106 19 109
rect -19 89 -13 106
rect 13 89 19 106
rect -19 86 19 89
rect 70 106 108 109
rect 70 89 76 106
rect 102 89 108 106
rect 70 86 108 89
rect 159 106 197 109
rect 159 89 165 106
rect 191 89 197 106
rect 159 86 197 89
rect 248 106 286 109
rect 248 89 254 106
rect 280 89 286 106
rect 248 86 286 89
rect 337 106 375 109
rect 337 89 343 106
rect 369 89 375 106
rect 337 86 375 89
rect 426 106 464 109
rect 426 89 432 106
rect 458 89 464 106
rect 426 86 464 89
rect 515 106 553 109
rect 515 89 521 106
rect 547 89 553 106
rect 515 86 553 89
rect 604 106 642 109
rect 604 89 610 106
rect 636 89 642 106
rect 604 86 642 89
rect 693 106 731 109
rect 693 89 699 106
rect 725 89 731 106
rect 693 86 731 89
rect 782 106 820 109
rect 782 89 788 106
rect 814 89 820 106
rect 782 86 820 89
rect 871 106 909 109
rect 871 89 877 106
rect 903 89 909 106
rect 871 86 909 89
rect 960 106 998 109
rect 960 89 966 106
rect 992 89 998 106
rect 960 86 998 89
rect 1049 106 1087 109
rect 1049 89 1055 106
rect 1081 89 1087 106
rect 1049 86 1087 89
rect -1087 -89 -1049 -86
rect -1087 -106 -1081 -89
rect -1055 -106 -1049 -89
rect -1087 -109 -1049 -106
rect -998 -89 -960 -86
rect -998 -106 -992 -89
rect -966 -106 -960 -89
rect -998 -109 -960 -106
rect -909 -89 -871 -86
rect -909 -106 -903 -89
rect -877 -106 -871 -89
rect -909 -109 -871 -106
rect -820 -89 -782 -86
rect -820 -106 -814 -89
rect -788 -106 -782 -89
rect -820 -109 -782 -106
rect -731 -89 -693 -86
rect -731 -106 -725 -89
rect -699 -106 -693 -89
rect -731 -109 -693 -106
rect -642 -89 -604 -86
rect -642 -106 -636 -89
rect -610 -106 -604 -89
rect -642 -109 -604 -106
rect -553 -89 -515 -86
rect -553 -106 -547 -89
rect -521 -106 -515 -89
rect -553 -109 -515 -106
rect -464 -89 -426 -86
rect -464 -106 -458 -89
rect -432 -106 -426 -89
rect -464 -109 -426 -106
rect -375 -89 -337 -86
rect -375 -106 -369 -89
rect -343 -106 -337 -89
rect -375 -109 -337 -106
rect -286 -89 -248 -86
rect -286 -106 -280 -89
rect -254 -106 -248 -89
rect -286 -109 -248 -106
rect -197 -89 -159 -86
rect -197 -106 -191 -89
rect -165 -106 -159 -89
rect -197 -109 -159 -106
rect -108 -89 -70 -86
rect -108 -106 -102 -89
rect -76 -106 -70 -89
rect -108 -109 -70 -106
rect -19 -89 19 -86
rect -19 -106 -13 -89
rect 13 -106 19 -89
rect -19 -109 19 -106
rect 70 -89 108 -86
rect 70 -106 76 -89
rect 102 -106 108 -89
rect 70 -109 108 -106
rect 159 -89 197 -86
rect 159 -106 165 -89
rect 191 -106 197 -89
rect 159 -109 197 -106
rect 248 -89 286 -86
rect 248 -106 254 -89
rect 280 -106 286 -89
rect 248 -109 286 -106
rect 337 -89 375 -86
rect 337 -106 343 -89
rect 369 -106 375 -89
rect 337 -109 375 -106
rect 426 -89 464 -86
rect 426 -106 432 -89
rect 458 -106 464 -89
rect 426 -109 464 -106
rect 515 -89 553 -86
rect 515 -106 521 -89
rect 547 -106 553 -89
rect 515 -109 553 -106
rect 604 -89 642 -86
rect 604 -106 610 -89
rect 636 -106 642 -89
rect 604 -109 642 -106
rect 693 -89 731 -86
rect 693 -106 699 -89
rect 725 -106 731 -89
rect 693 -109 731 -106
rect 782 -89 820 -86
rect 782 -106 788 -89
rect 814 -106 820 -89
rect 782 -109 820 -106
rect 871 -89 909 -86
rect 871 -106 877 -89
rect 903 -106 909 -89
rect 871 -109 909 -106
rect 960 -89 998 -86
rect 960 -106 966 -89
rect 992 -106 998 -89
rect 960 -109 998 -106
rect 1049 -89 1087 -86
rect 1049 -106 1055 -89
rect 1081 -106 1087 -89
rect 1049 -109 1087 -106
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 27 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
