* NGSPICE file created from ota_flat.ext - technology: sky130A

.subckt ota_flat ip in p1 p1_b p2 p2_b op on i_bias cm VDD VSS
X0 cm p2 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=1.1958e+13p pd=1.0498e+08u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X1 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=1.1368e+13p pd=9.464e+07u as=1.456e+13p ps=1.216e+08u w=1.4e+06u l=600000u
X2 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=1.582e+13p pd=1.318e+08u as=1.09496e+13p ps=9.46e+07u w=1.4e+06u l=600000u
X3 sc_cmfb_0/transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 sc_cmfb_0/transmission_gate_5/in p1_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=4.488e+12p pd=3.38e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X5 cm p2 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X6 a_12106_n11502# cm VSS VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=8.323e+13p ps=6.929e+08u w=1.4e+06u l=600000u
X7 op p2_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=1.01488e+13p pd=8.096e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X8 sc_cmfb_0/transmission_gate_5/out p2 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=8.212e+12p ps=7.108e+07u w=520000u l=150000u
X9 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=1.0556e+13p pd=8.788e+07u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_12398_n9962# cm cm VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.3884e+13p pd=1.9932e+08u as=0p ps=0u w=1.4e+06u l=600000u
X12 sc_cmfb_0/transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X13 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=1.624e+13p pd=1.352e+08u as=0p ps=0u w=1.4e+06u l=600000u
X14 op p2 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X15 VDD VDD a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.2152e+13p ps=1.0136e+08u w=1.4e+06u l=600000u
X17 a_n5928_n12940# ip a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+12p pd=2.98e+07u as=4.7212e+13p ps=3.9404e+08u w=1.2e+06u l=200000u
X18 cm p2 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X19 a_n6313_n3270# a_n6313_n3270# a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8_lvt ad=4.872e+12p pd=4.056e+07u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_n5580_n13620# in a_n5928_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.48e+12p ps=2.98e+07u w=1.2e+06u l=200000u
X22 sc_cmfb_0/transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X23 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n5580_n13620# a_n5580_n13620# a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 sc_cmfb_0/transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=1.06e+13p ps=8.112e+07u w=1.36e+06u l=150000u
X26 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=1.09496e+13p pd=9.46e+07u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.0556e+13p pd=8.788e+07u as=0p ps=0u w=1.4e+06u l=600000u
X31 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 sc_cmfb_0/transmission_gate_8/in p1 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=0p ps=0u w=520000u l=150000u
X33 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 c1_12802_1831# m3_12702_1731# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X35 on p1_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=1.01488e+13p pd=8.096e+07u as=4.8824e+12p ps=3.71e+07u w=1.36e+06u l=150000u
X36 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=1.624e+13p pd=1.352e+08u as=2.1112e+13p ps=1.7576e+08u w=1.4e+06u l=600000u
X37 op p1 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X38 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X40 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X41 VDD bias_b a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+12p ps=3.38e+07u w=1.4e+06u l=600000u
X42 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X43 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X44 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X45 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X46 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X47 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X48 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X49 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X50 a_n6313_n5010# a_n6313_n5010# a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8 ad=4.872e+12p pd=4.056e+07u as=0p ps=0u w=1.4e+06u l=600000u
X51 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X52 cm p1 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.8668e+12p ps=1.862e+07u w=520000u l=150000u
X53 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X54 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X55 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.872e+12p ps=4.056e+07u w=1.4e+06u l=600000u
X56 sc_cmfb_0/transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=1.8668e+12p pd=1.862e+07u as=0p ps=0u w=520000u l=150000u
X57 sc_cmfb_0/transmission_gate_5/out p2_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=4.8824e+12p pd=3.71e+07u as=0p ps=0u w=1.36e+06u l=150000u
X58 sc_cmfb_0/transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X59 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X60 sc_cmfb_0/transmission_gate_5/in p1 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X61 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X62 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X63 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X64 sc_cmfb_0/transmission_gate_5/out p2 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X65 sc_cmfb_0/transmission_gate_8/out p2_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=5.2768e+12p pd=4.04e+07u as=0p ps=0u w=1.36e+06u l=150000u
X66 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X67 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X68 op p2_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X69 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X70 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X71 sc_cmfb_0/transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X72 sc_cmfb_0/transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X73 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X74 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X75 op p2 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X76 sc_cmfb_0/transmission_gate_8/out p1_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X77 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X78 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X79 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X80 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X81 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X82 c1_16402_31# m3_16302_n69# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X83 c1_7402_n3569# m3_7302_n3669# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X84 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X85 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X86 cm p2_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X87 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X88 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X89 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X90 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X91 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X92 sc_cmfb_0/transmission_gate_8/in p2_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X93 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X94 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X95 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X96 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X97 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X98 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X99 sc_cmfb_0/transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X100 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X101 VSS VSS a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X102 on sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X103 VDD VDD op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X104 on p1_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X105 sc_cmfb_0/transmission_gate_8/in p1_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X106 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X107 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X108 a_n1110_n5852# bias_c a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8 ad=1.624e+12p pd=1.352e+07u as=0p ps=0u w=1.4e+06u l=600000u
X109 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X110 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X111 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X112 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X113 op p1_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X114 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X115 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X116 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X117 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X118 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X119 on VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X120 bias_d a_n1110_n5852# sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X121 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X122 a_n5928_n13620# in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X123 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X124 a_n5928_n12940# a_n5928_n12940# a_n5928_n12940# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X125 cm p1_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X126 a_n1651_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X127 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X128 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X129 a_n6313_n3270# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X130 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X131 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X132 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X133 sc_cmfb_0/transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X134 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X135 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X136 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X137 sc_cmfb_0/transmission_gate_5/in p2_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X138 a_n6313_n4140# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X139 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X140 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X141 sc_cmfb_0/transmission_gate_5/in p2 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X142 a_n1110_n5852# bias_c a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X143 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X144 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X145 sc_cmfb_0/transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X146 on p2_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X147 sc_cmfb_0/transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X148 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X149 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X150 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X151 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X152 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X153 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X154 sc_cmfb_0/transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X155 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X156 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X157 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X158 sc_cmfb_0/transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X159 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X160 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X161 on p2_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X162 a_n6313_n3270# a_n6313_n3270# a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X163 cm p2 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X164 sc_cmfb_0/transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X165 on VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X166 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X167 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X168 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X169 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X170 c1_14602_1831# m3_14502_1731# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X171 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X172 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X173 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X174 sc_cmfb_0/transmission_gate_8/in p2 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.0176e+12p ps=2.024e+07u w=520000u l=150000u
X175 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X176 sc_cmfb_0/transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X177 cm p1_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X178 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X179 on p2_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X180 c1_14602_n7169# m3_14502_n7269# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X181 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X182 sc_cmfb_0/transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X183 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X184 VSS VSS a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X185 sc_cmfb_0/transmission_gate_5/out p1_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X186 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X187 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X188 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X189 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X190 cm p2_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X191 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X192 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X193 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X194 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X195 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X196 VSS VSS a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X197 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X198 a_n5580_n13620# a_n5580_n13620# a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X199 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X200 c1_16402_n5369# m3_16302_n5469# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X201 a_12106_n9962# cm a_11928_n10732# VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=8.12e+11p ps=6.76e+06u w=1.4e+06u l=600000u
X202 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X203 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X204 on p2 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X205 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X206 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X207 sc_cmfb_0/transmission_gate_5/out p2_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X208 sc_cmfb_0/transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X209 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X210 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X211 a_n5928_n13620# a_n5928_n13620# a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X212 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X213 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X214 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X215 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X216 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X217 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X218 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X219 sc_cmfb_0/transmission_gate_5/out p2 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X220 VDD VDD a_n1110_n5852# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X221 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X222 op p2_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X223 sc_cmfb_0/transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X224 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X225 sc_cmfb_0/transmission_gate_5/in p1_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X226 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X227 sc_cmfb_0/transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X228 a_n5928_n12940# a_n5928_n12940# a_n5928_n12940# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X229 op p2 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X230 on p2 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X231 sc_cmfb_0/transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X232 sc_cmfb_0/transmission_gate_8/out p1 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X233 sc_cmfb_0/transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X234 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X235 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X236 a_n5580_n13620# in a_n5928_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X237 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X238 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X239 a_n6313_n3270# bias_c bias_b VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.624e+12p ps=1.352e+07u w=1.4e+06u l=600000u
X240 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X241 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X242 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X243 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X244 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X245 sc_cmfb_0/transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X246 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X247 VDD bias_b a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X248 on p2 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X249 a_n5580_n13620# a_n5580_n13620# a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X250 sc_cmfb_0/transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X251 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X252 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X253 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X254 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X255 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X256 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X257 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X258 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X259 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X260 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X261 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X262 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X263 VDD VDD a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X264 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X265 cm p2 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X266 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X267 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X268 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X269 cm p1 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X270 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X271 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X272 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X273 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X274 i_bias i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X275 VDD bias_b a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X276 sc_cmfb_0/transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X277 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X278 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X279 VSS VSS a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X280 sc_cmfb_0/transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X281 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X282 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X283 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X284 on sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X285 sc_cmfb_0/transmission_gate_8/out p2 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X286 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X287 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X288 sc_cmfb_0/transmission_gate_5/in p2_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X289 a_11230_n11502# cm VSS VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=0p ps=0u w=1.4e+06u l=600000u
X290 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X291 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X292 a_n6313_n3270# a_n6313_n3270# a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X293 VDD VDD op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X294 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X295 a_n6313_n4140# bias_c cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X296 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X297 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X298 sc_cmfb_0/transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X299 sc_cmfb_0/transmission_gate_5/in p2 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X300 cm p2 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X301 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X302 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X303 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X304 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X305 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X306 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X307 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X308 sc_cmfb_0/transmission_gate_8/in p2 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X309 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X310 sc_cmfb_0/transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X311 cm p1 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X312 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X313 c1_7402_31# m3_7302_n69# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X314 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X315 op sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X316 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X317 sc_cmfb_0/transmission_gate_5/out p1 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X318 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X319 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X320 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X321 sc_cmfb_0/transmission_gate_8/in p1 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X322 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X323 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X324 c1_16402_1831# m3_16302_1731# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X325 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X326 op p1 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X327 c1_7402_1831# m3_7302_1731# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X328 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X329 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X330 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X331 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X332 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X333 sc_cmfb_0/transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X334 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X335 a_11522_n11502# cm a_11344_n10732# VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=8.12e+11p ps=6.76e+06u w=1.4e+06u l=600000u
X336 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X337 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X338 on sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X339 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X340 sc_cmfb_0/transmission_gate_8/out p2 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X341 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X342 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X343 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X344 a_n6313_n3270# bias_c bias_b VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X345 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X346 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X347 a_n5928_n13620# in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X348 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X349 a_n5580_n13620# ip a_n5928_n12940# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X350 sc_cmfb_0/transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X351 a_n6313_n5010# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X352 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X353 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X354 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X355 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X356 sc_cmfb_0/transmission_gate_8/out p2_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X357 VDD VDD cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X358 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X359 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X360 bias_b bias_c a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X361 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X362 a_11522_n9962# cm cm VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=0p ps=0u w=1.4e+06u l=600000u
X363 c1_16402_n1769# m3_16302_n1869# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X364 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X365 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X366 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X367 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X368 VSS VSS a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X369 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X370 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X371 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X372 a_n6313_n4140# a_n6313_n4140# a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X373 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X374 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X375 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X376 sc_cmfb_0/transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X377 sc_cmfb_0/transmission_gate_5/out p2_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X378 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X379 op op op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X380 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X381 on p1 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X382 op p2_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X383 sc_cmfb_0/transmission_gate_5/out p2 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X384 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X385 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X386 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X387 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X388 op p2 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X389 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X390 cm p1_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X391 sc_cmfb_0/transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X392 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X393 cm p1 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X394 a_11814_n9962# cm cm VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=0p ps=0u w=1.4e+06u l=600000u
X395 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X396 bias_b bias_c a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X397 cm bias_c a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X398 sc_cmfb_0/transmission_gate_5/out p1_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X399 on p1_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X400 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X401 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X402 sc_cmfb_0/transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X403 VDD bias_b a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X404 sc_cmfb_0/transmission_gate_5/in p1 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X405 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X406 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X407 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X408 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X409 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X410 sc_cmfb_0/transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X411 sc_cmfb_0/transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X412 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X413 c1_9202_n7169# m3_9102_n7269# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X414 on p2_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X415 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X416 sc_cmfb_0/transmission_gate_8/out p2 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X417 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X418 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X419 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X420 sc_cmfb_0/transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X421 a_n1651_n11400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X422 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X423 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X424 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X425 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X426 sc_cmfb_0/transmission_gate_7/in p2_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X427 sc_cmfb_0/transmission_gate_8/out p1 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X428 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X429 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X430 sc_cmfb_0/transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X431 sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X432 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X433 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X434 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X435 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X436 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X437 on p1 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X438 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X439 cm p2_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X440 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X441 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X442 sc_cmfb_0/transmission_gate_6/in sc_cmfb_0/transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X443 sc_cmfb_0/transmission_gate_5/in p1_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X444 on on on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X445 sc_cmfb_0/transmission_gate_8/in p2_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X446 cm p2 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X447 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X448 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X449 VSS VSS a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X450 sc_cmfb_0/transmission_gate_5/in p2_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X451 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X452 bias_b bias_c a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X453 sc_cmfb_0/transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X454 a_11230_n9962# cm a_11052_n10732# VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=8.12e+11p ps=6.76e+06u w=1.4e+06u l=600000u
X455 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X456 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X457 sc_cmfb_0/transmission_gate_8/in p2 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X458 sc_cmfb_0/transmission_gate_5/in p2 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X459 a_n1651_n11400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X460 sc_cmfb_0/transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X461 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X462 on on on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X463 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X464 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X465 a_n1110_n5852# a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X466 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X467 cm bias_c a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X468 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X469 sc_cmfb_0/transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X470 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X471 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X472 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X473 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X474 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X475 VDD VDD bias_b VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X476 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X477 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X478 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X479 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X480 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X481 c1_9202_1831# m3_9102_1731# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X482 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X483 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X484 on p2 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X485 VDD bias_b a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X486 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X487 cm p1_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X488 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X489 a_n2185_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X490 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X491 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X492 a_12398_n9962# cm a_12220_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.12e+11p ps=6.76e+06u w=1.4e+06u l=600000u
X493 sc_cmfb_0/transmission_gate_7/in p2 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X494 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X495 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X496 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X497 sc_cmfb_0/transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X498 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X499 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X500 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X501 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X502 a_12398_n11502# cm a_12220_n10732# VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=0p ps=0u w=1.4e+06u l=600000u
X503 a_11814_n11502# cm VSS VSS sky130_fd_pr__nfet_01v8 ad=8.12e+11p pd=6.76e+06u as=0p ps=0u w=1.4e+06u l=600000u
X504 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X505 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X506 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X507 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X508 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X509 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X510 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X511 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X512 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X513 a_n1651_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X514 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X515 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X516 a_n6313_n4140# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X517 a_n6313_n3270# a_n6313_n3270# a_n6313_n3270# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X518 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X519 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X520 sc_cmfb_0/transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X521 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X522 sc_cmfb_0/transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X523 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X524 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X525 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X526 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X527 sc_cmfb_0/transmission_gate_8/out p1_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X528 on p1 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X529 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X530 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X531 op op op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X532 sc_cmfb_0/transmission_gate_8/in p1 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X533 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X534 op sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X535 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X536 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X537 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X538 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X539 VSS VSS op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X540 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X541 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X542 cm p1_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X543 op p1 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X544 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X545 a_n1651_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X546 VDD VDD on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X547 sc_cmfb_0/transmission_gate_5/out p1_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X548 a_12106_n11502# cm a_11928_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X549 a_n6313_n4140# bias_c cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X550 cm p1 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X551 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X552 VSS VSS a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X553 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X554 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X555 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X556 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X557 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X558 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X559 c1_7402_n5369# m3_7302_n5469# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X560 sc_cmfb_0/transmission_gate_5/out p1 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X561 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X562 a_n5580_n13620# ip a_n5928_n12940# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X563 cm p1 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X564 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X565 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X566 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X567 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X568 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X569 a_n5928_n13620# in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X570 sc_cmfb_0/transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X571 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X572 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X573 sc_cmfb_0/transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X574 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X575 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X576 sc_cmfb_0/transmission_gate_8/in p1_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X577 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X578 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X579 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X580 sc_cmfb_0/transmission_gate_8/out p2_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X581 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X582 sc_cmfb_0/transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X583 op p1_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X584 a_n6313_n5010# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X585 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X586 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X587 op sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X588 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X589 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X590 sc_cmfb_0/transmission_gate_8/out p1_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X591 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X592 sc_cmfb_0/transmission_gate_5/in a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X593 sc_cmfb_0/transmission_gate_5/in p1_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X594 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X595 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X596 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X597 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X598 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X599 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X600 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X601 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X602 sc_cmfb_0/transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X603 a_n6313_n5010# a_n6313_n5010# a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X604 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X605 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X606 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X607 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X608 a_n5928_n13620# a_n5928_n13620# a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X609 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X610 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X611 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X612 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X613 a_n6313_n5010# bias_c a_n1110_n5852# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X614 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X615 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X616 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X617 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X618 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X619 VDD VDD cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X620 sc_cmfb_0/transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X621 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X622 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X623 on p1_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X624 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X625 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X626 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X627 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X628 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X629 sc_cmfb_0/transmission_gate_8/in p1_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X630 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X631 VDD bias_b a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X632 op p1_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X633 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X634 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X635 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X636 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X637 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X638 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X639 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X640 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X641 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X642 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X643 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X644 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X645 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X646 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X647 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X648 sc_cmfb_0/transmission_gate_5/in p1 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X649 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X650 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X651 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X652 cm bias_c a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X653 sc_cmfb_0/transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X654 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X655 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X656 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X657 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X658 sc_cmfb_0/transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X659 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X660 sc_cmfb_0/transmission_gate_8/out p1_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X661 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X662 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X663 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X664 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X665 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X666 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X667 a_n2185_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X668 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X669 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X670 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X671 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X672 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X673 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X674 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X675 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X676 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X677 a_n5928_n13620# a_n5928_n13620# a_n5928_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X678 cm p2_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X679 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X680 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X681 a_n5580_n13620# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X682 a_n6313_n5010# a_n6313_n5010# a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X683 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X684 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X685 c1_16402_n7169# m3_16302_n7269# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X686 a_n5928_n12940# ip a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X687 sc_cmfb_0/transmission_gate_8/in p2_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X688 a_n6313_n3270# bias_c bias_b VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X689 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X690 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X691 cm p1_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X692 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X693 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X694 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X695 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X696 sc_cmfb_0/transmission_gate_5/out p1_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X697 VDD bias_b a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X698 sc_cmfb_0/transmission_gate_8/in p1_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X699 bias_c bias_c bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X700 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X701 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X702 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X703 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X704 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X705 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X706 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X707 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X708 op p1_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X709 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X710 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X711 a_n1110_n5852# bias_c a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X712 c1_7402_n1769# m3_7302_n1869# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X713 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X714 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X715 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X716 cm bias_c a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X717 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X718 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X719 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X720 sc_cmfb_0/transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X721 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X722 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X723 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X724 cm p1_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X725 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X726 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X727 sc_cmfb_0/transmission_gate_8/out p2 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X728 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X729 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X730 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X731 sc_cmfb_0/transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X732 sc_cmfb_0/transmission_gate_5/in p1_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X733 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X734 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X735 sc_cmfb_0/transmission_gate_4/out p1_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X736 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X737 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X738 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X739 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X740 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X741 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X742 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X743 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X744 a_n6313_n4140# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X745 c1_11002_n7169# m3_10902_n7269# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X746 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X747 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X748 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X749 cm p1 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X750 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X751 a_n6313_n5010# a_n6313_n5010# a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X752 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X753 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X754 on VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X755 sc_cmfb_0/transmission_gate_5/out p1 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X756 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X757 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X758 a_n5580_n13620# ip a_n5928_n12940# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X759 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X760 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X761 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X762 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X763 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X764 VSS VSS a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X765 a_n5928_n13620# a_n5928_n13620# a_n5928_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X766 sc_cmfb_0/transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X767 a_n6313_n4140# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X768 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X769 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X770 c1_12802_n7169# m3_12702_n7269# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X771 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X772 a_n2185_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X773 bias_b VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X774 VSS VSS on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X775 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X776 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X777 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X778 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X779 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X780 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X781 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X782 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X783 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X784 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X785 a_n5928_n12940# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X786 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X787 a_n6313_n5010# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X788 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X789 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X790 cm p2 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X791 a_12106_n9962# cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X792 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X793 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X794 sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X795 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X796 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X797 sc_cmfb_0/transmission_gate_8/in p2 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X798 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X799 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X800 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X801 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X802 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X803 sc_cmfb_0/transmission_gate_5/out p2_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X804 sc_cmfb_0/transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X805 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X806 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X807 sc_cmfb_0/transmission_gate_5/out p2 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X808 on p1 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X809 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X810 op p2_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X811 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X812 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X813 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X814 a_n5580_n13620# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X815 op p2 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X816 VDD bias_b a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X817 c1_16402_n3569# m3_16302_n3669# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X818 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X819 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X820 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X821 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X822 a_n5928_n12940# a_n5928_n12940# a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X823 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X824 a_11230_n11502# cm a_11052_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X825 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X826 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X827 a_n1110_n5852# a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X828 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X829 c1_11002_1831# m3_10902_1731# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X830 sc_cmfb_0/transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X831 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X832 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X833 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X834 op VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X835 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X836 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X837 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X838 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X839 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X840 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X841 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X842 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X843 a_11522_n9962# cm a_11344_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X844 sc_cmfb_0/transmission_gate_5/in p1 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X845 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X846 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X847 a_n2185_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X848 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X849 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X850 sc_cmfb_0/transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X851 VSS VSS a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X852 a_n5580_n13620# a_n5580_n13620# a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X853 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X854 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X855 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X856 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X857 a_n2185_n13400# a_n2185_n13400# a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X858 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X859 sc_cmfb_0/transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X860 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X861 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X862 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X863 sc_cmfb_0/transmission_gate_5/in bias_d a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X864 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X865 a_n1651_n13400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X866 sc_cmfb_0/transmission_gate_8/out p1 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X867 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X868 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X869 a_11522_n11502# cm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X870 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X871 VDD bias_b a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X872 op bias_c a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X873 a_n6313_n4140# a_n6313_n4140# a_n6313_n4140# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X874 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X875 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X876 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X877 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X878 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X879 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X880 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X881 a_11814_n9962# cm a_11636_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.12e+11p ps=6.76e+06u w=1.4e+06u l=600000u
X882 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X883 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X884 a_n5580_n13620# in a_n5928_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X885 cm p2_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X886 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X887 cm p1 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X888 a_n5928_n12940# ip a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+06u l=200000u
X889 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X890 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X891 sc_cmfb_0/transmission_gate_8/in p2_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X892 sc_cmfb_0/transmission_gate_5/out p1 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X893 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X894 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X895 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X896 sc_cmfb_0/transmission_gate_5/in p2_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X897 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X898 cm p1 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X899 VDD bias_b a_n6313_n5010# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X900 a_n5580_n13620# a_n5580_n13620# a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X901 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X902 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X903 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X904 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X905 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X906 sc_cmfb_0/transmission_gate_5/in p2 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X907 sc_cmfb_0/transmission_gate_3/out p1 on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X908 a_n2185_n13400# a_n2185_n13400# a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X909 sc_cmfb_0/transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X910 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X911 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X912 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X913 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X914 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X915 VDD bias_b a_n5928_n13620# VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X916 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X917 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X918 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X919 op bias_d a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X920 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X921 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X922 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X923 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X924 sc_cmfb_0/transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X925 sc_cmfb_0/transmission_gate_3/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X926 on sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X927 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X928 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X929 sc_cmfb_0/transmission_gate_8/out p2 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X930 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X931 sc_cmfb_0/transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X932 a_n1651_n13400# bias_d on VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X933 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X934 a_n6313_n5010# bias_c a_n1110_n5852# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X935 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X936 sc_cmfb_0/transmission_gate_8/out p1 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X937 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X938 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X939 a_n5580_n13620# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X940 sc_cmfb_0/transmission_gate_6/in sc_cmfb_0/transmission_gate_8/in sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X941 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X942 cm p1_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X943 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X944 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X945 VDD VDD on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X946 sc_cmfb_0/transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X947 i_bias i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X948 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X949 sc_cmfb_0/transmission_gate_6/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X950 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X951 VSS VSS a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X952 a_n5580_n13620# a_n5580_n13620# a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X953 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X954 a_n2185_n13400# a_n2185_n13400# a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X955 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X956 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X957 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X958 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X959 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X960 sc_cmfb_0/transmission_gate_8/out p1_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X961 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X962 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X963 a_n1651_n11400# VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X964 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X965 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X966 op sc_cmfb_0/transmission_gate_8/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X967 a_n5928_n13620# bias_c op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X968 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X969 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X970 VSS i_bias bias_c VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X971 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X972 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X973 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X974 bias_c i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X975 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X976 sc_cmfb_0/transmission_gate_8/in p1 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X977 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X978 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X979 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X980 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X981 op p1 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X982 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X983 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X984 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X985 a_n2185_n13400# a_n2185_n13400# a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X986 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X987 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X988 a_n6313_n3270# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X989 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X990 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X991 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X992 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X993 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X994 sc_cmfb_0/transmission_gate_8/in p1_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X995 sc_cmfb_0/transmission_gate_5/in p1 sc_cmfb_0/transmission_gate_8/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X996 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X997 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X998 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X999 op p1_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1000 sc_cmfb_0/transmission_gate_4/out p1 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1001 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1002 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1003 op VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1004 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1005 sc_cmfb_0/transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1006 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1007 cm p2_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1008 sc_cmfb_0/transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1009 op VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1010 a_n5928_n12940# bias_c on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1011 sc_cmfb_0/transmission_gate_6/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1012 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1013 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1014 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1015 c1_7402_n7169# m3_7302_n7269# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X1016 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1017 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1018 on p2_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1019 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1020 a_n6313_n4140# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1021 sc_cmfb_0/transmission_gate_8/out p2_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1022 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1023 sc_cmfb_0/transmission_gate_8/out p1 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1024 cm p2_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1025 a_n5928_n12940# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1026 sc_cmfb_0/transmission_gate_7/in p1 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1027 bias_b bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1028 a_n1651_n11400# bias_d op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1029 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1030 sc_cmfb_0/transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1031 a_n6313_n3270# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1032 cm p2_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1033 a_n2185_n13400# a_n2185_n13400# a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1034 on p1 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1035 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1036 cm p2_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1037 sc_cmfb_0/transmission_gate_8/in p1 sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1038 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1039 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1040 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1041 a_n1651_n11400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1042 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1043 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1044 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1045 sc_cmfb_0/transmission_gate_8/in p2_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1046 cm p2 sc_cmfb_0/transmission_gate_3/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1047 op p1 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1048 cm p2_b sc_cmfb_0/transmission_gate_4/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1049 sc_cmfb_0/transmission_gate_4/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1050 cm p1_b sc_cmfb_0/transmission_gate_6/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1051 VSS sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1052 a_n1110_n5852# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1053 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1054 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X1055 sc_cmfb_0/transmission_gate_8/in p2 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1056 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1057 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1058 sc_cmfb_0/transmission_gate_5/out p1_b sc_cmfb_0/transmission_gate_8/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1059 a_11814_n11502# cm a_11636_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1060 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1061 cm p1 sc_cmfb_0/transmission_gate_6/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1062 VSS sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1063 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_5/out sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
X1064 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1065 a_12398_n11502# cm VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1066 bias_b bias_b bias_c VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1067 a_11230_n9962# cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1068 on bias_c a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1069 sc_cmfb_0/transmission_gate_5/out p1 sc_cmfb_0/transmission_gate_8/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1070 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1071 sc_cmfb_0/transmission_gate_5/in p2_b sc_cmfb_0/transmission_gate_5/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1072 a_n5928_n13620# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1073 sc_cmfb_0/transmission_gate_7/in p1_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1074 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1075 cm cm cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1076 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1077 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1078 a_n2185_n13400# bias_d sc_cmfb_0/transmission_gate_5/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1079 sc_cmfb_0/transmission_gate_5/in p2 sc_cmfb_0/transmission_gate_5/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1080 a_n5928_n12940# a_n5928_n12940# a_n5928_n12940# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1081 on p1_b sc_cmfb_0/transmission_gate_3/out VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1082 a_n5580_n13620# sc_cmfb_0/transmission_gate_8/out VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1083 sc_cmfb_0/transmission_gate_6/in p2_b op VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1084 sc_cmfb_0/transmission_gate_3/out p2_b cm VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1085 a_n2185_n13400# a_n2185_n13400# a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1086 i_bias i_bias VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1087 VSS i_bias i_bias VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1088 sc_cmfb_0/transmission_gate_6/in p2 op VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1089 sc_cmfb_0/transmission_gate_4/out p2 cm VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1090 cm p2 sc_cmfb_0/transmission_gate_4/out VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1091 sc_cmfb_0/transmission_gate_8/out p2_b sc_cmfb_0/transmission_gate_8/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1092 bias_c bias_b bias_b VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1093 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1094 a_n1651_n13400# sc_cmfb_0/transmission_gate_5/in VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1095 VSS sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1096 on bias_d a_n1651_n13400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1097 a_n5928_n13620# bias_b VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1098 a_n6313_n5010# bias_c a_n1110_n5852# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1099 cm p1_b sc_cmfb_0/transmission_gate_7/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1100 a_n1110_n5852# a_n1110_n5852# bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1101 on p2 sc_cmfb_0/transmission_gate_7/in VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1102 bias_d a_n1110_n5852# a_n1110_n5852# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1103 bias_d bias_d bias_d VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X1104 sc_cmfb_0/transmission_gate_5/out p2_b sc_cmfb_0/transmission_gate_5/in VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1105 sc_cmfb_0/transmission_gate_3/out p1_b on VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X1106 VSS sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 c1_7402_31# sc_cmfb_0/transmission_gate_7/in 0.07fF
C1 sc_cmfb_0/transmission_gate_8/out sc_cmfb_0/transmission_gate_6/in 1.36fF
C2 sc_cmfb_0/transmission_gate_8/out m3_10902_n7269# 0.10fF
C3 a_n6313_n4140# cm 3.49fF
C4 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_8/in 6.67fF
C5 on cm 1.32fF
C6 c1_7402_n1769# c1_7402_31# 0.06fF
C7 a_11814_n11502# a_11230_n11502# 0.10fF
C8 m3_9102_1731# sc_cmfb_0/transmission_gate_6/in 0.39fF
C9 m3_7302_n7269# m3_7302_n5469# 0.10fF
C10 m3_7302_n3669# m3_7302_n5469# 0.10fF
C11 a_11522_n9962# a_11814_n9962# 0.22fF
C12 VDD op 9.84fF
C13 c1_7402_n7169# c1_7402_n5369# 0.06fF
C14 m3_16302_n3669# sc_cmfb_0/transmission_gate_6/in 0.79fF
C15 m3_9102_n7269# op 0.02fF
C16 p1 on 0.78fF
C17 c1_12802_1831# c1_14602_1831# 0.06fF
C18 sc_cmfb_0/transmission_gate_5/in m3_16302_1731# 0.99fF
C19 on a_n5580_n13620# 0.06fF
C20 sc_cmfb_0/transmission_gate_5/out cm 0.04fF
C21 bias_d on 14.35fF
C22 sc_cmfb_0/transmission_gate_8/out cm 0.85fF
C23 c1_11002_1831# c1_9202_1831# 0.06fF
C24 m3_10902_n7269# c1_11002_n7169# 2.67fF
C25 a_11522_n9962# a_12398_n9962# 0.07fF
C26 on m3_7302_n69# 0.87fF
C27 sc_cmfb_0/transmission_gate_4/out p1_b 1.18fF
C28 m3_7302_1731# c1_7402_1831# 2.73fF
C29 cm a_11814_n9962# 1.34fF
C30 a_11052_n10732# a_12220_n10732# 0.05fF
C31 bias_c op 5.28fF
C32 p1 sc_cmfb_0/transmission_gate_5/out 1.30fF
C33 a_11344_n10732# a_11052_n10732# 0.22fF
C34 m3_16302_n3669# cm 1.04fF
C35 sc_cmfb_0/transmission_gate_6/in p1_b 0.45fF
C36 m3_16302_n1869# cm 1.04fF
C37 p1 sc_cmfb_0/transmission_gate_8/out 0.60fF
C38 a_n2185_n13400# a_n1651_n11400# 11.80fF
C39 a_11814_n11502# cm 0.76fF
C40 sc_cmfb_0/transmission_gate_8/out a_n5580_n13620# 55.25fF
C41 m3_16302_n69# m3_16302_1731# 0.10fF
C42 bias_d sc_cmfb_0/transmission_gate_8/out 0.03fF
C43 a_12106_n11502# a_11928_n10732# 0.13fF
C44 a_11344_n10732# a_12220_n10732# 0.07fF
C45 a_12398_n9962# cm 1.57fF
C46 p1 m3_16302_n3669# 0.76fF
C47 i_bias ip 0.16fF
C48 sc_cmfb_0/transmission_gate_5/in a_n2185_n13400# 28.09fF
C49 p2 sc_cmfb_0/transmission_gate_7/in 1.30fF
C50 a_n6313_n3270# a_n6313_n5010# 4.77fF
C51 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_7/in 0.28fF
C52 p2_b p2 3.35fF
C53 cm p1_b 2.76fF
C54 a_n5928_n13620# i_bias 0.24fF
C55 m3_16302_n7269# p1_b 0.76fF
C56 sc_cmfb_0/transmission_gate_3/out p2_b 0.41fF
C57 a_n5928_n13620# a_n6313_n3270# 3.86fF
C58 m3_16302_n5469# sc_cmfb_0/transmission_gate_8/in 0.10fF
C59 c1_16402_31# c1_16402_n1769# 0.06fF
C60 a_11636_n10732# a_11814_n9962# 0.13fF
C61 in a_n5928_n12940# 1.60fF
C62 a_n2185_n13400# a_n1651_n13400# 12.32fF
C63 c1_11002_n7169# c1_12802_n7169# 0.06fF
C64 p1 p1_b 3.34fF
C65 a_11814_n11502# a_11636_n10732# 0.13fF
C66 a_12106_n11502# a_11230_n11502# 0.07fF
C67 a_11636_n10732# a_12398_n9962# 0.03fF
C68 sc_cmfb_0/transmission_gate_5/in a_n1110_n5852# 3.34fF
C69 on sc_cmfb_0/transmission_gate_7/in 9.74fF
C70 a_n6313_n4140# a_n6313_n3270# 0.56fF
C71 a_11052_n10732# a_11230_n9962# 0.13fF
C72 on a_n6313_n3270# 0.09fF
C73 sc_cmfb_0/transmission_gate_5/in a_n5928_n12940# 0.07fF
C74 on p2_b 0.52fF
C75 on c1_7402_n1769# 0.06fF
C76 m3_12702_1731# m3_14502_1731# 0.10fF
C77 a_11814_n11502# a_11522_n11502# 0.22fF
C78 VDD a_n6313_n5010# 10.33fF
C79 a_11230_n9962# a_12220_n10732# 0.02fF
C80 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_5/in 0.09fF
C81 VDD p2 0.40fF
C82 a_11344_n10732# a_11230_n9962# 0.25fF
C83 sc_cmfb_0/transmission_gate_5/out sc_cmfb_0/transmission_gate_7/in 0.02fF
C84 c1_7402_n1769# c1_7402_n3569# 0.06fF
C85 sc_cmfb_0/transmission_gate_8/out sc_cmfb_0/transmission_gate_7/in 0.06fF
C86 sc_cmfb_0/transmission_gate_3/out VDD 2.40fF
C87 a_n5928_n13620# VDD 22.54fF
C88 m3_7302_n1869# p2 0.76fF
C89 p2_b sc_cmfb_0/transmission_gate_5/out 0.44fF
C90 a_12106_n11502# cm 0.80fF
C91 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_6/in 0.05fF
C92 a_11052_n10732# a_12106_n9962# 0.02fF
C93 p2_b sc_cmfb_0/transmission_gate_8/out 0.45fF
C94 bias_b a_n1110_n5852# 0.39fF
C95 c1_7402_n5369# op 0.12fF
C96 a_12106_n9962# a_12220_n10732# 0.25fF
C97 op c1_16402_n1769# 0.06fF
C98 bias_b a_n5928_n12940# 10.81fF
C99 bias_c ip 0.11fF
C100 a_11344_n10732# a_12106_n9962# 0.03fF
C101 a_n5580_n13620# in 2.12fF
C102 bias_c a_n6313_n5010# 4.41fF
C103 p2_b m3_16302_n1869# 0.81fF
C104 sc_cmfb_0/transmission_gate_4/out m3_16302_n69# 0.77fF
C105 a_11814_n11502# a_12398_n11502# 0.10fF
C106 bias_c a_n5928_n13620# 8.60fF
C107 sc_cmfb_0/transmission_gate_5/in cm 1.53fF
C108 sc_cmfb_0/transmission_gate_4/out c1_9202_n7169# 0.06fF
C109 sc_cmfb_0/transmission_gate_5/in m3_16302_n7269# 0.99fF
C110 p1 m3_7302_n5469# 0.78fF
C111 a_n5580_n13620# a_n1651_n11400# 0.14fF
C112 a_12398_n9962# a_12398_n11502# 0.01fF
C113 m3_14502_1731# c1_14602_1831# 2.67fF
C114 bias_d a_n1651_n11400# 12.56fF
C115 a_n6313_n4140# VDD 6.60fF
C116 c1_9202_1831# sc_cmfb_0/transmission_gate_7/in 0.06fF
C117 on VDD 9.91fF
C118 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_8/in 0.23fF
C119 sc_cmfb_0/transmission_gate_7/in p1_b 0.44fF
C120 m3_16302_n5469# c1_16402_n5369# 2.66fF
C121 a_12106_n11502# a_11636_n10732# 0.04fF
C122 op a_n6313_n5010# 0.28fF
C123 p1 sc_cmfb_0/transmission_gate_5/in 1.41fF
C124 on c1_12802_1831# 0.06fF
C125 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/transmission_gate_6/in 6.06fF
C126 p2_b p1_b 0.01fF
C127 p2 op 0.60fF
C128 sc_cmfb_0/transmission_gate_5/in a_n5580_n13620# 21.74fF
C129 sc_cmfb_0/transmission_gate_3/out op 0.44fF
C130 a_n5928_n13620# op 7.39fF
C131 bias_d sc_cmfb_0/transmission_gate_5/in 9.24fF
C132 c1_16402_n5369# c1_16402_n3569# 0.06fF
C133 m3_16302_n69# cm 1.01fF
C134 sc_cmfb_0/transmission_gate_5/out VDD 2.30fF
C135 sc_cmfb_0/transmission_gate_4/out m3_7302_n7269# 0.89fF
C136 sc_cmfb_0/transmission_gate_8/out VDD 2.59fF
C137 m3_9102_n7269# sc_cmfb_0/transmission_gate_5/out 0.10fF
C138 sc_cmfb_0/transmission_gate_8/out m3_12702_1731# 0.10fF
C139 bias_c a_n6313_n4140# 3.58fF
C140 bias_b cm 0.36fF
C141 bias_c on 4.90fF
C142 sc_cmfb_0/transmission_gate_8/out m3_7302_n1869# 0.97fF
C143 a_n5580_n13620# a_n1651_n13400# 0.13fF
C144 m3_7302_1731# sc_cmfb_0/transmission_gate_6/in 0.95fF
C145 bias_d a_n1651_n13400# 16.52fF
C146 a_12106_n11502# a_11522_n11502# 0.10fF
C147 a_n1110_n5852# a_n2185_n13400# 0.00fF
C148 sc_cmfb_0/transmission_gate_8/in cm 0.07fF
C149 m3_16302_n3669# VDD 0.33fF
C150 sc_cmfb_0/transmission_gate_8/in m3_16302_n7269# 0.76fF
C151 VDD m3_16302_n1869# 0.34fF
C152 bias_b a_n5580_n13620# 0.11fF
C153 a_n2185_n13400# a_n5928_n12940# 0.11fF
C154 a_11230_n9962# a_12106_n9962# 0.07fF
C155 a_n6313_n4140# op 0.48fF
C156 bias_c sc_cmfb_0/transmission_gate_8/out 0.07fF
C157 on op 10.51fF
C158 p1 sc_cmfb_0/transmission_gate_8/in 0.58fF
C159 m3_16302_n5469# cm 1.04fF
C160 m3_16302_n5469# m3_16302_n7269# 0.10fF
C161 a_11052_n10732# a_11814_n9962# 0.03fF
C162 i_bias in 0.28fF
C163 VDD p1_b 7.40fF
C164 sc_cmfb_0/transmission_gate_8/in m3_7302_n69# 0.10fF
C165 op c1_7402_n3569# 0.07fF
C166 a_12106_n11502# a_12398_n11502# 0.22fF
C167 a_11928_n10732# a_11230_n11502# 0.03fF
C168 m3_12702_n7269# m3_10902_n7269# 0.10fF
C169 sc_cmfb_0/transmission_gate_5/out op 0.66fF
C170 p1 m3_7302_n7269# 0.82fF
C171 p1 m3_7302_n3669# 0.71fF
C172 a_11814_n11502# a_11052_n10732# 0.03fF
C173 sc_cmfb_0/transmission_gate_8/out op 17.23fF
C174 a_12220_n10732# a_11814_n9962# 0.05fF
C175 p1 m3_16302_n5469# 0.98fF
C176 a_11344_n10732# a_11814_n9962# 0.04fF
C177 m3_9102_1731# op 0.65fF
C178 a_n1110_n5852# a_n5928_n12940# 0.47fF
C179 a_11052_n10732# a_12398_n9962# 0.01fF
C180 a_11814_n11502# a_12220_n10732# 0.05fF
C181 m3_7302_1731# m3_7302_n69# 0.10fF
C182 a_11522_n9962# a_11928_n10732# 0.05fF
C183 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_7/in 0.09fF
C184 a_11814_n11502# a_11344_n10732# 0.04fF
C185 sc_cmfb_0/transmission_gate_4/out a_n1110_n5852# 0.01fF
C186 a_12398_n9962# a_12220_n10732# 0.13fF
C187 sc_cmfb_0/transmission_gate_5/in p2_b 1.25fF
C188 a_11344_n10732# a_12398_n9962# 0.02fF
C189 a_11928_n10732# cm 0.78fF
C190 c1_11002_1831# m3_10902_1731# 2.67fF
C191 a_n5580_n13620# a_n2185_n13400# 0.56fF
C192 bias_d a_n2185_n13400# 8.57fF
C193 a_n5928_n13620# ip 1.07fF
C194 op p1_b 0.52fF
C195 c1_7402_n7169# c1_9202_n7169# 0.06fF
C196 sc_cmfb_0/transmission_gate_6/in m3_10902_1731# 0.34fF
C197 m3_12702_n7269# c1_12802_n7169# 2.67fF
C198 a_n5928_n13620# a_n6313_n5010# 3.30fF
C199 m3_16302_n69# p2_b 0.91fF
C200 sc_cmfb_0/transmission_gate_3/out p2 0.59fF
C201 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_6/in 0.46fF
C202 bias_b a_n6313_n3270# 8.13fF
C203 a_n1110_n5852# cm 4.14fF
C204 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/transmission_gate_7/in 7.00fF
C205 VDD m3_7302_n5469# 0.33fF
C206 c1_7402_n5369# c1_7402_n3569# 0.06fF
C207 cm a_n5928_n12940# 1.56fF
C208 p2_b sc_cmfb_0/transmission_gate_8/in 1.17fF
C209 a_11230_n9962# a_11814_n9962# 0.10fF
C210 m3_7302_n7269# c1_7402_n7169# 2.73fF
C211 cm a_11230_n11502# 0.84fF
C212 bias_c in 0.43fF
C213 a_n5580_n13620# a_n1110_n5852# 0.08fF
C214 sc_cmfb_0/transmission_gate_5/in VDD 2.42fF
C215 a_11636_n10732# a_11928_n10732# 0.22fF
C216 sc_cmfb_0/transmission_gate_4/out cm 6.70fF
C217 bias_d a_n1110_n5852# 47.63fF
C218 a_n6313_n4140# a_n6313_n5010# 0.57fF
C219 a_12106_n11502# a_11052_n10732# 0.02fF
C220 on a_n6313_n5010# 0.42fF
C221 p2_b m3_16302_1731# 0.95fF
C222 a_n5580_n13620# a_n5928_n12940# 4.14fF
C223 m3_16302_n5469# sc_cmfb_0/transmission_gate_7/in 0.80fF
C224 sc_cmfb_0/transmission_gate_6/in cm 6.81fF
C225 on p2 0.83fF
C226 m3_16302_1731# c1_16402_1831# 2.73fF
C227 m3_16302_n69# c1_16402_31# 2.66fF
C228 m3_7302_1731# p2_b 0.91fF
C229 a_n5928_n13620# a_n6313_n4140# 4.04fF
C230 on sc_cmfb_0/transmission_gate_3/out 7.10fF
C231 a_12398_n9962# a_11230_n9962# 0.05fF
C232 a_11522_n9962# cm 1.35fF
C233 a_n5928_n13620# on 0.58fF
C234 m3_16302_n1869# c1_16402_n1769# 2.67fF
C235 a_12106_n9962# a_11814_n9962# 0.22fF
C236 p1 sc_cmfb_0/transmission_gate_4/out 1.32fF
C237 sc_cmfb_0/transmission_gate_5/out m3_14502_1731# 0.36fF
C238 a_12106_n11502# a_12220_n10732# 0.25fF
C239 a_11344_n10732# a_12106_n11502# 0.03fF
C240 p1 sc_cmfb_0/transmission_gate_6/in 0.56fF
C241 m3_16302_n69# VDD 0.33fF
C242 bias_c sc_cmfb_0/transmission_gate_5/in 0.00fF
C243 a_11928_n10732# a_11522_n11502# 0.05fF
C244 sc_cmfb_0/transmission_gate_5/out p2 0.58fF
C245 sc_cmfb_0/transmission_gate_8/out p2 1.11fF
C246 bias_b VDD 58.37fF
C247 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_5/out 8.24fF
C248 a_n1651_n11400# op 14.58fF
C249 a_12398_n9962# a_12106_n9962# 0.22fF
C250 a_11636_n10732# a_11230_n11502# 0.05fF
C251 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_8/out 1.22fF
C252 a_n5928_n13620# sc_cmfb_0/transmission_gate_8/out 0.14fF
C253 m3_9102_n7269# c1_9202_n7169# 2.59fF
C254 sc_cmfb_0/transmission_gate_8/in VDD 2.30fF
C255 on a_n6313_n4140# 0.39fF
C256 m3_16302_n1869# p2 0.96fF
C257 sc_cmfb_0/transmission_gate_8/in m3_7302_n1869# 0.91fF
C258 sc_cmfb_0/transmission_gate_5/in op 2.59fF
C259 sc_cmfb_0/transmission_gate_3/out m3_16302_n1869# 0.79fF
C260 p1 cm 2.90fF
C261 a_11522_n9962# a_11636_n10732# 0.25fF
C262 p1 m3_16302_n7269# 0.99fF
C263 a_n5580_n13620# cm 0.02fF
C264 bias_d cm 0.08fF
C265 bias_c bias_b 38.50fF
C266 VDD m3_16302_1731# 0.36fF
C267 m3_7302_n7269# VDD 0.31fF
C268 a_11522_n11502# a_11230_n11502# 0.22fF
C269 VDD m3_7302_n3669# 0.33fF
C270 a_11928_n10732# a_12398_n11502# 0.04fF
C271 m3_7302_1731# VDD 0.35fF
C272 m3_7302_n7269# m3_9102_n7269# 0.10fF
C273 a_n1651_n13400# op 2.21fF
C274 m3_16302_n5469# VDD 0.33fF
C275 m3_7302_n1869# m3_7302_n3669# 0.10fF
C276 on sc_cmfb_0/transmission_gate_5/out 1.21fF
C277 on sc_cmfb_0/transmission_gate_8/out 14.75fF
C278 p2 p1_b 0.24fF
C279 a_11636_n10732# cm 0.77fF
C280 sc_cmfb_0/transmission_gate_3/out p1_b 1.27fF
C281 c1_16402_n5369# sc_cmfb_0/transmission_gate_7/in 0.06fF
C282 a_11522_n9962# a_11522_n11502# 0.01fF
C283 a_n6313_n3270# a_n1110_n5852# 0.36fF
C284 bias_b op 0.30fF
C285 c1_14602_n7169# c1_12802_n7169# 0.06fF
C286 c1_9202_n7169# op 0.05fF
C287 i_bias a_n5928_n12940# 0.27fF
C288 a_n6313_n3270# a_n5928_n12940# 4.16fF
C289 sc_cmfb_0/transmission_gate_8/out sc_cmfb_0/transmission_gate_5/out 12.80fF
C290 sc_cmfb_0/transmission_gate_8/in op 0.85fF
C291 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_7/in 0.61fF
C292 a_12398_n11502# a_11230_n11502# 0.05fF
C293 on c1_11002_n7169# 0.06fF
C294 sc_cmfb_0/transmission_gate_4/out p2_b 0.44fF
C295 a_11522_n11502# cm 0.77fF
C296 c1_7402_n5369# m3_7302_n5469# 2.67fF
C297 c1_7402_1831# c1_7402_31# 0.06fF
C298 sc_cmfb_0/transmission_gate_6/in sc_cmfb_0/transmission_gate_7/in 0.44fF
C299 a_12106_n11502# a_12106_n9962# 0.01fF
C300 sc_cmfb_0/transmission_gate_8/out m3_16302_n3669# 0.10fF
C301 sc_cmfb_0/transmission_gate_8/out m3_16302_n1869# 0.10fF
C302 p2_b sc_cmfb_0/transmission_gate_6/in 1.21fF
C303 m3_7302_n7269# op 0.79fF
C304 on p1_b 0.53fF
C305 m3_7302_1731# op 0.93fF
C306 ip in 3.10fF
C307 a_11814_n11502# a_11814_n9962# 0.01fF
C308 m3_16302_n3669# m3_16302_n1869# 0.10fF
C309 bias_c a_n2185_n13400# 0.02fF
C310 a_12398_n9962# a_11814_n9962# 0.10fF
C311 cm sc_cmfb_0/transmission_gate_7/in 6.77fF
C312 a_n5928_n13620# in 3.26fF
C313 sc_cmfb_0/transmission_gate_5/out p1_b 1.19fF
C314 VDD a_n1110_n5852# 4.31fF
C315 sc_cmfb_0/transmission_gate_8/out p1_b 0.73fF
C316 p2_b cm 2.54fF
C317 m3_9102_1731# c1_9202_1831# 2.67fF
C318 a_n6313_n3270# cm 0.52fF
C319 a_12398_n11502# cm 1.27fF
C320 sc_cmfb_0/transmission_gate_4/out c1_16402_31# 0.06fF
C321 a_11636_n10732# a_11522_n11502# 0.25fF
C322 VDD a_n5928_n12940# 22.70fF
C323 sc_cmfb_0/transmission_gate_3/out m3_7302_n5469# 0.92fF
C324 p1 sc_cmfb_0/transmission_gate_7/in 0.58fF
C325 a_n2185_n13400# op 2.24fF
C326 a_11052_n10732# a_11928_n10732# 0.07fF
C327 m3_16302_n3669# p1_b 0.89fF
C328 m3_12702_1731# m3_10902_1731# 0.10fF
C329 c1_16402_n7169# c1_16402_n5369# 0.06fF
C330 sc_cmfb_0/transmission_gate_5/in a_n6313_n5010# 0.11fF
C331 i_bias a_n5580_n13620# 0.12fF
C332 sc_cmfb_0/transmission_gate_4/out VDD 2.35fF
C333 sc_cmfb_0/transmission_gate_5/in p2 1.35fF
C334 c1_14602_n7169# sc_cmfb_0/transmission_gate_7/in 0.06fF
C335 sc_cmfb_0/transmission_gate_4/out m3_9102_n7269# 0.53fF
C336 a_11928_n10732# a_12220_n10732# 0.22fF
C337 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_5/in 0.05fF
C338 m3_7302_n69# sc_cmfb_0/transmission_gate_7/in 0.94fF
C339 a_n5928_n13620# sc_cmfb_0/transmission_gate_5/in 0.04fF
C340 bias_c a_n1110_n5852# 1.61fF
C341 a_11344_n10732# a_11928_n10732# 0.10fF
C342 sc_cmfb_0/transmission_gate_6/in VDD 2.45fF
C343 p2_b m3_7302_n69# 0.84fF
C344 c1_11002_1831# c1_12802_1831# 0.06fF
C345 m3_9102_n7269# m3_10902_n7269# 0.10fF
C346 bias_c a_n5928_n12940# 7.44fF
C347 a_11636_n10732# a_12398_n11502# 0.03fF
C348 on a_n1651_n11400# 2.54fF
C349 bias_b ip 0.07fF
C350 a_11052_n10732# a_11230_n11502# 0.13fF
C351 on m3_7302_n5469# 0.96fF
C352 m3_16302_n69# p2 0.98fF
C353 a_n1110_n5852# op 2.51fF
C354 bias_b a_n6313_n5010# 3.89fF
C355 sc_cmfb_0/transmission_gate_8/in m3_14502_n7269# 0.51fF
C356 sc_cmfb_0/transmission_gate_8/out in 0.04fF
C357 VDD cm 8.94fF
C358 VDD m3_16302_n7269# 0.29fF
C359 a_12220_n10732# a_11230_n11502# 0.02fF
C360 op a_n5928_n12940# 0.96fF
C361 a_n5928_n13620# bias_b 9.36fF
C362 on sc_cmfb_0/transmission_gate_5/in 4.91fF
C363 a_11344_n10732# a_11230_n11502# 0.25fF
C364 m3_10902_1731# op 0.57fF
C365 a_11522_n9962# a_11052_n10732# 0.04fF
C366 sc_cmfb_0/transmission_gate_8/in p2 1.30fF
C367 sc_cmfb_0/transmission_gate_8/out a_n1651_n11400# 0.44fF
C368 sc_cmfb_0/transmission_gate_5/out m3_7302_n5469# 0.10fF
C369 c1_16402_n3569# c1_16402_n1769# 0.06fF
C370 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_8/in 0.23fF
C371 m3_14502_1731# m3_16302_1731# 0.10fF
C372 a_11522_n11502# a_12398_n11502# 0.07fF
C373 sc_cmfb_0/transmission_gate_4/out op 7.70fF
C374 sc_cmfb_0/transmission_gate_4/out c1_14602_1831# 0.06fF
C375 c1_16402_n7169# m3_16302_n7269# 2.73fF
C376 p1 VDD 0.36fF
C377 c1_11002_1831# op 0.06fF
C378 a_n5580_n13620# VDD 0.03fF
C379 a_11522_n9962# a_12220_n10732# 0.03fF
C380 a_11814_n11502# a_12106_n11502# 0.22fF
C381 sc_cmfb_0/transmission_gate_6/in op 7.21fF
C382 on a_n1651_n13400# 14.95fF
C383 a_11522_n9962# a_11344_n10732# 0.13fF
C384 bias_c cm 3.40fF
C385 m3_16302_1731# p2 0.74fF
C386 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_5/out 6.64fF
C387 VDD m3_7302_n69# 0.33fF
C388 sc_cmfb_0/transmission_gate_5/in sc_cmfb_0/transmission_gate_8/out 24.89fF
C389 m3_7302_1731# p2 0.71fF
C390 a_11052_n10732# cm 1.30fF
C391 m3_7302_n1869# m3_7302_n69# 0.10fF
C392 a_11928_n10732# a_11230_n9962# 0.03fF
C393 bias_b a_n6313_n4140# 2.96fF
C394 bias_b on 0.10fF
C395 c1_14602_n7169# c1_16402_n7169# 0.06fF
C396 p2_b sc_cmfb_0/transmission_gate_7/in 1.19fF
C397 cm a_12220_n10732# 0.86fF
C398 bias_c a_n5580_n13620# 0.50fF
C399 a_11344_n10732# cm 0.81fF
C400 sc_cmfb_0/transmission_gate_8/out a_n1651_n13400# 0.37fF
C401 cm op 1.07fF
C402 on sc_cmfb_0/transmission_gate_8/in 0.95fF
C403 m3_16302_n69# sc_cmfb_0/transmission_gate_5/out 0.10fF
C404 m3_7302_n5469# p1_b 0.84fF
C405 a_11928_n10732# a_12106_n9962# 0.13fF
C406 m3_12702_n7269# m3_14502_n7269# 0.10fF
C407 p1 op 0.66fF
C408 a_n5580_n13620# op 0.15fF
C409 a_n5928_n13620# a_n2185_n13400# 0.09fF
C410 m3_16302_n69# m3_16302_n1869# 0.10fF
C411 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/transmission_gate_5/out 3.09fF
C412 sc_cmfb_0/transmission_gate_5/in p1_b 1.25fF
C413 a_11052_n10732# a_11636_n10732# 0.10fF
C414 a_11230_n9962# a_11230_n11502# 0.01fF
C415 op c1_12802_n7169# 0.06fF
C416 bias_d op 12.81fF
C417 c1_7402_1831# c1_9202_1831# 0.06fF
C418 sc_cmfb_0/transmission_gate_8/out sc_cmfb_0/transmission_gate_8/in 14.62fF
C419 m3_9102_1731# sc_cmfb_0/transmission_gate_8/in 0.10fF
C420 a_11636_n10732# a_12220_n10732# 0.10fF
C421 sc_cmfb_0/transmission_gate_4/out c1_7402_n5369# 0.06fF
C422 on c1_16402_n3569# 0.06fF
C423 a_11344_n10732# a_11636_n10732# 0.22fF
C424 sc_cmfb_0/transmission_gate_5/out m3_16302_1731# 0.70fF
C425 a_11522_n9962# a_11230_n9962# 0.22fF
C426 m3_7302_n3669# c1_7402_n3569# 2.67fF
C427 c1_16402_31# c1_16402_1831# 0.06fF
C428 sc_cmfb_0/transmission_gate_5/out m3_7302_n3669# 0.91fF
C429 sc_cmfb_0/transmission_gate_8/out m3_7302_n3669# 1.00fF
C430 c1_9202_n7169# c1_11002_n7169# 0.06fF
C431 VDD sc_cmfb_0/transmission_gate_7/in 2.38fF
C432 a_n1110_n5852# a_n6313_n5010# 3.78fF
C433 a_11052_n10732# a_11522_n11502# 0.04fF
C434 m3_7302_1731# m3_9102_1731# 0.10fF
C435 a_n6313_n3270# VDD 11.02fF
C436 p2_b VDD 7.65fF
C437 ip a_n5928_n12940# 1.78fF
C438 on a_n2185_n13400# 9.23fF
C439 a_n5928_n13620# a_n1110_n5852# 0.10fF
C440 p2_b m3_7302_n1869# 0.77fF
C441 c1_7402_n1769# m3_7302_n1869# 2.67fF
C442 a_n6313_n5010# a_n5928_n12940# 4.84fF
C443 a_11522_n9962# a_12106_n9962# 0.10fF
C444 m3_16302_n5469# m3_16302_n3669# 0.10fF
C445 a_11230_n9962# cm 1.45fF
C446 a_11522_n11502# a_12220_n10732# 0.03fF
C447 sc_cmfb_0/transmission_gate_8/in p1_b 0.43fF
C448 a_n5928_n13620# a_n5928_n12940# 18.48fF
C449 a_11344_n10732# a_11522_n11502# 0.13fF
C450 m3_16302_n3669# c1_16402_n3569# 2.67fF
C451 sc_cmfb_0/transmission_gate_4/out p2 0.58fF
C452 c1_7402_31# m3_7302_n69# 2.67fF
C453 bias_c i_bias 13.86fF
C454 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_3/out 0.37fF
C455 sc_cmfb_0/transmission_gate_8/out a_n2185_n13400# 1.13fF
C456 bias_c a_n6313_n3270# 2.90fF
C457 sc_cmfb_0/transmission_gate_6/in p2 1.31fF
C458 a_12106_n9962# cm 1.34fF
C459 sc_cmfb_0/transmission_gate_8/out m3_12702_n7269# 0.10fF
C460 m3_7302_n7269# p1_b 0.76fF
C461 a_11052_n10732# a_12398_n11502# 0.01fF
C462 sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_6/in 0.76fF
C463 m3_7302_n3669# p1_b 0.84fF
C464 c1_7402_n7169# op 0.05fF
C465 sc_cmfb_0/transmission_gate_5/in a_n1651_n11400# 21.11fF
C466 m3_16302_n5469# p1_b 0.91fF
C467 on a_n1110_n5852# 1.83fF
C468 a_12398_n11502# a_12220_n10732# 0.13fF
C469 op sc_cmfb_0/transmission_gate_7/in 2.61fF
C470 m3_14502_n7269# m3_16302_n7269# 0.10fF
C471 a_n6313_n4140# a_n5928_n12940# 3.31fF
C472 a_11344_n10732# a_12398_n11502# 0.02fF
C473 a_11636_n10732# a_11230_n9962# 0.05fF
C474 on a_n5928_n12940# 6.91fF
C475 p2_b op 0.59fF
C476 a_n6313_n3270# op 0.40fF
C477 cm a_n6313_n5010# 1.44fF
C478 a_11928_n10732# a_11814_n9962# 0.25fF
C479 c1_14602_1831# c1_16402_1831# 0.06fF
C480 a_n1651_n13400# a_n1651_n11400# 11.78fF
C481 cm p2 2.82fF
C482 bias_b in 0.08fF
C483 sc_cmfb_0/transmission_gate_3/out cm 6.81fF
C484 VDD m3_7302_n1869# 0.33fF
C485 a_n5928_n13620# cm 0.39fF
C486 sc_cmfb_0/transmission_gate_4/out on 2.90fF
C487 sc_cmfb_0/transmission_gate_8/out a_n1110_n5852# 0.46fF
C488 a_11814_n11502# a_11928_n10732# 0.25fF
C489 c1_12802_1831# m3_12702_1731# 2.67fF
C490 a_n5580_n13620# ip 1.09fF
C491 on sc_cmfb_0/transmission_gate_6/in 0.39fF
C492 sc_cmfb_0/transmission_gate_5/in a_n1651_n13400# 22.42fF
C493 a_11636_n10732# a_12106_n9962# 0.04fF
C494 c1_14602_n7169# m3_14502_n7269# 2.67fF
C495 a_11928_n10732# a_12398_n9962# 0.04fF
C496 p1 p2 0.01fF
C497 sc_cmfb_0/transmission_gate_8/out a_n5928_n12940# 0.17fF
C498 p1 sc_cmfb_0/transmission_gate_3/out 1.30fF
C499 sc_cmfb_0/transmission_gate_8/out m3_10902_1731# 0.10fF
C500 a_n5928_n13620# a_n5580_n13620# 4.17fF
C501 bias_c VDD 30.03fF
C502 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_5/out 9.05fF
C503 m3_9102_1731# m3_10902_1731# 0.10fF
C504 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/transmission_gate_8/out 0.10fF
C505 p2 m3_7302_n69# 0.77fF
C506 sc_cmfb_0/transmission_gate_5/out sc_cmfb_0/transmission_gate_6/in 0.09fF
C507 i_bias VSS 33.90fF
C508 in VSS 2.99fF
C509 ip VSS 2.92fF
C510 m3_16302_n7269# VSS 0.75fF
C511 m3_14502_n7269# VSS 1.03fF
C512 m3_12702_n7269# VSS 1.07fF
C513 m3_10902_n7269# VSS 1.07fF
C514 m3_9102_n7269# VSS 1.01fF
C515 m3_7302_n7269# VSS 0.77fF
C516 m3_16302_n5469# VSS 0.70fF
C517 m3_16302_n3669# VSS 0.73fF
C518 m3_16302_n1869# VSS 0.70fF
C519 m3_7302_n5469# VSS 0.72fF
C520 m3_7302_n3669# VSS 0.73fF
C521 m3_7302_n1869# VSS 0.72fF
C522 m3_16302_n69# VSS 0.70fF
C523 m3_7302_n69# VSS 0.71fF
C524 m3_16302_1731# VSS 0.82fF
C525 m3_14502_1731# VSS 1.07fF
C526 m3_12702_1731# VSS 1.14fF
C527 m3_10902_1731# VSS 1.03fF
C528 m3_9102_1731# VSS 1.09fF
C529 m3_7302_1731# VSS 0.83fF
C530 a_n1651_n13400# VSS 29.40fF
C531 a_n1651_n11400# VSS 28.93fF
C532 a_n2185_n13400# VSS 24.97fF
C533 a_12398_n11502# VSS 0.32fF
C534 a_12106_n11502# VSS 0.57fF
C535 a_11814_n11502# VSS 0.62fF
C536 a_11522_n11502# VSS 0.65fF
C537 a_11230_n11502# VSS 0.64fF
C538 a_12220_n10732# VSS 0.12fF
C539 a_11928_n10732# VSS 0.12fF
C540 a_11636_n10732# VSS 0.14fF
C541 a_11344_n10732# VSS 0.15fF
C542 a_11052_n10732# VSS 0.16fF
C543 a_12398_n9962# VSS 0.09fF
C544 a_12106_n9962# VSS 0.11fF
C545 a_11814_n9962# VSS 0.12fF
C546 a_11522_n9962# VSS 0.15fF
C547 a_11230_n9962# VSS 0.16fF
C548 bias_d VSS 56.16fF
C549 a_n5580_n13620# VSS 110.90fF
C550 p1 VSS 11.82fF
C551 p1_b VSS 4.17fF
C552 a_n1110_n5852# VSS 23.20fF
C553 a_n6313_n5010# VSS 0.00fF
C554 bias_c VSS 18.47fF
C555 a_n6313_n3270# VSS 0.00fF
C556 a_n5928_n12940# VSS 4.89fF
C557 a_n5928_n13620# VSS 4.17fF
C558 bias_b VSS 19.59fF
C559 sc_cmfb_0/transmission_gate_3/out VSS 5.11fF
C560 sc_cmfb_0/transmission_gate_8/in VSS 10.71fF
C561 sc_cmfb_0/transmission_gate_8/out VSS 114.94fF
C562 cm VSS 24.55fF
C563 sc_cmfb_0/transmission_gate_4/out VSS 4.52fF
C564 sc_cmfb_0/transmission_gate_7/in VSS 4.36fF
C565 on VSS 25.08fF
C566 p2 VSS 11.67fF
C567 sc_cmfb_0/transmission_gate_5/in VSS 180.33fF
C568 sc_cmfb_0/transmission_gate_5/out VSS 11.54fF
C569 p2_b VSS 4.27fF
C570 sc_cmfb_0/transmission_gate_6/in VSS 6.83fF
C571 op VSS 27.64fF
C572 VDD VSS 253.65fF
.ends

