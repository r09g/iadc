magic
tech sky130A
magscale 1 2
timestamp 1653544574
<< nwell >>
rect -7664 -7309 3823 -1120
<< pwell >>
rect -7664 -17642 13838 -7439
<< nmos >>
rect -2127 -8400 -2007 -8120
rect -1949 -8400 -1829 -8120
rect -1771 -8400 -1651 -8120
rect -1593 -8400 -1473 -8120
rect -1415 -8400 -1295 -8120
rect -1237 -8400 -1117 -8120
rect -1059 -8400 -939 -8120
rect -881 -8400 -761 -8120
rect -703 -8400 -583 -8120
rect -525 -8400 -405 -8120
rect -347 -8400 -227 -8120
rect -169 -8400 -49 -8120
rect 9 -8400 129 -8120
rect 187 -8400 307 -8120
rect 365 -8400 485 -8120
rect 543 -8400 663 -8120
rect 721 -8400 841 -8120
rect 899 -8400 1019 -8120
rect 1077 -8400 1197 -8120
rect 1255 -8400 1375 -8120
rect 1433 -8400 1553 -8120
rect 1611 -8400 1731 -8120
rect 1789 -8400 1909 -8120
rect 1967 -8400 2087 -8120
rect 2145 -8400 2265 -8120
rect 2323 -8400 2443 -8120
rect 2501 -8400 2621 -8120
rect 2679 -8400 2799 -8120
rect 2857 -8400 2977 -8120
rect 3035 -8400 3155 -8120
rect 3213 -8400 3333 -8120
rect 3391 -8400 3511 -8120
rect 3569 -8400 3689 -8120
rect 3747 -8400 3867 -8120
rect 3925 -8400 4045 -8120
rect -2127 -9400 -2007 -9120
rect -1949 -9400 -1829 -9120
rect -1771 -9400 -1651 -9120
rect -1593 -9400 -1473 -9120
rect -1415 -9400 -1295 -9120
rect -1237 -9400 -1117 -9120
rect -1059 -9400 -939 -9120
rect -881 -9400 -761 -9120
rect -703 -9400 -583 -9120
rect -525 -9400 -405 -9120
rect -347 -9400 -227 -9120
rect -169 -9400 -49 -9120
rect 9 -9400 129 -9120
rect 187 -9400 307 -9120
rect 365 -9400 485 -9120
rect 543 -9400 663 -9120
rect 721 -9400 841 -9120
rect 899 -9400 1019 -9120
rect 1077 -9400 1197 -9120
rect 1255 -9400 1375 -9120
rect 1433 -9400 1553 -9120
rect 1611 -9400 1731 -9120
rect 1789 -9400 1909 -9120
rect 1967 -9400 2087 -9120
rect 2145 -9400 2265 -9120
rect 2323 -9400 2443 -9120
rect 2501 -9400 2621 -9120
rect 2679 -9400 2799 -9120
rect 2857 -9400 2977 -9120
rect 3035 -9400 3155 -9120
rect 3213 -9400 3333 -9120
rect 3391 -9400 3511 -9120
rect 3569 -9400 3689 -9120
rect 3747 -9400 3867 -9120
rect 3925 -9400 4045 -9120
rect 6558 -9162 6678 -8882
rect 6736 -9162 6856 -8882
rect 6914 -9162 7034 -8882
rect 7092 -9162 7212 -8882
rect 7270 -9162 7390 -8882
rect 7448 -9162 7568 -8882
rect 7626 -9162 7746 -8882
rect 7804 -9162 7924 -8882
rect 7982 -9162 8102 -8882
rect 8160 -9162 8280 -8882
rect 8338 -9162 8458 -8882
rect 8516 -9162 8636 -8882
rect 8694 -9162 8814 -8882
rect 8872 -9162 8992 -8882
rect 9050 -9162 9170 -8882
rect 9228 -9162 9348 -8882
rect 10818 -9192 10938 -8912
rect 11110 -9192 11230 -8912
rect 11402 -9192 11522 -8912
rect 11694 -9192 11814 -8912
rect 11986 -9192 12106 -8912
rect 12278 -9192 12398 -8912
rect 12570 -9192 12690 -8912
rect 6558 -10062 6678 -9782
rect 6736 -10062 6856 -9782
rect 6914 -10062 7034 -9782
rect 7092 -10062 7212 -9782
rect 7270 -10062 7390 -9782
rect 7448 -10062 7568 -9782
rect 7626 -10062 7746 -9782
rect 7804 -10062 7924 -9782
rect 7982 -10062 8102 -9782
rect 8160 -10062 8280 -9782
rect 8338 -10062 8458 -9782
rect 8516 -10062 8636 -9782
rect 8694 -10062 8814 -9782
rect 8872 -10062 8992 -9782
rect 9050 -10062 9170 -9782
rect 9228 -10062 9348 -9782
rect 10818 -9962 10938 -9682
rect 11110 -9962 11230 -9682
rect 11402 -9962 11522 -9682
rect 11694 -9962 11814 -9682
rect 11986 -9962 12106 -9682
rect 12278 -9962 12398 -9682
rect 12570 -9962 12690 -9682
rect -2127 -10400 -2007 -10120
rect -1949 -10400 -1829 -10120
rect -1771 -10400 -1651 -10120
rect -1593 -10400 -1473 -10120
rect -1415 -10400 -1295 -10120
rect -1237 -10400 -1117 -10120
rect -1059 -10400 -939 -10120
rect -881 -10400 -761 -10120
rect -703 -10400 -583 -10120
rect -525 -10400 -405 -10120
rect -347 -10400 -227 -10120
rect -169 -10400 -49 -10120
rect 9 -10400 129 -10120
rect 187 -10400 307 -10120
rect 365 -10400 485 -10120
rect 543 -10400 663 -10120
rect 721 -10400 841 -10120
rect 899 -10400 1019 -10120
rect 1077 -10400 1197 -10120
rect 1255 -10400 1375 -10120
rect 1433 -10400 1553 -10120
rect 1611 -10400 1731 -10120
rect 1789 -10400 1909 -10120
rect 1967 -10400 2087 -10120
rect 2145 -10400 2265 -10120
rect 2323 -10400 2443 -10120
rect 2501 -10400 2621 -10120
rect 2679 -10400 2799 -10120
rect 2857 -10400 2977 -10120
rect 3035 -10400 3155 -10120
rect 3213 -10400 3333 -10120
rect 3391 -10400 3511 -10120
rect 3569 -10400 3689 -10120
rect 3747 -10400 3867 -10120
rect 3925 -10400 4045 -10120
rect 6558 -10962 6678 -10682
rect 6736 -10962 6856 -10682
rect 6914 -10962 7034 -10682
rect 7092 -10962 7212 -10682
rect 7270 -10962 7390 -10682
rect 7448 -10962 7568 -10682
rect 7626 -10962 7746 -10682
rect 7804 -10962 7924 -10682
rect 7982 -10962 8102 -10682
rect 8160 -10962 8280 -10682
rect 8338 -10962 8458 -10682
rect 8516 -10962 8636 -10682
rect 8694 -10962 8814 -10682
rect 8872 -10962 8992 -10682
rect 9050 -10962 9170 -10682
rect 9228 -10962 9348 -10682
rect 10818 -10732 10938 -10452
rect 11110 -10732 11230 -10452
rect 11402 -10732 11522 -10452
rect 11694 -10732 11814 -10452
rect 11986 -10732 12106 -10452
rect 12278 -10732 12398 -10452
rect 12570 -10732 12690 -10452
rect -2127 -11400 -2007 -11120
rect -1949 -11400 -1829 -11120
rect -1771 -11400 -1651 -11120
rect -1593 -11400 -1473 -11120
rect -1415 -11400 -1295 -11120
rect -1237 -11400 -1117 -11120
rect -1059 -11400 -939 -11120
rect -881 -11400 -761 -11120
rect -703 -11400 -583 -11120
rect -525 -11400 -405 -11120
rect -347 -11400 -227 -11120
rect -169 -11400 -49 -11120
rect 9 -11400 129 -11120
rect 187 -11400 307 -11120
rect 365 -11400 485 -11120
rect 543 -11400 663 -11120
rect 721 -11400 841 -11120
rect 899 -11400 1019 -11120
rect 1077 -11400 1197 -11120
rect 1255 -11400 1375 -11120
rect 1433 -11400 1553 -11120
rect 1611 -11400 1731 -11120
rect 1789 -11400 1909 -11120
rect 1967 -11400 2087 -11120
rect 2145 -11400 2265 -11120
rect 2323 -11400 2443 -11120
rect 2501 -11400 2621 -11120
rect 2679 -11400 2799 -11120
rect 2857 -11400 2977 -11120
rect 3035 -11400 3155 -11120
rect 3213 -11400 3333 -11120
rect 3391 -11400 3511 -11120
rect 3569 -11400 3689 -11120
rect 3747 -11400 3867 -11120
rect 3925 -11400 4045 -11120
rect 10818 -11502 10938 -11222
rect 11110 -11502 11230 -11222
rect 11402 -11502 11522 -11222
rect 11694 -11502 11814 -11222
rect 11986 -11502 12106 -11222
rect 12278 -11502 12398 -11222
rect 12570 -11502 12690 -11222
rect 6558 -11862 6678 -11582
rect 6736 -11862 6856 -11582
rect 6914 -11862 7034 -11582
rect 7092 -11862 7212 -11582
rect 7270 -11862 7390 -11582
rect 7448 -11862 7568 -11582
rect 7626 -11862 7746 -11582
rect 7804 -11862 7924 -11582
rect 7982 -11862 8102 -11582
rect 8160 -11862 8280 -11582
rect 8338 -11862 8458 -11582
rect 8516 -11862 8636 -11582
rect 8694 -11862 8814 -11582
rect 8872 -11862 8992 -11582
rect 9050 -11862 9170 -11582
rect 9228 -11862 9348 -11582
rect -2127 -12400 -2007 -12120
rect -1949 -12400 -1829 -12120
rect -1771 -12400 -1651 -12120
rect -1593 -12400 -1473 -12120
rect -1415 -12400 -1295 -12120
rect -1237 -12400 -1117 -12120
rect -1059 -12400 -939 -12120
rect -881 -12400 -761 -12120
rect -703 -12400 -583 -12120
rect -525 -12400 -405 -12120
rect -347 -12400 -227 -12120
rect -169 -12400 -49 -12120
rect 9 -12400 129 -12120
rect 187 -12400 307 -12120
rect 365 -12400 485 -12120
rect 543 -12400 663 -12120
rect 721 -12400 841 -12120
rect 899 -12400 1019 -12120
rect 1077 -12400 1197 -12120
rect 1255 -12400 1375 -12120
rect 1433 -12400 1553 -12120
rect 1611 -12400 1731 -12120
rect 1789 -12400 1909 -12120
rect 1967 -12400 2087 -12120
rect 2145 -12400 2265 -12120
rect 2323 -12400 2443 -12120
rect 2501 -12400 2621 -12120
rect 2679 -12400 2799 -12120
rect 2857 -12400 2977 -12120
rect 3035 -12400 3155 -12120
rect 3213 -12400 3333 -12120
rect 3391 -12400 3511 -12120
rect 3569 -12400 3689 -12120
rect 3747 -12400 3867 -12120
rect 3925 -12400 4045 -12120
rect -2127 -13400 -2007 -13120
rect -1949 -13400 -1829 -13120
rect -1771 -13400 -1651 -13120
rect -1593 -13400 -1473 -13120
rect -1415 -13400 -1295 -13120
rect -1237 -13400 -1117 -13120
rect -1059 -13400 -939 -13120
rect -881 -13400 -761 -13120
rect -703 -13400 -583 -13120
rect -525 -13400 -405 -13120
rect -347 -13400 -227 -13120
rect -169 -13400 -49 -13120
rect 9 -13400 129 -13120
rect 187 -13400 307 -13120
rect 365 -13400 485 -13120
rect 543 -13400 663 -13120
rect 721 -13400 841 -13120
rect 899 -13400 1019 -13120
rect 1077 -13400 1197 -13120
rect 1255 -13400 1375 -13120
rect 1433 -13400 1553 -13120
rect 1611 -13400 1731 -13120
rect 1789 -13400 1909 -13120
rect 1967 -13400 2087 -13120
rect 2145 -13400 2265 -13120
rect 2323 -13400 2443 -13120
rect 2501 -13400 2621 -13120
rect 2679 -13400 2799 -13120
rect 2857 -13400 2977 -13120
rect 3035 -13400 3155 -13120
rect 3213 -13400 3333 -13120
rect 3391 -13400 3511 -13120
rect 3569 -13400 3689 -13120
rect 3747 -13400 3867 -13120
rect 3925 -13400 4045 -13120
rect -5982 -14662 -5862 -14382
rect -5804 -14662 -5684 -14382
rect -5626 -14662 -5506 -14382
rect -5448 -14662 -5328 -14382
rect -5270 -14662 -5150 -14382
rect -5092 -14662 -4972 -14382
rect -4914 -14662 -4794 -14382
rect -4736 -14662 -4616 -14382
rect -4558 -14662 -4438 -14382
rect -4380 -14662 -4260 -14382
rect -4202 -14662 -4082 -14382
rect -2127 -14400 -2007 -14120
rect -1949 -14400 -1829 -14120
rect -1771 -14400 -1651 -14120
rect -1593 -14400 -1473 -14120
rect -1415 -14400 -1295 -14120
rect -1237 -14400 -1117 -14120
rect -1059 -14400 -939 -14120
rect -881 -14400 -761 -14120
rect -703 -14400 -583 -14120
rect -525 -14400 -405 -14120
rect -347 -14400 -227 -14120
rect -169 -14400 -49 -14120
rect 9 -14400 129 -14120
rect 187 -14400 307 -14120
rect 365 -14400 485 -14120
rect 543 -14400 663 -14120
rect 721 -14400 841 -14120
rect 899 -14400 1019 -14120
rect 1077 -14400 1197 -14120
rect 1255 -14400 1375 -14120
rect 1433 -14400 1553 -14120
rect 1611 -14400 1731 -14120
rect 1789 -14400 1909 -14120
rect 1967 -14400 2087 -14120
rect 2145 -14400 2265 -14120
rect 2323 -14400 2443 -14120
rect 2501 -14400 2621 -14120
rect 2679 -14400 2799 -14120
rect 2857 -14400 2977 -14120
rect 3035 -14400 3155 -14120
rect 3213 -14400 3333 -14120
rect 3391 -14400 3511 -14120
rect 3569 -14400 3689 -14120
rect 3747 -14400 3867 -14120
rect 3925 -14400 4045 -14120
rect 5623 -14400 5743 -14120
rect 5801 -14400 5921 -14120
rect 5979 -14400 6099 -14120
rect 6157 -14400 6277 -14120
rect 6335 -14400 6455 -14120
rect 6513 -14400 6633 -14120
rect 6691 -14400 6811 -14120
rect 6869 -14400 6989 -14120
rect 7047 -14400 7167 -14120
rect 7225 -14400 7345 -14120
rect 7403 -14400 7523 -14120
rect 7581 -14400 7701 -14120
rect 7759 -14400 7879 -14120
rect 7937 -14400 8057 -14120
rect 8115 -14400 8235 -14120
rect 8293 -14400 8413 -14120
rect 8471 -14400 8591 -14120
rect 8649 -14400 8769 -14120
rect 8827 -14400 8947 -14120
rect 9005 -14400 9125 -14120
rect 9183 -14400 9303 -14120
rect 9361 -14400 9481 -14120
rect 9539 -14400 9659 -14120
rect 9717 -14400 9837 -14120
rect 9895 -14400 10015 -14120
rect 10073 -14400 10193 -14120
rect 10251 -14400 10371 -14120
rect 10429 -14400 10549 -14120
rect 10607 -14400 10727 -14120
rect 10785 -14400 10905 -14120
rect 10963 -14400 11083 -14120
rect 11141 -14400 11261 -14120
rect 11319 -14400 11439 -14120
rect 11497 -14400 11617 -14120
rect 11675 -14400 11795 -14120
rect 11853 -14400 11973 -14120
rect 12031 -14400 12151 -14120
rect 12209 -14400 12329 -14120
rect 12387 -14400 12507 -14120
rect 12565 -14400 12685 -14120
rect -5982 -15362 -5862 -15082
rect -5804 -15362 -5684 -15082
rect -5626 -15362 -5506 -15082
rect -5448 -15362 -5328 -15082
rect -5270 -15362 -5150 -15082
rect -5092 -15362 -4972 -15082
rect -4914 -15362 -4794 -15082
rect -4736 -15362 -4616 -15082
rect -4558 -15362 -4438 -15082
rect -4380 -15362 -4260 -15082
rect -4202 -15362 -4082 -15082
rect -2127 -15400 -2007 -15120
rect -1949 -15400 -1829 -15120
rect -1771 -15400 -1651 -15120
rect -1593 -15400 -1473 -15120
rect -1415 -15400 -1295 -15120
rect -1237 -15400 -1117 -15120
rect -1059 -15400 -939 -15120
rect -881 -15400 -761 -15120
rect -703 -15400 -583 -15120
rect -525 -15400 -405 -15120
rect -347 -15400 -227 -15120
rect -169 -15400 -49 -15120
rect 9 -15400 129 -15120
rect 187 -15400 307 -15120
rect 365 -15400 485 -15120
rect 543 -15400 663 -15120
rect 721 -15400 841 -15120
rect 899 -15400 1019 -15120
rect 1077 -15400 1197 -15120
rect 1255 -15400 1375 -15120
rect 1433 -15400 1553 -15120
rect 1611 -15400 1731 -15120
rect 1789 -15400 1909 -15120
rect 1967 -15400 2087 -15120
rect 2145 -15400 2265 -15120
rect 2323 -15400 2443 -15120
rect 2501 -15400 2621 -15120
rect 2679 -15400 2799 -15120
rect 2857 -15400 2977 -15120
rect 3035 -15400 3155 -15120
rect 3213 -15400 3333 -15120
rect 3391 -15400 3511 -15120
rect 3569 -15400 3689 -15120
rect 3747 -15400 3867 -15120
rect 3925 -15400 4045 -15120
rect 5623 -15400 5743 -15120
rect 5801 -15400 5921 -15120
rect 5979 -15400 6099 -15120
rect 6157 -15400 6277 -15120
rect 6335 -15400 6455 -15120
rect 6513 -15400 6633 -15120
rect 6691 -15400 6811 -15120
rect 6869 -15400 6989 -15120
rect 7047 -15400 7167 -15120
rect 7225 -15400 7345 -15120
rect 7403 -15400 7523 -15120
rect 7581 -15400 7701 -15120
rect 7759 -15400 7879 -15120
rect 7937 -15400 8057 -15120
rect 8115 -15400 8235 -15120
rect 8293 -15400 8413 -15120
rect 8471 -15400 8591 -15120
rect 8649 -15400 8769 -15120
rect 8827 -15400 8947 -15120
rect 9005 -15400 9125 -15120
rect 9183 -15400 9303 -15120
rect 9361 -15400 9481 -15120
rect 9539 -15400 9659 -15120
rect 9717 -15400 9837 -15120
rect 9895 -15400 10015 -15120
rect 10073 -15400 10193 -15120
rect 10251 -15400 10371 -15120
rect 10429 -15400 10549 -15120
rect 10607 -15400 10727 -15120
rect 10785 -15400 10905 -15120
rect 10963 -15400 11083 -15120
rect 11141 -15400 11261 -15120
rect 11319 -15400 11439 -15120
rect 11497 -15400 11617 -15120
rect 11675 -15400 11795 -15120
rect 11853 -15400 11973 -15120
rect 12031 -15400 12151 -15120
rect 12209 -15400 12329 -15120
rect 12387 -15400 12507 -15120
rect 12565 -15400 12685 -15120
rect -5982 -16062 -5862 -15782
rect -5804 -16062 -5684 -15782
rect -5626 -16062 -5506 -15782
rect -5448 -16062 -5328 -15782
rect -5270 -16062 -5150 -15782
rect -5092 -16062 -4972 -15782
rect -4914 -16062 -4794 -15782
rect -4736 -16062 -4616 -15782
rect -4558 -16062 -4438 -15782
rect -4380 -16062 -4260 -15782
rect -4202 -16062 -4082 -15782
rect -2127 -16400 -2007 -16120
rect -1949 -16400 -1829 -16120
rect -1771 -16400 -1651 -16120
rect -1593 -16400 -1473 -16120
rect -1415 -16400 -1295 -16120
rect -1237 -16400 -1117 -16120
rect -1059 -16400 -939 -16120
rect -881 -16400 -761 -16120
rect -703 -16400 -583 -16120
rect -525 -16400 -405 -16120
rect -347 -16400 -227 -16120
rect -169 -16400 -49 -16120
rect 9 -16400 129 -16120
rect 187 -16400 307 -16120
rect 365 -16400 485 -16120
rect 543 -16400 663 -16120
rect 721 -16400 841 -16120
rect 899 -16400 1019 -16120
rect 1077 -16400 1197 -16120
rect 1255 -16400 1375 -16120
rect 1433 -16400 1553 -16120
rect 1611 -16400 1731 -16120
rect 1789 -16400 1909 -16120
rect 1967 -16400 2087 -16120
rect 2145 -16400 2265 -16120
rect 2323 -16400 2443 -16120
rect 2501 -16400 2621 -16120
rect 2679 -16400 2799 -16120
rect 2857 -16400 2977 -16120
rect 3035 -16400 3155 -16120
rect 3213 -16400 3333 -16120
rect 3391 -16400 3511 -16120
rect 3569 -16400 3689 -16120
rect 3747 -16400 3867 -16120
rect 3925 -16400 4045 -16120
rect 5623 -16400 5743 -16120
rect 5801 -16400 5921 -16120
rect 5979 -16400 6099 -16120
rect 6157 -16400 6277 -16120
rect 6335 -16400 6455 -16120
rect 6513 -16400 6633 -16120
rect 6691 -16400 6811 -16120
rect 6869 -16400 6989 -16120
rect 7047 -16400 7167 -16120
rect 7225 -16400 7345 -16120
rect 7403 -16400 7523 -16120
rect 7581 -16400 7701 -16120
rect 7759 -16400 7879 -16120
rect 7937 -16400 8057 -16120
rect 8115 -16400 8235 -16120
rect 8293 -16400 8413 -16120
rect 8471 -16400 8591 -16120
rect 8649 -16400 8769 -16120
rect 8827 -16400 8947 -16120
rect 9005 -16400 9125 -16120
rect 9183 -16400 9303 -16120
rect 9361 -16400 9481 -16120
rect 9539 -16400 9659 -16120
rect 9717 -16400 9837 -16120
rect 9895 -16400 10015 -16120
rect 10073 -16400 10193 -16120
rect 10251 -16400 10371 -16120
rect 10429 -16400 10549 -16120
rect 10607 -16400 10727 -16120
rect 10785 -16400 10905 -16120
rect 10963 -16400 11083 -16120
rect 11141 -16400 11261 -16120
rect 11319 -16400 11439 -16120
rect 11497 -16400 11617 -16120
rect 11675 -16400 11795 -16120
rect 11853 -16400 11973 -16120
rect 12031 -16400 12151 -16120
rect 12209 -16400 12329 -16120
rect 12387 -16400 12507 -16120
rect 12565 -16400 12685 -16120
rect -5982 -16762 -5862 -16482
rect -5804 -16762 -5684 -16482
rect -5626 -16762 -5506 -16482
rect -5448 -16762 -5328 -16482
rect -5270 -16762 -5150 -16482
rect -5092 -16762 -4972 -16482
rect -4914 -16762 -4794 -16482
rect -4736 -16762 -4616 -16482
rect -4558 -16762 -4438 -16482
rect -4380 -16762 -4260 -16482
rect -4202 -16762 -4082 -16482
<< pmos >>
rect -1408 -3152 -1288 -2872
rect -1230 -3152 -1110 -2872
rect -1052 -3152 -932 -2872
rect -874 -3152 -754 -2872
rect -696 -3152 -576 -2872
rect -518 -3152 -398 -2872
rect -340 -3152 -220 -2872
rect -162 -3152 -42 -2872
rect 16 -3152 136 -2872
rect 194 -3152 314 -2872
rect 372 -3152 492 -2872
rect 550 -3152 670 -2872
rect 728 -3152 848 -2872
rect 906 -3152 1026 -2872
rect 1084 -3152 1204 -2872
rect 1262 -3152 1382 -2872
rect 1440 -3152 1560 -2872
rect 1618 -3152 1738 -2872
rect 1796 -3152 1916 -2872
rect 1974 -3152 2094 -2872
rect 2152 -3152 2272 -2872
rect 2330 -3152 2450 -2872
rect 2508 -3152 2628 -2872
rect -1408 -4052 -1288 -3772
rect -1230 -4052 -1110 -3772
rect -1052 -4052 -932 -3772
rect -874 -4052 -754 -3772
rect -696 -4052 -576 -3772
rect -518 -4052 -398 -3772
rect -340 -4052 -220 -3772
rect -162 -4052 -42 -3772
rect 16 -4052 136 -3772
rect 194 -4052 314 -3772
rect 372 -4052 492 -3772
rect 550 -4052 670 -3772
rect 728 -4052 848 -3772
rect 906 -4052 1026 -3772
rect 1084 -4052 1204 -3772
rect 1262 -4052 1382 -3772
rect 1440 -4052 1560 -3772
rect 1618 -4052 1738 -3772
rect 1796 -4052 1916 -3772
rect 1974 -4052 2094 -3772
rect 2152 -4052 2272 -3772
rect 2330 -4052 2450 -3772
rect 2508 -4052 2628 -3772
rect -1408 -4952 -1288 -4672
rect -1230 -4952 -1110 -4672
rect -1052 -4952 -932 -4672
rect -874 -4952 -754 -4672
rect -696 -4952 -576 -4672
rect -518 -4952 -398 -4672
rect -340 -4952 -220 -4672
rect -162 -4952 -42 -4672
rect 16 -4952 136 -4672
rect 194 -4952 314 -4672
rect 372 -4952 492 -4672
rect 550 -4952 670 -4672
rect 728 -4952 848 -4672
rect 906 -4952 1026 -4672
rect 1084 -4952 1204 -4672
rect 1262 -4952 1382 -4672
rect 1440 -4952 1560 -4672
rect 1618 -4952 1738 -4672
rect 1796 -4952 1916 -4672
rect 1974 -4952 2094 -4672
rect 2152 -4952 2272 -4672
rect 2330 -4952 2450 -4672
rect 2508 -4952 2628 -4672
rect -1408 -5852 -1288 -5572
rect -1230 -5852 -1110 -5572
rect -1052 -5852 -932 -5572
rect -874 -5852 -754 -5572
rect -696 -5852 -576 -5572
rect -518 -5852 -398 -5572
rect -340 -5852 -220 -5572
rect -162 -5852 -42 -5572
rect 16 -5852 136 -5572
rect 194 -5852 314 -5572
rect 372 -5852 492 -5572
rect 550 -5852 670 -5572
rect 728 -5852 848 -5572
rect 906 -5852 1026 -5572
rect 1084 -5852 1204 -5572
rect 1262 -5852 1382 -5572
rect 1440 -5852 1560 -5572
rect 1618 -5852 1738 -5572
rect 1796 -5852 1916 -5572
rect 1974 -5852 2094 -5572
rect 2152 -5852 2272 -5572
rect 2330 -5852 2450 -5572
rect 2508 -5852 2628 -5572
<< pmoslvt >>
rect -6256 -2400 -6136 -2120
rect -6078 -2400 -5958 -2120
rect -5900 -2400 -5780 -2120
rect -5722 -2400 -5602 -2120
rect -5544 -2400 -5424 -2120
rect -5366 -2400 -5246 -2120
rect -5188 -2400 -5068 -2120
rect -5010 -2400 -4890 -2120
rect -4832 -2400 -4712 -2120
rect -4654 -2400 -4534 -2120
rect -4476 -2400 -4356 -2120
rect -4298 -2400 -4178 -2120
rect -4120 -2400 -4000 -2120
rect -3942 -2400 -3822 -2120
rect -3764 -2400 -3644 -2120
rect -3586 -2400 -3466 -2120
rect -6256 -3270 -6136 -2990
rect -6078 -3270 -5958 -2990
rect -5900 -3270 -5780 -2990
rect -5722 -3270 -5602 -2990
rect -5544 -3270 -5424 -2990
rect -5366 -3270 -5246 -2990
rect -5188 -3270 -5068 -2990
rect -5010 -3270 -4890 -2990
rect -4832 -3270 -4712 -2990
rect -4654 -3270 -4534 -2990
rect -4476 -3270 -4356 -2990
rect -4298 -3270 -4178 -2990
rect -4120 -3270 -4000 -2990
rect -3942 -3270 -3822 -2990
rect -3764 -3270 -3644 -2990
rect -3586 -3270 -3466 -2990
rect -6256 -4140 -6136 -3860
rect -6078 -4140 -5958 -3860
rect -5900 -4140 -5780 -3860
rect -5722 -4140 -5602 -3860
rect -5544 -4140 -5424 -3860
rect -5366 -4140 -5246 -3860
rect -5188 -4140 -5068 -3860
rect -5010 -4140 -4890 -3860
rect -4832 -4140 -4712 -3860
rect -4654 -4140 -4534 -3860
rect -4476 -4140 -4356 -3860
rect -4298 -4140 -4178 -3860
rect -4120 -4140 -4000 -3860
rect -3942 -4140 -3822 -3860
rect -3764 -4140 -3644 -3860
rect -3586 -4140 -3466 -3860
rect -6256 -5010 -6136 -4730
rect -6078 -5010 -5958 -4730
rect -5900 -5010 -5780 -4730
rect -5722 -5010 -5602 -4730
rect -5544 -5010 -5424 -4730
rect -5366 -5010 -5246 -4730
rect -5188 -5010 -5068 -4730
rect -5010 -5010 -4890 -4730
rect -4832 -5010 -4712 -4730
rect -4654 -5010 -4534 -4730
rect -4476 -5010 -4356 -4730
rect -4298 -5010 -4178 -4730
rect -4120 -5010 -4000 -4730
rect -3942 -5010 -3822 -4730
rect -3764 -5010 -3644 -4730
rect -3586 -5010 -3466 -4730
rect -6256 -5880 -6136 -5600
rect -6078 -5880 -5958 -5600
rect -5900 -5880 -5780 -5600
rect -5722 -5880 -5602 -5600
rect -5544 -5880 -5424 -5600
rect -5366 -5880 -5246 -5600
rect -5188 -5880 -5068 -5600
rect -5010 -5880 -4890 -5600
rect -4832 -5880 -4712 -5600
rect -4654 -5880 -4534 -5600
rect -4476 -5880 -4356 -5600
rect -4298 -5880 -4178 -5600
rect -4120 -5880 -4000 -5600
rect -3942 -5880 -3822 -5600
rect -3764 -5880 -3644 -5600
rect -3586 -5880 -3466 -5600
<< nmoslvt >>
rect -5582 -8142 -5462 -7862
rect -5404 -8142 -5284 -7862
rect -5226 -8142 -5106 -7862
rect -5048 -8142 -4928 -7862
rect -4870 -8142 -4750 -7862
rect -4692 -8142 -4572 -7862
rect -4514 -8142 -4394 -7862
rect -4336 -8142 -4216 -7862
rect -4158 -8142 -4038 -7862
rect -5582 -8692 -5462 -8412
rect -5404 -8692 -5284 -8412
rect -5226 -8692 -5106 -8412
rect -5048 -8692 -4928 -8412
rect -4870 -8692 -4750 -8412
rect -4692 -8692 -4572 -8412
rect -4514 -8692 -4394 -8412
rect -4336 -8692 -4216 -8412
rect -4158 -8692 -4038 -8412
rect -5582 -9242 -5462 -8962
rect -5404 -9242 -5284 -8962
rect -5226 -9242 -5106 -8962
rect -5048 -9242 -4928 -8962
rect -4870 -9242 -4750 -8962
rect -4692 -9242 -4572 -8962
rect -4514 -9242 -4394 -8962
rect -4336 -9242 -4216 -8962
rect -4158 -9242 -4038 -8962
rect -5582 -9792 -5462 -9512
rect -5404 -9792 -5284 -9512
rect -5226 -9792 -5106 -9512
rect -5048 -9792 -4928 -9512
rect -4870 -9792 -4750 -9512
rect -4692 -9792 -4572 -9512
rect -4514 -9792 -4394 -9512
rect -4336 -9792 -4216 -9512
rect -4158 -9792 -4038 -9512
rect -5582 -10342 -5462 -10062
rect -5404 -10342 -5284 -10062
rect -5226 -10342 -5106 -10062
rect -5048 -10342 -4928 -10062
rect -4870 -10342 -4750 -10062
rect -4692 -10342 -4572 -10062
rect -4514 -10342 -4394 -10062
rect -4336 -10342 -4216 -10062
rect -4158 -10342 -4038 -10062
rect -5582 -10892 -5462 -10612
rect -5404 -10892 -5284 -10612
rect -5226 -10892 -5106 -10612
rect -5048 -10892 -4928 -10612
rect -4870 -10892 -4750 -10612
rect -4692 -10892 -4572 -10612
rect -4514 -10892 -4394 -10612
rect -4336 -10892 -4216 -10612
rect -4158 -10892 -4038 -10612
rect -5582 -11442 -5462 -11162
rect -5404 -11442 -5284 -11162
rect -5226 -11442 -5106 -11162
rect -5048 -11442 -4928 -11162
rect -4870 -11442 -4750 -11162
rect -4692 -11442 -4572 -11162
rect -4514 -11442 -4394 -11162
rect -4336 -11442 -4216 -11162
rect -4158 -11442 -4038 -11162
rect -5582 -11992 -5462 -11712
rect -5404 -11992 -5284 -11712
rect -5226 -11992 -5106 -11712
rect -5048 -11992 -4928 -11712
rect -4870 -11992 -4750 -11712
rect -4692 -11992 -4572 -11712
rect -4514 -11992 -4394 -11712
rect -4336 -11992 -4216 -11712
rect -4158 -11992 -4038 -11712
rect -5870 -12940 -5830 -12700
rect -5620 -12940 -5580 -12700
rect -5370 -12940 -5330 -12700
rect -5120 -12940 -5080 -12700
rect -4870 -12940 -4830 -12700
rect -4620 -12940 -4580 -12700
rect -4370 -12940 -4330 -12700
rect -4120 -12940 -4080 -12700
rect -5870 -13620 -5830 -13380
rect -5620 -13620 -5580 -13380
rect -5370 -13620 -5330 -13380
rect -5120 -13620 -5080 -13380
rect -4870 -13620 -4830 -13380
rect -4620 -13620 -4580 -13380
rect -4370 -13620 -4330 -13380
rect -4120 -13620 -4080 -13380
<< ndiff >>
rect -5640 -7874 -5582 -7862
rect -5640 -8130 -5628 -7874
rect -5594 -8130 -5582 -7874
rect -5640 -8142 -5582 -8130
rect -5462 -7874 -5404 -7862
rect -5462 -8130 -5450 -7874
rect -5416 -8130 -5404 -7874
rect -5462 -8142 -5404 -8130
rect -5284 -7874 -5226 -7862
rect -5284 -8130 -5272 -7874
rect -5238 -8130 -5226 -7874
rect -5284 -8142 -5226 -8130
rect -5106 -7874 -5048 -7862
rect -5106 -8130 -5094 -7874
rect -5060 -8130 -5048 -7874
rect -5106 -8142 -5048 -8130
rect -4928 -7874 -4870 -7862
rect -4928 -8130 -4916 -7874
rect -4882 -8130 -4870 -7874
rect -4928 -8142 -4870 -8130
rect -4750 -7874 -4692 -7862
rect -4750 -8130 -4738 -7874
rect -4704 -8130 -4692 -7874
rect -4750 -8142 -4692 -8130
rect -4572 -7874 -4514 -7862
rect -4572 -8130 -4560 -7874
rect -4526 -8130 -4514 -7874
rect -4572 -8142 -4514 -8130
rect -4394 -7874 -4336 -7862
rect -4394 -8130 -4382 -7874
rect -4348 -8130 -4336 -7874
rect -4394 -8142 -4336 -8130
rect -4216 -7874 -4158 -7862
rect -4216 -8130 -4204 -7874
rect -4170 -8130 -4158 -7874
rect -4216 -8142 -4158 -8130
rect -4038 -7874 -3980 -7862
rect -4038 -8130 -4026 -7874
rect -3992 -8130 -3980 -7874
rect -4038 -8142 -3980 -8130
rect -2185 -8132 -2127 -8120
rect -2185 -8388 -2173 -8132
rect -2139 -8388 -2127 -8132
rect -2185 -8400 -2127 -8388
rect -2007 -8132 -1949 -8120
rect -2007 -8388 -1995 -8132
rect -1961 -8388 -1949 -8132
rect -2007 -8400 -1949 -8388
rect -1829 -8132 -1771 -8120
rect -1829 -8388 -1817 -8132
rect -1783 -8388 -1771 -8132
rect -1829 -8400 -1771 -8388
rect -1651 -8132 -1593 -8120
rect -1651 -8388 -1639 -8132
rect -1605 -8388 -1593 -8132
rect -1651 -8400 -1593 -8388
rect -1473 -8132 -1415 -8120
rect -1473 -8388 -1461 -8132
rect -1427 -8388 -1415 -8132
rect -1473 -8400 -1415 -8388
rect -1295 -8132 -1237 -8120
rect -1295 -8388 -1283 -8132
rect -1249 -8388 -1237 -8132
rect -1295 -8400 -1237 -8388
rect -1117 -8132 -1059 -8120
rect -1117 -8388 -1105 -8132
rect -1071 -8388 -1059 -8132
rect -1117 -8400 -1059 -8388
rect -939 -8132 -881 -8120
rect -939 -8388 -927 -8132
rect -893 -8388 -881 -8132
rect -939 -8400 -881 -8388
rect -761 -8132 -703 -8120
rect -761 -8388 -749 -8132
rect -715 -8388 -703 -8132
rect -761 -8400 -703 -8388
rect -583 -8132 -525 -8120
rect -583 -8388 -571 -8132
rect -537 -8388 -525 -8132
rect -583 -8400 -525 -8388
rect -405 -8132 -347 -8120
rect -405 -8388 -393 -8132
rect -359 -8388 -347 -8132
rect -405 -8400 -347 -8388
rect -227 -8132 -169 -8120
rect -227 -8388 -215 -8132
rect -181 -8388 -169 -8132
rect -227 -8400 -169 -8388
rect -49 -8132 9 -8120
rect -49 -8388 -37 -8132
rect -3 -8388 9 -8132
rect -49 -8400 9 -8388
rect 129 -8132 187 -8120
rect 129 -8388 141 -8132
rect 175 -8388 187 -8132
rect 129 -8400 187 -8388
rect 307 -8132 365 -8120
rect 307 -8388 319 -8132
rect 353 -8388 365 -8132
rect 307 -8400 365 -8388
rect 485 -8132 543 -8120
rect 485 -8388 497 -8132
rect 531 -8388 543 -8132
rect 485 -8400 543 -8388
rect 663 -8132 721 -8120
rect 663 -8388 675 -8132
rect 709 -8388 721 -8132
rect 663 -8400 721 -8388
rect 841 -8132 899 -8120
rect 841 -8388 853 -8132
rect 887 -8388 899 -8132
rect 841 -8400 899 -8388
rect 1019 -8132 1077 -8120
rect 1019 -8388 1031 -8132
rect 1065 -8388 1077 -8132
rect 1019 -8400 1077 -8388
rect 1197 -8132 1255 -8120
rect 1197 -8388 1209 -8132
rect 1243 -8388 1255 -8132
rect 1197 -8400 1255 -8388
rect 1375 -8132 1433 -8120
rect 1375 -8388 1387 -8132
rect 1421 -8388 1433 -8132
rect 1375 -8400 1433 -8388
rect 1553 -8132 1611 -8120
rect 1553 -8388 1565 -8132
rect 1599 -8388 1611 -8132
rect 1553 -8400 1611 -8388
rect 1731 -8132 1789 -8120
rect 1731 -8388 1743 -8132
rect 1777 -8388 1789 -8132
rect 1731 -8400 1789 -8388
rect 1909 -8132 1967 -8120
rect 1909 -8388 1921 -8132
rect 1955 -8388 1967 -8132
rect 1909 -8400 1967 -8388
rect 2087 -8132 2145 -8120
rect 2087 -8388 2099 -8132
rect 2133 -8388 2145 -8132
rect 2087 -8400 2145 -8388
rect 2265 -8132 2323 -8120
rect 2265 -8388 2277 -8132
rect 2311 -8388 2323 -8132
rect 2265 -8400 2323 -8388
rect 2443 -8132 2501 -8120
rect 2443 -8388 2455 -8132
rect 2489 -8388 2501 -8132
rect 2443 -8400 2501 -8388
rect 2621 -8132 2679 -8120
rect 2621 -8388 2633 -8132
rect 2667 -8388 2679 -8132
rect 2621 -8400 2679 -8388
rect 2799 -8132 2857 -8120
rect 2799 -8388 2811 -8132
rect 2845 -8388 2857 -8132
rect 2799 -8400 2857 -8388
rect 2977 -8132 3035 -8120
rect 2977 -8388 2989 -8132
rect 3023 -8388 3035 -8132
rect 2977 -8400 3035 -8388
rect 3155 -8132 3213 -8120
rect 3155 -8388 3167 -8132
rect 3201 -8388 3213 -8132
rect 3155 -8400 3213 -8388
rect 3333 -8132 3391 -8120
rect 3333 -8388 3345 -8132
rect 3379 -8388 3391 -8132
rect 3333 -8400 3391 -8388
rect 3511 -8132 3569 -8120
rect 3511 -8388 3523 -8132
rect 3557 -8388 3569 -8132
rect 3511 -8400 3569 -8388
rect 3689 -8132 3747 -8120
rect 3689 -8388 3701 -8132
rect 3735 -8388 3747 -8132
rect 3689 -8400 3747 -8388
rect 3867 -8132 3925 -8120
rect 3867 -8388 3879 -8132
rect 3913 -8388 3925 -8132
rect 3867 -8400 3925 -8388
rect 4045 -8132 4103 -8120
rect 4045 -8388 4057 -8132
rect 4091 -8388 4103 -8132
rect 4045 -8400 4103 -8388
rect -5640 -8424 -5582 -8412
rect -5640 -8680 -5628 -8424
rect -5594 -8680 -5582 -8424
rect -5640 -8692 -5582 -8680
rect -5462 -8424 -5404 -8412
rect -5462 -8680 -5450 -8424
rect -5416 -8680 -5404 -8424
rect -5462 -8692 -5404 -8680
rect -5284 -8424 -5226 -8412
rect -5284 -8680 -5272 -8424
rect -5238 -8680 -5226 -8424
rect -5284 -8692 -5226 -8680
rect -5106 -8424 -5048 -8412
rect -5106 -8680 -5094 -8424
rect -5060 -8680 -5048 -8424
rect -5106 -8692 -5048 -8680
rect -4928 -8424 -4870 -8412
rect -4928 -8680 -4916 -8424
rect -4882 -8680 -4870 -8424
rect -4928 -8692 -4870 -8680
rect -4750 -8424 -4692 -8412
rect -4750 -8680 -4738 -8424
rect -4704 -8680 -4692 -8424
rect -4750 -8692 -4692 -8680
rect -4572 -8424 -4514 -8412
rect -4572 -8680 -4560 -8424
rect -4526 -8680 -4514 -8424
rect -4572 -8692 -4514 -8680
rect -4394 -8424 -4336 -8412
rect -4394 -8680 -4382 -8424
rect -4348 -8680 -4336 -8424
rect -4394 -8692 -4336 -8680
rect -4216 -8424 -4158 -8412
rect -4216 -8680 -4204 -8424
rect -4170 -8680 -4158 -8424
rect -4216 -8692 -4158 -8680
rect -4038 -8424 -3980 -8412
rect -4038 -8680 -4026 -8424
rect -3992 -8680 -3980 -8424
rect -4038 -8692 -3980 -8680
rect 6500 -8894 6558 -8882
rect -5640 -8974 -5582 -8962
rect -5640 -9230 -5628 -8974
rect -5594 -9230 -5582 -8974
rect -5640 -9242 -5582 -9230
rect -5462 -8974 -5404 -8962
rect -5462 -9230 -5450 -8974
rect -5416 -9230 -5404 -8974
rect -5462 -9242 -5404 -9230
rect -5284 -8974 -5226 -8962
rect -5284 -9230 -5272 -8974
rect -5238 -9230 -5226 -8974
rect -5284 -9242 -5226 -9230
rect -5106 -8974 -5048 -8962
rect -5106 -9230 -5094 -8974
rect -5060 -9230 -5048 -8974
rect -5106 -9242 -5048 -9230
rect -4928 -8974 -4870 -8962
rect -4928 -9230 -4916 -8974
rect -4882 -9230 -4870 -8974
rect -4928 -9242 -4870 -9230
rect -4750 -8974 -4692 -8962
rect -4750 -9230 -4738 -8974
rect -4704 -9230 -4692 -8974
rect -4750 -9242 -4692 -9230
rect -4572 -8974 -4514 -8962
rect -4572 -9230 -4560 -8974
rect -4526 -9230 -4514 -8974
rect -4572 -9242 -4514 -9230
rect -4394 -8974 -4336 -8962
rect -4394 -9230 -4382 -8974
rect -4348 -9230 -4336 -8974
rect -4394 -9242 -4336 -9230
rect -4216 -8974 -4158 -8962
rect -4216 -9230 -4204 -8974
rect -4170 -9230 -4158 -8974
rect -4216 -9242 -4158 -9230
rect -4038 -8974 -3980 -8962
rect -4038 -9230 -4026 -8974
rect -3992 -9230 -3980 -8974
rect -4038 -9242 -3980 -9230
rect -2185 -9132 -2127 -9120
rect -2185 -9388 -2173 -9132
rect -2139 -9388 -2127 -9132
rect -2185 -9400 -2127 -9388
rect -2007 -9132 -1949 -9120
rect -2007 -9388 -1995 -9132
rect -1961 -9388 -1949 -9132
rect -2007 -9400 -1949 -9388
rect -1829 -9132 -1771 -9120
rect -1829 -9388 -1817 -9132
rect -1783 -9388 -1771 -9132
rect -1829 -9400 -1771 -9388
rect -1651 -9132 -1593 -9120
rect -1651 -9388 -1639 -9132
rect -1605 -9388 -1593 -9132
rect -1651 -9400 -1593 -9388
rect -1473 -9132 -1415 -9120
rect -1473 -9388 -1461 -9132
rect -1427 -9388 -1415 -9132
rect -1473 -9400 -1415 -9388
rect -1295 -9132 -1237 -9120
rect -1295 -9388 -1283 -9132
rect -1249 -9388 -1237 -9132
rect -1295 -9400 -1237 -9388
rect -1117 -9132 -1059 -9120
rect -1117 -9388 -1105 -9132
rect -1071 -9388 -1059 -9132
rect -1117 -9400 -1059 -9388
rect -939 -9132 -881 -9120
rect -939 -9388 -927 -9132
rect -893 -9388 -881 -9132
rect -939 -9400 -881 -9388
rect -761 -9132 -703 -9120
rect -761 -9388 -749 -9132
rect -715 -9388 -703 -9132
rect -761 -9400 -703 -9388
rect -583 -9132 -525 -9120
rect -583 -9388 -571 -9132
rect -537 -9388 -525 -9132
rect -583 -9400 -525 -9388
rect -405 -9132 -347 -9120
rect -405 -9388 -393 -9132
rect -359 -9388 -347 -9132
rect -405 -9400 -347 -9388
rect -227 -9132 -169 -9120
rect -227 -9388 -215 -9132
rect -181 -9388 -169 -9132
rect -227 -9400 -169 -9388
rect -49 -9132 9 -9120
rect -49 -9388 -37 -9132
rect -3 -9388 9 -9132
rect -49 -9400 9 -9388
rect 129 -9132 187 -9120
rect 129 -9388 141 -9132
rect 175 -9388 187 -9132
rect 129 -9400 187 -9388
rect 307 -9132 365 -9120
rect 307 -9388 319 -9132
rect 353 -9388 365 -9132
rect 307 -9400 365 -9388
rect 485 -9132 543 -9120
rect 485 -9388 497 -9132
rect 531 -9388 543 -9132
rect 485 -9400 543 -9388
rect 663 -9132 721 -9120
rect 663 -9388 675 -9132
rect 709 -9388 721 -9132
rect 663 -9400 721 -9388
rect 841 -9132 899 -9120
rect 841 -9388 853 -9132
rect 887 -9388 899 -9132
rect 841 -9400 899 -9388
rect 1019 -9132 1077 -9120
rect 1019 -9388 1031 -9132
rect 1065 -9388 1077 -9132
rect 1019 -9400 1077 -9388
rect 1197 -9132 1255 -9120
rect 1197 -9388 1209 -9132
rect 1243 -9388 1255 -9132
rect 1197 -9400 1255 -9388
rect 1375 -9132 1433 -9120
rect 1375 -9388 1387 -9132
rect 1421 -9388 1433 -9132
rect 1375 -9400 1433 -9388
rect 1553 -9132 1611 -9120
rect 1553 -9388 1565 -9132
rect 1599 -9388 1611 -9132
rect 1553 -9400 1611 -9388
rect 1731 -9132 1789 -9120
rect 1731 -9388 1743 -9132
rect 1777 -9388 1789 -9132
rect 1731 -9400 1789 -9388
rect 1909 -9132 1967 -9120
rect 1909 -9388 1921 -9132
rect 1955 -9388 1967 -9132
rect 1909 -9400 1967 -9388
rect 2087 -9132 2145 -9120
rect 2087 -9388 2099 -9132
rect 2133 -9388 2145 -9132
rect 2087 -9400 2145 -9388
rect 2265 -9132 2323 -9120
rect 2265 -9388 2277 -9132
rect 2311 -9388 2323 -9132
rect 2265 -9400 2323 -9388
rect 2443 -9132 2501 -9120
rect 2443 -9388 2455 -9132
rect 2489 -9388 2501 -9132
rect 2443 -9400 2501 -9388
rect 2621 -9132 2679 -9120
rect 2621 -9388 2633 -9132
rect 2667 -9388 2679 -9132
rect 2621 -9400 2679 -9388
rect 2799 -9132 2857 -9120
rect 2799 -9388 2811 -9132
rect 2845 -9388 2857 -9132
rect 2799 -9400 2857 -9388
rect 2977 -9132 3035 -9120
rect 2977 -9388 2989 -9132
rect 3023 -9388 3035 -9132
rect 2977 -9400 3035 -9388
rect 3155 -9132 3213 -9120
rect 3155 -9388 3167 -9132
rect 3201 -9388 3213 -9132
rect 3155 -9400 3213 -9388
rect 3333 -9132 3391 -9120
rect 3333 -9388 3345 -9132
rect 3379 -9388 3391 -9132
rect 3333 -9400 3391 -9388
rect 3511 -9132 3569 -9120
rect 3511 -9388 3523 -9132
rect 3557 -9388 3569 -9132
rect 3511 -9400 3569 -9388
rect 3689 -9132 3747 -9120
rect 3689 -9388 3701 -9132
rect 3735 -9388 3747 -9132
rect 3689 -9400 3747 -9388
rect 3867 -9132 3925 -9120
rect 3867 -9388 3879 -9132
rect 3913 -9388 3925 -9132
rect 3867 -9400 3925 -9388
rect 4045 -9132 4103 -9120
rect 4045 -9388 4057 -9132
rect 4091 -9388 4103 -9132
rect 6500 -9150 6512 -8894
rect 6546 -9150 6558 -8894
rect 6500 -9162 6558 -9150
rect 6678 -8894 6736 -8882
rect 6678 -9150 6690 -8894
rect 6724 -9150 6736 -8894
rect 6678 -9162 6736 -9150
rect 6856 -8894 6914 -8882
rect 6856 -9150 6868 -8894
rect 6902 -9150 6914 -8894
rect 6856 -9162 6914 -9150
rect 7034 -8894 7092 -8882
rect 7034 -9150 7046 -8894
rect 7080 -9150 7092 -8894
rect 7034 -9162 7092 -9150
rect 7212 -8894 7270 -8882
rect 7212 -9150 7224 -8894
rect 7258 -9150 7270 -8894
rect 7212 -9162 7270 -9150
rect 7390 -8894 7448 -8882
rect 7390 -9150 7402 -8894
rect 7436 -9150 7448 -8894
rect 7390 -9162 7448 -9150
rect 7568 -8894 7626 -8882
rect 7568 -9150 7580 -8894
rect 7614 -9150 7626 -8894
rect 7568 -9162 7626 -9150
rect 7746 -8894 7804 -8882
rect 7746 -9150 7758 -8894
rect 7792 -9150 7804 -8894
rect 7746 -9162 7804 -9150
rect 7924 -8894 7982 -8882
rect 7924 -9150 7936 -8894
rect 7970 -9150 7982 -8894
rect 7924 -9162 7982 -9150
rect 8102 -8894 8160 -8882
rect 8102 -9150 8114 -8894
rect 8148 -9150 8160 -8894
rect 8102 -9162 8160 -9150
rect 8280 -8894 8338 -8882
rect 8280 -9150 8292 -8894
rect 8326 -9150 8338 -8894
rect 8280 -9162 8338 -9150
rect 8458 -8894 8516 -8882
rect 8458 -9150 8470 -8894
rect 8504 -9150 8516 -8894
rect 8458 -9162 8516 -9150
rect 8636 -8894 8694 -8882
rect 8636 -9150 8648 -8894
rect 8682 -9150 8694 -8894
rect 8636 -9162 8694 -9150
rect 8814 -8894 8872 -8882
rect 8814 -9150 8826 -8894
rect 8860 -9150 8872 -8894
rect 8814 -9162 8872 -9150
rect 8992 -8894 9050 -8882
rect 8992 -9150 9004 -8894
rect 9038 -9150 9050 -8894
rect 8992 -9162 9050 -9150
rect 9170 -8894 9228 -8882
rect 9170 -9150 9182 -8894
rect 9216 -9150 9228 -8894
rect 9170 -9162 9228 -9150
rect 9348 -8894 9406 -8882
rect 9348 -9150 9360 -8894
rect 9394 -9150 9406 -8894
rect 9348 -9162 9406 -9150
rect 10760 -8924 10818 -8912
rect 10760 -9180 10772 -8924
rect 10806 -9180 10818 -8924
rect 10760 -9192 10818 -9180
rect 10938 -8924 10996 -8912
rect 10938 -9180 10950 -8924
rect 10984 -9180 10996 -8924
rect 10938 -9192 10996 -9180
rect 11052 -8924 11110 -8912
rect 11052 -9180 11064 -8924
rect 11098 -9180 11110 -8924
rect 11052 -9192 11110 -9180
rect 11230 -8924 11288 -8912
rect 11230 -9180 11242 -8924
rect 11276 -9180 11288 -8924
rect 11230 -9192 11288 -9180
rect 11344 -8924 11402 -8912
rect 11344 -9180 11356 -8924
rect 11390 -9180 11402 -8924
rect 11344 -9192 11402 -9180
rect 11522 -8924 11580 -8912
rect 11522 -9180 11534 -8924
rect 11568 -9180 11580 -8924
rect 11522 -9192 11580 -9180
rect 11636 -8924 11694 -8912
rect 11636 -9180 11648 -8924
rect 11682 -9180 11694 -8924
rect 11636 -9192 11694 -9180
rect 11814 -8924 11872 -8912
rect 11814 -9180 11826 -8924
rect 11860 -9180 11872 -8924
rect 11814 -9192 11872 -9180
rect 11928 -8924 11986 -8912
rect 11928 -9180 11940 -8924
rect 11974 -9180 11986 -8924
rect 11928 -9192 11986 -9180
rect 12106 -8924 12164 -8912
rect 12106 -9180 12118 -8924
rect 12152 -9180 12164 -8924
rect 12106 -9192 12164 -9180
rect 12220 -8924 12278 -8912
rect 12220 -9180 12232 -8924
rect 12266 -9180 12278 -8924
rect 12220 -9192 12278 -9180
rect 12398 -8924 12456 -8912
rect 12398 -9180 12410 -8924
rect 12444 -9180 12456 -8924
rect 12398 -9192 12456 -9180
rect 12512 -8924 12570 -8912
rect 12512 -9180 12524 -8924
rect 12558 -9180 12570 -8924
rect 12512 -9192 12570 -9180
rect 12690 -8924 12748 -8912
rect 12690 -9180 12702 -8924
rect 12736 -9180 12748 -8924
rect 12690 -9192 12748 -9180
rect 4045 -9400 4103 -9388
rect -5640 -9524 -5582 -9512
rect -5640 -9780 -5628 -9524
rect -5594 -9780 -5582 -9524
rect -5640 -9792 -5582 -9780
rect -5462 -9524 -5404 -9512
rect -5462 -9780 -5450 -9524
rect -5416 -9780 -5404 -9524
rect -5462 -9792 -5404 -9780
rect -5284 -9524 -5226 -9512
rect -5284 -9780 -5272 -9524
rect -5238 -9780 -5226 -9524
rect -5284 -9792 -5226 -9780
rect -5106 -9524 -5048 -9512
rect -5106 -9780 -5094 -9524
rect -5060 -9780 -5048 -9524
rect -5106 -9792 -5048 -9780
rect -4928 -9524 -4870 -9512
rect -4928 -9780 -4916 -9524
rect -4882 -9780 -4870 -9524
rect -4928 -9792 -4870 -9780
rect -4750 -9524 -4692 -9512
rect -4750 -9780 -4738 -9524
rect -4704 -9780 -4692 -9524
rect -4750 -9792 -4692 -9780
rect -4572 -9524 -4514 -9512
rect -4572 -9780 -4560 -9524
rect -4526 -9780 -4514 -9524
rect -4572 -9792 -4514 -9780
rect -4394 -9524 -4336 -9512
rect -4394 -9780 -4382 -9524
rect -4348 -9780 -4336 -9524
rect -4394 -9792 -4336 -9780
rect -4216 -9524 -4158 -9512
rect -4216 -9780 -4204 -9524
rect -4170 -9780 -4158 -9524
rect -4216 -9792 -4158 -9780
rect -4038 -9524 -3980 -9512
rect -4038 -9780 -4026 -9524
rect -3992 -9780 -3980 -9524
rect 10760 -9694 10818 -9682
rect -4038 -9792 -3980 -9780
rect 6500 -9794 6558 -9782
rect -5640 -10074 -5582 -10062
rect -5640 -10330 -5628 -10074
rect -5594 -10330 -5582 -10074
rect -5640 -10342 -5582 -10330
rect -5462 -10074 -5404 -10062
rect -5462 -10330 -5450 -10074
rect -5416 -10330 -5404 -10074
rect -5462 -10342 -5404 -10330
rect -5284 -10074 -5226 -10062
rect -5284 -10330 -5272 -10074
rect -5238 -10330 -5226 -10074
rect -5284 -10342 -5226 -10330
rect -5106 -10074 -5048 -10062
rect -5106 -10330 -5094 -10074
rect -5060 -10330 -5048 -10074
rect -5106 -10342 -5048 -10330
rect -4928 -10074 -4870 -10062
rect -4928 -10330 -4916 -10074
rect -4882 -10330 -4870 -10074
rect -4928 -10342 -4870 -10330
rect -4750 -10074 -4692 -10062
rect -4750 -10330 -4738 -10074
rect -4704 -10330 -4692 -10074
rect -4750 -10342 -4692 -10330
rect -4572 -10074 -4514 -10062
rect -4572 -10330 -4560 -10074
rect -4526 -10330 -4514 -10074
rect -4572 -10342 -4514 -10330
rect -4394 -10074 -4336 -10062
rect -4394 -10330 -4382 -10074
rect -4348 -10330 -4336 -10074
rect -4394 -10342 -4336 -10330
rect -4216 -10074 -4158 -10062
rect -4216 -10330 -4204 -10074
rect -4170 -10330 -4158 -10074
rect -4216 -10342 -4158 -10330
rect -4038 -10074 -3980 -10062
rect -4038 -10330 -4026 -10074
rect -3992 -10330 -3980 -10074
rect 6500 -10050 6512 -9794
rect 6546 -10050 6558 -9794
rect 6500 -10062 6558 -10050
rect 6678 -9794 6736 -9782
rect 6678 -10050 6690 -9794
rect 6724 -10050 6736 -9794
rect 6678 -10062 6736 -10050
rect 6856 -9794 6914 -9782
rect 6856 -10050 6868 -9794
rect 6902 -10050 6914 -9794
rect 6856 -10062 6914 -10050
rect 7034 -9794 7092 -9782
rect 7034 -10050 7046 -9794
rect 7080 -10050 7092 -9794
rect 7034 -10062 7092 -10050
rect 7212 -9794 7270 -9782
rect 7212 -10050 7224 -9794
rect 7258 -10050 7270 -9794
rect 7212 -10062 7270 -10050
rect 7390 -9794 7448 -9782
rect 7390 -10050 7402 -9794
rect 7436 -10050 7448 -9794
rect 7390 -10062 7448 -10050
rect 7568 -9794 7626 -9782
rect 7568 -10050 7580 -9794
rect 7614 -10050 7626 -9794
rect 7568 -10062 7626 -10050
rect 7746 -9794 7804 -9782
rect 7746 -10050 7758 -9794
rect 7792 -10050 7804 -9794
rect 7746 -10062 7804 -10050
rect 7924 -9794 7982 -9782
rect 7924 -10050 7936 -9794
rect 7970 -10050 7982 -9794
rect 7924 -10062 7982 -10050
rect 8102 -9794 8160 -9782
rect 8102 -10050 8114 -9794
rect 8148 -10050 8160 -9794
rect 8102 -10062 8160 -10050
rect 8280 -9794 8338 -9782
rect 8280 -10050 8292 -9794
rect 8326 -10050 8338 -9794
rect 8280 -10062 8338 -10050
rect 8458 -9794 8516 -9782
rect 8458 -10050 8470 -9794
rect 8504 -10050 8516 -9794
rect 8458 -10062 8516 -10050
rect 8636 -9794 8694 -9782
rect 8636 -10050 8648 -9794
rect 8682 -10050 8694 -9794
rect 8636 -10062 8694 -10050
rect 8814 -9794 8872 -9782
rect 8814 -10050 8826 -9794
rect 8860 -10050 8872 -9794
rect 8814 -10062 8872 -10050
rect 8992 -9794 9050 -9782
rect 8992 -10050 9004 -9794
rect 9038 -10050 9050 -9794
rect 8992 -10062 9050 -10050
rect 9170 -9794 9228 -9782
rect 9170 -10050 9182 -9794
rect 9216 -10050 9228 -9794
rect 9170 -10062 9228 -10050
rect 9348 -9794 9406 -9782
rect 9348 -10050 9360 -9794
rect 9394 -10050 9406 -9794
rect 10760 -9950 10772 -9694
rect 10806 -9950 10818 -9694
rect 10760 -9962 10818 -9950
rect 10938 -9694 10996 -9682
rect 10938 -9950 10950 -9694
rect 10984 -9950 10996 -9694
rect 10938 -9962 10996 -9950
rect 11052 -9694 11110 -9682
rect 11052 -9950 11064 -9694
rect 11098 -9950 11110 -9694
rect 11052 -9962 11110 -9950
rect 11230 -9694 11288 -9682
rect 11230 -9950 11242 -9694
rect 11276 -9950 11288 -9694
rect 11230 -9962 11288 -9950
rect 11344 -9694 11402 -9682
rect 11344 -9950 11356 -9694
rect 11390 -9950 11402 -9694
rect 11344 -9962 11402 -9950
rect 11522 -9694 11580 -9682
rect 11522 -9950 11534 -9694
rect 11568 -9950 11580 -9694
rect 11522 -9962 11580 -9950
rect 11636 -9694 11694 -9682
rect 11636 -9950 11648 -9694
rect 11682 -9950 11694 -9694
rect 11636 -9962 11694 -9950
rect 11814 -9694 11872 -9682
rect 11814 -9950 11826 -9694
rect 11860 -9950 11872 -9694
rect 11814 -9962 11872 -9950
rect 11928 -9694 11986 -9682
rect 11928 -9950 11940 -9694
rect 11974 -9950 11986 -9694
rect 11928 -9962 11986 -9950
rect 12106 -9694 12164 -9682
rect 12106 -9950 12118 -9694
rect 12152 -9950 12164 -9694
rect 12106 -9962 12164 -9950
rect 12220 -9694 12278 -9682
rect 12220 -9950 12232 -9694
rect 12266 -9950 12278 -9694
rect 12220 -9962 12278 -9950
rect 12398 -9694 12456 -9682
rect 12398 -9950 12410 -9694
rect 12444 -9950 12456 -9694
rect 12398 -9962 12456 -9950
rect 12512 -9694 12570 -9682
rect 12512 -9950 12524 -9694
rect 12558 -9950 12570 -9694
rect 12512 -9962 12570 -9950
rect 12690 -9694 12748 -9682
rect 12690 -9950 12702 -9694
rect 12736 -9950 12748 -9694
rect 12690 -9962 12748 -9950
rect 9348 -10062 9406 -10050
rect -4038 -10342 -3980 -10330
rect -2185 -10132 -2127 -10120
rect -2185 -10388 -2173 -10132
rect -2139 -10388 -2127 -10132
rect -2185 -10400 -2127 -10388
rect -2007 -10132 -1949 -10120
rect -2007 -10388 -1995 -10132
rect -1961 -10388 -1949 -10132
rect -2007 -10400 -1949 -10388
rect -1829 -10132 -1771 -10120
rect -1829 -10388 -1817 -10132
rect -1783 -10388 -1771 -10132
rect -1829 -10400 -1771 -10388
rect -1651 -10132 -1593 -10120
rect -1651 -10388 -1639 -10132
rect -1605 -10388 -1593 -10132
rect -1651 -10400 -1593 -10388
rect -1473 -10132 -1415 -10120
rect -1473 -10388 -1461 -10132
rect -1427 -10388 -1415 -10132
rect -1473 -10400 -1415 -10388
rect -1295 -10132 -1237 -10120
rect -1295 -10388 -1283 -10132
rect -1249 -10388 -1237 -10132
rect -1295 -10400 -1237 -10388
rect -1117 -10132 -1059 -10120
rect -1117 -10388 -1105 -10132
rect -1071 -10388 -1059 -10132
rect -1117 -10400 -1059 -10388
rect -939 -10132 -881 -10120
rect -939 -10388 -927 -10132
rect -893 -10388 -881 -10132
rect -939 -10400 -881 -10388
rect -761 -10132 -703 -10120
rect -761 -10388 -749 -10132
rect -715 -10388 -703 -10132
rect -761 -10400 -703 -10388
rect -583 -10132 -525 -10120
rect -583 -10388 -571 -10132
rect -537 -10388 -525 -10132
rect -583 -10400 -525 -10388
rect -405 -10132 -347 -10120
rect -405 -10388 -393 -10132
rect -359 -10388 -347 -10132
rect -405 -10400 -347 -10388
rect -227 -10132 -169 -10120
rect -227 -10388 -215 -10132
rect -181 -10388 -169 -10132
rect -227 -10400 -169 -10388
rect -49 -10132 9 -10120
rect -49 -10388 -37 -10132
rect -3 -10388 9 -10132
rect -49 -10400 9 -10388
rect 129 -10132 187 -10120
rect 129 -10388 141 -10132
rect 175 -10388 187 -10132
rect 129 -10400 187 -10388
rect 307 -10132 365 -10120
rect 307 -10388 319 -10132
rect 353 -10388 365 -10132
rect 307 -10400 365 -10388
rect 485 -10132 543 -10120
rect 485 -10388 497 -10132
rect 531 -10388 543 -10132
rect 485 -10400 543 -10388
rect 663 -10132 721 -10120
rect 663 -10388 675 -10132
rect 709 -10388 721 -10132
rect 663 -10400 721 -10388
rect 841 -10132 899 -10120
rect 841 -10388 853 -10132
rect 887 -10388 899 -10132
rect 841 -10400 899 -10388
rect 1019 -10132 1077 -10120
rect 1019 -10388 1031 -10132
rect 1065 -10388 1077 -10132
rect 1019 -10400 1077 -10388
rect 1197 -10132 1255 -10120
rect 1197 -10388 1209 -10132
rect 1243 -10388 1255 -10132
rect 1197 -10400 1255 -10388
rect 1375 -10132 1433 -10120
rect 1375 -10388 1387 -10132
rect 1421 -10388 1433 -10132
rect 1375 -10400 1433 -10388
rect 1553 -10132 1611 -10120
rect 1553 -10388 1565 -10132
rect 1599 -10388 1611 -10132
rect 1553 -10400 1611 -10388
rect 1731 -10132 1789 -10120
rect 1731 -10388 1743 -10132
rect 1777 -10388 1789 -10132
rect 1731 -10400 1789 -10388
rect 1909 -10132 1967 -10120
rect 1909 -10388 1921 -10132
rect 1955 -10388 1967 -10132
rect 1909 -10400 1967 -10388
rect 2087 -10132 2145 -10120
rect 2087 -10388 2099 -10132
rect 2133 -10388 2145 -10132
rect 2087 -10400 2145 -10388
rect 2265 -10132 2323 -10120
rect 2265 -10388 2277 -10132
rect 2311 -10388 2323 -10132
rect 2265 -10400 2323 -10388
rect 2443 -10132 2501 -10120
rect 2443 -10388 2455 -10132
rect 2489 -10388 2501 -10132
rect 2443 -10400 2501 -10388
rect 2621 -10132 2679 -10120
rect 2621 -10388 2633 -10132
rect 2667 -10388 2679 -10132
rect 2621 -10400 2679 -10388
rect 2799 -10132 2857 -10120
rect 2799 -10388 2811 -10132
rect 2845 -10388 2857 -10132
rect 2799 -10400 2857 -10388
rect 2977 -10132 3035 -10120
rect 2977 -10388 2989 -10132
rect 3023 -10388 3035 -10132
rect 2977 -10400 3035 -10388
rect 3155 -10132 3213 -10120
rect 3155 -10388 3167 -10132
rect 3201 -10388 3213 -10132
rect 3155 -10400 3213 -10388
rect 3333 -10132 3391 -10120
rect 3333 -10388 3345 -10132
rect 3379 -10388 3391 -10132
rect 3333 -10400 3391 -10388
rect 3511 -10132 3569 -10120
rect 3511 -10388 3523 -10132
rect 3557 -10388 3569 -10132
rect 3511 -10400 3569 -10388
rect 3689 -10132 3747 -10120
rect 3689 -10388 3701 -10132
rect 3735 -10388 3747 -10132
rect 3689 -10400 3747 -10388
rect 3867 -10132 3925 -10120
rect 3867 -10388 3879 -10132
rect 3913 -10388 3925 -10132
rect 3867 -10400 3925 -10388
rect 4045 -10132 4103 -10120
rect 4045 -10388 4057 -10132
rect 4091 -10388 4103 -10132
rect 4045 -10400 4103 -10388
rect 10760 -10464 10818 -10452
rect -5640 -10624 -5582 -10612
rect -5640 -10880 -5628 -10624
rect -5594 -10880 -5582 -10624
rect -5640 -10892 -5582 -10880
rect -5462 -10624 -5404 -10612
rect -5462 -10880 -5450 -10624
rect -5416 -10880 -5404 -10624
rect -5462 -10892 -5404 -10880
rect -5284 -10624 -5226 -10612
rect -5284 -10880 -5272 -10624
rect -5238 -10880 -5226 -10624
rect -5284 -10892 -5226 -10880
rect -5106 -10624 -5048 -10612
rect -5106 -10880 -5094 -10624
rect -5060 -10880 -5048 -10624
rect -5106 -10892 -5048 -10880
rect -4928 -10624 -4870 -10612
rect -4928 -10880 -4916 -10624
rect -4882 -10880 -4870 -10624
rect -4928 -10892 -4870 -10880
rect -4750 -10624 -4692 -10612
rect -4750 -10880 -4738 -10624
rect -4704 -10880 -4692 -10624
rect -4750 -10892 -4692 -10880
rect -4572 -10624 -4514 -10612
rect -4572 -10880 -4560 -10624
rect -4526 -10880 -4514 -10624
rect -4572 -10892 -4514 -10880
rect -4394 -10624 -4336 -10612
rect -4394 -10880 -4382 -10624
rect -4348 -10880 -4336 -10624
rect -4394 -10892 -4336 -10880
rect -4216 -10624 -4158 -10612
rect -4216 -10880 -4204 -10624
rect -4170 -10880 -4158 -10624
rect -4216 -10892 -4158 -10880
rect -4038 -10624 -3980 -10612
rect -4038 -10880 -4026 -10624
rect -3992 -10880 -3980 -10624
rect -4038 -10892 -3980 -10880
rect 6500 -10694 6558 -10682
rect 6500 -10950 6512 -10694
rect 6546 -10950 6558 -10694
rect 6500 -10962 6558 -10950
rect 6678 -10694 6736 -10682
rect 6678 -10950 6690 -10694
rect 6724 -10950 6736 -10694
rect 6678 -10962 6736 -10950
rect 6856 -10694 6914 -10682
rect 6856 -10950 6868 -10694
rect 6902 -10950 6914 -10694
rect 6856 -10962 6914 -10950
rect 7034 -10694 7092 -10682
rect 7034 -10950 7046 -10694
rect 7080 -10950 7092 -10694
rect 7034 -10962 7092 -10950
rect 7212 -10694 7270 -10682
rect 7212 -10950 7224 -10694
rect 7258 -10950 7270 -10694
rect 7212 -10962 7270 -10950
rect 7390 -10694 7448 -10682
rect 7390 -10950 7402 -10694
rect 7436 -10950 7448 -10694
rect 7390 -10962 7448 -10950
rect 7568 -10694 7626 -10682
rect 7568 -10950 7580 -10694
rect 7614 -10950 7626 -10694
rect 7568 -10962 7626 -10950
rect 7746 -10694 7804 -10682
rect 7746 -10950 7758 -10694
rect 7792 -10950 7804 -10694
rect 7746 -10962 7804 -10950
rect 7924 -10694 7982 -10682
rect 7924 -10950 7936 -10694
rect 7970 -10950 7982 -10694
rect 7924 -10962 7982 -10950
rect 8102 -10694 8160 -10682
rect 8102 -10950 8114 -10694
rect 8148 -10950 8160 -10694
rect 8102 -10962 8160 -10950
rect 8280 -10694 8338 -10682
rect 8280 -10950 8292 -10694
rect 8326 -10950 8338 -10694
rect 8280 -10962 8338 -10950
rect 8458 -10694 8516 -10682
rect 8458 -10950 8470 -10694
rect 8504 -10950 8516 -10694
rect 8458 -10962 8516 -10950
rect 8636 -10694 8694 -10682
rect 8636 -10950 8648 -10694
rect 8682 -10950 8694 -10694
rect 8636 -10962 8694 -10950
rect 8814 -10694 8872 -10682
rect 8814 -10950 8826 -10694
rect 8860 -10950 8872 -10694
rect 8814 -10962 8872 -10950
rect 8992 -10694 9050 -10682
rect 8992 -10950 9004 -10694
rect 9038 -10950 9050 -10694
rect 8992 -10962 9050 -10950
rect 9170 -10694 9228 -10682
rect 9170 -10950 9182 -10694
rect 9216 -10950 9228 -10694
rect 9170 -10962 9228 -10950
rect 9348 -10694 9406 -10682
rect 9348 -10950 9360 -10694
rect 9394 -10950 9406 -10694
rect 10760 -10720 10772 -10464
rect 10806 -10720 10818 -10464
rect 10760 -10732 10818 -10720
rect 10938 -10464 10996 -10452
rect 10938 -10720 10950 -10464
rect 10984 -10720 10996 -10464
rect 10938 -10732 10996 -10720
rect 11052 -10464 11110 -10452
rect 11052 -10720 11064 -10464
rect 11098 -10720 11110 -10464
rect 11052 -10732 11110 -10720
rect 11230 -10464 11288 -10452
rect 11230 -10720 11242 -10464
rect 11276 -10720 11288 -10464
rect 11230 -10732 11288 -10720
rect 11344 -10464 11402 -10452
rect 11344 -10720 11356 -10464
rect 11390 -10720 11402 -10464
rect 11344 -10732 11402 -10720
rect 11522 -10464 11580 -10452
rect 11522 -10720 11534 -10464
rect 11568 -10720 11580 -10464
rect 11522 -10732 11580 -10720
rect 11636 -10464 11694 -10452
rect 11636 -10720 11648 -10464
rect 11682 -10720 11694 -10464
rect 11636 -10732 11694 -10720
rect 11814 -10464 11872 -10452
rect 11814 -10720 11826 -10464
rect 11860 -10720 11872 -10464
rect 11814 -10732 11872 -10720
rect 11928 -10464 11986 -10452
rect 11928 -10720 11940 -10464
rect 11974 -10720 11986 -10464
rect 11928 -10732 11986 -10720
rect 12106 -10464 12164 -10452
rect 12106 -10720 12118 -10464
rect 12152 -10720 12164 -10464
rect 12106 -10732 12164 -10720
rect 12220 -10464 12278 -10452
rect 12220 -10720 12232 -10464
rect 12266 -10720 12278 -10464
rect 12220 -10732 12278 -10720
rect 12398 -10464 12456 -10452
rect 12398 -10720 12410 -10464
rect 12444 -10720 12456 -10464
rect 12398 -10732 12456 -10720
rect 12512 -10464 12570 -10452
rect 12512 -10720 12524 -10464
rect 12558 -10720 12570 -10464
rect 12512 -10732 12570 -10720
rect 12690 -10464 12748 -10452
rect 12690 -10720 12702 -10464
rect 12736 -10720 12748 -10464
rect 12690 -10732 12748 -10720
rect 9348 -10962 9406 -10950
rect -2185 -11132 -2127 -11120
rect -5640 -11174 -5582 -11162
rect -5640 -11430 -5628 -11174
rect -5594 -11430 -5582 -11174
rect -5640 -11442 -5582 -11430
rect -5462 -11174 -5404 -11162
rect -5462 -11430 -5450 -11174
rect -5416 -11430 -5404 -11174
rect -5462 -11442 -5404 -11430
rect -5284 -11174 -5226 -11162
rect -5284 -11430 -5272 -11174
rect -5238 -11430 -5226 -11174
rect -5284 -11442 -5226 -11430
rect -5106 -11174 -5048 -11162
rect -5106 -11430 -5094 -11174
rect -5060 -11430 -5048 -11174
rect -5106 -11442 -5048 -11430
rect -4928 -11174 -4870 -11162
rect -4928 -11430 -4916 -11174
rect -4882 -11430 -4870 -11174
rect -4928 -11442 -4870 -11430
rect -4750 -11174 -4692 -11162
rect -4750 -11430 -4738 -11174
rect -4704 -11430 -4692 -11174
rect -4750 -11442 -4692 -11430
rect -4572 -11174 -4514 -11162
rect -4572 -11430 -4560 -11174
rect -4526 -11430 -4514 -11174
rect -4572 -11442 -4514 -11430
rect -4394 -11174 -4336 -11162
rect -4394 -11430 -4382 -11174
rect -4348 -11430 -4336 -11174
rect -4394 -11442 -4336 -11430
rect -4216 -11174 -4158 -11162
rect -4216 -11430 -4204 -11174
rect -4170 -11430 -4158 -11174
rect -4216 -11442 -4158 -11430
rect -4038 -11174 -3980 -11162
rect -4038 -11430 -4026 -11174
rect -3992 -11430 -3980 -11174
rect -2185 -11388 -2173 -11132
rect -2139 -11388 -2127 -11132
rect -2185 -11400 -2127 -11388
rect -2007 -11132 -1949 -11120
rect -2007 -11388 -1995 -11132
rect -1961 -11388 -1949 -11132
rect -2007 -11400 -1949 -11388
rect -1829 -11132 -1771 -11120
rect -1829 -11388 -1817 -11132
rect -1783 -11388 -1771 -11132
rect -1829 -11400 -1771 -11388
rect -1651 -11132 -1593 -11120
rect -1651 -11388 -1639 -11132
rect -1605 -11388 -1593 -11132
rect -1651 -11400 -1593 -11388
rect -1473 -11132 -1415 -11120
rect -1473 -11388 -1461 -11132
rect -1427 -11388 -1415 -11132
rect -1473 -11400 -1415 -11388
rect -1295 -11132 -1237 -11120
rect -1295 -11388 -1283 -11132
rect -1249 -11388 -1237 -11132
rect -1295 -11400 -1237 -11388
rect -1117 -11132 -1059 -11120
rect -1117 -11388 -1105 -11132
rect -1071 -11388 -1059 -11132
rect -1117 -11400 -1059 -11388
rect -939 -11132 -881 -11120
rect -939 -11388 -927 -11132
rect -893 -11388 -881 -11132
rect -939 -11400 -881 -11388
rect -761 -11132 -703 -11120
rect -761 -11388 -749 -11132
rect -715 -11388 -703 -11132
rect -761 -11400 -703 -11388
rect -583 -11132 -525 -11120
rect -583 -11388 -571 -11132
rect -537 -11388 -525 -11132
rect -583 -11400 -525 -11388
rect -405 -11132 -347 -11120
rect -405 -11388 -393 -11132
rect -359 -11388 -347 -11132
rect -405 -11400 -347 -11388
rect -227 -11132 -169 -11120
rect -227 -11388 -215 -11132
rect -181 -11388 -169 -11132
rect -227 -11400 -169 -11388
rect -49 -11132 9 -11120
rect -49 -11388 -37 -11132
rect -3 -11388 9 -11132
rect -49 -11400 9 -11388
rect 129 -11132 187 -11120
rect 129 -11388 141 -11132
rect 175 -11388 187 -11132
rect 129 -11400 187 -11388
rect 307 -11132 365 -11120
rect 307 -11388 319 -11132
rect 353 -11388 365 -11132
rect 307 -11400 365 -11388
rect 485 -11132 543 -11120
rect 485 -11388 497 -11132
rect 531 -11388 543 -11132
rect 485 -11400 543 -11388
rect 663 -11132 721 -11120
rect 663 -11388 675 -11132
rect 709 -11388 721 -11132
rect 663 -11400 721 -11388
rect 841 -11132 899 -11120
rect 841 -11388 853 -11132
rect 887 -11388 899 -11132
rect 841 -11400 899 -11388
rect 1019 -11132 1077 -11120
rect 1019 -11388 1031 -11132
rect 1065 -11388 1077 -11132
rect 1019 -11400 1077 -11388
rect 1197 -11132 1255 -11120
rect 1197 -11388 1209 -11132
rect 1243 -11388 1255 -11132
rect 1197 -11400 1255 -11388
rect 1375 -11132 1433 -11120
rect 1375 -11388 1387 -11132
rect 1421 -11388 1433 -11132
rect 1375 -11400 1433 -11388
rect 1553 -11132 1611 -11120
rect 1553 -11388 1565 -11132
rect 1599 -11388 1611 -11132
rect 1553 -11400 1611 -11388
rect 1731 -11132 1789 -11120
rect 1731 -11388 1743 -11132
rect 1777 -11388 1789 -11132
rect 1731 -11400 1789 -11388
rect 1909 -11132 1967 -11120
rect 1909 -11388 1921 -11132
rect 1955 -11388 1967 -11132
rect 1909 -11400 1967 -11388
rect 2087 -11132 2145 -11120
rect 2087 -11388 2099 -11132
rect 2133 -11388 2145 -11132
rect 2087 -11400 2145 -11388
rect 2265 -11132 2323 -11120
rect 2265 -11388 2277 -11132
rect 2311 -11388 2323 -11132
rect 2265 -11400 2323 -11388
rect 2443 -11132 2501 -11120
rect 2443 -11388 2455 -11132
rect 2489 -11388 2501 -11132
rect 2443 -11400 2501 -11388
rect 2621 -11132 2679 -11120
rect 2621 -11388 2633 -11132
rect 2667 -11388 2679 -11132
rect 2621 -11400 2679 -11388
rect 2799 -11132 2857 -11120
rect 2799 -11388 2811 -11132
rect 2845 -11388 2857 -11132
rect 2799 -11400 2857 -11388
rect 2977 -11132 3035 -11120
rect 2977 -11388 2989 -11132
rect 3023 -11388 3035 -11132
rect 2977 -11400 3035 -11388
rect 3155 -11132 3213 -11120
rect 3155 -11388 3167 -11132
rect 3201 -11388 3213 -11132
rect 3155 -11400 3213 -11388
rect 3333 -11132 3391 -11120
rect 3333 -11388 3345 -11132
rect 3379 -11388 3391 -11132
rect 3333 -11400 3391 -11388
rect 3511 -11132 3569 -11120
rect 3511 -11388 3523 -11132
rect 3557 -11388 3569 -11132
rect 3511 -11400 3569 -11388
rect 3689 -11132 3747 -11120
rect 3689 -11388 3701 -11132
rect 3735 -11388 3747 -11132
rect 3689 -11400 3747 -11388
rect 3867 -11132 3925 -11120
rect 3867 -11388 3879 -11132
rect 3913 -11388 3925 -11132
rect 3867 -11400 3925 -11388
rect 4045 -11132 4103 -11120
rect 4045 -11388 4057 -11132
rect 4091 -11388 4103 -11132
rect 4045 -11400 4103 -11388
rect 10760 -11234 10818 -11222
rect -4038 -11442 -3980 -11430
rect 10760 -11490 10772 -11234
rect 10806 -11490 10818 -11234
rect 10760 -11502 10818 -11490
rect 10938 -11234 10996 -11222
rect 10938 -11490 10950 -11234
rect 10984 -11490 10996 -11234
rect 10938 -11502 10996 -11490
rect 11052 -11234 11110 -11222
rect 11052 -11490 11064 -11234
rect 11098 -11490 11110 -11234
rect 11052 -11502 11110 -11490
rect 11230 -11234 11288 -11222
rect 11230 -11490 11242 -11234
rect 11276 -11490 11288 -11234
rect 11230 -11502 11288 -11490
rect 11344 -11234 11402 -11222
rect 11344 -11490 11356 -11234
rect 11390 -11490 11402 -11234
rect 11344 -11502 11402 -11490
rect 11522 -11234 11580 -11222
rect 11522 -11490 11534 -11234
rect 11568 -11490 11580 -11234
rect 11522 -11502 11580 -11490
rect 11636 -11234 11694 -11222
rect 11636 -11490 11648 -11234
rect 11682 -11490 11694 -11234
rect 11636 -11502 11694 -11490
rect 11814 -11234 11872 -11222
rect 11814 -11490 11826 -11234
rect 11860 -11490 11872 -11234
rect 11814 -11502 11872 -11490
rect 11928 -11234 11986 -11222
rect 11928 -11490 11940 -11234
rect 11974 -11490 11986 -11234
rect 11928 -11502 11986 -11490
rect 12106 -11234 12164 -11222
rect 12106 -11490 12118 -11234
rect 12152 -11490 12164 -11234
rect 12106 -11502 12164 -11490
rect 12220 -11234 12278 -11222
rect 12220 -11490 12232 -11234
rect 12266 -11490 12278 -11234
rect 12220 -11502 12278 -11490
rect 12398 -11234 12456 -11222
rect 12398 -11490 12410 -11234
rect 12444 -11490 12456 -11234
rect 12398 -11502 12456 -11490
rect 12512 -11234 12570 -11222
rect 12512 -11490 12524 -11234
rect 12558 -11490 12570 -11234
rect 12512 -11502 12570 -11490
rect 12690 -11234 12748 -11222
rect 12690 -11490 12702 -11234
rect 12736 -11490 12748 -11234
rect 12690 -11502 12748 -11490
rect 6500 -11594 6558 -11582
rect -5640 -11724 -5582 -11712
rect -5640 -11980 -5628 -11724
rect -5594 -11980 -5582 -11724
rect -5640 -11992 -5582 -11980
rect -5462 -11724 -5404 -11712
rect -5462 -11980 -5450 -11724
rect -5416 -11980 -5404 -11724
rect -5462 -11992 -5404 -11980
rect -5284 -11724 -5226 -11712
rect -5284 -11980 -5272 -11724
rect -5238 -11980 -5226 -11724
rect -5284 -11992 -5226 -11980
rect -5106 -11724 -5048 -11712
rect -5106 -11980 -5094 -11724
rect -5060 -11980 -5048 -11724
rect -5106 -11992 -5048 -11980
rect -4928 -11724 -4870 -11712
rect -4928 -11980 -4916 -11724
rect -4882 -11980 -4870 -11724
rect -4928 -11992 -4870 -11980
rect -4750 -11724 -4692 -11712
rect -4750 -11980 -4738 -11724
rect -4704 -11980 -4692 -11724
rect -4750 -11992 -4692 -11980
rect -4572 -11724 -4514 -11712
rect -4572 -11980 -4560 -11724
rect -4526 -11980 -4514 -11724
rect -4572 -11992 -4514 -11980
rect -4394 -11724 -4336 -11712
rect -4394 -11980 -4382 -11724
rect -4348 -11980 -4336 -11724
rect -4394 -11992 -4336 -11980
rect -4216 -11724 -4158 -11712
rect -4216 -11980 -4204 -11724
rect -4170 -11980 -4158 -11724
rect -4216 -11992 -4158 -11980
rect -4038 -11724 -3980 -11712
rect -4038 -11980 -4026 -11724
rect -3992 -11980 -3980 -11724
rect 6500 -11850 6512 -11594
rect 6546 -11850 6558 -11594
rect 6500 -11862 6558 -11850
rect 6678 -11594 6736 -11582
rect 6678 -11850 6690 -11594
rect 6724 -11850 6736 -11594
rect 6678 -11862 6736 -11850
rect 6856 -11594 6914 -11582
rect 6856 -11850 6868 -11594
rect 6902 -11850 6914 -11594
rect 6856 -11862 6914 -11850
rect 7034 -11594 7092 -11582
rect 7034 -11850 7046 -11594
rect 7080 -11850 7092 -11594
rect 7034 -11862 7092 -11850
rect 7212 -11594 7270 -11582
rect 7212 -11850 7224 -11594
rect 7258 -11850 7270 -11594
rect 7212 -11862 7270 -11850
rect 7390 -11594 7448 -11582
rect 7390 -11850 7402 -11594
rect 7436 -11850 7448 -11594
rect 7390 -11862 7448 -11850
rect 7568 -11594 7626 -11582
rect 7568 -11850 7580 -11594
rect 7614 -11850 7626 -11594
rect 7568 -11862 7626 -11850
rect 7746 -11594 7804 -11582
rect 7746 -11850 7758 -11594
rect 7792 -11850 7804 -11594
rect 7746 -11862 7804 -11850
rect 7924 -11594 7982 -11582
rect 7924 -11850 7936 -11594
rect 7970 -11850 7982 -11594
rect 7924 -11862 7982 -11850
rect 8102 -11594 8160 -11582
rect 8102 -11850 8114 -11594
rect 8148 -11850 8160 -11594
rect 8102 -11862 8160 -11850
rect 8280 -11594 8338 -11582
rect 8280 -11850 8292 -11594
rect 8326 -11850 8338 -11594
rect 8280 -11862 8338 -11850
rect 8458 -11594 8516 -11582
rect 8458 -11850 8470 -11594
rect 8504 -11850 8516 -11594
rect 8458 -11862 8516 -11850
rect 8636 -11594 8694 -11582
rect 8636 -11850 8648 -11594
rect 8682 -11850 8694 -11594
rect 8636 -11862 8694 -11850
rect 8814 -11594 8872 -11582
rect 8814 -11850 8826 -11594
rect 8860 -11850 8872 -11594
rect 8814 -11862 8872 -11850
rect 8992 -11594 9050 -11582
rect 8992 -11850 9004 -11594
rect 9038 -11850 9050 -11594
rect 8992 -11862 9050 -11850
rect 9170 -11594 9228 -11582
rect 9170 -11850 9182 -11594
rect 9216 -11850 9228 -11594
rect 9170 -11862 9228 -11850
rect 9348 -11594 9406 -11582
rect 9348 -11850 9360 -11594
rect 9394 -11850 9406 -11594
rect 9348 -11862 9406 -11850
rect -4038 -11992 -3980 -11980
rect -2185 -12132 -2127 -12120
rect -2185 -12388 -2173 -12132
rect -2139 -12388 -2127 -12132
rect -2185 -12400 -2127 -12388
rect -2007 -12132 -1949 -12120
rect -2007 -12388 -1995 -12132
rect -1961 -12388 -1949 -12132
rect -2007 -12400 -1949 -12388
rect -1829 -12132 -1771 -12120
rect -1829 -12388 -1817 -12132
rect -1783 -12388 -1771 -12132
rect -1829 -12400 -1771 -12388
rect -1651 -12132 -1593 -12120
rect -1651 -12388 -1639 -12132
rect -1605 -12388 -1593 -12132
rect -1651 -12400 -1593 -12388
rect -1473 -12132 -1415 -12120
rect -1473 -12388 -1461 -12132
rect -1427 -12388 -1415 -12132
rect -1473 -12400 -1415 -12388
rect -1295 -12132 -1237 -12120
rect -1295 -12388 -1283 -12132
rect -1249 -12388 -1237 -12132
rect -1295 -12400 -1237 -12388
rect -1117 -12132 -1059 -12120
rect -1117 -12388 -1105 -12132
rect -1071 -12388 -1059 -12132
rect -1117 -12400 -1059 -12388
rect -939 -12132 -881 -12120
rect -939 -12388 -927 -12132
rect -893 -12388 -881 -12132
rect -939 -12400 -881 -12388
rect -761 -12132 -703 -12120
rect -761 -12388 -749 -12132
rect -715 -12388 -703 -12132
rect -761 -12400 -703 -12388
rect -583 -12132 -525 -12120
rect -583 -12388 -571 -12132
rect -537 -12388 -525 -12132
rect -583 -12400 -525 -12388
rect -405 -12132 -347 -12120
rect -405 -12388 -393 -12132
rect -359 -12388 -347 -12132
rect -405 -12400 -347 -12388
rect -227 -12132 -169 -12120
rect -227 -12388 -215 -12132
rect -181 -12388 -169 -12132
rect -227 -12400 -169 -12388
rect -49 -12132 9 -12120
rect -49 -12388 -37 -12132
rect -3 -12388 9 -12132
rect -49 -12400 9 -12388
rect 129 -12132 187 -12120
rect 129 -12388 141 -12132
rect 175 -12388 187 -12132
rect 129 -12400 187 -12388
rect 307 -12132 365 -12120
rect 307 -12388 319 -12132
rect 353 -12388 365 -12132
rect 307 -12400 365 -12388
rect 485 -12132 543 -12120
rect 485 -12388 497 -12132
rect 531 -12388 543 -12132
rect 485 -12400 543 -12388
rect 663 -12132 721 -12120
rect 663 -12388 675 -12132
rect 709 -12388 721 -12132
rect 663 -12400 721 -12388
rect 841 -12132 899 -12120
rect 841 -12388 853 -12132
rect 887 -12388 899 -12132
rect 841 -12400 899 -12388
rect 1019 -12132 1077 -12120
rect 1019 -12388 1031 -12132
rect 1065 -12388 1077 -12132
rect 1019 -12400 1077 -12388
rect 1197 -12132 1255 -12120
rect 1197 -12388 1209 -12132
rect 1243 -12388 1255 -12132
rect 1197 -12400 1255 -12388
rect 1375 -12132 1433 -12120
rect 1375 -12388 1387 -12132
rect 1421 -12388 1433 -12132
rect 1375 -12400 1433 -12388
rect 1553 -12132 1611 -12120
rect 1553 -12388 1565 -12132
rect 1599 -12388 1611 -12132
rect 1553 -12400 1611 -12388
rect 1731 -12132 1789 -12120
rect 1731 -12388 1743 -12132
rect 1777 -12388 1789 -12132
rect 1731 -12400 1789 -12388
rect 1909 -12132 1967 -12120
rect 1909 -12388 1921 -12132
rect 1955 -12388 1967 -12132
rect 1909 -12400 1967 -12388
rect 2087 -12132 2145 -12120
rect 2087 -12388 2099 -12132
rect 2133 -12388 2145 -12132
rect 2087 -12400 2145 -12388
rect 2265 -12132 2323 -12120
rect 2265 -12388 2277 -12132
rect 2311 -12388 2323 -12132
rect 2265 -12400 2323 -12388
rect 2443 -12132 2501 -12120
rect 2443 -12388 2455 -12132
rect 2489 -12388 2501 -12132
rect 2443 -12400 2501 -12388
rect 2621 -12132 2679 -12120
rect 2621 -12388 2633 -12132
rect 2667 -12388 2679 -12132
rect 2621 -12400 2679 -12388
rect 2799 -12132 2857 -12120
rect 2799 -12388 2811 -12132
rect 2845 -12388 2857 -12132
rect 2799 -12400 2857 -12388
rect 2977 -12132 3035 -12120
rect 2977 -12388 2989 -12132
rect 3023 -12388 3035 -12132
rect 2977 -12400 3035 -12388
rect 3155 -12132 3213 -12120
rect 3155 -12388 3167 -12132
rect 3201 -12388 3213 -12132
rect 3155 -12400 3213 -12388
rect 3333 -12132 3391 -12120
rect 3333 -12388 3345 -12132
rect 3379 -12388 3391 -12132
rect 3333 -12400 3391 -12388
rect 3511 -12132 3569 -12120
rect 3511 -12388 3523 -12132
rect 3557 -12388 3569 -12132
rect 3511 -12400 3569 -12388
rect 3689 -12132 3747 -12120
rect 3689 -12388 3701 -12132
rect 3735 -12388 3747 -12132
rect 3689 -12400 3747 -12388
rect 3867 -12132 3925 -12120
rect 3867 -12388 3879 -12132
rect 3913 -12388 3925 -12132
rect 3867 -12400 3925 -12388
rect 4045 -12132 4103 -12120
rect 4045 -12388 4057 -12132
rect 4091 -12388 4103 -12132
rect 4045 -12400 4103 -12388
rect -5928 -12712 -5870 -12700
rect -5928 -12928 -5916 -12712
rect -5882 -12928 -5870 -12712
rect -5928 -12940 -5870 -12928
rect -5830 -12712 -5772 -12700
rect -5830 -12928 -5818 -12712
rect -5784 -12928 -5772 -12712
rect -5830 -12940 -5772 -12928
rect -5678 -12712 -5620 -12700
rect -5678 -12928 -5666 -12712
rect -5632 -12928 -5620 -12712
rect -5678 -12940 -5620 -12928
rect -5580 -12712 -5522 -12700
rect -5580 -12928 -5568 -12712
rect -5534 -12928 -5522 -12712
rect -5580 -12940 -5522 -12928
rect -5428 -12712 -5370 -12700
rect -5428 -12928 -5416 -12712
rect -5382 -12928 -5370 -12712
rect -5428 -12940 -5370 -12928
rect -5330 -12712 -5272 -12700
rect -5330 -12928 -5318 -12712
rect -5284 -12928 -5272 -12712
rect -5330 -12940 -5272 -12928
rect -5178 -12712 -5120 -12700
rect -5178 -12928 -5166 -12712
rect -5132 -12928 -5120 -12712
rect -5178 -12940 -5120 -12928
rect -5080 -12712 -5022 -12700
rect -5080 -12928 -5068 -12712
rect -5034 -12928 -5022 -12712
rect -5080 -12940 -5022 -12928
rect -4928 -12712 -4870 -12700
rect -4928 -12928 -4916 -12712
rect -4882 -12928 -4870 -12712
rect -4928 -12940 -4870 -12928
rect -4830 -12712 -4772 -12700
rect -4830 -12928 -4818 -12712
rect -4784 -12928 -4772 -12712
rect -4830 -12940 -4772 -12928
rect -4678 -12712 -4620 -12700
rect -4678 -12928 -4666 -12712
rect -4632 -12928 -4620 -12712
rect -4678 -12940 -4620 -12928
rect -4580 -12712 -4522 -12700
rect -4580 -12928 -4568 -12712
rect -4534 -12928 -4522 -12712
rect -4580 -12940 -4522 -12928
rect -4428 -12712 -4370 -12700
rect -4428 -12928 -4416 -12712
rect -4382 -12928 -4370 -12712
rect -4428 -12940 -4370 -12928
rect -4330 -12712 -4272 -12700
rect -4330 -12928 -4318 -12712
rect -4284 -12928 -4272 -12712
rect -4330 -12940 -4272 -12928
rect -4178 -12712 -4120 -12700
rect -4178 -12928 -4166 -12712
rect -4132 -12928 -4120 -12712
rect -4178 -12940 -4120 -12928
rect -4080 -12712 -4022 -12700
rect -4080 -12928 -4068 -12712
rect -4034 -12928 -4022 -12712
rect -4080 -12940 -4022 -12928
rect -2185 -13132 -2127 -13120
rect -5928 -13392 -5870 -13380
rect -5928 -13608 -5916 -13392
rect -5882 -13608 -5870 -13392
rect -5928 -13620 -5870 -13608
rect -5830 -13392 -5772 -13380
rect -5830 -13608 -5818 -13392
rect -5784 -13608 -5772 -13392
rect -5830 -13620 -5772 -13608
rect -5678 -13392 -5620 -13380
rect -5678 -13608 -5666 -13392
rect -5632 -13608 -5620 -13392
rect -5678 -13620 -5620 -13608
rect -5580 -13392 -5522 -13380
rect -5580 -13608 -5568 -13392
rect -5534 -13608 -5522 -13392
rect -5580 -13620 -5522 -13608
rect -5428 -13392 -5370 -13380
rect -5428 -13608 -5416 -13392
rect -5382 -13608 -5370 -13392
rect -5428 -13620 -5370 -13608
rect -5330 -13392 -5272 -13380
rect -5330 -13608 -5318 -13392
rect -5284 -13608 -5272 -13392
rect -5330 -13620 -5272 -13608
rect -5178 -13392 -5120 -13380
rect -5178 -13608 -5166 -13392
rect -5132 -13608 -5120 -13392
rect -5178 -13620 -5120 -13608
rect -5080 -13392 -5022 -13380
rect -5080 -13608 -5068 -13392
rect -5034 -13608 -5022 -13392
rect -5080 -13620 -5022 -13608
rect -4928 -13392 -4870 -13380
rect -4928 -13608 -4916 -13392
rect -4882 -13608 -4870 -13392
rect -4928 -13620 -4870 -13608
rect -4830 -13392 -4772 -13380
rect -4830 -13608 -4818 -13392
rect -4784 -13608 -4772 -13392
rect -4830 -13620 -4772 -13608
rect -4678 -13392 -4620 -13380
rect -4678 -13608 -4666 -13392
rect -4632 -13608 -4620 -13392
rect -4678 -13620 -4620 -13608
rect -4580 -13392 -4522 -13380
rect -4580 -13608 -4568 -13392
rect -4534 -13608 -4522 -13392
rect -4580 -13620 -4522 -13608
rect -4428 -13392 -4370 -13380
rect -4428 -13608 -4416 -13392
rect -4382 -13608 -4370 -13392
rect -4428 -13620 -4370 -13608
rect -4330 -13392 -4272 -13380
rect -4330 -13608 -4318 -13392
rect -4284 -13608 -4272 -13392
rect -4330 -13620 -4272 -13608
rect -4178 -13392 -4120 -13380
rect -4178 -13608 -4166 -13392
rect -4132 -13608 -4120 -13392
rect -4178 -13620 -4120 -13608
rect -4080 -13392 -4022 -13380
rect -4080 -13608 -4068 -13392
rect -4034 -13608 -4022 -13392
rect -2185 -13388 -2173 -13132
rect -2139 -13388 -2127 -13132
rect -2185 -13400 -2127 -13388
rect -2007 -13132 -1949 -13120
rect -2007 -13388 -1995 -13132
rect -1961 -13388 -1949 -13132
rect -2007 -13400 -1949 -13388
rect -1829 -13132 -1771 -13120
rect -1829 -13388 -1817 -13132
rect -1783 -13388 -1771 -13132
rect -1829 -13400 -1771 -13388
rect -1651 -13132 -1593 -13120
rect -1651 -13388 -1639 -13132
rect -1605 -13388 -1593 -13132
rect -1651 -13400 -1593 -13388
rect -1473 -13132 -1415 -13120
rect -1473 -13388 -1461 -13132
rect -1427 -13388 -1415 -13132
rect -1473 -13400 -1415 -13388
rect -1295 -13132 -1237 -13120
rect -1295 -13388 -1283 -13132
rect -1249 -13388 -1237 -13132
rect -1295 -13400 -1237 -13388
rect -1117 -13132 -1059 -13120
rect -1117 -13388 -1105 -13132
rect -1071 -13388 -1059 -13132
rect -1117 -13400 -1059 -13388
rect -939 -13132 -881 -13120
rect -939 -13388 -927 -13132
rect -893 -13388 -881 -13132
rect -939 -13400 -881 -13388
rect -761 -13132 -703 -13120
rect -761 -13388 -749 -13132
rect -715 -13388 -703 -13132
rect -761 -13400 -703 -13388
rect -583 -13132 -525 -13120
rect -583 -13388 -571 -13132
rect -537 -13388 -525 -13132
rect -583 -13400 -525 -13388
rect -405 -13132 -347 -13120
rect -405 -13388 -393 -13132
rect -359 -13388 -347 -13132
rect -405 -13400 -347 -13388
rect -227 -13132 -169 -13120
rect -227 -13388 -215 -13132
rect -181 -13388 -169 -13132
rect -227 -13400 -169 -13388
rect -49 -13132 9 -13120
rect -49 -13388 -37 -13132
rect -3 -13388 9 -13132
rect -49 -13400 9 -13388
rect 129 -13132 187 -13120
rect 129 -13388 141 -13132
rect 175 -13388 187 -13132
rect 129 -13400 187 -13388
rect 307 -13132 365 -13120
rect 307 -13388 319 -13132
rect 353 -13388 365 -13132
rect 307 -13400 365 -13388
rect 485 -13132 543 -13120
rect 485 -13388 497 -13132
rect 531 -13388 543 -13132
rect 485 -13400 543 -13388
rect 663 -13132 721 -13120
rect 663 -13388 675 -13132
rect 709 -13388 721 -13132
rect 663 -13400 721 -13388
rect 841 -13132 899 -13120
rect 841 -13388 853 -13132
rect 887 -13388 899 -13132
rect 841 -13400 899 -13388
rect 1019 -13132 1077 -13120
rect 1019 -13388 1031 -13132
rect 1065 -13388 1077 -13132
rect 1019 -13400 1077 -13388
rect 1197 -13132 1255 -13120
rect 1197 -13388 1209 -13132
rect 1243 -13388 1255 -13132
rect 1197 -13400 1255 -13388
rect 1375 -13132 1433 -13120
rect 1375 -13388 1387 -13132
rect 1421 -13388 1433 -13132
rect 1375 -13400 1433 -13388
rect 1553 -13132 1611 -13120
rect 1553 -13388 1565 -13132
rect 1599 -13388 1611 -13132
rect 1553 -13400 1611 -13388
rect 1731 -13132 1789 -13120
rect 1731 -13388 1743 -13132
rect 1777 -13388 1789 -13132
rect 1731 -13400 1789 -13388
rect 1909 -13132 1967 -13120
rect 1909 -13388 1921 -13132
rect 1955 -13388 1967 -13132
rect 1909 -13400 1967 -13388
rect 2087 -13132 2145 -13120
rect 2087 -13388 2099 -13132
rect 2133 -13388 2145 -13132
rect 2087 -13400 2145 -13388
rect 2265 -13132 2323 -13120
rect 2265 -13388 2277 -13132
rect 2311 -13388 2323 -13132
rect 2265 -13400 2323 -13388
rect 2443 -13132 2501 -13120
rect 2443 -13388 2455 -13132
rect 2489 -13388 2501 -13132
rect 2443 -13400 2501 -13388
rect 2621 -13132 2679 -13120
rect 2621 -13388 2633 -13132
rect 2667 -13388 2679 -13132
rect 2621 -13400 2679 -13388
rect 2799 -13132 2857 -13120
rect 2799 -13388 2811 -13132
rect 2845 -13388 2857 -13132
rect 2799 -13400 2857 -13388
rect 2977 -13132 3035 -13120
rect 2977 -13388 2989 -13132
rect 3023 -13388 3035 -13132
rect 2977 -13400 3035 -13388
rect 3155 -13132 3213 -13120
rect 3155 -13388 3167 -13132
rect 3201 -13388 3213 -13132
rect 3155 -13400 3213 -13388
rect 3333 -13132 3391 -13120
rect 3333 -13388 3345 -13132
rect 3379 -13388 3391 -13132
rect 3333 -13400 3391 -13388
rect 3511 -13132 3569 -13120
rect 3511 -13388 3523 -13132
rect 3557 -13388 3569 -13132
rect 3511 -13400 3569 -13388
rect 3689 -13132 3747 -13120
rect 3689 -13388 3701 -13132
rect 3735 -13388 3747 -13132
rect 3689 -13400 3747 -13388
rect 3867 -13132 3925 -13120
rect 3867 -13388 3879 -13132
rect 3913 -13388 3925 -13132
rect 3867 -13400 3925 -13388
rect 4045 -13132 4103 -13120
rect 4045 -13388 4057 -13132
rect 4091 -13388 4103 -13132
rect 4045 -13400 4103 -13388
rect -4080 -13620 -4022 -13608
rect -2185 -14132 -2127 -14120
rect -6040 -14394 -5982 -14382
rect -6040 -14650 -6028 -14394
rect -5994 -14650 -5982 -14394
rect -6040 -14662 -5982 -14650
rect -5862 -14394 -5804 -14382
rect -5862 -14650 -5850 -14394
rect -5816 -14650 -5804 -14394
rect -5862 -14662 -5804 -14650
rect -5684 -14394 -5626 -14382
rect -5684 -14650 -5672 -14394
rect -5638 -14650 -5626 -14394
rect -5684 -14662 -5626 -14650
rect -5506 -14394 -5448 -14382
rect -5506 -14650 -5494 -14394
rect -5460 -14650 -5448 -14394
rect -5506 -14662 -5448 -14650
rect -5328 -14394 -5270 -14382
rect -5328 -14650 -5316 -14394
rect -5282 -14650 -5270 -14394
rect -5328 -14662 -5270 -14650
rect -5150 -14394 -5092 -14382
rect -5150 -14650 -5138 -14394
rect -5104 -14650 -5092 -14394
rect -5150 -14662 -5092 -14650
rect -4972 -14394 -4914 -14382
rect -4972 -14650 -4960 -14394
rect -4926 -14650 -4914 -14394
rect -4972 -14662 -4914 -14650
rect -4794 -14394 -4736 -14382
rect -4794 -14650 -4782 -14394
rect -4748 -14650 -4736 -14394
rect -4794 -14662 -4736 -14650
rect -4616 -14394 -4558 -14382
rect -4616 -14650 -4604 -14394
rect -4570 -14650 -4558 -14394
rect -4616 -14662 -4558 -14650
rect -4438 -14394 -4380 -14382
rect -4438 -14650 -4426 -14394
rect -4392 -14650 -4380 -14394
rect -4438 -14662 -4380 -14650
rect -4260 -14394 -4202 -14382
rect -4260 -14650 -4248 -14394
rect -4214 -14650 -4202 -14394
rect -4260 -14662 -4202 -14650
rect -4082 -14394 -4024 -14382
rect -4082 -14650 -4070 -14394
rect -4036 -14650 -4024 -14394
rect -2185 -14388 -2173 -14132
rect -2139 -14388 -2127 -14132
rect -2185 -14400 -2127 -14388
rect -2007 -14132 -1949 -14120
rect -2007 -14388 -1995 -14132
rect -1961 -14388 -1949 -14132
rect -2007 -14400 -1949 -14388
rect -1829 -14132 -1771 -14120
rect -1829 -14388 -1817 -14132
rect -1783 -14388 -1771 -14132
rect -1829 -14400 -1771 -14388
rect -1651 -14132 -1593 -14120
rect -1651 -14388 -1639 -14132
rect -1605 -14388 -1593 -14132
rect -1651 -14400 -1593 -14388
rect -1473 -14132 -1415 -14120
rect -1473 -14388 -1461 -14132
rect -1427 -14388 -1415 -14132
rect -1473 -14400 -1415 -14388
rect -1295 -14132 -1237 -14120
rect -1295 -14388 -1283 -14132
rect -1249 -14388 -1237 -14132
rect -1295 -14400 -1237 -14388
rect -1117 -14132 -1059 -14120
rect -1117 -14388 -1105 -14132
rect -1071 -14388 -1059 -14132
rect -1117 -14400 -1059 -14388
rect -939 -14132 -881 -14120
rect -939 -14388 -927 -14132
rect -893 -14388 -881 -14132
rect -939 -14400 -881 -14388
rect -761 -14132 -703 -14120
rect -761 -14388 -749 -14132
rect -715 -14388 -703 -14132
rect -761 -14400 -703 -14388
rect -583 -14132 -525 -14120
rect -583 -14388 -571 -14132
rect -537 -14388 -525 -14132
rect -583 -14400 -525 -14388
rect -405 -14132 -347 -14120
rect -405 -14388 -393 -14132
rect -359 -14388 -347 -14132
rect -405 -14400 -347 -14388
rect -227 -14132 -169 -14120
rect -227 -14388 -215 -14132
rect -181 -14388 -169 -14132
rect -227 -14400 -169 -14388
rect -49 -14132 9 -14120
rect -49 -14388 -37 -14132
rect -3 -14388 9 -14132
rect -49 -14400 9 -14388
rect 129 -14132 187 -14120
rect 129 -14388 141 -14132
rect 175 -14388 187 -14132
rect 129 -14400 187 -14388
rect 307 -14132 365 -14120
rect 307 -14388 319 -14132
rect 353 -14388 365 -14132
rect 307 -14400 365 -14388
rect 485 -14132 543 -14120
rect 485 -14388 497 -14132
rect 531 -14388 543 -14132
rect 485 -14400 543 -14388
rect 663 -14132 721 -14120
rect 663 -14388 675 -14132
rect 709 -14388 721 -14132
rect 663 -14400 721 -14388
rect 841 -14132 899 -14120
rect 841 -14388 853 -14132
rect 887 -14388 899 -14132
rect 841 -14400 899 -14388
rect 1019 -14132 1077 -14120
rect 1019 -14388 1031 -14132
rect 1065 -14388 1077 -14132
rect 1019 -14400 1077 -14388
rect 1197 -14132 1255 -14120
rect 1197 -14388 1209 -14132
rect 1243 -14388 1255 -14132
rect 1197 -14400 1255 -14388
rect 1375 -14132 1433 -14120
rect 1375 -14388 1387 -14132
rect 1421 -14388 1433 -14132
rect 1375 -14400 1433 -14388
rect 1553 -14132 1611 -14120
rect 1553 -14388 1565 -14132
rect 1599 -14388 1611 -14132
rect 1553 -14400 1611 -14388
rect 1731 -14132 1789 -14120
rect 1731 -14388 1743 -14132
rect 1777 -14388 1789 -14132
rect 1731 -14400 1789 -14388
rect 1909 -14132 1967 -14120
rect 1909 -14388 1921 -14132
rect 1955 -14388 1967 -14132
rect 1909 -14400 1967 -14388
rect 2087 -14132 2145 -14120
rect 2087 -14388 2099 -14132
rect 2133 -14388 2145 -14132
rect 2087 -14400 2145 -14388
rect 2265 -14132 2323 -14120
rect 2265 -14388 2277 -14132
rect 2311 -14388 2323 -14132
rect 2265 -14400 2323 -14388
rect 2443 -14132 2501 -14120
rect 2443 -14388 2455 -14132
rect 2489 -14388 2501 -14132
rect 2443 -14400 2501 -14388
rect 2621 -14132 2679 -14120
rect 2621 -14388 2633 -14132
rect 2667 -14388 2679 -14132
rect 2621 -14400 2679 -14388
rect 2799 -14132 2857 -14120
rect 2799 -14388 2811 -14132
rect 2845 -14388 2857 -14132
rect 2799 -14400 2857 -14388
rect 2977 -14132 3035 -14120
rect 2977 -14388 2989 -14132
rect 3023 -14388 3035 -14132
rect 2977 -14400 3035 -14388
rect 3155 -14132 3213 -14120
rect 3155 -14388 3167 -14132
rect 3201 -14388 3213 -14132
rect 3155 -14400 3213 -14388
rect 3333 -14132 3391 -14120
rect 3333 -14388 3345 -14132
rect 3379 -14388 3391 -14132
rect 3333 -14400 3391 -14388
rect 3511 -14132 3569 -14120
rect 3511 -14388 3523 -14132
rect 3557 -14388 3569 -14132
rect 3511 -14400 3569 -14388
rect 3689 -14132 3747 -14120
rect 3689 -14388 3701 -14132
rect 3735 -14388 3747 -14132
rect 3689 -14400 3747 -14388
rect 3867 -14132 3925 -14120
rect 3867 -14388 3879 -14132
rect 3913 -14388 3925 -14132
rect 3867 -14400 3925 -14388
rect 4045 -14132 4103 -14120
rect 4045 -14388 4057 -14132
rect 4091 -14388 4103 -14132
rect 4045 -14400 4103 -14388
rect 5565 -14132 5623 -14120
rect 5565 -14388 5577 -14132
rect 5611 -14388 5623 -14132
rect 5565 -14400 5623 -14388
rect 5743 -14132 5801 -14120
rect 5743 -14388 5755 -14132
rect 5789 -14388 5801 -14132
rect 5743 -14400 5801 -14388
rect 5921 -14132 5979 -14120
rect 5921 -14388 5933 -14132
rect 5967 -14388 5979 -14132
rect 5921 -14400 5979 -14388
rect 6099 -14132 6157 -14120
rect 6099 -14388 6111 -14132
rect 6145 -14388 6157 -14132
rect 6099 -14400 6157 -14388
rect 6277 -14132 6335 -14120
rect 6277 -14388 6289 -14132
rect 6323 -14388 6335 -14132
rect 6277 -14400 6335 -14388
rect 6455 -14132 6513 -14120
rect 6455 -14388 6467 -14132
rect 6501 -14388 6513 -14132
rect 6455 -14400 6513 -14388
rect 6633 -14132 6691 -14120
rect 6633 -14388 6645 -14132
rect 6679 -14388 6691 -14132
rect 6633 -14400 6691 -14388
rect 6811 -14132 6869 -14120
rect 6811 -14388 6823 -14132
rect 6857 -14388 6869 -14132
rect 6811 -14400 6869 -14388
rect 6989 -14132 7047 -14120
rect 6989 -14388 7001 -14132
rect 7035 -14388 7047 -14132
rect 6989 -14400 7047 -14388
rect 7167 -14132 7225 -14120
rect 7167 -14388 7179 -14132
rect 7213 -14388 7225 -14132
rect 7167 -14400 7225 -14388
rect 7345 -14132 7403 -14120
rect 7345 -14388 7357 -14132
rect 7391 -14388 7403 -14132
rect 7345 -14400 7403 -14388
rect 7523 -14132 7581 -14120
rect 7523 -14388 7535 -14132
rect 7569 -14388 7581 -14132
rect 7523 -14400 7581 -14388
rect 7701 -14132 7759 -14120
rect 7701 -14388 7713 -14132
rect 7747 -14388 7759 -14132
rect 7701 -14400 7759 -14388
rect 7879 -14132 7937 -14120
rect 7879 -14388 7891 -14132
rect 7925 -14388 7937 -14132
rect 7879 -14400 7937 -14388
rect 8057 -14132 8115 -14120
rect 8057 -14388 8069 -14132
rect 8103 -14388 8115 -14132
rect 8057 -14400 8115 -14388
rect 8235 -14132 8293 -14120
rect 8235 -14388 8247 -14132
rect 8281 -14388 8293 -14132
rect 8235 -14400 8293 -14388
rect 8413 -14132 8471 -14120
rect 8413 -14388 8425 -14132
rect 8459 -14388 8471 -14132
rect 8413 -14400 8471 -14388
rect 8591 -14132 8649 -14120
rect 8591 -14388 8603 -14132
rect 8637 -14388 8649 -14132
rect 8591 -14400 8649 -14388
rect 8769 -14132 8827 -14120
rect 8769 -14388 8781 -14132
rect 8815 -14388 8827 -14132
rect 8769 -14400 8827 -14388
rect 8947 -14132 9005 -14120
rect 8947 -14388 8959 -14132
rect 8993 -14388 9005 -14132
rect 8947 -14400 9005 -14388
rect 9125 -14132 9183 -14120
rect 9125 -14388 9137 -14132
rect 9171 -14388 9183 -14132
rect 9125 -14400 9183 -14388
rect 9303 -14132 9361 -14120
rect 9303 -14388 9315 -14132
rect 9349 -14388 9361 -14132
rect 9303 -14400 9361 -14388
rect 9481 -14132 9539 -14120
rect 9481 -14388 9493 -14132
rect 9527 -14388 9539 -14132
rect 9481 -14400 9539 -14388
rect 9659 -14132 9717 -14120
rect 9659 -14388 9671 -14132
rect 9705 -14388 9717 -14132
rect 9659 -14400 9717 -14388
rect 9837 -14132 9895 -14120
rect 9837 -14388 9849 -14132
rect 9883 -14388 9895 -14132
rect 9837 -14400 9895 -14388
rect 10015 -14132 10073 -14120
rect 10015 -14388 10027 -14132
rect 10061 -14388 10073 -14132
rect 10015 -14400 10073 -14388
rect 10193 -14132 10251 -14120
rect 10193 -14388 10205 -14132
rect 10239 -14388 10251 -14132
rect 10193 -14400 10251 -14388
rect 10371 -14132 10429 -14120
rect 10371 -14388 10383 -14132
rect 10417 -14388 10429 -14132
rect 10371 -14400 10429 -14388
rect 10549 -14132 10607 -14120
rect 10549 -14388 10561 -14132
rect 10595 -14388 10607 -14132
rect 10549 -14400 10607 -14388
rect 10727 -14132 10785 -14120
rect 10727 -14388 10739 -14132
rect 10773 -14388 10785 -14132
rect 10727 -14400 10785 -14388
rect 10905 -14132 10963 -14120
rect 10905 -14388 10917 -14132
rect 10951 -14388 10963 -14132
rect 10905 -14400 10963 -14388
rect 11083 -14132 11141 -14120
rect 11083 -14388 11095 -14132
rect 11129 -14388 11141 -14132
rect 11083 -14400 11141 -14388
rect 11261 -14132 11319 -14120
rect 11261 -14388 11273 -14132
rect 11307 -14388 11319 -14132
rect 11261 -14400 11319 -14388
rect 11439 -14132 11497 -14120
rect 11439 -14388 11451 -14132
rect 11485 -14388 11497 -14132
rect 11439 -14400 11497 -14388
rect 11617 -14132 11675 -14120
rect 11617 -14388 11629 -14132
rect 11663 -14388 11675 -14132
rect 11617 -14400 11675 -14388
rect 11795 -14132 11853 -14120
rect 11795 -14388 11807 -14132
rect 11841 -14388 11853 -14132
rect 11795 -14400 11853 -14388
rect 11973 -14132 12031 -14120
rect 11973 -14388 11985 -14132
rect 12019 -14388 12031 -14132
rect 11973 -14400 12031 -14388
rect 12151 -14132 12209 -14120
rect 12151 -14388 12163 -14132
rect 12197 -14388 12209 -14132
rect 12151 -14400 12209 -14388
rect 12329 -14132 12387 -14120
rect 12329 -14388 12341 -14132
rect 12375 -14388 12387 -14132
rect 12329 -14400 12387 -14388
rect 12507 -14132 12565 -14120
rect 12507 -14388 12519 -14132
rect 12553 -14388 12565 -14132
rect 12507 -14400 12565 -14388
rect 12685 -14132 12743 -14120
rect 12685 -14388 12697 -14132
rect 12731 -14388 12743 -14132
rect 12685 -14400 12743 -14388
rect -4082 -14662 -4024 -14650
rect -6040 -15094 -5982 -15082
rect -6040 -15350 -6028 -15094
rect -5994 -15350 -5982 -15094
rect -6040 -15362 -5982 -15350
rect -5862 -15094 -5804 -15082
rect -5862 -15350 -5850 -15094
rect -5816 -15350 -5804 -15094
rect -5862 -15362 -5804 -15350
rect -5684 -15094 -5626 -15082
rect -5684 -15350 -5672 -15094
rect -5638 -15350 -5626 -15094
rect -5684 -15362 -5626 -15350
rect -5506 -15094 -5448 -15082
rect -5506 -15350 -5494 -15094
rect -5460 -15350 -5448 -15094
rect -5506 -15362 -5448 -15350
rect -5328 -15094 -5270 -15082
rect -5328 -15350 -5316 -15094
rect -5282 -15350 -5270 -15094
rect -5328 -15362 -5270 -15350
rect -5150 -15094 -5092 -15082
rect -5150 -15350 -5138 -15094
rect -5104 -15350 -5092 -15094
rect -5150 -15362 -5092 -15350
rect -4972 -15094 -4914 -15082
rect -4972 -15350 -4960 -15094
rect -4926 -15350 -4914 -15094
rect -4972 -15362 -4914 -15350
rect -4794 -15094 -4736 -15082
rect -4794 -15350 -4782 -15094
rect -4748 -15350 -4736 -15094
rect -4794 -15362 -4736 -15350
rect -4616 -15094 -4558 -15082
rect -4616 -15350 -4604 -15094
rect -4570 -15350 -4558 -15094
rect -4616 -15362 -4558 -15350
rect -4438 -15094 -4380 -15082
rect -4438 -15350 -4426 -15094
rect -4392 -15350 -4380 -15094
rect -4438 -15362 -4380 -15350
rect -4260 -15094 -4202 -15082
rect -4260 -15350 -4248 -15094
rect -4214 -15350 -4202 -15094
rect -4260 -15362 -4202 -15350
rect -4082 -15094 -4024 -15082
rect -4082 -15350 -4070 -15094
rect -4036 -15350 -4024 -15094
rect -4082 -15362 -4024 -15350
rect -2185 -15132 -2127 -15120
rect -2185 -15388 -2173 -15132
rect -2139 -15388 -2127 -15132
rect -2185 -15400 -2127 -15388
rect -2007 -15132 -1949 -15120
rect -2007 -15388 -1995 -15132
rect -1961 -15388 -1949 -15132
rect -2007 -15400 -1949 -15388
rect -1829 -15132 -1771 -15120
rect -1829 -15388 -1817 -15132
rect -1783 -15388 -1771 -15132
rect -1829 -15400 -1771 -15388
rect -1651 -15132 -1593 -15120
rect -1651 -15388 -1639 -15132
rect -1605 -15388 -1593 -15132
rect -1651 -15400 -1593 -15388
rect -1473 -15132 -1415 -15120
rect -1473 -15388 -1461 -15132
rect -1427 -15388 -1415 -15132
rect -1473 -15400 -1415 -15388
rect -1295 -15132 -1237 -15120
rect -1295 -15388 -1283 -15132
rect -1249 -15388 -1237 -15132
rect -1295 -15400 -1237 -15388
rect -1117 -15132 -1059 -15120
rect -1117 -15388 -1105 -15132
rect -1071 -15388 -1059 -15132
rect -1117 -15400 -1059 -15388
rect -939 -15132 -881 -15120
rect -939 -15388 -927 -15132
rect -893 -15388 -881 -15132
rect -939 -15400 -881 -15388
rect -761 -15132 -703 -15120
rect -761 -15388 -749 -15132
rect -715 -15388 -703 -15132
rect -761 -15400 -703 -15388
rect -583 -15132 -525 -15120
rect -583 -15388 -571 -15132
rect -537 -15388 -525 -15132
rect -583 -15400 -525 -15388
rect -405 -15132 -347 -15120
rect -405 -15388 -393 -15132
rect -359 -15388 -347 -15132
rect -405 -15400 -347 -15388
rect -227 -15132 -169 -15120
rect -227 -15388 -215 -15132
rect -181 -15388 -169 -15132
rect -227 -15400 -169 -15388
rect -49 -15132 9 -15120
rect -49 -15388 -37 -15132
rect -3 -15388 9 -15132
rect -49 -15400 9 -15388
rect 129 -15132 187 -15120
rect 129 -15388 141 -15132
rect 175 -15388 187 -15132
rect 129 -15400 187 -15388
rect 307 -15132 365 -15120
rect 307 -15388 319 -15132
rect 353 -15388 365 -15132
rect 307 -15400 365 -15388
rect 485 -15132 543 -15120
rect 485 -15388 497 -15132
rect 531 -15388 543 -15132
rect 485 -15400 543 -15388
rect 663 -15132 721 -15120
rect 663 -15388 675 -15132
rect 709 -15388 721 -15132
rect 663 -15400 721 -15388
rect 841 -15132 899 -15120
rect 841 -15388 853 -15132
rect 887 -15388 899 -15132
rect 841 -15400 899 -15388
rect 1019 -15132 1077 -15120
rect 1019 -15388 1031 -15132
rect 1065 -15388 1077 -15132
rect 1019 -15400 1077 -15388
rect 1197 -15132 1255 -15120
rect 1197 -15388 1209 -15132
rect 1243 -15388 1255 -15132
rect 1197 -15400 1255 -15388
rect 1375 -15132 1433 -15120
rect 1375 -15388 1387 -15132
rect 1421 -15388 1433 -15132
rect 1375 -15400 1433 -15388
rect 1553 -15132 1611 -15120
rect 1553 -15388 1565 -15132
rect 1599 -15388 1611 -15132
rect 1553 -15400 1611 -15388
rect 1731 -15132 1789 -15120
rect 1731 -15388 1743 -15132
rect 1777 -15388 1789 -15132
rect 1731 -15400 1789 -15388
rect 1909 -15132 1967 -15120
rect 1909 -15388 1921 -15132
rect 1955 -15388 1967 -15132
rect 1909 -15400 1967 -15388
rect 2087 -15132 2145 -15120
rect 2087 -15388 2099 -15132
rect 2133 -15388 2145 -15132
rect 2087 -15400 2145 -15388
rect 2265 -15132 2323 -15120
rect 2265 -15388 2277 -15132
rect 2311 -15388 2323 -15132
rect 2265 -15400 2323 -15388
rect 2443 -15132 2501 -15120
rect 2443 -15388 2455 -15132
rect 2489 -15388 2501 -15132
rect 2443 -15400 2501 -15388
rect 2621 -15132 2679 -15120
rect 2621 -15388 2633 -15132
rect 2667 -15388 2679 -15132
rect 2621 -15400 2679 -15388
rect 2799 -15132 2857 -15120
rect 2799 -15388 2811 -15132
rect 2845 -15388 2857 -15132
rect 2799 -15400 2857 -15388
rect 2977 -15132 3035 -15120
rect 2977 -15388 2989 -15132
rect 3023 -15388 3035 -15132
rect 2977 -15400 3035 -15388
rect 3155 -15132 3213 -15120
rect 3155 -15388 3167 -15132
rect 3201 -15388 3213 -15132
rect 3155 -15400 3213 -15388
rect 3333 -15132 3391 -15120
rect 3333 -15388 3345 -15132
rect 3379 -15388 3391 -15132
rect 3333 -15400 3391 -15388
rect 3511 -15132 3569 -15120
rect 3511 -15388 3523 -15132
rect 3557 -15388 3569 -15132
rect 3511 -15400 3569 -15388
rect 3689 -15132 3747 -15120
rect 3689 -15388 3701 -15132
rect 3735 -15388 3747 -15132
rect 3689 -15400 3747 -15388
rect 3867 -15132 3925 -15120
rect 3867 -15388 3879 -15132
rect 3913 -15388 3925 -15132
rect 3867 -15400 3925 -15388
rect 4045 -15132 4103 -15120
rect 4045 -15388 4057 -15132
rect 4091 -15388 4103 -15132
rect 4045 -15400 4103 -15388
rect 5565 -15132 5623 -15120
rect 5565 -15388 5577 -15132
rect 5611 -15388 5623 -15132
rect 5565 -15400 5623 -15388
rect 5743 -15132 5801 -15120
rect 5743 -15388 5755 -15132
rect 5789 -15388 5801 -15132
rect 5743 -15400 5801 -15388
rect 5921 -15132 5979 -15120
rect 5921 -15388 5933 -15132
rect 5967 -15388 5979 -15132
rect 5921 -15400 5979 -15388
rect 6099 -15132 6157 -15120
rect 6099 -15388 6111 -15132
rect 6145 -15388 6157 -15132
rect 6099 -15400 6157 -15388
rect 6277 -15132 6335 -15120
rect 6277 -15388 6289 -15132
rect 6323 -15388 6335 -15132
rect 6277 -15400 6335 -15388
rect 6455 -15132 6513 -15120
rect 6455 -15388 6467 -15132
rect 6501 -15388 6513 -15132
rect 6455 -15400 6513 -15388
rect 6633 -15132 6691 -15120
rect 6633 -15388 6645 -15132
rect 6679 -15388 6691 -15132
rect 6633 -15400 6691 -15388
rect 6811 -15132 6869 -15120
rect 6811 -15388 6823 -15132
rect 6857 -15388 6869 -15132
rect 6811 -15400 6869 -15388
rect 6989 -15132 7047 -15120
rect 6989 -15388 7001 -15132
rect 7035 -15388 7047 -15132
rect 6989 -15400 7047 -15388
rect 7167 -15132 7225 -15120
rect 7167 -15388 7179 -15132
rect 7213 -15388 7225 -15132
rect 7167 -15400 7225 -15388
rect 7345 -15132 7403 -15120
rect 7345 -15388 7357 -15132
rect 7391 -15388 7403 -15132
rect 7345 -15400 7403 -15388
rect 7523 -15132 7581 -15120
rect 7523 -15388 7535 -15132
rect 7569 -15388 7581 -15132
rect 7523 -15400 7581 -15388
rect 7701 -15132 7759 -15120
rect 7701 -15388 7713 -15132
rect 7747 -15388 7759 -15132
rect 7701 -15400 7759 -15388
rect 7879 -15132 7937 -15120
rect 7879 -15388 7891 -15132
rect 7925 -15388 7937 -15132
rect 7879 -15400 7937 -15388
rect 8057 -15132 8115 -15120
rect 8057 -15388 8069 -15132
rect 8103 -15388 8115 -15132
rect 8057 -15400 8115 -15388
rect 8235 -15132 8293 -15120
rect 8235 -15388 8247 -15132
rect 8281 -15388 8293 -15132
rect 8235 -15400 8293 -15388
rect 8413 -15132 8471 -15120
rect 8413 -15388 8425 -15132
rect 8459 -15388 8471 -15132
rect 8413 -15400 8471 -15388
rect 8591 -15132 8649 -15120
rect 8591 -15388 8603 -15132
rect 8637 -15388 8649 -15132
rect 8591 -15400 8649 -15388
rect 8769 -15132 8827 -15120
rect 8769 -15388 8781 -15132
rect 8815 -15388 8827 -15132
rect 8769 -15400 8827 -15388
rect 8947 -15132 9005 -15120
rect 8947 -15388 8959 -15132
rect 8993 -15388 9005 -15132
rect 8947 -15400 9005 -15388
rect 9125 -15132 9183 -15120
rect 9125 -15388 9137 -15132
rect 9171 -15388 9183 -15132
rect 9125 -15400 9183 -15388
rect 9303 -15132 9361 -15120
rect 9303 -15388 9315 -15132
rect 9349 -15388 9361 -15132
rect 9303 -15400 9361 -15388
rect 9481 -15132 9539 -15120
rect 9481 -15388 9493 -15132
rect 9527 -15388 9539 -15132
rect 9481 -15400 9539 -15388
rect 9659 -15132 9717 -15120
rect 9659 -15388 9671 -15132
rect 9705 -15388 9717 -15132
rect 9659 -15400 9717 -15388
rect 9837 -15132 9895 -15120
rect 9837 -15388 9849 -15132
rect 9883 -15388 9895 -15132
rect 9837 -15400 9895 -15388
rect 10015 -15132 10073 -15120
rect 10015 -15388 10027 -15132
rect 10061 -15388 10073 -15132
rect 10015 -15400 10073 -15388
rect 10193 -15132 10251 -15120
rect 10193 -15388 10205 -15132
rect 10239 -15388 10251 -15132
rect 10193 -15400 10251 -15388
rect 10371 -15132 10429 -15120
rect 10371 -15388 10383 -15132
rect 10417 -15388 10429 -15132
rect 10371 -15400 10429 -15388
rect 10549 -15132 10607 -15120
rect 10549 -15388 10561 -15132
rect 10595 -15388 10607 -15132
rect 10549 -15400 10607 -15388
rect 10727 -15132 10785 -15120
rect 10727 -15388 10739 -15132
rect 10773 -15388 10785 -15132
rect 10727 -15400 10785 -15388
rect 10905 -15132 10963 -15120
rect 10905 -15388 10917 -15132
rect 10951 -15388 10963 -15132
rect 10905 -15400 10963 -15388
rect 11083 -15132 11141 -15120
rect 11083 -15388 11095 -15132
rect 11129 -15388 11141 -15132
rect 11083 -15400 11141 -15388
rect 11261 -15132 11319 -15120
rect 11261 -15388 11273 -15132
rect 11307 -15388 11319 -15132
rect 11261 -15400 11319 -15388
rect 11439 -15132 11497 -15120
rect 11439 -15388 11451 -15132
rect 11485 -15388 11497 -15132
rect 11439 -15400 11497 -15388
rect 11617 -15132 11675 -15120
rect 11617 -15388 11629 -15132
rect 11663 -15388 11675 -15132
rect 11617 -15400 11675 -15388
rect 11795 -15132 11853 -15120
rect 11795 -15388 11807 -15132
rect 11841 -15388 11853 -15132
rect 11795 -15400 11853 -15388
rect 11973 -15132 12031 -15120
rect 11973 -15388 11985 -15132
rect 12019 -15388 12031 -15132
rect 11973 -15400 12031 -15388
rect 12151 -15132 12209 -15120
rect 12151 -15388 12163 -15132
rect 12197 -15388 12209 -15132
rect 12151 -15400 12209 -15388
rect 12329 -15132 12387 -15120
rect 12329 -15388 12341 -15132
rect 12375 -15388 12387 -15132
rect 12329 -15400 12387 -15388
rect 12507 -15132 12565 -15120
rect 12507 -15388 12519 -15132
rect 12553 -15388 12565 -15132
rect 12507 -15400 12565 -15388
rect 12685 -15132 12743 -15120
rect 12685 -15388 12697 -15132
rect 12731 -15388 12743 -15132
rect 12685 -15400 12743 -15388
rect -6040 -15794 -5982 -15782
rect -6040 -16050 -6028 -15794
rect -5994 -16050 -5982 -15794
rect -6040 -16062 -5982 -16050
rect -5862 -15794 -5804 -15782
rect -5862 -16050 -5850 -15794
rect -5816 -16050 -5804 -15794
rect -5862 -16062 -5804 -16050
rect -5684 -15794 -5626 -15782
rect -5684 -16050 -5672 -15794
rect -5638 -16050 -5626 -15794
rect -5684 -16062 -5626 -16050
rect -5506 -15794 -5448 -15782
rect -5506 -16050 -5494 -15794
rect -5460 -16050 -5448 -15794
rect -5506 -16062 -5448 -16050
rect -5328 -15794 -5270 -15782
rect -5328 -16050 -5316 -15794
rect -5282 -16050 -5270 -15794
rect -5328 -16062 -5270 -16050
rect -5150 -15794 -5092 -15782
rect -5150 -16050 -5138 -15794
rect -5104 -16050 -5092 -15794
rect -5150 -16062 -5092 -16050
rect -4972 -15794 -4914 -15782
rect -4972 -16050 -4960 -15794
rect -4926 -16050 -4914 -15794
rect -4972 -16062 -4914 -16050
rect -4794 -15794 -4736 -15782
rect -4794 -16050 -4782 -15794
rect -4748 -16050 -4736 -15794
rect -4794 -16062 -4736 -16050
rect -4616 -15794 -4558 -15782
rect -4616 -16050 -4604 -15794
rect -4570 -16050 -4558 -15794
rect -4616 -16062 -4558 -16050
rect -4438 -15794 -4380 -15782
rect -4438 -16050 -4426 -15794
rect -4392 -16050 -4380 -15794
rect -4438 -16062 -4380 -16050
rect -4260 -15794 -4202 -15782
rect -4260 -16050 -4248 -15794
rect -4214 -16050 -4202 -15794
rect -4260 -16062 -4202 -16050
rect -4082 -15794 -4024 -15782
rect -4082 -16050 -4070 -15794
rect -4036 -16050 -4024 -15794
rect -4082 -16062 -4024 -16050
rect -2185 -16132 -2127 -16120
rect -2185 -16388 -2173 -16132
rect -2139 -16388 -2127 -16132
rect -2185 -16400 -2127 -16388
rect -2007 -16132 -1949 -16120
rect -2007 -16388 -1995 -16132
rect -1961 -16388 -1949 -16132
rect -2007 -16400 -1949 -16388
rect -1829 -16132 -1771 -16120
rect -1829 -16388 -1817 -16132
rect -1783 -16388 -1771 -16132
rect -1829 -16400 -1771 -16388
rect -1651 -16132 -1593 -16120
rect -1651 -16388 -1639 -16132
rect -1605 -16388 -1593 -16132
rect -1651 -16400 -1593 -16388
rect -1473 -16132 -1415 -16120
rect -1473 -16388 -1461 -16132
rect -1427 -16388 -1415 -16132
rect -1473 -16400 -1415 -16388
rect -1295 -16132 -1237 -16120
rect -1295 -16388 -1283 -16132
rect -1249 -16388 -1237 -16132
rect -1295 -16400 -1237 -16388
rect -1117 -16132 -1059 -16120
rect -1117 -16388 -1105 -16132
rect -1071 -16388 -1059 -16132
rect -1117 -16400 -1059 -16388
rect -939 -16132 -881 -16120
rect -939 -16388 -927 -16132
rect -893 -16388 -881 -16132
rect -939 -16400 -881 -16388
rect -761 -16132 -703 -16120
rect -761 -16388 -749 -16132
rect -715 -16388 -703 -16132
rect -761 -16400 -703 -16388
rect -583 -16132 -525 -16120
rect -583 -16388 -571 -16132
rect -537 -16388 -525 -16132
rect -583 -16400 -525 -16388
rect -405 -16132 -347 -16120
rect -405 -16388 -393 -16132
rect -359 -16388 -347 -16132
rect -405 -16400 -347 -16388
rect -227 -16132 -169 -16120
rect -227 -16388 -215 -16132
rect -181 -16388 -169 -16132
rect -227 -16400 -169 -16388
rect -49 -16132 9 -16120
rect -49 -16388 -37 -16132
rect -3 -16388 9 -16132
rect -49 -16400 9 -16388
rect 129 -16132 187 -16120
rect 129 -16388 141 -16132
rect 175 -16388 187 -16132
rect 129 -16400 187 -16388
rect 307 -16132 365 -16120
rect 307 -16388 319 -16132
rect 353 -16388 365 -16132
rect 307 -16400 365 -16388
rect 485 -16132 543 -16120
rect 485 -16388 497 -16132
rect 531 -16388 543 -16132
rect 485 -16400 543 -16388
rect 663 -16132 721 -16120
rect 663 -16388 675 -16132
rect 709 -16388 721 -16132
rect 663 -16400 721 -16388
rect 841 -16132 899 -16120
rect 841 -16388 853 -16132
rect 887 -16388 899 -16132
rect 841 -16400 899 -16388
rect 1019 -16132 1077 -16120
rect 1019 -16388 1031 -16132
rect 1065 -16388 1077 -16132
rect 1019 -16400 1077 -16388
rect 1197 -16132 1255 -16120
rect 1197 -16388 1209 -16132
rect 1243 -16388 1255 -16132
rect 1197 -16400 1255 -16388
rect 1375 -16132 1433 -16120
rect 1375 -16388 1387 -16132
rect 1421 -16388 1433 -16132
rect 1375 -16400 1433 -16388
rect 1553 -16132 1611 -16120
rect 1553 -16388 1565 -16132
rect 1599 -16388 1611 -16132
rect 1553 -16400 1611 -16388
rect 1731 -16132 1789 -16120
rect 1731 -16388 1743 -16132
rect 1777 -16388 1789 -16132
rect 1731 -16400 1789 -16388
rect 1909 -16132 1967 -16120
rect 1909 -16388 1921 -16132
rect 1955 -16388 1967 -16132
rect 1909 -16400 1967 -16388
rect 2087 -16132 2145 -16120
rect 2087 -16388 2099 -16132
rect 2133 -16388 2145 -16132
rect 2087 -16400 2145 -16388
rect 2265 -16132 2323 -16120
rect 2265 -16388 2277 -16132
rect 2311 -16388 2323 -16132
rect 2265 -16400 2323 -16388
rect 2443 -16132 2501 -16120
rect 2443 -16388 2455 -16132
rect 2489 -16388 2501 -16132
rect 2443 -16400 2501 -16388
rect 2621 -16132 2679 -16120
rect 2621 -16388 2633 -16132
rect 2667 -16388 2679 -16132
rect 2621 -16400 2679 -16388
rect 2799 -16132 2857 -16120
rect 2799 -16388 2811 -16132
rect 2845 -16388 2857 -16132
rect 2799 -16400 2857 -16388
rect 2977 -16132 3035 -16120
rect 2977 -16388 2989 -16132
rect 3023 -16388 3035 -16132
rect 2977 -16400 3035 -16388
rect 3155 -16132 3213 -16120
rect 3155 -16388 3167 -16132
rect 3201 -16388 3213 -16132
rect 3155 -16400 3213 -16388
rect 3333 -16132 3391 -16120
rect 3333 -16388 3345 -16132
rect 3379 -16388 3391 -16132
rect 3333 -16400 3391 -16388
rect 3511 -16132 3569 -16120
rect 3511 -16388 3523 -16132
rect 3557 -16388 3569 -16132
rect 3511 -16400 3569 -16388
rect 3689 -16132 3747 -16120
rect 3689 -16388 3701 -16132
rect 3735 -16388 3747 -16132
rect 3689 -16400 3747 -16388
rect 3867 -16132 3925 -16120
rect 3867 -16388 3879 -16132
rect 3913 -16388 3925 -16132
rect 3867 -16400 3925 -16388
rect 4045 -16132 4103 -16120
rect 4045 -16388 4057 -16132
rect 4091 -16388 4103 -16132
rect 4045 -16400 4103 -16388
rect 5565 -16132 5623 -16120
rect 5565 -16388 5577 -16132
rect 5611 -16388 5623 -16132
rect 5565 -16400 5623 -16388
rect 5743 -16132 5801 -16120
rect 5743 -16388 5755 -16132
rect 5789 -16388 5801 -16132
rect 5743 -16400 5801 -16388
rect 5921 -16132 5979 -16120
rect 5921 -16388 5933 -16132
rect 5967 -16388 5979 -16132
rect 5921 -16400 5979 -16388
rect 6099 -16132 6157 -16120
rect 6099 -16388 6111 -16132
rect 6145 -16388 6157 -16132
rect 6099 -16400 6157 -16388
rect 6277 -16132 6335 -16120
rect 6277 -16388 6289 -16132
rect 6323 -16388 6335 -16132
rect 6277 -16400 6335 -16388
rect 6455 -16132 6513 -16120
rect 6455 -16388 6467 -16132
rect 6501 -16388 6513 -16132
rect 6455 -16400 6513 -16388
rect 6633 -16132 6691 -16120
rect 6633 -16388 6645 -16132
rect 6679 -16388 6691 -16132
rect 6633 -16400 6691 -16388
rect 6811 -16132 6869 -16120
rect 6811 -16388 6823 -16132
rect 6857 -16388 6869 -16132
rect 6811 -16400 6869 -16388
rect 6989 -16132 7047 -16120
rect 6989 -16388 7001 -16132
rect 7035 -16388 7047 -16132
rect 6989 -16400 7047 -16388
rect 7167 -16132 7225 -16120
rect 7167 -16388 7179 -16132
rect 7213 -16388 7225 -16132
rect 7167 -16400 7225 -16388
rect 7345 -16132 7403 -16120
rect 7345 -16388 7357 -16132
rect 7391 -16388 7403 -16132
rect 7345 -16400 7403 -16388
rect 7523 -16132 7581 -16120
rect 7523 -16388 7535 -16132
rect 7569 -16388 7581 -16132
rect 7523 -16400 7581 -16388
rect 7701 -16132 7759 -16120
rect 7701 -16388 7713 -16132
rect 7747 -16388 7759 -16132
rect 7701 -16400 7759 -16388
rect 7879 -16132 7937 -16120
rect 7879 -16388 7891 -16132
rect 7925 -16388 7937 -16132
rect 7879 -16400 7937 -16388
rect 8057 -16132 8115 -16120
rect 8057 -16388 8069 -16132
rect 8103 -16388 8115 -16132
rect 8057 -16400 8115 -16388
rect 8235 -16132 8293 -16120
rect 8235 -16388 8247 -16132
rect 8281 -16388 8293 -16132
rect 8235 -16400 8293 -16388
rect 8413 -16132 8471 -16120
rect 8413 -16388 8425 -16132
rect 8459 -16388 8471 -16132
rect 8413 -16400 8471 -16388
rect 8591 -16132 8649 -16120
rect 8591 -16388 8603 -16132
rect 8637 -16388 8649 -16132
rect 8591 -16400 8649 -16388
rect 8769 -16132 8827 -16120
rect 8769 -16388 8781 -16132
rect 8815 -16388 8827 -16132
rect 8769 -16400 8827 -16388
rect 8947 -16132 9005 -16120
rect 8947 -16388 8959 -16132
rect 8993 -16388 9005 -16132
rect 8947 -16400 9005 -16388
rect 9125 -16132 9183 -16120
rect 9125 -16388 9137 -16132
rect 9171 -16388 9183 -16132
rect 9125 -16400 9183 -16388
rect 9303 -16132 9361 -16120
rect 9303 -16388 9315 -16132
rect 9349 -16388 9361 -16132
rect 9303 -16400 9361 -16388
rect 9481 -16132 9539 -16120
rect 9481 -16388 9493 -16132
rect 9527 -16388 9539 -16132
rect 9481 -16400 9539 -16388
rect 9659 -16132 9717 -16120
rect 9659 -16388 9671 -16132
rect 9705 -16388 9717 -16132
rect 9659 -16400 9717 -16388
rect 9837 -16132 9895 -16120
rect 9837 -16388 9849 -16132
rect 9883 -16388 9895 -16132
rect 9837 -16400 9895 -16388
rect 10015 -16132 10073 -16120
rect 10015 -16388 10027 -16132
rect 10061 -16388 10073 -16132
rect 10015 -16400 10073 -16388
rect 10193 -16132 10251 -16120
rect 10193 -16388 10205 -16132
rect 10239 -16388 10251 -16132
rect 10193 -16400 10251 -16388
rect 10371 -16132 10429 -16120
rect 10371 -16388 10383 -16132
rect 10417 -16388 10429 -16132
rect 10371 -16400 10429 -16388
rect 10549 -16132 10607 -16120
rect 10549 -16388 10561 -16132
rect 10595 -16388 10607 -16132
rect 10549 -16400 10607 -16388
rect 10727 -16132 10785 -16120
rect 10727 -16388 10739 -16132
rect 10773 -16388 10785 -16132
rect 10727 -16400 10785 -16388
rect 10905 -16132 10963 -16120
rect 10905 -16388 10917 -16132
rect 10951 -16388 10963 -16132
rect 10905 -16400 10963 -16388
rect 11083 -16132 11141 -16120
rect 11083 -16388 11095 -16132
rect 11129 -16388 11141 -16132
rect 11083 -16400 11141 -16388
rect 11261 -16132 11319 -16120
rect 11261 -16388 11273 -16132
rect 11307 -16388 11319 -16132
rect 11261 -16400 11319 -16388
rect 11439 -16132 11497 -16120
rect 11439 -16388 11451 -16132
rect 11485 -16388 11497 -16132
rect 11439 -16400 11497 -16388
rect 11617 -16132 11675 -16120
rect 11617 -16388 11629 -16132
rect 11663 -16388 11675 -16132
rect 11617 -16400 11675 -16388
rect 11795 -16132 11853 -16120
rect 11795 -16388 11807 -16132
rect 11841 -16388 11853 -16132
rect 11795 -16400 11853 -16388
rect 11973 -16132 12031 -16120
rect 11973 -16388 11985 -16132
rect 12019 -16388 12031 -16132
rect 11973 -16400 12031 -16388
rect 12151 -16132 12209 -16120
rect 12151 -16388 12163 -16132
rect 12197 -16388 12209 -16132
rect 12151 -16400 12209 -16388
rect 12329 -16132 12387 -16120
rect 12329 -16388 12341 -16132
rect 12375 -16388 12387 -16132
rect 12329 -16400 12387 -16388
rect 12507 -16132 12565 -16120
rect 12507 -16388 12519 -16132
rect 12553 -16388 12565 -16132
rect 12507 -16400 12565 -16388
rect 12685 -16132 12743 -16120
rect 12685 -16388 12697 -16132
rect 12731 -16388 12743 -16132
rect 12685 -16400 12743 -16388
rect -6040 -16494 -5982 -16482
rect -6040 -16750 -6028 -16494
rect -5994 -16750 -5982 -16494
rect -6040 -16762 -5982 -16750
rect -5862 -16494 -5804 -16482
rect -5862 -16750 -5850 -16494
rect -5816 -16750 -5804 -16494
rect -5862 -16762 -5804 -16750
rect -5684 -16494 -5626 -16482
rect -5684 -16750 -5672 -16494
rect -5638 -16750 -5626 -16494
rect -5684 -16762 -5626 -16750
rect -5506 -16494 -5448 -16482
rect -5506 -16750 -5494 -16494
rect -5460 -16750 -5448 -16494
rect -5506 -16762 -5448 -16750
rect -5328 -16494 -5270 -16482
rect -5328 -16750 -5316 -16494
rect -5282 -16750 -5270 -16494
rect -5328 -16762 -5270 -16750
rect -5150 -16494 -5092 -16482
rect -5150 -16750 -5138 -16494
rect -5104 -16750 -5092 -16494
rect -5150 -16762 -5092 -16750
rect -4972 -16494 -4914 -16482
rect -4972 -16750 -4960 -16494
rect -4926 -16750 -4914 -16494
rect -4972 -16762 -4914 -16750
rect -4794 -16494 -4736 -16482
rect -4794 -16750 -4782 -16494
rect -4748 -16750 -4736 -16494
rect -4794 -16762 -4736 -16750
rect -4616 -16494 -4558 -16482
rect -4616 -16750 -4604 -16494
rect -4570 -16750 -4558 -16494
rect -4616 -16762 -4558 -16750
rect -4438 -16494 -4380 -16482
rect -4438 -16750 -4426 -16494
rect -4392 -16750 -4380 -16494
rect -4438 -16762 -4380 -16750
rect -4260 -16494 -4202 -16482
rect -4260 -16750 -4248 -16494
rect -4214 -16750 -4202 -16494
rect -4260 -16762 -4202 -16750
rect -4082 -16494 -4024 -16482
rect -4082 -16750 -4070 -16494
rect -4036 -16750 -4024 -16494
rect -4082 -16762 -4024 -16750
<< pdiff >>
rect -6314 -2132 -6256 -2120
rect -6314 -2388 -6302 -2132
rect -6268 -2388 -6256 -2132
rect -6314 -2400 -6256 -2388
rect -6136 -2132 -6078 -2120
rect -6136 -2388 -6124 -2132
rect -6090 -2388 -6078 -2132
rect -6136 -2400 -6078 -2388
rect -5958 -2132 -5900 -2120
rect -5958 -2388 -5946 -2132
rect -5912 -2388 -5900 -2132
rect -5958 -2400 -5900 -2388
rect -5780 -2132 -5722 -2120
rect -5780 -2388 -5768 -2132
rect -5734 -2388 -5722 -2132
rect -5780 -2400 -5722 -2388
rect -5602 -2132 -5544 -2120
rect -5602 -2388 -5590 -2132
rect -5556 -2388 -5544 -2132
rect -5602 -2400 -5544 -2388
rect -5424 -2132 -5366 -2120
rect -5424 -2388 -5412 -2132
rect -5378 -2388 -5366 -2132
rect -5424 -2400 -5366 -2388
rect -5246 -2132 -5188 -2120
rect -5246 -2388 -5234 -2132
rect -5200 -2388 -5188 -2132
rect -5246 -2400 -5188 -2388
rect -5068 -2132 -5010 -2120
rect -5068 -2388 -5056 -2132
rect -5022 -2388 -5010 -2132
rect -5068 -2400 -5010 -2388
rect -4890 -2132 -4832 -2120
rect -4890 -2388 -4878 -2132
rect -4844 -2388 -4832 -2132
rect -4890 -2400 -4832 -2388
rect -4712 -2132 -4654 -2120
rect -4712 -2388 -4700 -2132
rect -4666 -2388 -4654 -2132
rect -4712 -2400 -4654 -2388
rect -4534 -2132 -4476 -2120
rect -4534 -2388 -4522 -2132
rect -4488 -2388 -4476 -2132
rect -4534 -2400 -4476 -2388
rect -4356 -2132 -4298 -2120
rect -4356 -2388 -4344 -2132
rect -4310 -2388 -4298 -2132
rect -4356 -2400 -4298 -2388
rect -4178 -2132 -4120 -2120
rect -4178 -2388 -4166 -2132
rect -4132 -2388 -4120 -2132
rect -4178 -2400 -4120 -2388
rect -4000 -2132 -3942 -2120
rect -4000 -2388 -3988 -2132
rect -3954 -2388 -3942 -2132
rect -4000 -2400 -3942 -2388
rect -3822 -2132 -3764 -2120
rect -3822 -2388 -3810 -2132
rect -3776 -2388 -3764 -2132
rect -3822 -2400 -3764 -2388
rect -3644 -2132 -3586 -2120
rect -3644 -2388 -3632 -2132
rect -3598 -2388 -3586 -2132
rect -3644 -2400 -3586 -2388
rect -3466 -2132 -3408 -2120
rect -3466 -2388 -3454 -2132
rect -3420 -2388 -3408 -2132
rect -3466 -2400 -3408 -2388
rect -1466 -2884 -1408 -2872
rect -6314 -3002 -6256 -2990
rect -6314 -3258 -6302 -3002
rect -6268 -3258 -6256 -3002
rect -6314 -3270 -6256 -3258
rect -6136 -3002 -6078 -2990
rect -6136 -3258 -6124 -3002
rect -6090 -3258 -6078 -3002
rect -6136 -3270 -6078 -3258
rect -5958 -3002 -5900 -2990
rect -5958 -3258 -5946 -3002
rect -5912 -3258 -5900 -3002
rect -5958 -3270 -5900 -3258
rect -5780 -3002 -5722 -2990
rect -5780 -3258 -5768 -3002
rect -5734 -3258 -5722 -3002
rect -5780 -3270 -5722 -3258
rect -5602 -3002 -5544 -2990
rect -5602 -3258 -5590 -3002
rect -5556 -3258 -5544 -3002
rect -5602 -3270 -5544 -3258
rect -5424 -3002 -5366 -2990
rect -5424 -3258 -5412 -3002
rect -5378 -3258 -5366 -3002
rect -5424 -3270 -5366 -3258
rect -5246 -3002 -5188 -2990
rect -5246 -3258 -5234 -3002
rect -5200 -3258 -5188 -3002
rect -5246 -3270 -5188 -3258
rect -5068 -3002 -5010 -2990
rect -5068 -3258 -5056 -3002
rect -5022 -3258 -5010 -3002
rect -5068 -3270 -5010 -3258
rect -4890 -3002 -4832 -2990
rect -4890 -3258 -4878 -3002
rect -4844 -3258 -4832 -3002
rect -4890 -3270 -4832 -3258
rect -4712 -3002 -4654 -2990
rect -4712 -3258 -4700 -3002
rect -4666 -3258 -4654 -3002
rect -4712 -3270 -4654 -3258
rect -4534 -3002 -4476 -2990
rect -4534 -3258 -4522 -3002
rect -4488 -3258 -4476 -3002
rect -4534 -3270 -4476 -3258
rect -4356 -3002 -4298 -2990
rect -4356 -3258 -4344 -3002
rect -4310 -3258 -4298 -3002
rect -4356 -3270 -4298 -3258
rect -4178 -3002 -4120 -2990
rect -4178 -3258 -4166 -3002
rect -4132 -3258 -4120 -3002
rect -4178 -3270 -4120 -3258
rect -4000 -3002 -3942 -2990
rect -4000 -3258 -3988 -3002
rect -3954 -3258 -3942 -3002
rect -4000 -3270 -3942 -3258
rect -3822 -3002 -3764 -2990
rect -3822 -3258 -3810 -3002
rect -3776 -3258 -3764 -3002
rect -3822 -3270 -3764 -3258
rect -3644 -3002 -3586 -2990
rect -3644 -3258 -3632 -3002
rect -3598 -3258 -3586 -3002
rect -3644 -3270 -3586 -3258
rect -3466 -3002 -3408 -2990
rect -3466 -3258 -3454 -3002
rect -3420 -3258 -3408 -3002
rect -1466 -3140 -1454 -2884
rect -1420 -3140 -1408 -2884
rect -1466 -3152 -1408 -3140
rect -1288 -2884 -1230 -2872
rect -1288 -3140 -1276 -2884
rect -1242 -3140 -1230 -2884
rect -1288 -3152 -1230 -3140
rect -1110 -2884 -1052 -2872
rect -1110 -3140 -1098 -2884
rect -1064 -3140 -1052 -2884
rect -1110 -3152 -1052 -3140
rect -932 -2884 -874 -2872
rect -932 -3140 -920 -2884
rect -886 -3140 -874 -2884
rect -932 -3152 -874 -3140
rect -754 -2884 -696 -2872
rect -754 -3140 -742 -2884
rect -708 -3140 -696 -2884
rect -754 -3152 -696 -3140
rect -576 -2884 -518 -2872
rect -576 -3140 -564 -2884
rect -530 -3140 -518 -2884
rect -576 -3152 -518 -3140
rect -398 -2884 -340 -2872
rect -398 -3140 -386 -2884
rect -352 -3140 -340 -2884
rect -398 -3152 -340 -3140
rect -220 -2884 -162 -2872
rect -220 -3140 -208 -2884
rect -174 -3140 -162 -2884
rect -220 -3152 -162 -3140
rect -42 -2884 16 -2872
rect -42 -3140 -30 -2884
rect 4 -3140 16 -2884
rect -42 -3152 16 -3140
rect 136 -2884 194 -2872
rect 136 -3140 148 -2884
rect 182 -3140 194 -2884
rect 136 -3152 194 -3140
rect 314 -2884 372 -2872
rect 314 -3140 326 -2884
rect 360 -3140 372 -2884
rect 314 -3152 372 -3140
rect 492 -2884 550 -2872
rect 492 -3140 504 -2884
rect 538 -3140 550 -2884
rect 492 -3152 550 -3140
rect 670 -2884 728 -2872
rect 670 -3140 682 -2884
rect 716 -3140 728 -2884
rect 670 -3152 728 -3140
rect 848 -2884 906 -2872
rect 848 -3140 860 -2884
rect 894 -3140 906 -2884
rect 848 -3152 906 -3140
rect 1026 -2884 1084 -2872
rect 1026 -3140 1038 -2884
rect 1072 -3140 1084 -2884
rect 1026 -3152 1084 -3140
rect 1204 -2884 1262 -2872
rect 1204 -3140 1216 -2884
rect 1250 -3140 1262 -2884
rect 1204 -3152 1262 -3140
rect 1382 -2884 1440 -2872
rect 1382 -3140 1394 -2884
rect 1428 -3140 1440 -2884
rect 1382 -3152 1440 -3140
rect 1560 -2884 1618 -2872
rect 1560 -3140 1572 -2884
rect 1606 -3140 1618 -2884
rect 1560 -3152 1618 -3140
rect 1738 -2884 1796 -2872
rect 1738 -3140 1750 -2884
rect 1784 -3140 1796 -2884
rect 1738 -3152 1796 -3140
rect 1916 -2884 1974 -2872
rect 1916 -3140 1928 -2884
rect 1962 -3140 1974 -2884
rect 1916 -3152 1974 -3140
rect 2094 -2884 2152 -2872
rect 2094 -3140 2106 -2884
rect 2140 -3140 2152 -2884
rect 2094 -3152 2152 -3140
rect 2272 -2884 2330 -2872
rect 2272 -3140 2284 -2884
rect 2318 -3140 2330 -2884
rect 2272 -3152 2330 -3140
rect 2450 -2884 2508 -2872
rect 2450 -3140 2462 -2884
rect 2496 -3140 2508 -2884
rect 2450 -3152 2508 -3140
rect 2628 -2884 2686 -2872
rect 2628 -3140 2640 -2884
rect 2674 -3140 2686 -2884
rect 2628 -3152 2686 -3140
rect -3466 -3270 -3408 -3258
rect -1466 -3784 -1408 -3772
rect -6314 -3872 -6256 -3860
rect -6314 -4128 -6302 -3872
rect -6268 -4128 -6256 -3872
rect -6314 -4140 -6256 -4128
rect -6136 -3872 -6078 -3860
rect -6136 -4128 -6124 -3872
rect -6090 -4128 -6078 -3872
rect -6136 -4140 -6078 -4128
rect -5958 -3872 -5900 -3860
rect -5958 -4128 -5946 -3872
rect -5912 -4128 -5900 -3872
rect -5958 -4140 -5900 -4128
rect -5780 -3872 -5722 -3860
rect -5780 -4128 -5768 -3872
rect -5734 -4128 -5722 -3872
rect -5780 -4140 -5722 -4128
rect -5602 -3872 -5544 -3860
rect -5602 -4128 -5590 -3872
rect -5556 -4128 -5544 -3872
rect -5602 -4140 -5544 -4128
rect -5424 -3872 -5366 -3860
rect -5424 -4128 -5412 -3872
rect -5378 -4128 -5366 -3872
rect -5424 -4140 -5366 -4128
rect -5246 -3872 -5188 -3860
rect -5246 -4128 -5234 -3872
rect -5200 -4128 -5188 -3872
rect -5246 -4140 -5188 -4128
rect -5068 -3872 -5010 -3860
rect -5068 -4128 -5056 -3872
rect -5022 -4128 -5010 -3872
rect -5068 -4140 -5010 -4128
rect -4890 -3872 -4832 -3860
rect -4890 -4128 -4878 -3872
rect -4844 -4128 -4832 -3872
rect -4890 -4140 -4832 -4128
rect -4712 -3872 -4654 -3860
rect -4712 -4128 -4700 -3872
rect -4666 -4128 -4654 -3872
rect -4712 -4140 -4654 -4128
rect -4534 -3872 -4476 -3860
rect -4534 -4128 -4522 -3872
rect -4488 -4128 -4476 -3872
rect -4534 -4140 -4476 -4128
rect -4356 -3872 -4298 -3860
rect -4356 -4128 -4344 -3872
rect -4310 -4128 -4298 -3872
rect -4356 -4140 -4298 -4128
rect -4178 -3872 -4120 -3860
rect -4178 -4128 -4166 -3872
rect -4132 -4128 -4120 -3872
rect -4178 -4140 -4120 -4128
rect -4000 -3872 -3942 -3860
rect -4000 -4128 -3988 -3872
rect -3954 -4128 -3942 -3872
rect -4000 -4140 -3942 -4128
rect -3822 -3872 -3764 -3860
rect -3822 -4128 -3810 -3872
rect -3776 -4128 -3764 -3872
rect -3822 -4140 -3764 -4128
rect -3644 -3872 -3586 -3860
rect -3644 -4128 -3632 -3872
rect -3598 -4128 -3586 -3872
rect -3644 -4140 -3586 -4128
rect -3466 -3872 -3408 -3860
rect -3466 -4128 -3454 -3872
rect -3420 -4128 -3408 -3872
rect -1466 -4040 -1454 -3784
rect -1420 -4040 -1408 -3784
rect -1466 -4052 -1408 -4040
rect -1288 -3784 -1230 -3772
rect -1288 -4040 -1276 -3784
rect -1242 -4040 -1230 -3784
rect -1288 -4052 -1230 -4040
rect -1110 -3784 -1052 -3772
rect -1110 -4040 -1098 -3784
rect -1064 -4040 -1052 -3784
rect -1110 -4052 -1052 -4040
rect -932 -3784 -874 -3772
rect -932 -4040 -920 -3784
rect -886 -4040 -874 -3784
rect -932 -4052 -874 -4040
rect -754 -3784 -696 -3772
rect -754 -4040 -742 -3784
rect -708 -4040 -696 -3784
rect -754 -4052 -696 -4040
rect -576 -3784 -518 -3772
rect -576 -4040 -564 -3784
rect -530 -4040 -518 -3784
rect -576 -4052 -518 -4040
rect -398 -3784 -340 -3772
rect -398 -4040 -386 -3784
rect -352 -4040 -340 -3784
rect -398 -4052 -340 -4040
rect -220 -3784 -162 -3772
rect -220 -4040 -208 -3784
rect -174 -4040 -162 -3784
rect -220 -4052 -162 -4040
rect -42 -3784 16 -3772
rect -42 -4040 -30 -3784
rect 4 -4040 16 -3784
rect -42 -4052 16 -4040
rect 136 -3784 194 -3772
rect 136 -4040 148 -3784
rect 182 -4040 194 -3784
rect 136 -4052 194 -4040
rect 314 -3784 372 -3772
rect 314 -4040 326 -3784
rect 360 -4040 372 -3784
rect 314 -4052 372 -4040
rect 492 -3784 550 -3772
rect 492 -4040 504 -3784
rect 538 -4040 550 -3784
rect 492 -4052 550 -4040
rect 670 -3784 728 -3772
rect 670 -4040 682 -3784
rect 716 -4040 728 -3784
rect 670 -4052 728 -4040
rect 848 -3784 906 -3772
rect 848 -4040 860 -3784
rect 894 -4040 906 -3784
rect 848 -4052 906 -4040
rect 1026 -3784 1084 -3772
rect 1026 -4040 1038 -3784
rect 1072 -4040 1084 -3784
rect 1026 -4052 1084 -4040
rect 1204 -3784 1262 -3772
rect 1204 -4040 1216 -3784
rect 1250 -4040 1262 -3784
rect 1204 -4052 1262 -4040
rect 1382 -3784 1440 -3772
rect 1382 -4040 1394 -3784
rect 1428 -4040 1440 -3784
rect 1382 -4052 1440 -4040
rect 1560 -3784 1618 -3772
rect 1560 -4040 1572 -3784
rect 1606 -4040 1618 -3784
rect 1560 -4052 1618 -4040
rect 1738 -3784 1796 -3772
rect 1738 -4040 1750 -3784
rect 1784 -4040 1796 -3784
rect 1738 -4052 1796 -4040
rect 1916 -3784 1974 -3772
rect 1916 -4040 1928 -3784
rect 1962 -4040 1974 -3784
rect 1916 -4052 1974 -4040
rect 2094 -3784 2152 -3772
rect 2094 -4040 2106 -3784
rect 2140 -4040 2152 -3784
rect 2094 -4052 2152 -4040
rect 2272 -3784 2330 -3772
rect 2272 -4040 2284 -3784
rect 2318 -4040 2330 -3784
rect 2272 -4052 2330 -4040
rect 2450 -3784 2508 -3772
rect 2450 -4040 2462 -3784
rect 2496 -4040 2508 -3784
rect 2450 -4052 2508 -4040
rect 2628 -3784 2686 -3772
rect 2628 -4040 2640 -3784
rect 2674 -4040 2686 -3784
rect 2628 -4052 2686 -4040
rect -3466 -4140 -3408 -4128
rect -1466 -4684 -1408 -4672
rect -6314 -4742 -6256 -4730
rect -6314 -4998 -6302 -4742
rect -6268 -4998 -6256 -4742
rect -6314 -5010 -6256 -4998
rect -6136 -4742 -6078 -4730
rect -6136 -4998 -6124 -4742
rect -6090 -4998 -6078 -4742
rect -6136 -5010 -6078 -4998
rect -5958 -4742 -5900 -4730
rect -5958 -4998 -5946 -4742
rect -5912 -4998 -5900 -4742
rect -5958 -5010 -5900 -4998
rect -5780 -4742 -5722 -4730
rect -5780 -4998 -5768 -4742
rect -5734 -4998 -5722 -4742
rect -5780 -5010 -5722 -4998
rect -5602 -4742 -5544 -4730
rect -5602 -4998 -5590 -4742
rect -5556 -4998 -5544 -4742
rect -5602 -5010 -5544 -4998
rect -5424 -4742 -5366 -4730
rect -5424 -4998 -5412 -4742
rect -5378 -4998 -5366 -4742
rect -5424 -5010 -5366 -4998
rect -5246 -4742 -5188 -4730
rect -5246 -4998 -5234 -4742
rect -5200 -4998 -5188 -4742
rect -5246 -5010 -5188 -4998
rect -5068 -4742 -5010 -4730
rect -5068 -4998 -5056 -4742
rect -5022 -4998 -5010 -4742
rect -5068 -5010 -5010 -4998
rect -4890 -4742 -4832 -4730
rect -4890 -4998 -4878 -4742
rect -4844 -4998 -4832 -4742
rect -4890 -5010 -4832 -4998
rect -4712 -4742 -4654 -4730
rect -4712 -4998 -4700 -4742
rect -4666 -4998 -4654 -4742
rect -4712 -5010 -4654 -4998
rect -4534 -4742 -4476 -4730
rect -4534 -4998 -4522 -4742
rect -4488 -4998 -4476 -4742
rect -4534 -5010 -4476 -4998
rect -4356 -4742 -4298 -4730
rect -4356 -4998 -4344 -4742
rect -4310 -4998 -4298 -4742
rect -4356 -5010 -4298 -4998
rect -4178 -4742 -4120 -4730
rect -4178 -4998 -4166 -4742
rect -4132 -4998 -4120 -4742
rect -4178 -5010 -4120 -4998
rect -4000 -4742 -3942 -4730
rect -4000 -4998 -3988 -4742
rect -3954 -4998 -3942 -4742
rect -4000 -5010 -3942 -4998
rect -3822 -4742 -3764 -4730
rect -3822 -4998 -3810 -4742
rect -3776 -4998 -3764 -4742
rect -3822 -5010 -3764 -4998
rect -3644 -4742 -3586 -4730
rect -3644 -4998 -3632 -4742
rect -3598 -4998 -3586 -4742
rect -3644 -5010 -3586 -4998
rect -3466 -4742 -3408 -4730
rect -3466 -4998 -3454 -4742
rect -3420 -4998 -3408 -4742
rect -1466 -4940 -1454 -4684
rect -1420 -4940 -1408 -4684
rect -1466 -4952 -1408 -4940
rect -1288 -4684 -1230 -4672
rect -1288 -4940 -1276 -4684
rect -1242 -4940 -1230 -4684
rect -1288 -4952 -1230 -4940
rect -1110 -4684 -1052 -4672
rect -1110 -4940 -1098 -4684
rect -1064 -4940 -1052 -4684
rect -1110 -4952 -1052 -4940
rect -932 -4684 -874 -4672
rect -932 -4940 -920 -4684
rect -886 -4940 -874 -4684
rect -932 -4952 -874 -4940
rect -754 -4684 -696 -4672
rect -754 -4940 -742 -4684
rect -708 -4940 -696 -4684
rect -754 -4952 -696 -4940
rect -576 -4684 -518 -4672
rect -576 -4940 -564 -4684
rect -530 -4940 -518 -4684
rect -576 -4952 -518 -4940
rect -398 -4684 -340 -4672
rect -398 -4940 -386 -4684
rect -352 -4940 -340 -4684
rect -398 -4952 -340 -4940
rect -220 -4684 -162 -4672
rect -220 -4940 -208 -4684
rect -174 -4940 -162 -4684
rect -220 -4952 -162 -4940
rect -42 -4684 16 -4672
rect -42 -4940 -30 -4684
rect 4 -4940 16 -4684
rect -42 -4952 16 -4940
rect 136 -4684 194 -4672
rect 136 -4940 148 -4684
rect 182 -4940 194 -4684
rect 136 -4952 194 -4940
rect 314 -4684 372 -4672
rect 314 -4940 326 -4684
rect 360 -4940 372 -4684
rect 314 -4952 372 -4940
rect 492 -4684 550 -4672
rect 492 -4940 504 -4684
rect 538 -4940 550 -4684
rect 492 -4952 550 -4940
rect 670 -4684 728 -4672
rect 670 -4940 682 -4684
rect 716 -4940 728 -4684
rect 670 -4952 728 -4940
rect 848 -4684 906 -4672
rect 848 -4940 860 -4684
rect 894 -4940 906 -4684
rect 848 -4952 906 -4940
rect 1026 -4684 1084 -4672
rect 1026 -4940 1038 -4684
rect 1072 -4940 1084 -4684
rect 1026 -4952 1084 -4940
rect 1204 -4684 1262 -4672
rect 1204 -4940 1216 -4684
rect 1250 -4940 1262 -4684
rect 1204 -4952 1262 -4940
rect 1382 -4684 1440 -4672
rect 1382 -4940 1394 -4684
rect 1428 -4940 1440 -4684
rect 1382 -4952 1440 -4940
rect 1560 -4684 1618 -4672
rect 1560 -4940 1572 -4684
rect 1606 -4940 1618 -4684
rect 1560 -4952 1618 -4940
rect 1738 -4684 1796 -4672
rect 1738 -4940 1750 -4684
rect 1784 -4940 1796 -4684
rect 1738 -4952 1796 -4940
rect 1916 -4684 1974 -4672
rect 1916 -4940 1928 -4684
rect 1962 -4940 1974 -4684
rect 1916 -4952 1974 -4940
rect 2094 -4684 2152 -4672
rect 2094 -4940 2106 -4684
rect 2140 -4940 2152 -4684
rect 2094 -4952 2152 -4940
rect 2272 -4684 2330 -4672
rect 2272 -4940 2284 -4684
rect 2318 -4940 2330 -4684
rect 2272 -4952 2330 -4940
rect 2450 -4684 2508 -4672
rect 2450 -4940 2462 -4684
rect 2496 -4940 2508 -4684
rect 2450 -4952 2508 -4940
rect 2628 -4684 2686 -4672
rect 2628 -4940 2640 -4684
rect 2674 -4940 2686 -4684
rect 2628 -4952 2686 -4940
rect -3466 -5010 -3408 -4998
rect -1466 -5584 -1408 -5572
rect -6314 -5612 -6256 -5600
rect -6314 -5868 -6302 -5612
rect -6268 -5868 -6256 -5612
rect -6314 -5880 -6256 -5868
rect -6136 -5612 -6078 -5600
rect -6136 -5868 -6124 -5612
rect -6090 -5868 -6078 -5612
rect -6136 -5880 -6078 -5868
rect -5958 -5612 -5900 -5600
rect -5958 -5868 -5946 -5612
rect -5912 -5868 -5900 -5612
rect -5958 -5880 -5900 -5868
rect -5780 -5612 -5722 -5600
rect -5780 -5868 -5768 -5612
rect -5734 -5868 -5722 -5612
rect -5780 -5880 -5722 -5868
rect -5602 -5612 -5544 -5600
rect -5602 -5868 -5590 -5612
rect -5556 -5868 -5544 -5612
rect -5602 -5880 -5544 -5868
rect -5424 -5612 -5366 -5600
rect -5424 -5868 -5412 -5612
rect -5378 -5868 -5366 -5612
rect -5424 -5880 -5366 -5868
rect -5246 -5612 -5188 -5600
rect -5246 -5868 -5234 -5612
rect -5200 -5868 -5188 -5612
rect -5246 -5880 -5188 -5868
rect -5068 -5612 -5010 -5600
rect -5068 -5868 -5056 -5612
rect -5022 -5868 -5010 -5612
rect -5068 -5880 -5010 -5868
rect -4890 -5612 -4832 -5600
rect -4890 -5868 -4878 -5612
rect -4844 -5868 -4832 -5612
rect -4890 -5880 -4832 -5868
rect -4712 -5612 -4654 -5600
rect -4712 -5868 -4700 -5612
rect -4666 -5868 -4654 -5612
rect -4712 -5880 -4654 -5868
rect -4534 -5612 -4476 -5600
rect -4534 -5868 -4522 -5612
rect -4488 -5868 -4476 -5612
rect -4534 -5880 -4476 -5868
rect -4356 -5612 -4298 -5600
rect -4356 -5868 -4344 -5612
rect -4310 -5868 -4298 -5612
rect -4356 -5880 -4298 -5868
rect -4178 -5612 -4120 -5600
rect -4178 -5868 -4166 -5612
rect -4132 -5868 -4120 -5612
rect -4178 -5880 -4120 -5868
rect -4000 -5612 -3942 -5600
rect -4000 -5868 -3988 -5612
rect -3954 -5868 -3942 -5612
rect -4000 -5880 -3942 -5868
rect -3822 -5612 -3764 -5600
rect -3822 -5868 -3810 -5612
rect -3776 -5868 -3764 -5612
rect -3822 -5880 -3764 -5868
rect -3644 -5612 -3586 -5600
rect -3644 -5868 -3632 -5612
rect -3598 -5868 -3586 -5612
rect -3644 -5880 -3586 -5868
rect -3466 -5612 -3408 -5600
rect -3466 -5868 -3454 -5612
rect -3420 -5868 -3408 -5612
rect -1466 -5840 -1454 -5584
rect -1420 -5840 -1408 -5584
rect -1466 -5852 -1408 -5840
rect -1288 -5584 -1230 -5572
rect -1288 -5840 -1276 -5584
rect -1242 -5840 -1230 -5584
rect -1288 -5852 -1230 -5840
rect -1110 -5584 -1052 -5572
rect -1110 -5840 -1098 -5584
rect -1064 -5840 -1052 -5584
rect -1110 -5852 -1052 -5840
rect -932 -5584 -874 -5572
rect -932 -5840 -920 -5584
rect -886 -5840 -874 -5584
rect -932 -5852 -874 -5840
rect -754 -5584 -696 -5572
rect -754 -5840 -742 -5584
rect -708 -5840 -696 -5584
rect -754 -5852 -696 -5840
rect -576 -5584 -518 -5572
rect -576 -5840 -564 -5584
rect -530 -5840 -518 -5584
rect -576 -5852 -518 -5840
rect -398 -5584 -340 -5572
rect -398 -5840 -386 -5584
rect -352 -5840 -340 -5584
rect -398 -5852 -340 -5840
rect -220 -5584 -162 -5572
rect -220 -5840 -208 -5584
rect -174 -5840 -162 -5584
rect -220 -5852 -162 -5840
rect -42 -5584 16 -5572
rect -42 -5840 -30 -5584
rect 4 -5840 16 -5584
rect -42 -5852 16 -5840
rect 136 -5584 194 -5572
rect 136 -5840 148 -5584
rect 182 -5840 194 -5584
rect 136 -5852 194 -5840
rect 314 -5584 372 -5572
rect 314 -5840 326 -5584
rect 360 -5840 372 -5584
rect 314 -5852 372 -5840
rect 492 -5584 550 -5572
rect 492 -5840 504 -5584
rect 538 -5840 550 -5584
rect 492 -5852 550 -5840
rect 670 -5584 728 -5572
rect 670 -5840 682 -5584
rect 716 -5840 728 -5584
rect 670 -5852 728 -5840
rect 848 -5584 906 -5572
rect 848 -5840 860 -5584
rect 894 -5840 906 -5584
rect 848 -5852 906 -5840
rect 1026 -5584 1084 -5572
rect 1026 -5840 1038 -5584
rect 1072 -5840 1084 -5584
rect 1026 -5852 1084 -5840
rect 1204 -5584 1262 -5572
rect 1204 -5840 1216 -5584
rect 1250 -5840 1262 -5584
rect 1204 -5852 1262 -5840
rect 1382 -5584 1440 -5572
rect 1382 -5840 1394 -5584
rect 1428 -5840 1440 -5584
rect 1382 -5852 1440 -5840
rect 1560 -5584 1618 -5572
rect 1560 -5840 1572 -5584
rect 1606 -5840 1618 -5584
rect 1560 -5852 1618 -5840
rect 1738 -5584 1796 -5572
rect 1738 -5840 1750 -5584
rect 1784 -5840 1796 -5584
rect 1738 -5852 1796 -5840
rect 1916 -5584 1974 -5572
rect 1916 -5840 1928 -5584
rect 1962 -5840 1974 -5584
rect 1916 -5852 1974 -5840
rect 2094 -5584 2152 -5572
rect 2094 -5840 2106 -5584
rect 2140 -5840 2152 -5584
rect 2094 -5852 2152 -5840
rect 2272 -5584 2330 -5572
rect 2272 -5840 2284 -5584
rect 2318 -5840 2330 -5584
rect 2272 -5852 2330 -5840
rect 2450 -5584 2508 -5572
rect 2450 -5840 2462 -5584
rect 2496 -5840 2508 -5584
rect 2450 -5852 2508 -5840
rect 2628 -5584 2686 -5572
rect 2628 -5840 2640 -5584
rect 2674 -5840 2686 -5584
rect 2628 -5852 2686 -5840
rect -3466 -5880 -3408 -5868
<< ndiffc >>
rect -5628 -8130 -5594 -7874
rect -5450 -8130 -5416 -7874
rect -5272 -8130 -5238 -7874
rect -5094 -8130 -5060 -7874
rect -4916 -8130 -4882 -7874
rect -4738 -8130 -4704 -7874
rect -4560 -8130 -4526 -7874
rect -4382 -8130 -4348 -7874
rect -4204 -8130 -4170 -7874
rect -4026 -8130 -3992 -7874
rect -2173 -8388 -2139 -8132
rect -1995 -8388 -1961 -8132
rect -1817 -8388 -1783 -8132
rect -1639 -8388 -1605 -8132
rect -1461 -8388 -1427 -8132
rect -1283 -8388 -1249 -8132
rect -1105 -8388 -1071 -8132
rect -927 -8388 -893 -8132
rect -749 -8388 -715 -8132
rect -571 -8388 -537 -8132
rect -393 -8388 -359 -8132
rect -215 -8388 -181 -8132
rect -37 -8388 -3 -8132
rect 141 -8388 175 -8132
rect 319 -8388 353 -8132
rect 497 -8388 531 -8132
rect 675 -8388 709 -8132
rect 853 -8388 887 -8132
rect 1031 -8388 1065 -8132
rect 1209 -8388 1243 -8132
rect 1387 -8388 1421 -8132
rect 1565 -8388 1599 -8132
rect 1743 -8388 1777 -8132
rect 1921 -8388 1955 -8132
rect 2099 -8388 2133 -8132
rect 2277 -8388 2311 -8132
rect 2455 -8388 2489 -8132
rect 2633 -8388 2667 -8132
rect 2811 -8388 2845 -8132
rect 2989 -8388 3023 -8132
rect 3167 -8388 3201 -8132
rect 3345 -8388 3379 -8132
rect 3523 -8388 3557 -8132
rect 3701 -8388 3735 -8132
rect 3879 -8388 3913 -8132
rect 4057 -8388 4091 -8132
rect -5628 -8680 -5594 -8424
rect -5450 -8680 -5416 -8424
rect -5272 -8680 -5238 -8424
rect -5094 -8680 -5060 -8424
rect -4916 -8680 -4882 -8424
rect -4738 -8680 -4704 -8424
rect -4560 -8680 -4526 -8424
rect -4382 -8680 -4348 -8424
rect -4204 -8680 -4170 -8424
rect -4026 -8680 -3992 -8424
rect -5628 -9230 -5594 -8974
rect -5450 -9230 -5416 -8974
rect -5272 -9230 -5238 -8974
rect -5094 -9230 -5060 -8974
rect -4916 -9230 -4882 -8974
rect -4738 -9230 -4704 -8974
rect -4560 -9230 -4526 -8974
rect -4382 -9230 -4348 -8974
rect -4204 -9230 -4170 -8974
rect -4026 -9230 -3992 -8974
rect -2173 -9388 -2139 -9132
rect -1995 -9388 -1961 -9132
rect -1817 -9388 -1783 -9132
rect -1639 -9388 -1605 -9132
rect -1461 -9388 -1427 -9132
rect -1283 -9388 -1249 -9132
rect -1105 -9388 -1071 -9132
rect -927 -9388 -893 -9132
rect -749 -9388 -715 -9132
rect -571 -9388 -537 -9132
rect -393 -9388 -359 -9132
rect -215 -9388 -181 -9132
rect -37 -9388 -3 -9132
rect 141 -9388 175 -9132
rect 319 -9388 353 -9132
rect 497 -9388 531 -9132
rect 675 -9388 709 -9132
rect 853 -9388 887 -9132
rect 1031 -9388 1065 -9132
rect 1209 -9388 1243 -9132
rect 1387 -9388 1421 -9132
rect 1565 -9388 1599 -9132
rect 1743 -9388 1777 -9132
rect 1921 -9388 1955 -9132
rect 2099 -9388 2133 -9132
rect 2277 -9388 2311 -9132
rect 2455 -9388 2489 -9132
rect 2633 -9388 2667 -9132
rect 2811 -9388 2845 -9132
rect 2989 -9388 3023 -9132
rect 3167 -9388 3201 -9132
rect 3345 -9388 3379 -9132
rect 3523 -9388 3557 -9132
rect 3701 -9388 3735 -9132
rect 3879 -9388 3913 -9132
rect 4057 -9388 4091 -9132
rect 6512 -9150 6546 -8894
rect 6690 -9150 6724 -8894
rect 6868 -9150 6902 -8894
rect 7046 -9150 7080 -8894
rect 7224 -9150 7258 -8894
rect 7402 -9150 7436 -8894
rect 7580 -9150 7614 -8894
rect 7758 -9150 7792 -8894
rect 7936 -9150 7970 -8894
rect 8114 -9150 8148 -8894
rect 8292 -9150 8326 -8894
rect 8470 -9150 8504 -8894
rect 8648 -9150 8682 -8894
rect 8826 -9150 8860 -8894
rect 9004 -9150 9038 -8894
rect 9182 -9150 9216 -8894
rect 9360 -9150 9394 -8894
rect 10772 -9180 10806 -8924
rect 10950 -9180 10984 -8924
rect 11064 -9180 11098 -8924
rect 11242 -9180 11276 -8924
rect 11356 -9180 11390 -8924
rect 11534 -9180 11568 -8924
rect 11648 -9180 11682 -8924
rect 11826 -9180 11860 -8924
rect 11940 -9180 11974 -8924
rect 12118 -9180 12152 -8924
rect 12232 -9180 12266 -8924
rect 12410 -9180 12444 -8924
rect 12524 -9180 12558 -8924
rect 12702 -9180 12736 -8924
rect -5628 -9780 -5594 -9524
rect -5450 -9780 -5416 -9524
rect -5272 -9780 -5238 -9524
rect -5094 -9780 -5060 -9524
rect -4916 -9780 -4882 -9524
rect -4738 -9780 -4704 -9524
rect -4560 -9780 -4526 -9524
rect -4382 -9780 -4348 -9524
rect -4204 -9780 -4170 -9524
rect -4026 -9780 -3992 -9524
rect -5628 -10330 -5594 -10074
rect -5450 -10330 -5416 -10074
rect -5272 -10330 -5238 -10074
rect -5094 -10330 -5060 -10074
rect -4916 -10330 -4882 -10074
rect -4738 -10330 -4704 -10074
rect -4560 -10330 -4526 -10074
rect -4382 -10330 -4348 -10074
rect -4204 -10330 -4170 -10074
rect -4026 -10330 -3992 -10074
rect 6512 -10050 6546 -9794
rect 6690 -10050 6724 -9794
rect 6868 -10050 6902 -9794
rect 7046 -10050 7080 -9794
rect 7224 -10050 7258 -9794
rect 7402 -10050 7436 -9794
rect 7580 -10050 7614 -9794
rect 7758 -10050 7792 -9794
rect 7936 -10050 7970 -9794
rect 8114 -10050 8148 -9794
rect 8292 -10050 8326 -9794
rect 8470 -10050 8504 -9794
rect 8648 -10050 8682 -9794
rect 8826 -10050 8860 -9794
rect 9004 -10050 9038 -9794
rect 9182 -10050 9216 -9794
rect 9360 -10050 9394 -9794
rect 10772 -9950 10806 -9694
rect 10950 -9950 10984 -9694
rect 11064 -9950 11098 -9694
rect 11242 -9950 11276 -9694
rect 11356 -9950 11390 -9694
rect 11534 -9950 11568 -9694
rect 11648 -9950 11682 -9694
rect 11826 -9950 11860 -9694
rect 11940 -9950 11974 -9694
rect 12118 -9950 12152 -9694
rect 12232 -9950 12266 -9694
rect 12410 -9950 12444 -9694
rect 12524 -9950 12558 -9694
rect 12702 -9950 12736 -9694
rect -2173 -10388 -2139 -10132
rect -1995 -10388 -1961 -10132
rect -1817 -10388 -1783 -10132
rect -1639 -10388 -1605 -10132
rect -1461 -10388 -1427 -10132
rect -1283 -10388 -1249 -10132
rect -1105 -10388 -1071 -10132
rect -927 -10388 -893 -10132
rect -749 -10388 -715 -10132
rect -571 -10388 -537 -10132
rect -393 -10388 -359 -10132
rect -215 -10388 -181 -10132
rect -37 -10388 -3 -10132
rect 141 -10388 175 -10132
rect 319 -10388 353 -10132
rect 497 -10388 531 -10132
rect 675 -10388 709 -10132
rect 853 -10388 887 -10132
rect 1031 -10388 1065 -10132
rect 1209 -10388 1243 -10132
rect 1387 -10388 1421 -10132
rect 1565 -10388 1599 -10132
rect 1743 -10388 1777 -10132
rect 1921 -10388 1955 -10132
rect 2099 -10388 2133 -10132
rect 2277 -10388 2311 -10132
rect 2455 -10388 2489 -10132
rect 2633 -10388 2667 -10132
rect 2811 -10388 2845 -10132
rect 2989 -10388 3023 -10132
rect 3167 -10388 3201 -10132
rect 3345 -10388 3379 -10132
rect 3523 -10388 3557 -10132
rect 3701 -10388 3735 -10132
rect 3879 -10388 3913 -10132
rect 4057 -10388 4091 -10132
rect -5628 -10880 -5594 -10624
rect -5450 -10880 -5416 -10624
rect -5272 -10880 -5238 -10624
rect -5094 -10880 -5060 -10624
rect -4916 -10880 -4882 -10624
rect -4738 -10880 -4704 -10624
rect -4560 -10880 -4526 -10624
rect -4382 -10880 -4348 -10624
rect -4204 -10880 -4170 -10624
rect -4026 -10880 -3992 -10624
rect 6512 -10950 6546 -10694
rect 6690 -10950 6724 -10694
rect 6868 -10950 6902 -10694
rect 7046 -10950 7080 -10694
rect 7224 -10950 7258 -10694
rect 7402 -10950 7436 -10694
rect 7580 -10950 7614 -10694
rect 7758 -10950 7792 -10694
rect 7936 -10950 7970 -10694
rect 8114 -10950 8148 -10694
rect 8292 -10950 8326 -10694
rect 8470 -10950 8504 -10694
rect 8648 -10950 8682 -10694
rect 8826 -10950 8860 -10694
rect 9004 -10950 9038 -10694
rect 9182 -10950 9216 -10694
rect 9360 -10950 9394 -10694
rect 10772 -10720 10806 -10464
rect 10950 -10720 10984 -10464
rect 11064 -10720 11098 -10464
rect 11242 -10720 11276 -10464
rect 11356 -10720 11390 -10464
rect 11534 -10720 11568 -10464
rect 11648 -10720 11682 -10464
rect 11826 -10720 11860 -10464
rect 11940 -10720 11974 -10464
rect 12118 -10720 12152 -10464
rect 12232 -10720 12266 -10464
rect 12410 -10720 12444 -10464
rect 12524 -10720 12558 -10464
rect 12702 -10720 12736 -10464
rect -5628 -11430 -5594 -11174
rect -5450 -11430 -5416 -11174
rect -5272 -11430 -5238 -11174
rect -5094 -11430 -5060 -11174
rect -4916 -11430 -4882 -11174
rect -4738 -11430 -4704 -11174
rect -4560 -11430 -4526 -11174
rect -4382 -11430 -4348 -11174
rect -4204 -11430 -4170 -11174
rect -4026 -11430 -3992 -11174
rect -2173 -11388 -2139 -11132
rect -1995 -11388 -1961 -11132
rect -1817 -11388 -1783 -11132
rect -1639 -11388 -1605 -11132
rect -1461 -11388 -1427 -11132
rect -1283 -11388 -1249 -11132
rect -1105 -11388 -1071 -11132
rect -927 -11388 -893 -11132
rect -749 -11388 -715 -11132
rect -571 -11388 -537 -11132
rect -393 -11388 -359 -11132
rect -215 -11388 -181 -11132
rect -37 -11388 -3 -11132
rect 141 -11388 175 -11132
rect 319 -11388 353 -11132
rect 497 -11388 531 -11132
rect 675 -11388 709 -11132
rect 853 -11388 887 -11132
rect 1031 -11388 1065 -11132
rect 1209 -11388 1243 -11132
rect 1387 -11388 1421 -11132
rect 1565 -11388 1599 -11132
rect 1743 -11388 1777 -11132
rect 1921 -11388 1955 -11132
rect 2099 -11388 2133 -11132
rect 2277 -11388 2311 -11132
rect 2455 -11388 2489 -11132
rect 2633 -11388 2667 -11132
rect 2811 -11388 2845 -11132
rect 2989 -11388 3023 -11132
rect 3167 -11388 3201 -11132
rect 3345 -11388 3379 -11132
rect 3523 -11388 3557 -11132
rect 3701 -11388 3735 -11132
rect 3879 -11388 3913 -11132
rect 4057 -11388 4091 -11132
rect 10772 -11490 10806 -11234
rect 10950 -11490 10984 -11234
rect 11064 -11490 11098 -11234
rect 11242 -11490 11276 -11234
rect 11356 -11490 11390 -11234
rect 11534 -11490 11568 -11234
rect 11648 -11490 11682 -11234
rect 11826 -11490 11860 -11234
rect 11940 -11490 11974 -11234
rect 12118 -11490 12152 -11234
rect 12232 -11490 12266 -11234
rect 12410 -11490 12444 -11234
rect 12524 -11490 12558 -11234
rect 12702 -11490 12736 -11234
rect -5628 -11980 -5594 -11724
rect -5450 -11980 -5416 -11724
rect -5272 -11980 -5238 -11724
rect -5094 -11980 -5060 -11724
rect -4916 -11980 -4882 -11724
rect -4738 -11980 -4704 -11724
rect -4560 -11980 -4526 -11724
rect -4382 -11980 -4348 -11724
rect -4204 -11980 -4170 -11724
rect -4026 -11980 -3992 -11724
rect 6512 -11850 6546 -11594
rect 6690 -11850 6724 -11594
rect 6868 -11850 6902 -11594
rect 7046 -11850 7080 -11594
rect 7224 -11850 7258 -11594
rect 7402 -11850 7436 -11594
rect 7580 -11850 7614 -11594
rect 7758 -11850 7792 -11594
rect 7936 -11850 7970 -11594
rect 8114 -11850 8148 -11594
rect 8292 -11850 8326 -11594
rect 8470 -11850 8504 -11594
rect 8648 -11850 8682 -11594
rect 8826 -11850 8860 -11594
rect 9004 -11850 9038 -11594
rect 9182 -11850 9216 -11594
rect 9360 -11850 9394 -11594
rect -2173 -12388 -2139 -12132
rect -1995 -12388 -1961 -12132
rect -1817 -12388 -1783 -12132
rect -1639 -12388 -1605 -12132
rect -1461 -12388 -1427 -12132
rect -1283 -12388 -1249 -12132
rect -1105 -12388 -1071 -12132
rect -927 -12388 -893 -12132
rect -749 -12388 -715 -12132
rect -571 -12388 -537 -12132
rect -393 -12388 -359 -12132
rect -215 -12388 -181 -12132
rect -37 -12388 -3 -12132
rect 141 -12388 175 -12132
rect 319 -12388 353 -12132
rect 497 -12388 531 -12132
rect 675 -12388 709 -12132
rect 853 -12388 887 -12132
rect 1031 -12388 1065 -12132
rect 1209 -12388 1243 -12132
rect 1387 -12388 1421 -12132
rect 1565 -12388 1599 -12132
rect 1743 -12388 1777 -12132
rect 1921 -12388 1955 -12132
rect 2099 -12388 2133 -12132
rect 2277 -12388 2311 -12132
rect 2455 -12388 2489 -12132
rect 2633 -12388 2667 -12132
rect 2811 -12388 2845 -12132
rect 2989 -12388 3023 -12132
rect 3167 -12388 3201 -12132
rect 3345 -12388 3379 -12132
rect 3523 -12388 3557 -12132
rect 3701 -12388 3735 -12132
rect 3879 -12388 3913 -12132
rect 4057 -12388 4091 -12132
rect -5916 -12928 -5882 -12712
rect -5818 -12928 -5784 -12712
rect -5666 -12928 -5632 -12712
rect -5568 -12928 -5534 -12712
rect -5416 -12928 -5382 -12712
rect -5318 -12928 -5284 -12712
rect -5166 -12928 -5132 -12712
rect -5068 -12928 -5034 -12712
rect -4916 -12928 -4882 -12712
rect -4818 -12928 -4784 -12712
rect -4666 -12928 -4632 -12712
rect -4568 -12928 -4534 -12712
rect -4416 -12928 -4382 -12712
rect -4318 -12928 -4284 -12712
rect -4166 -12928 -4132 -12712
rect -4068 -12928 -4034 -12712
rect -5916 -13608 -5882 -13392
rect -5818 -13608 -5784 -13392
rect -5666 -13608 -5632 -13392
rect -5568 -13608 -5534 -13392
rect -5416 -13608 -5382 -13392
rect -5318 -13608 -5284 -13392
rect -5166 -13608 -5132 -13392
rect -5068 -13608 -5034 -13392
rect -4916 -13608 -4882 -13392
rect -4818 -13608 -4784 -13392
rect -4666 -13608 -4632 -13392
rect -4568 -13608 -4534 -13392
rect -4416 -13608 -4382 -13392
rect -4318 -13608 -4284 -13392
rect -4166 -13608 -4132 -13392
rect -4068 -13608 -4034 -13392
rect -2173 -13388 -2139 -13132
rect -1995 -13388 -1961 -13132
rect -1817 -13388 -1783 -13132
rect -1639 -13388 -1605 -13132
rect -1461 -13388 -1427 -13132
rect -1283 -13388 -1249 -13132
rect -1105 -13388 -1071 -13132
rect -927 -13388 -893 -13132
rect -749 -13388 -715 -13132
rect -571 -13388 -537 -13132
rect -393 -13388 -359 -13132
rect -215 -13388 -181 -13132
rect -37 -13388 -3 -13132
rect 141 -13388 175 -13132
rect 319 -13388 353 -13132
rect 497 -13388 531 -13132
rect 675 -13388 709 -13132
rect 853 -13388 887 -13132
rect 1031 -13388 1065 -13132
rect 1209 -13388 1243 -13132
rect 1387 -13388 1421 -13132
rect 1565 -13388 1599 -13132
rect 1743 -13388 1777 -13132
rect 1921 -13388 1955 -13132
rect 2099 -13388 2133 -13132
rect 2277 -13388 2311 -13132
rect 2455 -13388 2489 -13132
rect 2633 -13388 2667 -13132
rect 2811 -13388 2845 -13132
rect 2989 -13388 3023 -13132
rect 3167 -13388 3201 -13132
rect 3345 -13388 3379 -13132
rect 3523 -13388 3557 -13132
rect 3701 -13388 3735 -13132
rect 3879 -13388 3913 -13132
rect 4057 -13388 4091 -13132
rect -6028 -14650 -5994 -14394
rect -5850 -14650 -5816 -14394
rect -5672 -14650 -5638 -14394
rect -5494 -14650 -5460 -14394
rect -5316 -14650 -5282 -14394
rect -5138 -14650 -5104 -14394
rect -4960 -14650 -4926 -14394
rect -4782 -14650 -4748 -14394
rect -4604 -14650 -4570 -14394
rect -4426 -14650 -4392 -14394
rect -4248 -14650 -4214 -14394
rect -4070 -14650 -4036 -14394
rect -2173 -14388 -2139 -14132
rect -1995 -14388 -1961 -14132
rect -1817 -14388 -1783 -14132
rect -1639 -14388 -1605 -14132
rect -1461 -14388 -1427 -14132
rect -1283 -14388 -1249 -14132
rect -1105 -14388 -1071 -14132
rect -927 -14388 -893 -14132
rect -749 -14388 -715 -14132
rect -571 -14388 -537 -14132
rect -393 -14388 -359 -14132
rect -215 -14388 -181 -14132
rect -37 -14388 -3 -14132
rect 141 -14388 175 -14132
rect 319 -14388 353 -14132
rect 497 -14388 531 -14132
rect 675 -14388 709 -14132
rect 853 -14388 887 -14132
rect 1031 -14388 1065 -14132
rect 1209 -14388 1243 -14132
rect 1387 -14388 1421 -14132
rect 1565 -14388 1599 -14132
rect 1743 -14388 1777 -14132
rect 1921 -14388 1955 -14132
rect 2099 -14388 2133 -14132
rect 2277 -14388 2311 -14132
rect 2455 -14388 2489 -14132
rect 2633 -14388 2667 -14132
rect 2811 -14388 2845 -14132
rect 2989 -14388 3023 -14132
rect 3167 -14388 3201 -14132
rect 3345 -14388 3379 -14132
rect 3523 -14388 3557 -14132
rect 3701 -14388 3735 -14132
rect 3879 -14388 3913 -14132
rect 4057 -14388 4091 -14132
rect 5577 -14388 5611 -14132
rect 5755 -14388 5789 -14132
rect 5933 -14388 5967 -14132
rect 6111 -14388 6145 -14132
rect 6289 -14388 6323 -14132
rect 6467 -14388 6501 -14132
rect 6645 -14388 6679 -14132
rect 6823 -14388 6857 -14132
rect 7001 -14388 7035 -14132
rect 7179 -14388 7213 -14132
rect 7357 -14388 7391 -14132
rect 7535 -14388 7569 -14132
rect 7713 -14388 7747 -14132
rect 7891 -14388 7925 -14132
rect 8069 -14388 8103 -14132
rect 8247 -14388 8281 -14132
rect 8425 -14388 8459 -14132
rect 8603 -14388 8637 -14132
rect 8781 -14388 8815 -14132
rect 8959 -14388 8993 -14132
rect 9137 -14388 9171 -14132
rect 9315 -14388 9349 -14132
rect 9493 -14388 9527 -14132
rect 9671 -14388 9705 -14132
rect 9849 -14388 9883 -14132
rect 10027 -14388 10061 -14132
rect 10205 -14388 10239 -14132
rect 10383 -14388 10417 -14132
rect 10561 -14388 10595 -14132
rect 10739 -14388 10773 -14132
rect 10917 -14388 10951 -14132
rect 11095 -14388 11129 -14132
rect 11273 -14388 11307 -14132
rect 11451 -14388 11485 -14132
rect 11629 -14388 11663 -14132
rect 11807 -14388 11841 -14132
rect 11985 -14388 12019 -14132
rect 12163 -14388 12197 -14132
rect 12341 -14388 12375 -14132
rect 12519 -14388 12553 -14132
rect 12697 -14388 12731 -14132
rect -6028 -15350 -5994 -15094
rect -5850 -15350 -5816 -15094
rect -5672 -15350 -5638 -15094
rect -5494 -15350 -5460 -15094
rect -5316 -15350 -5282 -15094
rect -5138 -15350 -5104 -15094
rect -4960 -15350 -4926 -15094
rect -4782 -15350 -4748 -15094
rect -4604 -15350 -4570 -15094
rect -4426 -15350 -4392 -15094
rect -4248 -15350 -4214 -15094
rect -4070 -15350 -4036 -15094
rect -2173 -15388 -2139 -15132
rect -1995 -15388 -1961 -15132
rect -1817 -15388 -1783 -15132
rect -1639 -15388 -1605 -15132
rect -1461 -15388 -1427 -15132
rect -1283 -15388 -1249 -15132
rect -1105 -15388 -1071 -15132
rect -927 -15388 -893 -15132
rect -749 -15388 -715 -15132
rect -571 -15388 -537 -15132
rect -393 -15388 -359 -15132
rect -215 -15388 -181 -15132
rect -37 -15388 -3 -15132
rect 141 -15388 175 -15132
rect 319 -15388 353 -15132
rect 497 -15388 531 -15132
rect 675 -15388 709 -15132
rect 853 -15388 887 -15132
rect 1031 -15388 1065 -15132
rect 1209 -15388 1243 -15132
rect 1387 -15388 1421 -15132
rect 1565 -15388 1599 -15132
rect 1743 -15388 1777 -15132
rect 1921 -15388 1955 -15132
rect 2099 -15388 2133 -15132
rect 2277 -15388 2311 -15132
rect 2455 -15388 2489 -15132
rect 2633 -15388 2667 -15132
rect 2811 -15388 2845 -15132
rect 2989 -15388 3023 -15132
rect 3167 -15388 3201 -15132
rect 3345 -15388 3379 -15132
rect 3523 -15388 3557 -15132
rect 3701 -15388 3735 -15132
rect 3879 -15388 3913 -15132
rect 4057 -15388 4091 -15132
rect 5577 -15388 5611 -15132
rect 5755 -15388 5789 -15132
rect 5933 -15388 5967 -15132
rect 6111 -15388 6145 -15132
rect 6289 -15388 6323 -15132
rect 6467 -15388 6501 -15132
rect 6645 -15388 6679 -15132
rect 6823 -15388 6857 -15132
rect 7001 -15388 7035 -15132
rect 7179 -15388 7213 -15132
rect 7357 -15388 7391 -15132
rect 7535 -15388 7569 -15132
rect 7713 -15388 7747 -15132
rect 7891 -15388 7925 -15132
rect 8069 -15388 8103 -15132
rect 8247 -15388 8281 -15132
rect 8425 -15388 8459 -15132
rect 8603 -15388 8637 -15132
rect 8781 -15388 8815 -15132
rect 8959 -15388 8993 -15132
rect 9137 -15388 9171 -15132
rect 9315 -15388 9349 -15132
rect 9493 -15388 9527 -15132
rect 9671 -15388 9705 -15132
rect 9849 -15388 9883 -15132
rect 10027 -15388 10061 -15132
rect 10205 -15388 10239 -15132
rect 10383 -15388 10417 -15132
rect 10561 -15388 10595 -15132
rect 10739 -15388 10773 -15132
rect 10917 -15388 10951 -15132
rect 11095 -15388 11129 -15132
rect 11273 -15388 11307 -15132
rect 11451 -15388 11485 -15132
rect 11629 -15388 11663 -15132
rect 11807 -15388 11841 -15132
rect 11985 -15388 12019 -15132
rect 12163 -15388 12197 -15132
rect 12341 -15388 12375 -15132
rect 12519 -15388 12553 -15132
rect 12697 -15388 12731 -15132
rect -6028 -16050 -5994 -15794
rect -5850 -16050 -5816 -15794
rect -5672 -16050 -5638 -15794
rect -5494 -16050 -5460 -15794
rect -5316 -16050 -5282 -15794
rect -5138 -16050 -5104 -15794
rect -4960 -16050 -4926 -15794
rect -4782 -16050 -4748 -15794
rect -4604 -16050 -4570 -15794
rect -4426 -16050 -4392 -15794
rect -4248 -16050 -4214 -15794
rect -4070 -16050 -4036 -15794
rect -2173 -16388 -2139 -16132
rect -1995 -16388 -1961 -16132
rect -1817 -16388 -1783 -16132
rect -1639 -16388 -1605 -16132
rect -1461 -16388 -1427 -16132
rect -1283 -16388 -1249 -16132
rect -1105 -16388 -1071 -16132
rect -927 -16388 -893 -16132
rect -749 -16388 -715 -16132
rect -571 -16388 -537 -16132
rect -393 -16388 -359 -16132
rect -215 -16388 -181 -16132
rect -37 -16388 -3 -16132
rect 141 -16388 175 -16132
rect 319 -16388 353 -16132
rect 497 -16388 531 -16132
rect 675 -16388 709 -16132
rect 853 -16388 887 -16132
rect 1031 -16388 1065 -16132
rect 1209 -16388 1243 -16132
rect 1387 -16388 1421 -16132
rect 1565 -16388 1599 -16132
rect 1743 -16388 1777 -16132
rect 1921 -16388 1955 -16132
rect 2099 -16388 2133 -16132
rect 2277 -16388 2311 -16132
rect 2455 -16388 2489 -16132
rect 2633 -16388 2667 -16132
rect 2811 -16388 2845 -16132
rect 2989 -16388 3023 -16132
rect 3167 -16388 3201 -16132
rect 3345 -16388 3379 -16132
rect 3523 -16388 3557 -16132
rect 3701 -16388 3735 -16132
rect 3879 -16388 3913 -16132
rect 4057 -16388 4091 -16132
rect 5577 -16388 5611 -16132
rect 5755 -16388 5789 -16132
rect 5933 -16388 5967 -16132
rect 6111 -16388 6145 -16132
rect 6289 -16388 6323 -16132
rect 6467 -16388 6501 -16132
rect 6645 -16388 6679 -16132
rect 6823 -16388 6857 -16132
rect 7001 -16388 7035 -16132
rect 7179 -16388 7213 -16132
rect 7357 -16388 7391 -16132
rect 7535 -16388 7569 -16132
rect 7713 -16388 7747 -16132
rect 7891 -16388 7925 -16132
rect 8069 -16388 8103 -16132
rect 8247 -16388 8281 -16132
rect 8425 -16388 8459 -16132
rect 8603 -16388 8637 -16132
rect 8781 -16388 8815 -16132
rect 8959 -16388 8993 -16132
rect 9137 -16388 9171 -16132
rect 9315 -16388 9349 -16132
rect 9493 -16388 9527 -16132
rect 9671 -16388 9705 -16132
rect 9849 -16388 9883 -16132
rect 10027 -16388 10061 -16132
rect 10205 -16388 10239 -16132
rect 10383 -16388 10417 -16132
rect 10561 -16388 10595 -16132
rect 10739 -16388 10773 -16132
rect 10917 -16388 10951 -16132
rect 11095 -16388 11129 -16132
rect 11273 -16388 11307 -16132
rect 11451 -16388 11485 -16132
rect 11629 -16388 11663 -16132
rect 11807 -16388 11841 -16132
rect 11985 -16388 12019 -16132
rect 12163 -16388 12197 -16132
rect 12341 -16388 12375 -16132
rect 12519 -16388 12553 -16132
rect 12697 -16388 12731 -16132
rect -6028 -16750 -5994 -16494
rect -5850 -16750 -5816 -16494
rect -5672 -16750 -5638 -16494
rect -5494 -16750 -5460 -16494
rect -5316 -16750 -5282 -16494
rect -5138 -16750 -5104 -16494
rect -4960 -16750 -4926 -16494
rect -4782 -16750 -4748 -16494
rect -4604 -16750 -4570 -16494
rect -4426 -16750 -4392 -16494
rect -4248 -16750 -4214 -16494
rect -4070 -16750 -4036 -16494
<< pdiffc >>
rect -6302 -2388 -6268 -2132
rect -6124 -2388 -6090 -2132
rect -5946 -2388 -5912 -2132
rect -5768 -2388 -5734 -2132
rect -5590 -2388 -5556 -2132
rect -5412 -2388 -5378 -2132
rect -5234 -2388 -5200 -2132
rect -5056 -2388 -5022 -2132
rect -4878 -2388 -4844 -2132
rect -4700 -2388 -4666 -2132
rect -4522 -2388 -4488 -2132
rect -4344 -2388 -4310 -2132
rect -4166 -2388 -4132 -2132
rect -3988 -2388 -3954 -2132
rect -3810 -2388 -3776 -2132
rect -3632 -2388 -3598 -2132
rect -3454 -2388 -3420 -2132
rect -6302 -3258 -6268 -3002
rect -6124 -3258 -6090 -3002
rect -5946 -3258 -5912 -3002
rect -5768 -3258 -5734 -3002
rect -5590 -3258 -5556 -3002
rect -5412 -3258 -5378 -3002
rect -5234 -3258 -5200 -3002
rect -5056 -3258 -5022 -3002
rect -4878 -3258 -4844 -3002
rect -4700 -3258 -4666 -3002
rect -4522 -3258 -4488 -3002
rect -4344 -3258 -4310 -3002
rect -4166 -3258 -4132 -3002
rect -3988 -3258 -3954 -3002
rect -3810 -3258 -3776 -3002
rect -3632 -3258 -3598 -3002
rect -3454 -3258 -3420 -3002
rect -1454 -3140 -1420 -2884
rect -1276 -3140 -1242 -2884
rect -1098 -3140 -1064 -2884
rect -920 -3140 -886 -2884
rect -742 -3140 -708 -2884
rect -564 -3140 -530 -2884
rect -386 -3140 -352 -2884
rect -208 -3140 -174 -2884
rect -30 -3140 4 -2884
rect 148 -3140 182 -2884
rect 326 -3140 360 -2884
rect 504 -3140 538 -2884
rect 682 -3140 716 -2884
rect 860 -3140 894 -2884
rect 1038 -3140 1072 -2884
rect 1216 -3140 1250 -2884
rect 1394 -3140 1428 -2884
rect 1572 -3140 1606 -2884
rect 1750 -3140 1784 -2884
rect 1928 -3140 1962 -2884
rect 2106 -3140 2140 -2884
rect 2284 -3140 2318 -2884
rect 2462 -3140 2496 -2884
rect 2640 -3140 2674 -2884
rect -6302 -4128 -6268 -3872
rect -6124 -4128 -6090 -3872
rect -5946 -4128 -5912 -3872
rect -5768 -4128 -5734 -3872
rect -5590 -4128 -5556 -3872
rect -5412 -4128 -5378 -3872
rect -5234 -4128 -5200 -3872
rect -5056 -4128 -5022 -3872
rect -4878 -4128 -4844 -3872
rect -4700 -4128 -4666 -3872
rect -4522 -4128 -4488 -3872
rect -4344 -4128 -4310 -3872
rect -4166 -4128 -4132 -3872
rect -3988 -4128 -3954 -3872
rect -3810 -4128 -3776 -3872
rect -3632 -4128 -3598 -3872
rect -3454 -4128 -3420 -3872
rect -1454 -4040 -1420 -3784
rect -1276 -4040 -1242 -3784
rect -1098 -4040 -1064 -3784
rect -920 -4040 -886 -3784
rect -742 -4040 -708 -3784
rect -564 -4040 -530 -3784
rect -386 -4040 -352 -3784
rect -208 -4040 -174 -3784
rect -30 -4040 4 -3784
rect 148 -4040 182 -3784
rect 326 -4040 360 -3784
rect 504 -4040 538 -3784
rect 682 -4040 716 -3784
rect 860 -4040 894 -3784
rect 1038 -4040 1072 -3784
rect 1216 -4040 1250 -3784
rect 1394 -4040 1428 -3784
rect 1572 -4040 1606 -3784
rect 1750 -4040 1784 -3784
rect 1928 -4040 1962 -3784
rect 2106 -4040 2140 -3784
rect 2284 -4040 2318 -3784
rect 2462 -4040 2496 -3784
rect 2640 -4040 2674 -3784
rect -6302 -4998 -6268 -4742
rect -6124 -4998 -6090 -4742
rect -5946 -4998 -5912 -4742
rect -5768 -4998 -5734 -4742
rect -5590 -4998 -5556 -4742
rect -5412 -4998 -5378 -4742
rect -5234 -4998 -5200 -4742
rect -5056 -4998 -5022 -4742
rect -4878 -4998 -4844 -4742
rect -4700 -4998 -4666 -4742
rect -4522 -4998 -4488 -4742
rect -4344 -4998 -4310 -4742
rect -4166 -4998 -4132 -4742
rect -3988 -4998 -3954 -4742
rect -3810 -4998 -3776 -4742
rect -3632 -4998 -3598 -4742
rect -3454 -4998 -3420 -4742
rect -1454 -4940 -1420 -4684
rect -1276 -4940 -1242 -4684
rect -1098 -4940 -1064 -4684
rect -920 -4940 -886 -4684
rect -742 -4940 -708 -4684
rect -564 -4940 -530 -4684
rect -386 -4940 -352 -4684
rect -208 -4940 -174 -4684
rect -30 -4940 4 -4684
rect 148 -4940 182 -4684
rect 326 -4940 360 -4684
rect 504 -4940 538 -4684
rect 682 -4940 716 -4684
rect 860 -4940 894 -4684
rect 1038 -4940 1072 -4684
rect 1216 -4940 1250 -4684
rect 1394 -4940 1428 -4684
rect 1572 -4940 1606 -4684
rect 1750 -4940 1784 -4684
rect 1928 -4940 1962 -4684
rect 2106 -4940 2140 -4684
rect 2284 -4940 2318 -4684
rect 2462 -4940 2496 -4684
rect 2640 -4940 2674 -4684
rect -6302 -5868 -6268 -5612
rect -6124 -5868 -6090 -5612
rect -5946 -5868 -5912 -5612
rect -5768 -5868 -5734 -5612
rect -5590 -5868 -5556 -5612
rect -5412 -5868 -5378 -5612
rect -5234 -5868 -5200 -5612
rect -5056 -5868 -5022 -5612
rect -4878 -5868 -4844 -5612
rect -4700 -5868 -4666 -5612
rect -4522 -5868 -4488 -5612
rect -4344 -5868 -4310 -5612
rect -4166 -5868 -4132 -5612
rect -3988 -5868 -3954 -5612
rect -3810 -5868 -3776 -5612
rect -3632 -5868 -3598 -5612
rect -3454 -5868 -3420 -5612
rect -1454 -5840 -1420 -5584
rect -1276 -5840 -1242 -5584
rect -1098 -5840 -1064 -5584
rect -920 -5840 -886 -5584
rect -742 -5840 -708 -5584
rect -564 -5840 -530 -5584
rect -386 -5840 -352 -5584
rect -208 -5840 -174 -5584
rect -30 -5840 4 -5584
rect 148 -5840 182 -5584
rect 326 -5840 360 -5584
rect 504 -5840 538 -5584
rect 682 -5840 716 -5584
rect 860 -5840 894 -5584
rect 1038 -5840 1072 -5584
rect 1216 -5840 1250 -5584
rect 1394 -5840 1428 -5584
rect 1572 -5840 1606 -5584
rect 1750 -5840 1784 -5584
rect 1928 -5840 1962 -5584
rect 2106 -5840 2140 -5584
rect 2284 -5840 2318 -5584
rect 2462 -5840 2496 -5584
rect 2640 -5840 2674 -5584
<< psubdiff >>
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect 13619 -7731 13719 -7621
rect -7605 -17459 -7505 -17268
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< nsubdiff >>
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect 3610 -1520 3703 -1353
rect -7605 -7140 -7512 -6976
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
<< psubdiffcont >>
rect -7264 -7621 13443 -7521
rect -7605 -17268 -7505 -7850
rect 13619 -17149 13719 -7731
rect -7323 -17559 13384 -17459
<< nsubdiffcont >>
rect -7379 -1353 3329 -1260
rect -7605 -6976 -7512 -1507
rect 3610 -6989 3703 -1520
rect -7282 -7233 3426 -7140
<< poly >>
rect -6234 -2039 -6158 -2023
rect -6234 -2056 -6218 -2039
rect -6256 -2073 -6218 -2056
rect -6174 -2056 -6158 -2039
rect -6056 -2039 -5980 -2023
rect -6056 -2056 -6040 -2039
rect -6174 -2073 -6136 -2056
rect -6256 -2120 -6136 -2073
rect -6078 -2073 -6040 -2056
rect -5996 -2056 -5980 -2039
rect -5878 -2039 -5802 -2023
rect -5878 -2056 -5862 -2039
rect -5996 -2073 -5958 -2056
rect -6078 -2120 -5958 -2073
rect -5900 -2073 -5862 -2056
rect -5818 -2056 -5802 -2039
rect -5700 -2039 -5624 -2023
rect -5700 -2056 -5684 -2039
rect -5818 -2073 -5780 -2056
rect -5900 -2120 -5780 -2073
rect -5722 -2073 -5684 -2056
rect -5640 -2056 -5624 -2039
rect -5522 -2039 -5446 -2023
rect -5522 -2056 -5506 -2039
rect -5640 -2073 -5602 -2056
rect -5722 -2120 -5602 -2073
rect -5544 -2073 -5506 -2056
rect -5462 -2056 -5446 -2039
rect -5344 -2039 -5268 -2023
rect -5344 -2056 -5328 -2039
rect -5462 -2073 -5424 -2056
rect -5544 -2120 -5424 -2073
rect -5366 -2073 -5328 -2056
rect -5284 -2056 -5268 -2039
rect -5166 -2039 -5090 -2023
rect -5166 -2056 -5150 -2039
rect -5284 -2073 -5246 -2056
rect -5366 -2120 -5246 -2073
rect -5188 -2073 -5150 -2056
rect -5106 -2056 -5090 -2039
rect -4988 -2039 -4912 -2023
rect -4988 -2056 -4972 -2039
rect -5106 -2073 -5068 -2056
rect -5188 -2120 -5068 -2073
rect -5010 -2073 -4972 -2056
rect -4928 -2056 -4912 -2039
rect -4810 -2039 -4734 -2023
rect -4810 -2056 -4794 -2039
rect -4928 -2073 -4890 -2056
rect -5010 -2120 -4890 -2073
rect -4832 -2073 -4794 -2056
rect -4750 -2056 -4734 -2039
rect -4632 -2039 -4556 -2023
rect -4632 -2056 -4616 -2039
rect -4750 -2073 -4712 -2056
rect -4832 -2120 -4712 -2073
rect -4654 -2073 -4616 -2056
rect -4572 -2056 -4556 -2039
rect -4454 -2039 -4378 -2023
rect -4454 -2056 -4438 -2039
rect -4572 -2073 -4534 -2056
rect -4654 -2120 -4534 -2073
rect -4476 -2073 -4438 -2056
rect -4394 -2056 -4378 -2039
rect -4276 -2039 -4200 -2023
rect -4276 -2056 -4260 -2039
rect -4394 -2073 -4356 -2056
rect -4476 -2120 -4356 -2073
rect -4298 -2073 -4260 -2056
rect -4216 -2056 -4200 -2039
rect -4098 -2039 -4022 -2023
rect -4098 -2056 -4082 -2039
rect -4216 -2073 -4178 -2056
rect -4298 -2120 -4178 -2073
rect -4120 -2073 -4082 -2056
rect -4038 -2056 -4022 -2039
rect -3920 -2039 -3844 -2023
rect -3920 -2056 -3904 -2039
rect -4038 -2073 -4000 -2056
rect -4120 -2120 -4000 -2073
rect -3942 -2073 -3904 -2056
rect -3860 -2056 -3844 -2039
rect -3742 -2039 -3666 -2023
rect -3742 -2056 -3726 -2039
rect -3860 -2073 -3822 -2056
rect -3942 -2120 -3822 -2073
rect -3764 -2073 -3726 -2056
rect -3682 -2056 -3666 -2039
rect -3564 -2039 -3488 -2023
rect -3564 -2056 -3548 -2039
rect -3682 -2073 -3644 -2056
rect -3764 -2120 -3644 -2073
rect -3586 -2073 -3548 -2056
rect -3504 -2056 -3488 -2039
rect -3504 -2073 -3466 -2056
rect -3586 -2120 -3466 -2073
rect -6256 -2447 -6136 -2400
rect -6256 -2464 -6218 -2447
rect -6234 -2481 -6218 -2464
rect -6174 -2464 -6136 -2447
rect -6078 -2447 -5958 -2400
rect -6078 -2464 -6040 -2447
rect -6174 -2481 -6158 -2464
rect -6234 -2497 -6158 -2481
rect -6056 -2481 -6040 -2464
rect -5996 -2464 -5958 -2447
rect -5900 -2447 -5780 -2400
rect -5900 -2464 -5862 -2447
rect -5996 -2481 -5980 -2464
rect -6056 -2497 -5980 -2481
rect -5878 -2481 -5862 -2464
rect -5818 -2464 -5780 -2447
rect -5722 -2447 -5602 -2400
rect -5722 -2464 -5684 -2447
rect -5818 -2481 -5802 -2464
rect -5878 -2497 -5802 -2481
rect -5700 -2481 -5684 -2464
rect -5640 -2464 -5602 -2447
rect -5544 -2447 -5424 -2400
rect -5544 -2464 -5506 -2447
rect -5640 -2481 -5624 -2464
rect -5700 -2497 -5624 -2481
rect -5522 -2481 -5506 -2464
rect -5462 -2464 -5424 -2447
rect -5366 -2447 -5246 -2400
rect -5366 -2464 -5328 -2447
rect -5462 -2481 -5446 -2464
rect -5522 -2497 -5446 -2481
rect -5344 -2481 -5328 -2464
rect -5284 -2464 -5246 -2447
rect -5188 -2447 -5068 -2400
rect -5188 -2464 -5150 -2447
rect -5284 -2481 -5268 -2464
rect -5344 -2497 -5268 -2481
rect -5166 -2481 -5150 -2464
rect -5106 -2464 -5068 -2447
rect -5010 -2447 -4890 -2400
rect -5010 -2464 -4972 -2447
rect -5106 -2481 -5090 -2464
rect -5166 -2497 -5090 -2481
rect -4988 -2481 -4972 -2464
rect -4928 -2464 -4890 -2447
rect -4832 -2447 -4712 -2400
rect -4832 -2464 -4794 -2447
rect -4928 -2481 -4912 -2464
rect -4988 -2497 -4912 -2481
rect -4810 -2481 -4794 -2464
rect -4750 -2464 -4712 -2447
rect -4654 -2447 -4534 -2400
rect -4654 -2464 -4616 -2447
rect -4750 -2481 -4734 -2464
rect -4810 -2497 -4734 -2481
rect -4632 -2481 -4616 -2464
rect -4572 -2464 -4534 -2447
rect -4476 -2447 -4356 -2400
rect -4476 -2464 -4438 -2447
rect -4572 -2481 -4556 -2464
rect -4632 -2497 -4556 -2481
rect -4454 -2481 -4438 -2464
rect -4394 -2464 -4356 -2447
rect -4298 -2447 -4178 -2400
rect -4298 -2464 -4260 -2447
rect -4394 -2481 -4378 -2464
rect -4454 -2497 -4378 -2481
rect -4276 -2481 -4260 -2464
rect -4216 -2464 -4178 -2447
rect -4120 -2447 -4000 -2400
rect -4120 -2464 -4082 -2447
rect -4216 -2481 -4200 -2464
rect -4276 -2497 -4200 -2481
rect -4098 -2481 -4082 -2464
rect -4038 -2464 -4000 -2447
rect -3942 -2447 -3822 -2400
rect -3942 -2464 -3904 -2447
rect -4038 -2481 -4022 -2464
rect -4098 -2497 -4022 -2481
rect -3920 -2481 -3904 -2464
rect -3860 -2464 -3822 -2447
rect -3764 -2447 -3644 -2400
rect -3764 -2464 -3726 -2447
rect -3860 -2481 -3844 -2464
rect -3920 -2497 -3844 -2481
rect -3742 -2481 -3726 -2464
rect -3682 -2464 -3644 -2447
rect -3586 -2447 -3466 -2400
rect -3586 -2464 -3548 -2447
rect -3682 -2481 -3666 -2464
rect -3742 -2497 -3666 -2481
rect -3564 -2481 -3548 -2464
rect -3504 -2464 -3466 -2447
rect -3504 -2481 -3488 -2464
rect -3564 -2497 -3488 -2481
rect -1386 -2791 -1310 -2775
rect -1386 -2808 -1370 -2791
rect -1408 -2825 -1370 -2808
rect -1326 -2808 -1310 -2791
rect -1208 -2791 -1132 -2775
rect -1208 -2808 -1192 -2791
rect -1326 -2825 -1288 -2808
rect -1408 -2872 -1288 -2825
rect -1230 -2825 -1192 -2808
rect -1148 -2808 -1132 -2791
rect -1030 -2791 -954 -2775
rect -1030 -2808 -1014 -2791
rect -1148 -2825 -1110 -2808
rect -1230 -2872 -1110 -2825
rect -1052 -2825 -1014 -2808
rect -970 -2808 -954 -2791
rect -852 -2791 -776 -2775
rect -852 -2808 -836 -2791
rect -970 -2825 -932 -2808
rect -1052 -2872 -932 -2825
rect -874 -2825 -836 -2808
rect -792 -2808 -776 -2791
rect -674 -2791 -598 -2775
rect -674 -2808 -658 -2791
rect -792 -2825 -754 -2808
rect -874 -2872 -754 -2825
rect -696 -2825 -658 -2808
rect -614 -2808 -598 -2791
rect -496 -2791 -420 -2775
rect -496 -2808 -480 -2791
rect -614 -2825 -576 -2808
rect -696 -2872 -576 -2825
rect -518 -2825 -480 -2808
rect -436 -2808 -420 -2791
rect -318 -2791 -242 -2775
rect -318 -2808 -302 -2791
rect -436 -2825 -398 -2808
rect -518 -2872 -398 -2825
rect -340 -2825 -302 -2808
rect -258 -2808 -242 -2791
rect -140 -2791 -64 -2775
rect -140 -2808 -124 -2791
rect -258 -2825 -220 -2808
rect -340 -2872 -220 -2825
rect -162 -2825 -124 -2808
rect -80 -2808 -64 -2791
rect 38 -2791 114 -2775
rect 38 -2808 54 -2791
rect -80 -2825 -42 -2808
rect -162 -2872 -42 -2825
rect 16 -2825 54 -2808
rect 98 -2808 114 -2791
rect 216 -2791 292 -2775
rect 216 -2808 232 -2791
rect 98 -2825 136 -2808
rect 16 -2872 136 -2825
rect 194 -2825 232 -2808
rect 276 -2808 292 -2791
rect 394 -2791 470 -2775
rect 394 -2808 410 -2791
rect 276 -2825 314 -2808
rect 194 -2872 314 -2825
rect 372 -2825 410 -2808
rect 454 -2808 470 -2791
rect 572 -2791 648 -2775
rect 572 -2808 588 -2791
rect 454 -2825 492 -2808
rect 372 -2872 492 -2825
rect 550 -2825 588 -2808
rect 632 -2808 648 -2791
rect 750 -2791 826 -2775
rect 750 -2808 766 -2791
rect 632 -2825 670 -2808
rect 550 -2872 670 -2825
rect 728 -2825 766 -2808
rect 810 -2808 826 -2791
rect 928 -2791 1004 -2775
rect 928 -2808 944 -2791
rect 810 -2825 848 -2808
rect 728 -2872 848 -2825
rect 906 -2825 944 -2808
rect 988 -2808 1004 -2791
rect 1106 -2791 1182 -2775
rect 1106 -2808 1122 -2791
rect 988 -2825 1026 -2808
rect 906 -2872 1026 -2825
rect 1084 -2825 1122 -2808
rect 1166 -2808 1182 -2791
rect 1284 -2791 1360 -2775
rect 1284 -2808 1300 -2791
rect 1166 -2825 1204 -2808
rect 1084 -2872 1204 -2825
rect 1262 -2825 1300 -2808
rect 1344 -2808 1360 -2791
rect 1462 -2791 1538 -2775
rect 1462 -2808 1478 -2791
rect 1344 -2825 1382 -2808
rect 1262 -2872 1382 -2825
rect 1440 -2825 1478 -2808
rect 1522 -2808 1538 -2791
rect 1640 -2791 1716 -2775
rect 1640 -2808 1656 -2791
rect 1522 -2825 1560 -2808
rect 1440 -2872 1560 -2825
rect 1618 -2825 1656 -2808
rect 1700 -2808 1716 -2791
rect 1818 -2791 1894 -2775
rect 1818 -2808 1834 -2791
rect 1700 -2825 1738 -2808
rect 1618 -2872 1738 -2825
rect 1796 -2825 1834 -2808
rect 1878 -2808 1894 -2791
rect 1996 -2791 2072 -2775
rect 1996 -2808 2012 -2791
rect 1878 -2825 1916 -2808
rect 1796 -2872 1916 -2825
rect 1974 -2825 2012 -2808
rect 2056 -2808 2072 -2791
rect 2174 -2791 2250 -2775
rect 2174 -2808 2190 -2791
rect 2056 -2825 2094 -2808
rect 1974 -2872 2094 -2825
rect 2152 -2825 2190 -2808
rect 2234 -2808 2250 -2791
rect 2352 -2791 2428 -2775
rect 2352 -2808 2368 -2791
rect 2234 -2825 2272 -2808
rect 2152 -2872 2272 -2825
rect 2330 -2825 2368 -2808
rect 2412 -2808 2428 -2791
rect 2530 -2791 2606 -2775
rect 2530 -2808 2546 -2791
rect 2412 -2825 2450 -2808
rect 2330 -2872 2450 -2825
rect 2508 -2825 2546 -2808
rect 2590 -2808 2606 -2791
rect 2590 -2825 2628 -2808
rect 2508 -2872 2628 -2825
rect -6234 -2909 -6158 -2893
rect -6234 -2926 -6218 -2909
rect -6256 -2943 -6218 -2926
rect -6174 -2926 -6158 -2909
rect -6056 -2909 -5980 -2893
rect -6056 -2926 -6040 -2909
rect -6174 -2943 -6136 -2926
rect -6256 -2990 -6136 -2943
rect -6078 -2943 -6040 -2926
rect -5996 -2926 -5980 -2909
rect -5878 -2909 -5802 -2893
rect -5878 -2926 -5862 -2909
rect -5996 -2943 -5958 -2926
rect -6078 -2990 -5958 -2943
rect -5900 -2943 -5862 -2926
rect -5818 -2926 -5802 -2909
rect -5700 -2909 -5624 -2893
rect -5700 -2926 -5684 -2909
rect -5818 -2943 -5780 -2926
rect -5900 -2990 -5780 -2943
rect -5722 -2943 -5684 -2926
rect -5640 -2926 -5624 -2909
rect -5522 -2909 -5446 -2893
rect -5522 -2926 -5506 -2909
rect -5640 -2943 -5602 -2926
rect -5722 -2990 -5602 -2943
rect -5544 -2943 -5506 -2926
rect -5462 -2926 -5446 -2909
rect -5344 -2909 -5268 -2893
rect -5344 -2926 -5328 -2909
rect -5462 -2943 -5424 -2926
rect -5544 -2990 -5424 -2943
rect -5366 -2943 -5328 -2926
rect -5284 -2926 -5268 -2909
rect -5166 -2909 -5090 -2893
rect -5166 -2926 -5150 -2909
rect -5284 -2943 -5246 -2926
rect -5366 -2990 -5246 -2943
rect -5188 -2943 -5150 -2926
rect -5106 -2926 -5090 -2909
rect -4988 -2909 -4912 -2893
rect -4988 -2926 -4972 -2909
rect -5106 -2943 -5068 -2926
rect -5188 -2990 -5068 -2943
rect -5010 -2943 -4972 -2926
rect -4928 -2926 -4912 -2909
rect -4810 -2909 -4734 -2893
rect -4810 -2926 -4794 -2909
rect -4928 -2943 -4890 -2926
rect -5010 -2990 -4890 -2943
rect -4832 -2943 -4794 -2926
rect -4750 -2926 -4734 -2909
rect -4632 -2909 -4556 -2893
rect -4632 -2926 -4616 -2909
rect -4750 -2943 -4712 -2926
rect -4832 -2990 -4712 -2943
rect -4654 -2943 -4616 -2926
rect -4572 -2926 -4556 -2909
rect -4454 -2909 -4378 -2893
rect -4454 -2926 -4438 -2909
rect -4572 -2943 -4534 -2926
rect -4654 -2990 -4534 -2943
rect -4476 -2943 -4438 -2926
rect -4394 -2926 -4378 -2909
rect -4276 -2909 -4200 -2893
rect -4276 -2926 -4260 -2909
rect -4394 -2943 -4356 -2926
rect -4476 -2990 -4356 -2943
rect -4298 -2943 -4260 -2926
rect -4216 -2926 -4200 -2909
rect -4098 -2909 -4022 -2893
rect -4098 -2926 -4082 -2909
rect -4216 -2943 -4178 -2926
rect -4298 -2990 -4178 -2943
rect -4120 -2943 -4082 -2926
rect -4038 -2926 -4022 -2909
rect -3920 -2909 -3844 -2893
rect -3920 -2926 -3904 -2909
rect -4038 -2943 -4000 -2926
rect -4120 -2990 -4000 -2943
rect -3942 -2943 -3904 -2926
rect -3860 -2926 -3844 -2909
rect -3742 -2909 -3666 -2893
rect -3742 -2926 -3726 -2909
rect -3860 -2943 -3822 -2926
rect -3942 -2990 -3822 -2943
rect -3764 -2943 -3726 -2926
rect -3682 -2926 -3666 -2909
rect -3564 -2909 -3488 -2893
rect -3564 -2926 -3548 -2909
rect -3682 -2943 -3644 -2926
rect -3764 -2990 -3644 -2943
rect -3586 -2943 -3548 -2926
rect -3504 -2926 -3488 -2909
rect -3504 -2943 -3466 -2926
rect -3586 -2990 -3466 -2943
rect -1408 -3199 -1288 -3152
rect -1408 -3216 -1370 -3199
rect -1386 -3233 -1370 -3216
rect -1326 -3216 -1288 -3199
rect -1230 -3199 -1110 -3152
rect -1230 -3216 -1192 -3199
rect -1326 -3233 -1310 -3216
rect -1386 -3249 -1310 -3233
rect -1208 -3233 -1192 -3216
rect -1148 -3216 -1110 -3199
rect -1052 -3199 -932 -3152
rect -1052 -3216 -1014 -3199
rect -1148 -3233 -1132 -3216
rect -1208 -3249 -1132 -3233
rect -1030 -3233 -1014 -3216
rect -970 -3216 -932 -3199
rect -874 -3199 -754 -3152
rect -874 -3216 -836 -3199
rect -970 -3233 -954 -3216
rect -1030 -3249 -954 -3233
rect -852 -3233 -836 -3216
rect -792 -3216 -754 -3199
rect -696 -3199 -576 -3152
rect -696 -3216 -658 -3199
rect -792 -3233 -776 -3216
rect -852 -3249 -776 -3233
rect -674 -3233 -658 -3216
rect -614 -3216 -576 -3199
rect -518 -3199 -398 -3152
rect -518 -3216 -480 -3199
rect -614 -3233 -598 -3216
rect -674 -3249 -598 -3233
rect -496 -3233 -480 -3216
rect -436 -3216 -398 -3199
rect -340 -3199 -220 -3152
rect -340 -3216 -302 -3199
rect -436 -3233 -420 -3216
rect -496 -3249 -420 -3233
rect -318 -3233 -302 -3216
rect -258 -3216 -220 -3199
rect -162 -3199 -42 -3152
rect -162 -3216 -124 -3199
rect -258 -3233 -242 -3216
rect -318 -3249 -242 -3233
rect -140 -3233 -124 -3216
rect -80 -3216 -42 -3199
rect 16 -3199 136 -3152
rect 16 -3216 54 -3199
rect -80 -3233 -64 -3216
rect -140 -3249 -64 -3233
rect 38 -3233 54 -3216
rect 98 -3216 136 -3199
rect 194 -3199 314 -3152
rect 194 -3216 232 -3199
rect 98 -3233 114 -3216
rect 38 -3249 114 -3233
rect 216 -3233 232 -3216
rect 276 -3216 314 -3199
rect 372 -3199 492 -3152
rect 372 -3216 410 -3199
rect 276 -3233 292 -3216
rect 216 -3249 292 -3233
rect 394 -3233 410 -3216
rect 454 -3216 492 -3199
rect 550 -3199 670 -3152
rect 550 -3216 588 -3199
rect 454 -3233 470 -3216
rect 394 -3249 470 -3233
rect 572 -3233 588 -3216
rect 632 -3216 670 -3199
rect 728 -3199 848 -3152
rect 728 -3216 766 -3199
rect 632 -3233 648 -3216
rect 572 -3249 648 -3233
rect 750 -3233 766 -3216
rect 810 -3216 848 -3199
rect 906 -3199 1026 -3152
rect 906 -3216 944 -3199
rect 810 -3233 826 -3216
rect 750 -3249 826 -3233
rect 928 -3233 944 -3216
rect 988 -3216 1026 -3199
rect 1084 -3199 1204 -3152
rect 1084 -3216 1122 -3199
rect 988 -3233 1004 -3216
rect 928 -3249 1004 -3233
rect 1106 -3233 1122 -3216
rect 1166 -3216 1204 -3199
rect 1262 -3199 1382 -3152
rect 1262 -3216 1300 -3199
rect 1166 -3233 1182 -3216
rect 1106 -3249 1182 -3233
rect 1284 -3233 1300 -3216
rect 1344 -3216 1382 -3199
rect 1440 -3199 1560 -3152
rect 1440 -3216 1478 -3199
rect 1344 -3233 1360 -3216
rect 1284 -3249 1360 -3233
rect 1462 -3233 1478 -3216
rect 1522 -3216 1560 -3199
rect 1618 -3199 1738 -3152
rect 1618 -3216 1656 -3199
rect 1522 -3233 1538 -3216
rect 1462 -3249 1538 -3233
rect 1640 -3233 1656 -3216
rect 1700 -3216 1738 -3199
rect 1796 -3199 1916 -3152
rect 1796 -3216 1834 -3199
rect 1700 -3233 1716 -3216
rect 1640 -3249 1716 -3233
rect 1818 -3233 1834 -3216
rect 1878 -3216 1916 -3199
rect 1974 -3199 2094 -3152
rect 1974 -3216 2012 -3199
rect 1878 -3233 1894 -3216
rect 1818 -3249 1894 -3233
rect 1996 -3233 2012 -3216
rect 2056 -3216 2094 -3199
rect 2152 -3199 2272 -3152
rect 2152 -3216 2190 -3199
rect 2056 -3233 2072 -3216
rect 1996 -3249 2072 -3233
rect 2174 -3233 2190 -3216
rect 2234 -3216 2272 -3199
rect 2330 -3199 2450 -3152
rect 2330 -3216 2368 -3199
rect 2234 -3233 2250 -3216
rect 2174 -3249 2250 -3233
rect 2352 -3233 2368 -3216
rect 2412 -3216 2450 -3199
rect 2508 -3199 2628 -3152
rect 2508 -3216 2546 -3199
rect 2412 -3233 2428 -3216
rect 2352 -3249 2428 -3233
rect 2530 -3233 2546 -3216
rect 2590 -3216 2628 -3199
rect 2590 -3233 2606 -3216
rect 2530 -3249 2606 -3233
rect -6256 -3317 -6136 -3270
rect -6256 -3334 -6218 -3317
rect -6234 -3351 -6218 -3334
rect -6174 -3334 -6136 -3317
rect -6078 -3317 -5958 -3270
rect -6078 -3334 -6040 -3317
rect -6174 -3351 -6158 -3334
rect -6234 -3367 -6158 -3351
rect -6056 -3351 -6040 -3334
rect -5996 -3334 -5958 -3317
rect -5900 -3317 -5780 -3270
rect -5900 -3334 -5862 -3317
rect -5996 -3351 -5980 -3334
rect -6056 -3367 -5980 -3351
rect -5878 -3351 -5862 -3334
rect -5818 -3334 -5780 -3317
rect -5722 -3317 -5602 -3270
rect -5722 -3334 -5684 -3317
rect -5818 -3351 -5802 -3334
rect -5878 -3367 -5802 -3351
rect -5700 -3351 -5684 -3334
rect -5640 -3334 -5602 -3317
rect -5544 -3317 -5424 -3270
rect -5544 -3334 -5506 -3317
rect -5640 -3351 -5624 -3334
rect -5700 -3367 -5624 -3351
rect -5522 -3351 -5506 -3334
rect -5462 -3334 -5424 -3317
rect -5366 -3317 -5246 -3270
rect -5366 -3334 -5328 -3317
rect -5462 -3351 -5446 -3334
rect -5522 -3367 -5446 -3351
rect -5344 -3351 -5328 -3334
rect -5284 -3334 -5246 -3317
rect -5188 -3317 -5068 -3270
rect -5188 -3334 -5150 -3317
rect -5284 -3351 -5268 -3334
rect -5344 -3367 -5268 -3351
rect -5166 -3351 -5150 -3334
rect -5106 -3334 -5068 -3317
rect -5010 -3317 -4890 -3270
rect -5010 -3334 -4972 -3317
rect -5106 -3351 -5090 -3334
rect -5166 -3367 -5090 -3351
rect -4988 -3351 -4972 -3334
rect -4928 -3334 -4890 -3317
rect -4832 -3317 -4712 -3270
rect -4832 -3334 -4794 -3317
rect -4928 -3351 -4912 -3334
rect -4988 -3367 -4912 -3351
rect -4810 -3351 -4794 -3334
rect -4750 -3334 -4712 -3317
rect -4654 -3317 -4534 -3270
rect -4654 -3334 -4616 -3317
rect -4750 -3351 -4734 -3334
rect -4810 -3367 -4734 -3351
rect -4632 -3351 -4616 -3334
rect -4572 -3334 -4534 -3317
rect -4476 -3317 -4356 -3270
rect -4476 -3334 -4438 -3317
rect -4572 -3351 -4556 -3334
rect -4632 -3367 -4556 -3351
rect -4454 -3351 -4438 -3334
rect -4394 -3334 -4356 -3317
rect -4298 -3317 -4178 -3270
rect -4298 -3334 -4260 -3317
rect -4394 -3351 -4378 -3334
rect -4454 -3367 -4378 -3351
rect -4276 -3351 -4260 -3334
rect -4216 -3334 -4178 -3317
rect -4120 -3317 -4000 -3270
rect -4120 -3334 -4082 -3317
rect -4216 -3351 -4200 -3334
rect -4276 -3367 -4200 -3351
rect -4098 -3351 -4082 -3334
rect -4038 -3334 -4000 -3317
rect -3942 -3317 -3822 -3270
rect -3942 -3334 -3904 -3317
rect -4038 -3351 -4022 -3334
rect -4098 -3367 -4022 -3351
rect -3920 -3351 -3904 -3334
rect -3860 -3334 -3822 -3317
rect -3764 -3317 -3644 -3270
rect -3764 -3334 -3726 -3317
rect -3860 -3351 -3844 -3334
rect -3920 -3367 -3844 -3351
rect -3742 -3351 -3726 -3334
rect -3682 -3334 -3644 -3317
rect -3586 -3317 -3466 -3270
rect -3586 -3334 -3548 -3317
rect -3682 -3351 -3666 -3334
rect -3742 -3367 -3666 -3351
rect -3564 -3351 -3548 -3334
rect -3504 -3334 -3466 -3317
rect -3504 -3351 -3488 -3334
rect -3564 -3367 -3488 -3351
rect -1386 -3691 -1310 -3675
rect -1386 -3708 -1370 -3691
rect -1408 -3725 -1370 -3708
rect -1326 -3708 -1310 -3691
rect -1208 -3691 -1132 -3675
rect -1208 -3708 -1192 -3691
rect -1326 -3725 -1288 -3708
rect -6234 -3779 -6158 -3763
rect -6234 -3796 -6218 -3779
rect -6256 -3813 -6218 -3796
rect -6174 -3796 -6158 -3779
rect -6056 -3779 -5980 -3763
rect -6056 -3796 -6040 -3779
rect -6174 -3813 -6136 -3796
rect -6256 -3860 -6136 -3813
rect -6078 -3813 -6040 -3796
rect -5996 -3796 -5980 -3779
rect -5878 -3779 -5802 -3763
rect -5878 -3796 -5862 -3779
rect -5996 -3813 -5958 -3796
rect -6078 -3860 -5958 -3813
rect -5900 -3813 -5862 -3796
rect -5818 -3796 -5802 -3779
rect -5700 -3779 -5624 -3763
rect -5700 -3796 -5684 -3779
rect -5818 -3813 -5780 -3796
rect -5900 -3860 -5780 -3813
rect -5722 -3813 -5684 -3796
rect -5640 -3796 -5624 -3779
rect -5522 -3779 -5446 -3763
rect -5522 -3796 -5506 -3779
rect -5640 -3813 -5602 -3796
rect -5722 -3860 -5602 -3813
rect -5544 -3813 -5506 -3796
rect -5462 -3796 -5446 -3779
rect -5344 -3779 -5268 -3763
rect -5344 -3796 -5328 -3779
rect -5462 -3813 -5424 -3796
rect -5544 -3860 -5424 -3813
rect -5366 -3813 -5328 -3796
rect -5284 -3796 -5268 -3779
rect -5166 -3779 -5090 -3763
rect -5166 -3796 -5150 -3779
rect -5284 -3813 -5246 -3796
rect -5366 -3860 -5246 -3813
rect -5188 -3813 -5150 -3796
rect -5106 -3796 -5090 -3779
rect -4988 -3779 -4912 -3763
rect -4988 -3796 -4972 -3779
rect -5106 -3813 -5068 -3796
rect -5188 -3860 -5068 -3813
rect -5010 -3813 -4972 -3796
rect -4928 -3796 -4912 -3779
rect -4810 -3779 -4734 -3763
rect -4810 -3796 -4794 -3779
rect -4928 -3813 -4890 -3796
rect -5010 -3860 -4890 -3813
rect -4832 -3813 -4794 -3796
rect -4750 -3796 -4734 -3779
rect -4632 -3779 -4556 -3763
rect -4632 -3796 -4616 -3779
rect -4750 -3813 -4712 -3796
rect -4832 -3860 -4712 -3813
rect -4654 -3813 -4616 -3796
rect -4572 -3796 -4556 -3779
rect -4454 -3779 -4378 -3763
rect -4454 -3796 -4438 -3779
rect -4572 -3813 -4534 -3796
rect -4654 -3860 -4534 -3813
rect -4476 -3813 -4438 -3796
rect -4394 -3796 -4378 -3779
rect -4276 -3779 -4200 -3763
rect -4276 -3796 -4260 -3779
rect -4394 -3813 -4356 -3796
rect -4476 -3860 -4356 -3813
rect -4298 -3813 -4260 -3796
rect -4216 -3796 -4200 -3779
rect -4098 -3779 -4022 -3763
rect -4098 -3796 -4082 -3779
rect -4216 -3813 -4178 -3796
rect -4298 -3860 -4178 -3813
rect -4120 -3813 -4082 -3796
rect -4038 -3796 -4022 -3779
rect -3920 -3779 -3844 -3763
rect -3920 -3796 -3904 -3779
rect -4038 -3813 -4000 -3796
rect -4120 -3860 -4000 -3813
rect -3942 -3813 -3904 -3796
rect -3860 -3796 -3844 -3779
rect -3742 -3779 -3666 -3763
rect -3742 -3796 -3726 -3779
rect -3860 -3813 -3822 -3796
rect -3942 -3860 -3822 -3813
rect -3764 -3813 -3726 -3796
rect -3682 -3796 -3666 -3779
rect -3564 -3779 -3488 -3763
rect -1408 -3772 -1288 -3725
rect -1230 -3725 -1192 -3708
rect -1148 -3708 -1132 -3691
rect -1030 -3691 -954 -3675
rect -1030 -3708 -1014 -3691
rect -1148 -3725 -1110 -3708
rect -1230 -3772 -1110 -3725
rect -1052 -3725 -1014 -3708
rect -970 -3708 -954 -3691
rect -852 -3691 -776 -3675
rect -852 -3708 -836 -3691
rect -970 -3725 -932 -3708
rect -1052 -3772 -932 -3725
rect -874 -3725 -836 -3708
rect -792 -3708 -776 -3691
rect -674 -3691 -598 -3675
rect -674 -3708 -658 -3691
rect -792 -3725 -754 -3708
rect -874 -3772 -754 -3725
rect -696 -3725 -658 -3708
rect -614 -3708 -598 -3691
rect -496 -3691 -420 -3675
rect -496 -3708 -480 -3691
rect -614 -3725 -576 -3708
rect -696 -3772 -576 -3725
rect -518 -3725 -480 -3708
rect -436 -3708 -420 -3691
rect -318 -3691 -242 -3675
rect -318 -3708 -302 -3691
rect -436 -3725 -398 -3708
rect -518 -3772 -398 -3725
rect -340 -3725 -302 -3708
rect -258 -3708 -242 -3691
rect -140 -3691 -64 -3675
rect -140 -3708 -124 -3691
rect -258 -3725 -220 -3708
rect -340 -3772 -220 -3725
rect -162 -3725 -124 -3708
rect -80 -3708 -64 -3691
rect 38 -3691 114 -3675
rect 38 -3708 54 -3691
rect -80 -3725 -42 -3708
rect -162 -3772 -42 -3725
rect 16 -3725 54 -3708
rect 98 -3708 114 -3691
rect 216 -3691 292 -3675
rect 216 -3708 232 -3691
rect 98 -3725 136 -3708
rect 16 -3772 136 -3725
rect 194 -3725 232 -3708
rect 276 -3708 292 -3691
rect 394 -3691 470 -3675
rect 394 -3708 410 -3691
rect 276 -3725 314 -3708
rect 194 -3772 314 -3725
rect 372 -3725 410 -3708
rect 454 -3708 470 -3691
rect 572 -3691 648 -3675
rect 572 -3708 588 -3691
rect 454 -3725 492 -3708
rect 372 -3772 492 -3725
rect 550 -3725 588 -3708
rect 632 -3708 648 -3691
rect 750 -3691 826 -3675
rect 750 -3708 766 -3691
rect 632 -3725 670 -3708
rect 550 -3772 670 -3725
rect 728 -3725 766 -3708
rect 810 -3708 826 -3691
rect 928 -3691 1004 -3675
rect 928 -3708 944 -3691
rect 810 -3725 848 -3708
rect 728 -3772 848 -3725
rect 906 -3725 944 -3708
rect 988 -3708 1004 -3691
rect 1106 -3691 1182 -3675
rect 1106 -3708 1122 -3691
rect 988 -3725 1026 -3708
rect 906 -3772 1026 -3725
rect 1084 -3725 1122 -3708
rect 1166 -3708 1182 -3691
rect 1284 -3691 1360 -3675
rect 1284 -3708 1300 -3691
rect 1166 -3725 1204 -3708
rect 1084 -3772 1204 -3725
rect 1262 -3725 1300 -3708
rect 1344 -3708 1360 -3691
rect 1462 -3691 1538 -3675
rect 1462 -3708 1478 -3691
rect 1344 -3725 1382 -3708
rect 1262 -3772 1382 -3725
rect 1440 -3725 1478 -3708
rect 1522 -3708 1538 -3691
rect 1640 -3691 1716 -3675
rect 1640 -3708 1656 -3691
rect 1522 -3725 1560 -3708
rect 1440 -3772 1560 -3725
rect 1618 -3725 1656 -3708
rect 1700 -3708 1716 -3691
rect 1818 -3691 1894 -3675
rect 1818 -3708 1834 -3691
rect 1700 -3725 1738 -3708
rect 1618 -3772 1738 -3725
rect 1796 -3725 1834 -3708
rect 1878 -3708 1894 -3691
rect 1996 -3691 2072 -3675
rect 1996 -3708 2012 -3691
rect 1878 -3725 1916 -3708
rect 1796 -3772 1916 -3725
rect 1974 -3725 2012 -3708
rect 2056 -3708 2072 -3691
rect 2174 -3691 2250 -3675
rect 2174 -3708 2190 -3691
rect 2056 -3725 2094 -3708
rect 1974 -3772 2094 -3725
rect 2152 -3725 2190 -3708
rect 2234 -3708 2250 -3691
rect 2352 -3691 2428 -3675
rect 2352 -3708 2368 -3691
rect 2234 -3725 2272 -3708
rect 2152 -3772 2272 -3725
rect 2330 -3725 2368 -3708
rect 2412 -3708 2428 -3691
rect 2530 -3691 2606 -3675
rect 2530 -3708 2546 -3691
rect 2412 -3725 2450 -3708
rect 2330 -3772 2450 -3725
rect 2508 -3725 2546 -3708
rect 2590 -3708 2606 -3691
rect 2590 -3725 2628 -3708
rect 2508 -3772 2628 -3725
rect -3564 -3796 -3548 -3779
rect -3682 -3813 -3644 -3796
rect -3764 -3860 -3644 -3813
rect -3586 -3813 -3548 -3796
rect -3504 -3796 -3488 -3779
rect -3504 -3813 -3466 -3796
rect -3586 -3860 -3466 -3813
rect -1408 -4099 -1288 -4052
rect -1408 -4116 -1370 -4099
rect -1386 -4133 -1370 -4116
rect -1326 -4116 -1288 -4099
rect -1230 -4099 -1110 -4052
rect -1230 -4116 -1192 -4099
rect -1326 -4133 -1310 -4116
rect -6256 -4187 -6136 -4140
rect -6256 -4204 -6218 -4187
rect -6234 -4221 -6218 -4204
rect -6174 -4204 -6136 -4187
rect -6078 -4187 -5958 -4140
rect -6078 -4204 -6040 -4187
rect -6174 -4221 -6158 -4204
rect -6234 -4237 -6158 -4221
rect -6056 -4221 -6040 -4204
rect -5996 -4204 -5958 -4187
rect -5900 -4187 -5780 -4140
rect -5900 -4204 -5862 -4187
rect -5996 -4221 -5980 -4204
rect -6056 -4237 -5980 -4221
rect -5878 -4221 -5862 -4204
rect -5818 -4204 -5780 -4187
rect -5722 -4187 -5602 -4140
rect -5722 -4204 -5684 -4187
rect -5818 -4221 -5802 -4204
rect -5878 -4237 -5802 -4221
rect -5700 -4221 -5684 -4204
rect -5640 -4204 -5602 -4187
rect -5544 -4187 -5424 -4140
rect -5544 -4204 -5506 -4187
rect -5640 -4221 -5624 -4204
rect -5700 -4237 -5624 -4221
rect -5522 -4221 -5506 -4204
rect -5462 -4204 -5424 -4187
rect -5366 -4187 -5246 -4140
rect -5366 -4204 -5328 -4187
rect -5462 -4221 -5446 -4204
rect -5522 -4237 -5446 -4221
rect -5344 -4221 -5328 -4204
rect -5284 -4204 -5246 -4187
rect -5188 -4187 -5068 -4140
rect -5188 -4204 -5150 -4187
rect -5284 -4221 -5268 -4204
rect -5344 -4237 -5268 -4221
rect -5166 -4221 -5150 -4204
rect -5106 -4204 -5068 -4187
rect -5010 -4187 -4890 -4140
rect -5010 -4204 -4972 -4187
rect -5106 -4221 -5090 -4204
rect -5166 -4237 -5090 -4221
rect -4988 -4221 -4972 -4204
rect -4928 -4204 -4890 -4187
rect -4832 -4187 -4712 -4140
rect -4832 -4204 -4794 -4187
rect -4928 -4221 -4912 -4204
rect -4988 -4237 -4912 -4221
rect -4810 -4221 -4794 -4204
rect -4750 -4204 -4712 -4187
rect -4654 -4187 -4534 -4140
rect -4654 -4204 -4616 -4187
rect -4750 -4221 -4734 -4204
rect -4810 -4237 -4734 -4221
rect -4632 -4221 -4616 -4204
rect -4572 -4204 -4534 -4187
rect -4476 -4187 -4356 -4140
rect -4476 -4204 -4438 -4187
rect -4572 -4221 -4556 -4204
rect -4632 -4237 -4556 -4221
rect -4454 -4221 -4438 -4204
rect -4394 -4204 -4356 -4187
rect -4298 -4187 -4178 -4140
rect -4298 -4204 -4260 -4187
rect -4394 -4221 -4378 -4204
rect -4454 -4237 -4378 -4221
rect -4276 -4221 -4260 -4204
rect -4216 -4204 -4178 -4187
rect -4120 -4187 -4000 -4140
rect -4120 -4204 -4082 -4187
rect -4216 -4221 -4200 -4204
rect -4276 -4237 -4200 -4221
rect -4098 -4221 -4082 -4204
rect -4038 -4204 -4000 -4187
rect -3942 -4187 -3822 -4140
rect -3942 -4204 -3904 -4187
rect -4038 -4221 -4022 -4204
rect -4098 -4237 -4022 -4221
rect -3920 -4221 -3904 -4204
rect -3860 -4204 -3822 -4187
rect -3764 -4187 -3644 -4140
rect -3764 -4204 -3726 -4187
rect -3860 -4221 -3844 -4204
rect -3920 -4237 -3844 -4221
rect -3742 -4221 -3726 -4204
rect -3682 -4204 -3644 -4187
rect -3586 -4187 -3466 -4140
rect -1386 -4149 -1310 -4133
rect -1208 -4133 -1192 -4116
rect -1148 -4116 -1110 -4099
rect -1052 -4099 -932 -4052
rect -1052 -4116 -1014 -4099
rect -1148 -4133 -1132 -4116
rect -1208 -4149 -1132 -4133
rect -1030 -4133 -1014 -4116
rect -970 -4116 -932 -4099
rect -874 -4099 -754 -4052
rect -874 -4116 -836 -4099
rect -970 -4133 -954 -4116
rect -1030 -4149 -954 -4133
rect -852 -4133 -836 -4116
rect -792 -4116 -754 -4099
rect -696 -4099 -576 -4052
rect -696 -4116 -658 -4099
rect -792 -4133 -776 -4116
rect -852 -4149 -776 -4133
rect -674 -4133 -658 -4116
rect -614 -4116 -576 -4099
rect -518 -4099 -398 -4052
rect -518 -4116 -480 -4099
rect -614 -4133 -598 -4116
rect -674 -4149 -598 -4133
rect -496 -4133 -480 -4116
rect -436 -4116 -398 -4099
rect -340 -4099 -220 -4052
rect -340 -4116 -302 -4099
rect -436 -4133 -420 -4116
rect -496 -4149 -420 -4133
rect -318 -4133 -302 -4116
rect -258 -4116 -220 -4099
rect -162 -4099 -42 -4052
rect -162 -4116 -124 -4099
rect -258 -4133 -242 -4116
rect -318 -4149 -242 -4133
rect -140 -4133 -124 -4116
rect -80 -4116 -42 -4099
rect 16 -4099 136 -4052
rect 16 -4116 54 -4099
rect -80 -4133 -64 -4116
rect -140 -4149 -64 -4133
rect 38 -4133 54 -4116
rect 98 -4116 136 -4099
rect 194 -4099 314 -4052
rect 194 -4116 232 -4099
rect 98 -4133 114 -4116
rect 38 -4149 114 -4133
rect 216 -4133 232 -4116
rect 276 -4116 314 -4099
rect 372 -4099 492 -4052
rect 372 -4116 410 -4099
rect 276 -4133 292 -4116
rect 216 -4149 292 -4133
rect 394 -4133 410 -4116
rect 454 -4116 492 -4099
rect 550 -4099 670 -4052
rect 550 -4116 588 -4099
rect 454 -4133 470 -4116
rect 394 -4149 470 -4133
rect 572 -4133 588 -4116
rect 632 -4116 670 -4099
rect 728 -4099 848 -4052
rect 728 -4116 766 -4099
rect 632 -4133 648 -4116
rect 572 -4149 648 -4133
rect 750 -4133 766 -4116
rect 810 -4116 848 -4099
rect 906 -4099 1026 -4052
rect 906 -4116 944 -4099
rect 810 -4133 826 -4116
rect 750 -4149 826 -4133
rect 928 -4133 944 -4116
rect 988 -4116 1026 -4099
rect 1084 -4099 1204 -4052
rect 1084 -4116 1122 -4099
rect 988 -4133 1004 -4116
rect 928 -4149 1004 -4133
rect 1106 -4133 1122 -4116
rect 1166 -4116 1204 -4099
rect 1262 -4099 1382 -4052
rect 1262 -4116 1300 -4099
rect 1166 -4133 1182 -4116
rect 1106 -4149 1182 -4133
rect 1284 -4133 1300 -4116
rect 1344 -4116 1382 -4099
rect 1440 -4099 1560 -4052
rect 1440 -4116 1478 -4099
rect 1344 -4133 1360 -4116
rect 1284 -4149 1360 -4133
rect 1462 -4133 1478 -4116
rect 1522 -4116 1560 -4099
rect 1618 -4099 1738 -4052
rect 1618 -4116 1656 -4099
rect 1522 -4133 1538 -4116
rect 1462 -4149 1538 -4133
rect 1640 -4133 1656 -4116
rect 1700 -4116 1738 -4099
rect 1796 -4099 1916 -4052
rect 1796 -4116 1834 -4099
rect 1700 -4133 1716 -4116
rect 1640 -4149 1716 -4133
rect 1818 -4133 1834 -4116
rect 1878 -4116 1916 -4099
rect 1974 -4099 2094 -4052
rect 1974 -4116 2012 -4099
rect 1878 -4133 1894 -4116
rect 1818 -4149 1894 -4133
rect 1996 -4133 2012 -4116
rect 2056 -4116 2094 -4099
rect 2152 -4099 2272 -4052
rect 2152 -4116 2190 -4099
rect 2056 -4133 2072 -4116
rect 1996 -4149 2072 -4133
rect 2174 -4133 2190 -4116
rect 2234 -4116 2272 -4099
rect 2330 -4099 2450 -4052
rect 2330 -4116 2368 -4099
rect 2234 -4133 2250 -4116
rect 2174 -4149 2250 -4133
rect 2352 -4133 2368 -4116
rect 2412 -4116 2450 -4099
rect 2508 -4099 2628 -4052
rect 2508 -4116 2546 -4099
rect 2412 -4133 2428 -4116
rect 2352 -4149 2428 -4133
rect 2530 -4133 2546 -4116
rect 2590 -4116 2628 -4099
rect 2590 -4133 2606 -4116
rect 2530 -4149 2606 -4133
rect -3586 -4204 -3548 -4187
rect -3682 -4221 -3666 -4204
rect -3742 -4237 -3666 -4221
rect -3564 -4221 -3548 -4204
rect -3504 -4204 -3466 -4187
rect -3504 -4221 -3488 -4204
rect -3564 -4237 -3488 -4221
rect -1386 -4591 -1310 -4575
rect -1386 -4608 -1370 -4591
rect -1408 -4625 -1370 -4608
rect -1326 -4608 -1310 -4591
rect -1208 -4591 -1132 -4575
rect -1208 -4608 -1192 -4591
rect -1326 -4625 -1288 -4608
rect -6234 -4649 -6158 -4633
rect -6234 -4666 -6218 -4649
rect -6256 -4683 -6218 -4666
rect -6174 -4666 -6158 -4649
rect -6056 -4649 -5980 -4633
rect -6056 -4666 -6040 -4649
rect -6174 -4683 -6136 -4666
rect -6256 -4730 -6136 -4683
rect -6078 -4683 -6040 -4666
rect -5996 -4666 -5980 -4649
rect -5878 -4649 -5802 -4633
rect -5878 -4666 -5862 -4649
rect -5996 -4683 -5958 -4666
rect -6078 -4730 -5958 -4683
rect -5900 -4683 -5862 -4666
rect -5818 -4666 -5802 -4649
rect -5700 -4649 -5624 -4633
rect -5700 -4666 -5684 -4649
rect -5818 -4683 -5780 -4666
rect -5900 -4730 -5780 -4683
rect -5722 -4683 -5684 -4666
rect -5640 -4666 -5624 -4649
rect -5522 -4649 -5446 -4633
rect -5522 -4666 -5506 -4649
rect -5640 -4683 -5602 -4666
rect -5722 -4730 -5602 -4683
rect -5544 -4683 -5506 -4666
rect -5462 -4666 -5446 -4649
rect -5344 -4649 -5268 -4633
rect -5344 -4666 -5328 -4649
rect -5462 -4683 -5424 -4666
rect -5544 -4730 -5424 -4683
rect -5366 -4683 -5328 -4666
rect -5284 -4666 -5268 -4649
rect -5166 -4649 -5090 -4633
rect -5166 -4666 -5150 -4649
rect -5284 -4683 -5246 -4666
rect -5366 -4730 -5246 -4683
rect -5188 -4683 -5150 -4666
rect -5106 -4666 -5090 -4649
rect -4988 -4649 -4912 -4633
rect -4988 -4666 -4972 -4649
rect -5106 -4683 -5068 -4666
rect -5188 -4730 -5068 -4683
rect -5010 -4683 -4972 -4666
rect -4928 -4666 -4912 -4649
rect -4810 -4649 -4734 -4633
rect -4810 -4666 -4794 -4649
rect -4928 -4683 -4890 -4666
rect -5010 -4730 -4890 -4683
rect -4832 -4683 -4794 -4666
rect -4750 -4666 -4734 -4649
rect -4632 -4649 -4556 -4633
rect -4632 -4666 -4616 -4649
rect -4750 -4683 -4712 -4666
rect -4832 -4730 -4712 -4683
rect -4654 -4683 -4616 -4666
rect -4572 -4666 -4556 -4649
rect -4454 -4649 -4378 -4633
rect -4454 -4666 -4438 -4649
rect -4572 -4683 -4534 -4666
rect -4654 -4730 -4534 -4683
rect -4476 -4683 -4438 -4666
rect -4394 -4666 -4378 -4649
rect -4276 -4649 -4200 -4633
rect -4276 -4666 -4260 -4649
rect -4394 -4683 -4356 -4666
rect -4476 -4730 -4356 -4683
rect -4298 -4683 -4260 -4666
rect -4216 -4666 -4200 -4649
rect -4098 -4649 -4022 -4633
rect -4098 -4666 -4082 -4649
rect -4216 -4683 -4178 -4666
rect -4298 -4730 -4178 -4683
rect -4120 -4683 -4082 -4666
rect -4038 -4666 -4022 -4649
rect -3920 -4649 -3844 -4633
rect -3920 -4666 -3904 -4649
rect -4038 -4683 -4000 -4666
rect -4120 -4730 -4000 -4683
rect -3942 -4683 -3904 -4666
rect -3860 -4666 -3844 -4649
rect -3742 -4649 -3666 -4633
rect -3742 -4666 -3726 -4649
rect -3860 -4683 -3822 -4666
rect -3942 -4730 -3822 -4683
rect -3764 -4683 -3726 -4666
rect -3682 -4666 -3666 -4649
rect -3564 -4649 -3488 -4633
rect -3564 -4666 -3548 -4649
rect -3682 -4683 -3644 -4666
rect -3764 -4730 -3644 -4683
rect -3586 -4683 -3548 -4666
rect -3504 -4666 -3488 -4649
rect -3504 -4683 -3466 -4666
rect -1408 -4672 -1288 -4625
rect -1230 -4625 -1192 -4608
rect -1148 -4608 -1132 -4591
rect -1030 -4591 -954 -4575
rect -1030 -4608 -1014 -4591
rect -1148 -4625 -1110 -4608
rect -1230 -4672 -1110 -4625
rect -1052 -4625 -1014 -4608
rect -970 -4608 -954 -4591
rect -852 -4591 -776 -4575
rect -852 -4608 -836 -4591
rect -970 -4625 -932 -4608
rect -1052 -4672 -932 -4625
rect -874 -4625 -836 -4608
rect -792 -4608 -776 -4591
rect -674 -4591 -598 -4575
rect -674 -4608 -658 -4591
rect -792 -4625 -754 -4608
rect -874 -4672 -754 -4625
rect -696 -4625 -658 -4608
rect -614 -4608 -598 -4591
rect -496 -4591 -420 -4575
rect -496 -4608 -480 -4591
rect -614 -4625 -576 -4608
rect -696 -4672 -576 -4625
rect -518 -4625 -480 -4608
rect -436 -4608 -420 -4591
rect -318 -4591 -242 -4575
rect -318 -4608 -302 -4591
rect -436 -4625 -398 -4608
rect -518 -4672 -398 -4625
rect -340 -4625 -302 -4608
rect -258 -4608 -242 -4591
rect -140 -4591 -64 -4575
rect -140 -4608 -124 -4591
rect -258 -4625 -220 -4608
rect -340 -4672 -220 -4625
rect -162 -4625 -124 -4608
rect -80 -4608 -64 -4591
rect 38 -4591 114 -4575
rect 38 -4608 54 -4591
rect -80 -4625 -42 -4608
rect -162 -4672 -42 -4625
rect 16 -4625 54 -4608
rect 98 -4608 114 -4591
rect 216 -4591 292 -4575
rect 216 -4608 232 -4591
rect 98 -4625 136 -4608
rect 16 -4672 136 -4625
rect 194 -4625 232 -4608
rect 276 -4608 292 -4591
rect 394 -4591 470 -4575
rect 394 -4608 410 -4591
rect 276 -4625 314 -4608
rect 194 -4672 314 -4625
rect 372 -4625 410 -4608
rect 454 -4608 470 -4591
rect 572 -4591 648 -4575
rect 572 -4608 588 -4591
rect 454 -4625 492 -4608
rect 372 -4672 492 -4625
rect 550 -4625 588 -4608
rect 632 -4608 648 -4591
rect 750 -4591 826 -4575
rect 750 -4608 766 -4591
rect 632 -4625 670 -4608
rect 550 -4672 670 -4625
rect 728 -4625 766 -4608
rect 810 -4608 826 -4591
rect 928 -4591 1004 -4575
rect 928 -4608 944 -4591
rect 810 -4625 848 -4608
rect 728 -4672 848 -4625
rect 906 -4625 944 -4608
rect 988 -4608 1004 -4591
rect 1106 -4591 1182 -4575
rect 1106 -4608 1122 -4591
rect 988 -4625 1026 -4608
rect 906 -4672 1026 -4625
rect 1084 -4625 1122 -4608
rect 1166 -4608 1182 -4591
rect 1284 -4591 1360 -4575
rect 1284 -4608 1300 -4591
rect 1166 -4625 1204 -4608
rect 1084 -4672 1204 -4625
rect 1262 -4625 1300 -4608
rect 1344 -4608 1360 -4591
rect 1462 -4591 1538 -4575
rect 1462 -4608 1478 -4591
rect 1344 -4625 1382 -4608
rect 1262 -4672 1382 -4625
rect 1440 -4625 1478 -4608
rect 1522 -4608 1538 -4591
rect 1640 -4591 1716 -4575
rect 1640 -4608 1656 -4591
rect 1522 -4625 1560 -4608
rect 1440 -4672 1560 -4625
rect 1618 -4625 1656 -4608
rect 1700 -4608 1716 -4591
rect 1818 -4591 1894 -4575
rect 1818 -4608 1834 -4591
rect 1700 -4625 1738 -4608
rect 1618 -4672 1738 -4625
rect 1796 -4625 1834 -4608
rect 1878 -4608 1894 -4591
rect 1996 -4591 2072 -4575
rect 1996 -4608 2012 -4591
rect 1878 -4625 1916 -4608
rect 1796 -4672 1916 -4625
rect 1974 -4625 2012 -4608
rect 2056 -4608 2072 -4591
rect 2174 -4591 2250 -4575
rect 2174 -4608 2190 -4591
rect 2056 -4625 2094 -4608
rect 1974 -4672 2094 -4625
rect 2152 -4625 2190 -4608
rect 2234 -4608 2250 -4591
rect 2352 -4591 2428 -4575
rect 2352 -4608 2368 -4591
rect 2234 -4625 2272 -4608
rect 2152 -4672 2272 -4625
rect 2330 -4625 2368 -4608
rect 2412 -4608 2428 -4591
rect 2530 -4591 2606 -4575
rect 2530 -4608 2546 -4591
rect 2412 -4625 2450 -4608
rect 2330 -4672 2450 -4625
rect 2508 -4625 2546 -4608
rect 2590 -4608 2606 -4591
rect 2590 -4625 2628 -4608
rect 2508 -4672 2628 -4625
rect -3586 -4730 -3466 -4683
rect -1408 -4999 -1288 -4952
rect -6256 -5057 -6136 -5010
rect -6256 -5074 -6218 -5057
rect -6234 -5091 -6218 -5074
rect -6174 -5074 -6136 -5057
rect -6078 -5057 -5958 -5010
rect -6078 -5074 -6040 -5057
rect -6174 -5091 -6158 -5074
rect -6234 -5107 -6158 -5091
rect -6056 -5091 -6040 -5074
rect -5996 -5074 -5958 -5057
rect -5900 -5057 -5780 -5010
rect -5900 -5074 -5862 -5057
rect -5996 -5091 -5980 -5074
rect -6056 -5107 -5980 -5091
rect -5878 -5091 -5862 -5074
rect -5818 -5074 -5780 -5057
rect -5722 -5057 -5602 -5010
rect -5722 -5074 -5684 -5057
rect -5818 -5091 -5802 -5074
rect -5878 -5107 -5802 -5091
rect -5700 -5091 -5684 -5074
rect -5640 -5074 -5602 -5057
rect -5544 -5057 -5424 -5010
rect -5544 -5074 -5506 -5057
rect -5640 -5091 -5624 -5074
rect -5700 -5107 -5624 -5091
rect -5522 -5091 -5506 -5074
rect -5462 -5074 -5424 -5057
rect -5366 -5057 -5246 -5010
rect -5366 -5074 -5328 -5057
rect -5462 -5091 -5446 -5074
rect -5522 -5107 -5446 -5091
rect -5344 -5091 -5328 -5074
rect -5284 -5074 -5246 -5057
rect -5188 -5057 -5068 -5010
rect -5188 -5074 -5150 -5057
rect -5284 -5091 -5268 -5074
rect -5344 -5107 -5268 -5091
rect -5166 -5091 -5150 -5074
rect -5106 -5074 -5068 -5057
rect -5010 -5057 -4890 -5010
rect -5010 -5074 -4972 -5057
rect -5106 -5091 -5090 -5074
rect -5166 -5107 -5090 -5091
rect -4988 -5091 -4972 -5074
rect -4928 -5074 -4890 -5057
rect -4832 -5057 -4712 -5010
rect -4832 -5074 -4794 -5057
rect -4928 -5091 -4912 -5074
rect -4988 -5107 -4912 -5091
rect -4810 -5091 -4794 -5074
rect -4750 -5074 -4712 -5057
rect -4654 -5057 -4534 -5010
rect -4654 -5074 -4616 -5057
rect -4750 -5091 -4734 -5074
rect -4810 -5107 -4734 -5091
rect -4632 -5091 -4616 -5074
rect -4572 -5074 -4534 -5057
rect -4476 -5057 -4356 -5010
rect -4476 -5074 -4438 -5057
rect -4572 -5091 -4556 -5074
rect -4632 -5107 -4556 -5091
rect -4454 -5091 -4438 -5074
rect -4394 -5074 -4356 -5057
rect -4298 -5057 -4178 -5010
rect -4298 -5074 -4260 -5057
rect -4394 -5091 -4378 -5074
rect -4454 -5107 -4378 -5091
rect -4276 -5091 -4260 -5074
rect -4216 -5074 -4178 -5057
rect -4120 -5057 -4000 -5010
rect -4120 -5074 -4082 -5057
rect -4216 -5091 -4200 -5074
rect -4276 -5107 -4200 -5091
rect -4098 -5091 -4082 -5074
rect -4038 -5074 -4000 -5057
rect -3942 -5057 -3822 -5010
rect -3942 -5074 -3904 -5057
rect -4038 -5091 -4022 -5074
rect -4098 -5107 -4022 -5091
rect -3920 -5091 -3904 -5074
rect -3860 -5074 -3822 -5057
rect -3764 -5057 -3644 -5010
rect -3764 -5074 -3726 -5057
rect -3860 -5091 -3844 -5074
rect -3920 -5107 -3844 -5091
rect -3742 -5091 -3726 -5074
rect -3682 -5074 -3644 -5057
rect -3586 -5057 -3466 -5010
rect -1408 -5016 -1370 -4999
rect -1386 -5033 -1370 -5016
rect -1326 -5016 -1288 -4999
rect -1230 -4999 -1110 -4952
rect -1230 -5016 -1192 -4999
rect -1326 -5033 -1310 -5016
rect -1386 -5049 -1310 -5033
rect -1208 -5033 -1192 -5016
rect -1148 -5016 -1110 -4999
rect -1052 -4999 -932 -4952
rect -1052 -5016 -1014 -4999
rect -1148 -5033 -1132 -5016
rect -1208 -5049 -1132 -5033
rect -1030 -5033 -1014 -5016
rect -970 -5016 -932 -4999
rect -874 -4999 -754 -4952
rect -874 -5016 -836 -4999
rect -970 -5033 -954 -5016
rect -1030 -5049 -954 -5033
rect -852 -5033 -836 -5016
rect -792 -5016 -754 -4999
rect -696 -4999 -576 -4952
rect -696 -5016 -658 -4999
rect -792 -5033 -776 -5016
rect -852 -5049 -776 -5033
rect -674 -5033 -658 -5016
rect -614 -5016 -576 -4999
rect -518 -4999 -398 -4952
rect -518 -5016 -480 -4999
rect -614 -5033 -598 -5016
rect -674 -5049 -598 -5033
rect -496 -5033 -480 -5016
rect -436 -5016 -398 -4999
rect -340 -4999 -220 -4952
rect -340 -5016 -302 -4999
rect -436 -5033 -420 -5016
rect -496 -5049 -420 -5033
rect -318 -5033 -302 -5016
rect -258 -5016 -220 -4999
rect -162 -4999 -42 -4952
rect -162 -5016 -124 -4999
rect -258 -5033 -242 -5016
rect -318 -5049 -242 -5033
rect -140 -5033 -124 -5016
rect -80 -5016 -42 -4999
rect 16 -4999 136 -4952
rect 16 -5016 54 -4999
rect -80 -5033 -64 -5016
rect -140 -5049 -64 -5033
rect 38 -5033 54 -5016
rect 98 -5016 136 -4999
rect 194 -4999 314 -4952
rect 194 -5016 232 -4999
rect 98 -5033 114 -5016
rect 38 -5049 114 -5033
rect 216 -5033 232 -5016
rect 276 -5016 314 -4999
rect 372 -4999 492 -4952
rect 372 -5016 410 -4999
rect 276 -5033 292 -5016
rect 216 -5049 292 -5033
rect 394 -5033 410 -5016
rect 454 -5016 492 -4999
rect 550 -4999 670 -4952
rect 550 -5016 588 -4999
rect 454 -5033 470 -5016
rect 394 -5049 470 -5033
rect 572 -5033 588 -5016
rect 632 -5016 670 -4999
rect 728 -4999 848 -4952
rect 728 -5016 766 -4999
rect 632 -5033 648 -5016
rect 572 -5049 648 -5033
rect 750 -5033 766 -5016
rect 810 -5016 848 -4999
rect 906 -4999 1026 -4952
rect 906 -5016 944 -4999
rect 810 -5033 826 -5016
rect 750 -5049 826 -5033
rect 928 -5033 944 -5016
rect 988 -5016 1026 -4999
rect 1084 -4999 1204 -4952
rect 1084 -5016 1122 -4999
rect 988 -5033 1004 -5016
rect 928 -5049 1004 -5033
rect 1106 -5033 1122 -5016
rect 1166 -5016 1204 -4999
rect 1262 -4999 1382 -4952
rect 1262 -5016 1300 -4999
rect 1166 -5033 1182 -5016
rect 1106 -5049 1182 -5033
rect 1284 -5033 1300 -5016
rect 1344 -5016 1382 -4999
rect 1440 -4999 1560 -4952
rect 1440 -5016 1478 -4999
rect 1344 -5033 1360 -5016
rect 1284 -5049 1360 -5033
rect 1462 -5033 1478 -5016
rect 1522 -5016 1560 -4999
rect 1618 -4999 1738 -4952
rect 1618 -5016 1656 -4999
rect 1522 -5033 1538 -5016
rect 1462 -5049 1538 -5033
rect 1640 -5033 1656 -5016
rect 1700 -5016 1738 -4999
rect 1796 -4999 1916 -4952
rect 1796 -5016 1834 -4999
rect 1700 -5033 1716 -5016
rect 1640 -5049 1716 -5033
rect 1818 -5033 1834 -5016
rect 1878 -5016 1916 -4999
rect 1974 -4999 2094 -4952
rect 1974 -5016 2012 -4999
rect 1878 -5033 1894 -5016
rect 1818 -5049 1894 -5033
rect 1996 -5033 2012 -5016
rect 2056 -5016 2094 -4999
rect 2152 -4999 2272 -4952
rect 2152 -5016 2190 -4999
rect 2056 -5033 2072 -5016
rect 1996 -5049 2072 -5033
rect 2174 -5033 2190 -5016
rect 2234 -5016 2272 -4999
rect 2330 -4999 2450 -4952
rect 2330 -5016 2368 -4999
rect 2234 -5033 2250 -5016
rect 2174 -5049 2250 -5033
rect 2352 -5033 2368 -5016
rect 2412 -5016 2450 -4999
rect 2508 -4999 2628 -4952
rect 2508 -5016 2546 -4999
rect 2412 -5033 2428 -5016
rect 2352 -5049 2428 -5033
rect 2530 -5033 2546 -5016
rect 2590 -5016 2628 -4999
rect 2590 -5033 2606 -5016
rect 2530 -5049 2606 -5033
rect -3586 -5074 -3548 -5057
rect -3682 -5091 -3666 -5074
rect -3742 -5107 -3666 -5091
rect -3564 -5091 -3548 -5074
rect -3504 -5074 -3466 -5057
rect -3504 -5091 -3488 -5074
rect -3564 -5107 -3488 -5091
rect -1386 -5491 -1310 -5475
rect -6234 -5519 -6158 -5503
rect -6234 -5536 -6218 -5519
rect -6256 -5553 -6218 -5536
rect -6174 -5536 -6158 -5519
rect -6056 -5519 -5980 -5503
rect -6056 -5536 -6040 -5519
rect -6174 -5553 -6136 -5536
rect -6256 -5600 -6136 -5553
rect -6078 -5553 -6040 -5536
rect -5996 -5536 -5980 -5519
rect -5878 -5519 -5802 -5503
rect -5878 -5536 -5862 -5519
rect -5996 -5553 -5958 -5536
rect -6078 -5600 -5958 -5553
rect -5900 -5553 -5862 -5536
rect -5818 -5536 -5802 -5519
rect -5700 -5519 -5624 -5503
rect -5700 -5536 -5684 -5519
rect -5818 -5553 -5780 -5536
rect -5900 -5600 -5780 -5553
rect -5722 -5553 -5684 -5536
rect -5640 -5536 -5624 -5519
rect -5522 -5519 -5446 -5503
rect -5522 -5536 -5506 -5519
rect -5640 -5553 -5602 -5536
rect -5722 -5600 -5602 -5553
rect -5544 -5553 -5506 -5536
rect -5462 -5536 -5446 -5519
rect -5344 -5519 -5268 -5503
rect -5344 -5536 -5328 -5519
rect -5462 -5553 -5424 -5536
rect -5544 -5600 -5424 -5553
rect -5366 -5553 -5328 -5536
rect -5284 -5536 -5268 -5519
rect -5166 -5519 -5090 -5503
rect -5166 -5536 -5150 -5519
rect -5284 -5553 -5246 -5536
rect -5366 -5600 -5246 -5553
rect -5188 -5553 -5150 -5536
rect -5106 -5536 -5090 -5519
rect -4988 -5519 -4912 -5503
rect -4988 -5536 -4972 -5519
rect -5106 -5553 -5068 -5536
rect -5188 -5600 -5068 -5553
rect -5010 -5553 -4972 -5536
rect -4928 -5536 -4912 -5519
rect -4810 -5519 -4734 -5503
rect -4810 -5536 -4794 -5519
rect -4928 -5553 -4890 -5536
rect -5010 -5600 -4890 -5553
rect -4832 -5553 -4794 -5536
rect -4750 -5536 -4734 -5519
rect -4632 -5519 -4556 -5503
rect -4632 -5536 -4616 -5519
rect -4750 -5553 -4712 -5536
rect -4832 -5600 -4712 -5553
rect -4654 -5553 -4616 -5536
rect -4572 -5536 -4556 -5519
rect -4454 -5519 -4378 -5503
rect -4454 -5536 -4438 -5519
rect -4572 -5553 -4534 -5536
rect -4654 -5600 -4534 -5553
rect -4476 -5553 -4438 -5536
rect -4394 -5536 -4378 -5519
rect -4276 -5519 -4200 -5503
rect -4276 -5536 -4260 -5519
rect -4394 -5553 -4356 -5536
rect -4476 -5600 -4356 -5553
rect -4298 -5553 -4260 -5536
rect -4216 -5536 -4200 -5519
rect -4098 -5519 -4022 -5503
rect -4098 -5536 -4082 -5519
rect -4216 -5553 -4178 -5536
rect -4298 -5600 -4178 -5553
rect -4120 -5553 -4082 -5536
rect -4038 -5536 -4022 -5519
rect -3920 -5519 -3844 -5503
rect -3920 -5536 -3904 -5519
rect -4038 -5553 -4000 -5536
rect -4120 -5600 -4000 -5553
rect -3942 -5553 -3904 -5536
rect -3860 -5536 -3844 -5519
rect -3742 -5519 -3666 -5503
rect -3742 -5536 -3726 -5519
rect -3860 -5553 -3822 -5536
rect -3942 -5600 -3822 -5553
rect -3764 -5553 -3726 -5536
rect -3682 -5536 -3666 -5519
rect -3564 -5519 -3488 -5503
rect -1386 -5508 -1370 -5491
rect -3564 -5536 -3548 -5519
rect -3682 -5553 -3644 -5536
rect -3764 -5600 -3644 -5553
rect -3586 -5553 -3548 -5536
rect -3504 -5536 -3488 -5519
rect -1408 -5525 -1370 -5508
rect -1326 -5508 -1310 -5491
rect -1208 -5491 -1132 -5475
rect -1208 -5508 -1192 -5491
rect -1326 -5525 -1288 -5508
rect -3504 -5553 -3466 -5536
rect -3586 -5600 -3466 -5553
rect -1408 -5572 -1288 -5525
rect -1230 -5525 -1192 -5508
rect -1148 -5508 -1132 -5491
rect -1030 -5491 -954 -5475
rect -1030 -5508 -1014 -5491
rect -1148 -5525 -1110 -5508
rect -1230 -5572 -1110 -5525
rect -1052 -5525 -1014 -5508
rect -970 -5508 -954 -5491
rect -852 -5491 -776 -5475
rect -852 -5508 -836 -5491
rect -970 -5525 -932 -5508
rect -1052 -5572 -932 -5525
rect -874 -5525 -836 -5508
rect -792 -5508 -776 -5491
rect -674 -5491 -598 -5475
rect -674 -5508 -658 -5491
rect -792 -5525 -754 -5508
rect -874 -5572 -754 -5525
rect -696 -5525 -658 -5508
rect -614 -5508 -598 -5491
rect -496 -5491 -420 -5475
rect -496 -5508 -480 -5491
rect -614 -5525 -576 -5508
rect -696 -5572 -576 -5525
rect -518 -5525 -480 -5508
rect -436 -5508 -420 -5491
rect -318 -5491 -242 -5475
rect -318 -5508 -302 -5491
rect -436 -5525 -398 -5508
rect -518 -5572 -398 -5525
rect -340 -5525 -302 -5508
rect -258 -5508 -242 -5491
rect -140 -5491 -64 -5475
rect -140 -5508 -124 -5491
rect -258 -5525 -220 -5508
rect -340 -5572 -220 -5525
rect -162 -5525 -124 -5508
rect -80 -5508 -64 -5491
rect 38 -5491 114 -5475
rect 38 -5508 54 -5491
rect -80 -5525 -42 -5508
rect -162 -5572 -42 -5525
rect 16 -5525 54 -5508
rect 98 -5508 114 -5491
rect 216 -5491 292 -5475
rect 216 -5508 232 -5491
rect 98 -5525 136 -5508
rect 16 -5572 136 -5525
rect 194 -5525 232 -5508
rect 276 -5508 292 -5491
rect 394 -5491 470 -5475
rect 394 -5508 410 -5491
rect 276 -5525 314 -5508
rect 194 -5572 314 -5525
rect 372 -5525 410 -5508
rect 454 -5508 470 -5491
rect 572 -5491 648 -5475
rect 572 -5508 588 -5491
rect 454 -5525 492 -5508
rect 372 -5572 492 -5525
rect 550 -5525 588 -5508
rect 632 -5508 648 -5491
rect 750 -5491 826 -5475
rect 750 -5508 766 -5491
rect 632 -5525 670 -5508
rect 550 -5572 670 -5525
rect 728 -5525 766 -5508
rect 810 -5508 826 -5491
rect 928 -5491 1004 -5475
rect 928 -5508 944 -5491
rect 810 -5525 848 -5508
rect 728 -5572 848 -5525
rect 906 -5525 944 -5508
rect 988 -5508 1004 -5491
rect 1106 -5491 1182 -5475
rect 1106 -5508 1122 -5491
rect 988 -5525 1026 -5508
rect 906 -5572 1026 -5525
rect 1084 -5525 1122 -5508
rect 1166 -5508 1182 -5491
rect 1284 -5491 1360 -5475
rect 1284 -5508 1300 -5491
rect 1166 -5525 1204 -5508
rect 1084 -5572 1204 -5525
rect 1262 -5525 1300 -5508
rect 1344 -5508 1360 -5491
rect 1462 -5491 1538 -5475
rect 1462 -5508 1478 -5491
rect 1344 -5525 1382 -5508
rect 1262 -5572 1382 -5525
rect 1440 -5525 1478 -5508
rect 1522 -5508 1538 -5491
rect 1640 -5491 1716 -5475
rect 1640 -5508 1656 -5491
rect 1522 -5525 1560 -5508
rect 1440 -5572 1560 -5525
rect 1618 -5525 1656 -5508
rect 1700 -5508 1716 -5491
rect 1818 -5491 1894 -5475
rect 1818 -5508 1834 -5491
rect 1700 -5525 1738 -5508
rect 1618 -5572 1738 -5525
rect 1796 -5525 1834 -5508
rect 1878 -5508 1894 -5491
rect 1996 -5491 2072 -5475
rect 1996 -5508 2012 -5491
rect 1878 -5525 1916 -5508
rect 1796 -5572 1916 -5525
rect 1974 -5525 2012 -5508
rect 2056 -5508 2072 -5491
rect 2174 -5491 2250 -5475
rect 2174 -5508 2190 -5491
rect 2056 -5525 2094 -5508
rect 1974 -5572 2094 -5525
rect 2152 -5525 2190 -5508
rect 2234 -5508 2250 -5491
rect 2352 -5491 2428 -5475
rect 2352 -5508 2368 -5491
rect 2234 -5525 2272 -5508
rect 2152 -5572 2272 -5525
rect 2330 -5525 2368 -5508
rect 2412 -5508 2428 -5491
rect 2530 -5491 2606 -5475
rect 2530 -5508 2546 -5491
rect 2412 -5525 2450 -5508
rect 2330 -5572 2450 -5525
rect 2508 -5525 2546 -5508
rect 2590 -5508 2606 -5491
rect 2590 -5525 2628 -5508
rect 2508 -5572 2628 -5525
rect -6256 -5927 -6136 -5880
rect -6256 -5944 -6218 -5927
rect -6234 -5961 -6218 -5944
rect -6174 -5944 -6136 -5927
rect -6078 -5927 -5958 -5880
rect -6078 -5944 -6040 -5927
rect -6174 -5961 -6158 -5944
rect -6234 -5977 -6158 -5961
rect -6056 -5961 -6040 -5944
rect -5996 -5944 -5958 -5927
rect -5900 -5927 -5780 -5880
rect -5900 -5944 -5862 -5927
rect -5996 -5961 -5980 -5944
rect -6056 -5977 -5980 -5961
rect -5878 -5961 -5862 -5944
rect -5818 -5944 -5780 -5927
rect -5722 -5927 -5602 -5880
rect -5722 -5944 -5684 -5927
rect -5818 -5961 -5802 -5944
rect -5878 -5977 -5802 -5961
rect -5700 -5961 -5684 -5944
rect -5640 -5944 -5602 -5927
rect -5544 -5927 -5424 -5880
rect -5544 -5944 -5506 -5927
rect -5640 -5961 -5624 -5944
rect -5700 -5977 -5624 -5961
rect -5522 -5961 -5506 -5944
rect -5462 -5944 -5424 -5927
rect -5366 -5927 -5246 -5880
rect -5366 -5944 -5328 -5927
rect -5462 -5961 -5446 -5944
rect -5522 -5977 -5446 -5961
rect -5344 -5961 -5328 -5944
rect -5284 -5944 -5246 -5927
rect -5188 -5927 -5068 -5880
rect -5188 -5944 -5150 -5927
rect -5284 -5961 -5268 -5944
rect -5344 -5977 -5268 -5961
rect -5166 -5961 -5150 -5944
rect -5106 -5944 -5068 -5927
rect -5010 -5927 -4890 -5880
rect -5010 -5944 -4972 -5927
rect -5106 -5961 -5090 -5944
rect -5166 -5977 -5090 -5961
rect -4988 -5961 -4972 -5944
rect -4928 -5944 -4890 -5927
rect -4832 -5927 -4712 -5880
rect -4832 -5944 -4794 -5927
rect -4928 -5961 -4912 -5944
rect -4988 -5977 -4912 -5961
rect -4810 -5961 -4794 -5944
rect -4750 -5944 -4712 -5927
rect -4654 -5927 -4534 -5880
rect -4654 -5944 -4616 -5927
rect -4750 -5961 -4734 -5944
rect -4810 -5977 -4734 -5961
rect -4632 -5961 -4616 -5944
rect -4572 -5944 -4534 -5927
rect -4476 -5927 -4356 -5880
rect -4476 -5944 -4438 -5927
rect -4572 -5961 -4556 -5944
rect -4632 -5977 -4556 -5961
rect -4454 -5961 -4438 -5944
rect -4394 -5944 -4356 -5927
rect -4298 -5927 -4178 -5880
rect -4298 -5944 -4260 -5927
rect -4394 -5961 -4378 -5944
rect -4454 -5977 -4378 -5961
rect -4276 -5961 -4260 -5944
rect -4216 -5944 -4178 -5927
rect -4120 -5927 -4000 -5880
rect -4120 -5944 -4082 -5927
rect -4216 -5961 -4200 -5944
rect -4276 -5977 -4200 -5961
rect -4098 -5961 -4082 -5944
rect -4038 -5944 -4000 -5927
rect -3942 -5927 -3822 -5880
rect -3942 -5944 -3904 -5927
rect -4038 -5961 -4022 -5944
rect -4098 -5977 -4022 -5961
rect -3920 -5961 -3904 -5944
rect -3860 -5944 -3822 -5927
rect -3764 -5927 -3644 -5880
rect -3764 -5944 -3726 -5927
rect -3860 -5961 -3844 -5944
rect -3920 -5977 -3844 -5961
rect -3742 -5961 -3726 -5944
rect -3682 -5944 -3644 -5927
rect -3586 -5927 -3466 -5880
rect -1408 -5899 -1288 -5852
rect -1408 -5916 -1370 -5899
rect -3586 -5944 -3548 -5927
rect -3682 -5961 -3666 -5944
rect -3742 -5977 -3666 -5961
rect -3564 -5961 -3548 -5944
rect -3504 -5944 -3466 -5927
rect -1386 -5933 -1370 -5916
rect -1326 -5916 -1288 -5899
rect -1230 -5899 -1110 -5852
rect -1230 -5916 -1192 -5899
rect -1326 -5933 -1310 -5916
rect -3504 -5961 -3488 -5944
rect -1386 -5949 -1310 -5933
rect -1208 -5933 -1192 -5916
rect -1148 -5916 -1110 -5899
rect -1052 -5899 -932 -5852
rect -1052 -5916 -1014 -5899
rect -1148 -5933 -1132 -5916
rect -1208 -5949 -1132 -5933
rect -1030 -5933 -1014 -5916
rect -970 -5916 -932 -5899
rect -874 -5899 -754 -5852
rect -874 -5916 -836 -5899
rect -970 -5933 -954 -5916
rect -1030 -5949 -954 -5933
rect -852 -5933 -836 -5916
rect -792 -5916 -754 -5899
rect -696 -5899 -576 -5852
rect -696 -5916 -658 -5899
rect -792 -5933 -776 -5916
rect -852 -5949 -776 -5933
rect -674 -5933 -658 -5916
rect -614 -5916 -576 -5899
rect -518 -5899 -398 -5852
rect -518 -5916 -480 -5899
rect -614 -5933 -598 -5916
rect -674 -5949 -598 -5933
rect -496 -5933 -480 -5916
rect -436 -5916 -398 -5899
rect -340 -5899 -220 -5852
rect -340 -5916 -302 -5899
rect -436 -5933 -420 -5916
rect -496 -5949 -420 -5933
rect -318 -5933 -302 -5916
rect -258 -5916 -220 -5899
rect -162 -5899 -42 -5852
rect -162 -5916 -124 -5899
rect -258 -5933 -242 -5916
rect -318 -5949 -242 -5933
rect -140 -5933 -124 -5916
rect -80 -5916 -42 -5899
rect 16 -5899 136 -5852
rect 16 -5916 54 -5899
rect -80 -5933 -64 -5916
rect -140 -5949 -64 -5933
rect 38 -5933 54 -5916
rect 98 -5916 136 -5899
rect 194 -5899 314 -5852
rect 194 -5916 232 -5899
rect 98 -5933 114 -5916
rect 38 -5949 114 -5933
rect 216 -5933 232 -5916
rect 276 -5916 314 -5899
rect 372 -5899 492 -5852
rect 372 -5916 410 -5899
rect 276 -5933 292 -5916
rect 216 -5949 292 -5933
rect 394 -5933 410 -5916
rect 454 -5916 492 -5899
rect 550 -5899 670 -5852
rect 550 -5916 588 -5899
rect 454 -5933 470 -5916
rect 394 -5949 470 -5933
rect 572 -5933 588 -5916
rect 632 -5916 670 -5899
rect 728 -5899 848 -5852
rect 728 -5916 766 -5899
rect 632 -5933 648 -5916
rect 572 -5949 648 -5933
rect 750 -5933 766 -5916
rect 810 -5916 848 -5899
rect 906 -5899 1026 -5852
rect 906 -5916 944 -5899
rect 810 -5933 826 -5916
rect 750 -5949 826 -5933
rect 928 -5933 944 -5916
rect 988 -5916 1026 -5899
rect 1084 -5899 1204 -5852
rect 1084 -5916 1122 -5899
rect 988 -5933 1004 -5916
rect 928 -5949 1004 -5933
rect 1106 -5933 1122 -5916
rect 1166 -5916 1204 -5899
rect 1262 -5899 1382 -5852
rect 1262 -5916 1300 -5899
rect 1166 -5933 1182 -5916
rect 1106 -5949 1182 -5933
rect 1284 -5933 1300 -5916
rect 1344 -5916 1382 -5899
rect 1440 -5899 1560 -5852
rect 1440 -5916 1478 -5899
rect 1344 -5933 1360 -5916
rect 1284 -5949 1360 -5933
rect 1462 -5933 1478 -5916
rect 1522 -5916 1560 -5899
rect 1618 -5899 1738 -5852
rect 1618 -5916 1656 -5899
rect 1522 -5933 1538 -5916
rect 1462 -5949 1538 -5933
rect 1640 -5933 1656 -5916
rect 1700 -5916 1738 -5899
rect 1796 -5899 1916 -5852
rect 1796 -5916 1834 -5899
rect 1700 -5933 1716 -5916
rect 1640 -5949 1716 -5933
rect 1818 -5933 1834 -5916
rect 1878 -5916 1916 -5899
rect 1974 -5899 2094 -5852
rect 1974 -5916 2012 -5899
rect 1878 -5933 1894 -5916
rect 1818 -5949 1894 -5933
rect 1996 -5933 2012 -5916
rect 2056 -5916 2094 -5899
rect 2152 -5899 2272 -5852
rect 2152 -5916 2190 -5899
rect 2056 -5933 2072 -5916
rect 1996 -5949 2072 -5933
rect 2174 -5933 2190 -5916
rect 2234 -5916 2272 -5899
rect 2330 -5899 2450 -5852
rect 2330 -5916 2368 -5899
rect 2234 -5933 2250 -5916
rect 2174 -5949 2250 -5933
rect 2352 -5933 2368 -5916
rect 2412 -5916 2450 -5899
rect 2508 -5899 2628 -5852
rect 2508 -5916 2546 -5899
rect 2412 -5933 2428 -5916
rect 2352 -5949 2428 -5933
rect 2530 -5933 2546 -5916
rect 2590 -5916 2628 -5899
rect 2590 -5933 2606 -5916
rect 2530 -5949 2606 -5933
rect -3564 -5977 -3488 -5961
rect -5560 -7790 -5484 -7774
rect -5560 -7807 -5544 -7790
rect -5582 -7824 -5544 -7807
rect -5500 -7807 -5484 -7790
rect -5382 -7790 -5306 -7774
rect -5382 -7807 -5366 -7790
rect -5500 -7824 -5462 -7807
rect -5582 -7862 -5462 -7824
rect -5404 -7824 -5366 -7807
rect -5322 -7807 -5306 -7790
rect -5204 -7790 -5128 -7774
rect -5204 -7807 -5188 -7790
rect -5322 -7824 -5284 -7807
rect -5404 -7862 -5284 -7824
rect -5226 -7824 -5188 -7807
rect -5144 -7807 -5128 -7790
rect -5026 -7790 -4950 -7774
rect -5026 -7807 -5010 -7790
rect -5144 -7824 -5106 -7807
rect -5226 -7862 -5106 -7824
rect -5048 -7824 -5010 -7807
rect -4966 -7807 -4950 -7790
rect -4848 -7790 -4772 -7774
rect -4848 -7807 -4832 -7790
rect -4966 -7824 -4928 -7807
rect -5048 -7862 -4928 -7824
rect -4870 -7824 -4832 -7807
rect -4788 -7807 -4772 -7790
rect -4670 -7790 -4594 -7774
rect -4670 -7807 -4654 -7790
rect -4788 -7824 -4750 -7807
rect -4870 -7862 -4750 -7824
rect -4692 -7824 -4654 -7807
rect -4610 -7807 -4594 -7790
rect -4492 -7790 -4416 -7774
rect -4492 -7807 -4476 -7790
rect -4610 -7824 -4572 -7807
rect -4692 -7862 -4572 -7824
rect -4514 -7824 -4476 -7807
rect -4432 -7807 -4416 -7790
rect -4314 -7790 -4238 -7774
rect -4314 -7807 -4298 -7790
rect -4432 -7824 -4394 -7807
rect -4514 -7862 -4394 -7824
rect -4336 -7824 -4298 -7807
rect -4254 -7807 -4238 -7790
rect -4136 -7790 -4060 -7774
rect -4136 -7807 -4120 -7790
rect -4254 -7824 -4216 -7807
rect -4336 -7862 -4216 -7824
rect -4158 -7824 -4120 -7807
rect -4076 -7807 -4060 -7790
rect -4076 -7824 -4038 -7807
rect -4158 -7862 -4038 -7824
rect -2105 -8048 -2029 -8032
rect -2105 -8065 -2089 -8048
rect -2127 -8082 -2089 -8065
rect -2045 -8065 -2029 -8048
rect -1927 -8048 -1851 -8032
rect -1927 -8065 -1911 -8048
rect -2045 -8082 -2007 -8065
rect -2127 -8120 -2007 -8082
rect -1949 -8082 -1911 -8065
rect -1867 -8065 -1851 -8048
rect -1749 -8048 -1673 -8032
rect -1749 -8065 -1733 -8048
rect -1867 -8082 -1829 -8065
rect -1949 -8120 -1829 -8082
rect -1771 -8082 -1733 -8065
rect -1689 -8065 -1673 -8048
rect -1571 -8048 -1495 -8032
rect -1571 -8065 -1555 -8048
rect -1689 -8082 -1651 -8065
rect -1771 -8120 -1651 -8082
rect -1593 -8082 -1555 -8065
rect -1511 -8065 -1495 -8048
rect -1393 -8048 -1317 -8032
rect -1393 -8065 -1377 -8048
rect -1511 -8082 -1473 -8065
rect -1593 -8120 -1473 -8082
rect -1415 -8082 -1377 -8065
rect -1333 -8065 -1317 -8048
rect -1215 -8048 -1139 -8032
rect -1215 -8065 -1199 -8048
rect -1333 -8082 -1295 -8065
rect -1415 -8120 -1295 -8082
rect -1237 -8082 -1199 -8065
rect -1155 -8065 -1139 -8048
rect -1037 -8048 -961 -8032
rect -1037 -8065 -1021 -8048
rect -1155 -8082 -1117 -8065
rect -1237 -8120 -1117 -8082
rect -1059 -8082 -1021 -8065
rect -977 -8065 -961 -8048
rect -859 -8048 -783 -8032
rect -859 -8065 -843 -8048
rect -977 -8082 -939 -8065
rect -1059 -8120 -939 -8082
rect -881 -8082 -843 -8065
rect -799 -8065 -783 -8048
rect -681 -8048 -605 -8032
rect -681 -8065 -665 -8048
rect -799 -8082 -761 -8065
rect -881 -8120 -761 -8082
rect -703 -8082 -665 -8065
rect -621 -8065 -605 -8048
rect -503 -8048 -427 -8032
rect -503 -8065 -487 -8048
rect -621 -8082 -583 -8065
rect -703 -8120 -583 -8082
rect -525 -8082 -487 -8065
rect -443 -8065 -427 -8048
rect -325 -8048 -249 -8032
rect -325 -8065 -309 -8048
rect -443 -8082 -405 -8065
rect -525 -8120 -405 -8082
rect -347 -8082 -309 -8065
rect -265 -8065 -249 -8048
rect -147 -8048 -71 -8032
rect -147 -8065 -131 -8048
rect -265 -8082 -227 -8065
rect -347 -8120 -227 -8082
rect -169 -8082 -131 -8065
rect -87 -8065 -71 -8048
rect 31 -8048 107 -8032
rect 31 -8065 47 -8048
rect -87 -8082 -49 -8065
rect -169 -8120 -49 -8082
rect 9 -8082 47 -8065
rect 91 -8065 107 -8048
rect 209 -8048 285 -8032
rect 209 -8065 225 -8048
rect 91 -8082 129 -8065
rect 9 -8120 129 -8082
rect 187 -8082 225 -8065
rect 269 -8065 285 -8048
rect 387 -8048 463 -8032
rect 387 -8065 403 -8048
rect 269 -8082 307 -8065
rect 187 -8120 307 -8082
rect 365 -8082 403 -8065
rect 447 -8065 463 -8048
rect 565 -8048 641 -8032
rect 565 -8065 581 -8048
rect 447 -8082 485 -8065
rect 365 -8120 485 -8082
rect 543 -8082 581 -8065
rect 625 -8065 641 -8048
rect 743 -8048 819 -8032
rect 743 -8065 759 -8048
rect 625 -8082 663 -8065
rect 543 -8120 663 -8082
rect 721 -8082 759 -8065
rect 803 -8065 819 -8048
rect 921 -8048 997 -8032
rect 921 -8065 937 -8048
rect 803 -8082 841 -8065
rect 721 -8120 841 -8082
rect 899 -8082 937 -8065
rect 981 -8065 997 -8048
rect 1099 -8048 1175 -8032
rect 1099 -8065 1115 -8048
rect 981 -8082 1019 -8065
rect 899 -8120 1019 -8082
rect 1077 -8082 1115 -8065
rect 1159 -8065 1175 -8048
rect 1277 -8048 1353 -8032
rect 1277 -8065 1293 -8048
rect 1159 -8082 1197 -8065
rect 1077 -8120 1197 -8082
rect 1255 -8082 1293 -8065
rect 1337 -8065 1353 -8048
rect 1455 -8048 1531 -8032
rect 1455 -8065 1471 -8048
rect 1337 -8082 1375 -8065
rect 1255 -8120 1375 -8082
rect 1433 -8082 1471 -8065
rect 1515 -8065 1531 -8048
rect 1633 -8048 1709 -8032
rect 1633 -8065 1649 -8048
rect 1515 -8082 1553 -8065
rect 1433 -8120 1553 -8082
rect 1611 -8082 1649 -8065
rect 1693 -8065 1709 -8048
rect 1811 -8048 1887 -8032
rect 1811 -8065 1827 -8048
rect 1693 -8082 1731 -8065
rect 1611 -8120 1731 -8082
rect 1789 -8082 1827 -8065
rect 1871 -8065 1887 -8048
rect 1989 -8048 2065 -8032
rect 1989 -8065 2005 -8048
rect 1871 -8082 1909 -8065
rect 1789 -8120 1909 -8082
rect 1967 -8082 2005 -8065
rect 2049 -8065 2065 -8048
rect 2167 -8048 2243 -8032
rect 2167 -8065 2183 -8048
rect 2049 -8082 2087 -8065
rect 1967 -8120 2087 -8082
rect 2145 -8082 2183 -8065
rect 2227 -8065 2243 -8048
rect 2345 -8048 2421 -8032
rect 2345 -8065 2361 -8048
rect 2227 -8082 2265 -8065
rect 2145 -8120 2265 -8082
rect 2323 -8082 2361 -8065
rect 2405 -8065 2421 -8048
rect 2523 -8048 2599 -8032
rect 2523 -8065 2539 -8048
rect 2405 -8082 2443 -8065
rect 2323 -8120 2443 -8082
rect 2501 -8082 2539 -8065
rect 2583 -8065 2599 -8048
rect 2701 -8048 2777 -8032
rect 2701 -8065 2717 -8048
rect 2583 -8082 2621 -8065
rect 2501 -8120 2621 -8082
rect 2679 -8082 2717 -8065
rect 2761 -8065 2777 -8048
rect 2879 -8048 2955 -8032
rect 2879 -8065 2895 -8048
rect 2761 -8082 2799 -8065
rect 2679 -8120 2799 -8082
rect 2857 -8082 2895 -8065
rect 2939 -8065 2955 -8048
rect 3057 -8048 3133 -8032
rect 3057 -8065 3073 -8048
rect 2939 -8082 2977 -8065
rect 2857 -8120 2977 -8082
rect 3035 -8082 3073 -8065
rect 3117 -8065 3133 -8048
rect 3235 -8048 3311 -8032
rect 3235 -8065 3251 -8048
rect 3117 -8082 3155 -8065
rect 3035 -8120 3155 -8082
rect 3213 -8082 3251 -8065
rect 3295 -8065 3311 -8048
rect 3413 -8048 3489 -8032
rect 3413 -8065 3429 -8048
rect 3295 -8082 3333 -8065
rect 3213 -8120 3333 -8082
rect 3391 -8082 3429 -8065
rect 3473 -8065 3489 -8048
rect 3591 -8048 3667 -8032
rect 3591 -8065 3607 -8048
rect 3473 -8082 3511 -8065
rect 3391 -8120 3511 -8082
rect 3569 -8082 3607 -8065
rect 3651 -8065 3667 -8048
rect 3769 -8048 3845 -8032
rect 3769 -8065 3785 -8048
rect 3651 -8082 3689 -8065
rect 3569 -8120 3689 -8082
rect 3747 -8082 3785 -8065
rect 3829 -8065 3845 -8048
rect 3947 -8048 4023 -8032
rect 3947 -8065 3963 -8048
rect 3829 -8082 3867 -8065
rect 3747 -8120 3867 -8082
rect 3925 -8082 3963 -8065
rect 4007 -8065 4023 -8048
rect 4007 -8082 4045 -8065
rect 3925 -8120 4045 -8082
rect -5582 -8180 -5462 -8142
rect -5582 -8197 -5544 -8180
rect -5560 -8214 -5544 -8197
rect -5500 -8197 -5462 -8180
rect -5404 -8180 -5284 -8142
rect -5404 -8197 -5366 -8180
rect -5500 -8214 -5484 -8197
rect -5560 -8230 -5484 -8214
rect -5382 -8214 -5366 -8197
rect -5322 -8197 -5284 -8180
rect -5226 -8180 -5106 -8142
rect -5226 -8197 -5188 -8180
rect -5322 -8214 -5306 -8197
rect -5382 -8230 -5306 -8214
rect -5204 -8214 -5188 -8197
rect -5144 -8197 -5106 -8180
rect -5048 -8180 -4928 -8142
rect -5048 -8197 -5010 -8180
rect -5144 -8214 -5128 -8197
rect -5204 -8230 -5128 -8214
rect -5026 -8214 -5010 -8197
rect -4966 -8197 -4928 -8180
rect -4870 -8180 -4750 -8142
rect -4870 -8197 -4832 -8180
rect -4966 -8214 -4950 -8197
rect -5026 -8230 -4950 -8214
rect -4848 -8214 -4832 -8197
rect -4788 -8197 -4750 -8180
rect -4692 -8180 -4572 -8142
rect -4692 -8197 -4654 -8180
rect -4788 -8214 -4772 -8197
rect -4848 -8230 -4772 -8214
rect -4670 -8214 -4654 -8197
rect -4610 -8197 -4572 -8180
rect -4514 -8180 -4394 -8142
rect -4514 -8197 -4476 -8180
rect -4610 -8214 -4594 -8197
rect -4670 -8230 -4594 -8214
rect -4492 -8214 -4476 -8197
rect -4432 -8197 -4394 -8180
rect -4336 -8180 -4216 -8142
rect -4336 -8197 -4298 -8180
rect -4432 -8214 -4416 -8197
rect -4492 -8230 -4416 -8214
rect -4314 -8214 -4298 -8197
rect -4254 -8197 -4216 -8180
rect -4158 -8180 -4038 -8142
rect -4158 -8197 -4120 -8180
rect -4254 -8214 -4238 -8197
rect -4314 -8230 -4238 -8214
rect -4136 -8214 -4120 -8197
rect -4076 -8197 -4038 -8180
rect -4076 -8214 -4060 -8197
rect -4136 -8230 -4060 -8214
rect -5560 -8340 -5484 -8324
rect -5560 -8357 -5544 -8340
rect -5582 -8374 -5544 -8357
rect -5500 -8357 -5484 -8340
rect -5382 -8340 -5306 -8324
rect -5382 -8357 -5366 -8340
rect -5500 -8374 -5462 -8357
rect -5582 -8412 -5462 -8374
rect -5404 -8374 -5366 -8357
rect -5322 -8357 -5306 -8340
rect -5204 -8340 -5128 -8324
rect -5204 -8357 -5188 -8340
rect -5322 -8374 -5284 -8357
rect -5404 -8412 -5284 -8374
rect -5226 -8374 -5188 -8357
rect -5144 -8357 -5128 -8340
rect -5026 -8340 -4950 -8324
rect -5026 -8357 -5010 -8340
rect -5144 -8374 -5106 -8357
rect -5226 -8412 -5106 -8374
rect -5048 -8374 -5010 -8357
rect -4966 -8357 -4950 -8340
rect -4848 -8340 -4772 -8324
rect -4848 -8357 -4832 -8340
rect -4966 -8374 -4928 -8357
rect -5048 -8412 -4928 -8374
rect -4870 -8374 -4832 -8357
rect -4788 -8357 -4772 -8340
rect -4670 -8340 -4594 -8324
rect -4670 -8357 -4654 -8340
rect -4788 -8374 -4750 -8357
rect -4870 -8412 -4750 -8374
rect -4692 -8374 -4654 -8357
rect -4610 -8357 -4594 -8340
rect -4492 -8340 -4416 -8324
rect -4492 -8357 -4476 -8340
rect -4610 -8374 -4572 -8357
rect -4692 -8412 -4572 -8374
rect -4514 -8374 -4476 -8357
rect -4432 -8357 -4416 -8340
rect -4314 -8340 -4238 -8324
rect -4314 -8357 -4298 -8340
rect -4432 -8374 -4394 -8357
rect -4514 -8412 -4394 -8374
rect -4336 -8374 -4298 -8357
rect -4254 -8357 -4238 -8340
rect -4136 -8340 -4060 -8324
rect -4136 -8357 -4120 -8340
rect -4254 -8374 -4216 -8357
rect -4336 -8412 -4216 -8374
rect -4158 -8374 -4120 -8357
rect -4076 -8357 -4060 -8340
rect -4076 -8374 -4038 -8357
rect -4158 -8412 -4038 -8374
rect -2127 -8438 -2007 -8400
rect -2127 -8455 -2089 -8438
rect -2105 -8472 -2089 -8455
rect -2045 -8455 -2007 -8438
rect -1949 -8438 -1829 -8400
rect -1949 -8455 -1911 -8438
rect -2045 -8472 -2029 -8455
rect -2105 -8488 -2029 -8472
rect -1927 -8472 -1911 -8455
rect -1867 -8455 -1829 -8438
rect -1771 -8438 -1651 -8400
rect -1771 -8455 -1733 -8438
rect -1867 -8472 -1851 -8455
rect -1927 -8488 -1851 -8472
rect -1749 -8472 -1733 -8455
rect -1689 -8455 -1651 -8438
rect -1593 -8438 -1473 -8400
rect -1593 -8455 -1555 -8438
rect -1689 -8472 -1673 -8455
rect -1749 -8488 -1673 -8472
rect -1571 -8472 -1555 -8455
rect -1511 -8455 -1473 -8438
rect -1415 -8438 -1295 -8400
rect -1415 -8455 -1377 -8438
rect -1511 -8472 -1495 -8455
rect -1571 -8488 -1495 -8472
rect -1393 -8472 -1377 -8455
rect -1333 -8455 -1295 -8438
rect -1237 -8438 -1117 -8400
rect -1237 -8455 -1199 -8438
rect -1333 -8472 -1317 -8455
rect -1393 -8488 -1317 -8472
rect -1215 -8472 -1199 -8455
rect -1155 -8455 -1117 -8438
rect -1059 -8438 -939 -8400
rect -1059 -8455 -1021 -8438
rect -1155 -8472 -1139 -8455
rect -1215 -8488 -1139 -8472
rect -1037 -8472 -1021 -8455
rect -977 -8455 -939 -8438
rect -881 -8438 -761 -8400
rect -881 -8455 -843 -8438
rect -977 -8472 -961 -8455
rect -1037 -8488 -961 -8472
rect -859 -8472 -843 -8455
rect -799 -8455 -761 -8438
rect -703 -8438 -583 -8400
rect -703 -8455 -665 -8438
rect -799 -8472 -783 -8455
rect -859 -8488 -783 -8472
rect -681 -8472 -665 -8455
rect -621 -8455 -583 -8438
rect -525 -8438 -405 -8400
rect -525 -8455 -487 -8438
rect -621 -8472 -605 -8455
rect -681 -8488 -605 -8472
rect -503 -8472 -487 -8455
rect -443 -8455 -405 -8438
rect -347 -8438 -227 -8400
rect -347 -8455 -309 -8438
rect -443 -8472 -427 -8455
rect -503 -8488 -427 -8472
rect -325 -8472 -309 -8455
rect -265 -8455 -227 -8438
rect -169 -8438 -49 -8400
rect -169 -8455 -131 -8438
rect -265 -8472 -249 -8455
rect -325 -8488 -249 -8472
rect -147 -8472 -131 -8455
rect -87 -8455 -49 -8438
rect 9 -8438 129 -8400
rect 9 -8455 47 -8438
rect -87 -8472 -71 -8455
rect -147 -8488 -71 -8472
rect 31 -8472 47 -8455
rect 91 -8455 129 -8438
rect 187 -8438 307 -8400
rect 187 -8455 225 -8438
rect 91 -8472 107 -8455
rect 31 -8488 107 -8472
rect 209 -8472 225 -8455
rect 269 -8455 307 -8438
rect 365 -8438 485 -8400
rect 365 -8455 403 -8438
rect 269 -8472 285 -8455
rect 209 -8488 285 -8472
rect 387 -8472 403 -8455
rect 447 -8455 485 -8438
rect 543 -8438 663 -8400
rect 543 -8455 581 -8438
rect 447 -8472 463 -8455
rect 387 -8488 463 -8472
rect 565 -8472 581 -8455
rect 625 -8455 663 -8438
rect 721 -8438 841 -8400
rect 721 -8455 759 -8438
rect 625 -8472 641 -8455
rect 565 -8488 641 -8472
rect 743 -8472 759 -8455
rect 803 -8455 841 -8438
rect 899 -8438 1019 -8400
rect 899 -8455 937 -8438
rect 803 -8472 819 -8455
rect 743 -8488 819 -8472
rect 921 -8472 937 -8455
rect 981 -8455 1019 -8438
rect 1077 -8438 1197 -8400
rect 1077 -8455 1115 -8438
rect 981 -8472 997 -8455
rect 921 -8488 997 -8472
rect 1099 -8472 1115 -8455
rect 1159 -8455 1197 -8438
rect 1255 -8438 1375 -8400
rect 1255 -8455 1293 -8438
rect 1159 -8472 1175 -8455
rect 1099 -8488 1175 -8472
rect 1277 -8472 1293 -8455
rect 1337 -8455 1375 -8438
rect 1433 -8438 1553 -8400
rect 1433 -8455 1471 -8438
rect 1337 -8472 1353 -8455
rect 1277 -8488 1353 -8472
rect 1455 -8472 1471 -8455
rect 1515 -8455 1553 -8438
rect 1611 -8438 1731 -8400
rect 1611 -8455 1649 -8438
rect 1515 -8472 1531 -8455
rect 1455 -8488 1531 -8472
rect 1633 -8472 1649 -8455
rect 1693 -8455 1731 -8438
rect 1789 -8438 1909 -8400
rect 1789 -8455 1827 -8438
rect 1693 -8472 1709 -8455
rect 1633 -8488 1709 -8472
rect 1811 -8472 1827 -8455
rect 1871 -8455 1909 -8438
rect 1967 -8438 2087 -8400
rect 1967 -8455 2005 -8438
rect 1871 -8472 1887 -8455
rect 1811 -8488 1887 -8472
rect 1989 -8472 2005 -8455
rect 2049 -8455 2087 -8438
rect 2145 -8438 2265 -8400
rect 2145 -8455 2183 -8438
rect 2049 -8472 2065 -8455
rect 1989 -8488 2065 -8472
rect 2167 -8472 2183 -8455
rect 2227 -8455 2265 -8438
rect 2323 -8438 2443 -8400
rect 2323 -8455 2361 -8438
rect 2227 -8472 2243 -8455
rect 2167 -8488 2243 -8472
rect 2345 -8472 2361 -8455
rect 2405 -8455 2443 -8438
rect 2501 -8438 2621 -8400
rect 2501 -8455 2539 -8438
rect 2405 -8472 2421 -8455
rect 2345 -8488 2421 -8472
rect 2523 -8472 2539 -8455
rect 2583 -8455 2621 -8438
rect 2679 -8438 2799 -8400
rect 2679 -8455 2717 -8438
rect 2583 -8472 2599 -8455
rect 2523 -8488 2599 -8472
rect 2701 -8472 2717 -8455
rect 2761 -8455 2799 -8438
rect 2857 -8438 2977 -8400
rect 2857 -8455 2895 -8438
rect 2761 -8472 2777 -8455
rect 2701 -8488 2777 -8472
rect 2879 -8472 2895 -8455
rect 2939 -8455 2977 -8438
rect 3035 -8438 3155 -8400
rect 3035 -8455 3073 -8438
rect 2939 -8472 2955 -8455
rect 2879 -8488 2955 -8472
rect 3057 -8472 3073 -8455
rect 3117 -8455 3155 -8438
rect 3213 -8438 3333 -8400
rect 3213 -8455 3251 -8438
rect 3117 -8472 3133 -8455
rect 3057 -8488 3133 -8472
rect 3235 -8472 3251 -8455
rect 3295 -8455 3333 -8438
rect 3391 -8438 3511 -8400
rect 3391 -8455 3429 -8438
rect 3295 -8472 3311 -8455
rect 3235 -8488 3311 -8472
rect 3413 -8472 3429 -8455
rect 3473 -8455 3511 -8438
rect 3569 -8438 3689 -8400
rect 3569 -8455 3607 -8438
rect 3473 -8472 3489 -8455
rect 3413 -8488 3489 -8472
rect 3591 -8472 3607 -8455
rect 3651 -8455 3689 -8438
rect 3747 -8438 3867 -8400
rect 3747 -8455 3785 -8438
rect 3651 -8472 3667 -8455
rect 3591 -8488 3667 -8472
rect 3769 -8472 3785 -8455
rect 3829 -8455 3867 -8438
rect 3925 -8438 4045 -8400
rect 3925 -8455 3963 -8438
rect 3829 -8472 3845 -8455
rect 3769 -8488 3845 -8472
rect 3947 -8472 3963 -8455
rect 4007 -8455 4045 -8438
rect 4007 -8472 4023 -8455
rect 3947 -8488 4023 -8472
rect -5582 -8730 -5462 -8692
rect -5582 -8747 -5544 -8730
rect -5560 -8764 -5544 -8747
rect -5500 -8747 -5462 -8730
rect -5404 -8730 -5284 -8692
rect -5404 -8747 -5366 -8730
rect -5500 -8764 -5484 -8747
rect -5560 -8780 -5484 -8764
rect -5382 -8764 -5366 -8747
rect -5322 -8747 -5284 -8730
rect -5226 -8730 -5106 -8692
rect -5226 -8747 -5188 -8730
rect -5322 -8764 -5306 -8747
rect -5382 -8780 -5306 -8764
rect -5204 -8764 -5188 -8747
rect -5144 -8747 -5106 -8730
rect -5048 -8730 -4928 -8692
rect -5048 -8747 -5010 -8730
rect -5144 -8764 -5128 -8747
rect -5204 -8780 -5128 -8764
rect -5026 -8764 -5010 -8747
rect -4966 -8747 -4928 -8730
rect -4870 -8730 -4750 -8692
rect -4870 -8747 -4832 -8730
rect -4966 -8764 -4950 -8747
rect -5026 -8780 -4950 -8764
rect -4848 -8764 -4832 -8747
rect -4788 -8747 -4750 -8730
rect -4692 -8730 -4572 -8692
rect -4692 -8747 -4654 -8730
rect -4788 -8764 -4772 -8747
rect -4848 -8780 -4772 -8764
rect -4670 -8764 -4654 -8747
rect -4610 -8747 -4572 -8730
rect -4514 -8730 -4394 -8692
rect -4514 -8747 -4476 -8730
rect -4610 -8764 -4594 -8747
rect -4670 -8780 -4594 -8764
rect -4492 -8764 -4476 -8747
rect -4432 -8747 -4394 -8730
rect -4336 -8730 -4216 -8692
rect -4336 -8747 -4298 -8730
rect -4432 -8764 -4416 -8747
rect -4492 -8780 -4416 -8764
rect -4314 -8764 -4298 -8747
rect -4254 -8747 -4216 -8730
rect -4158 -8730 -4038 -8692
rect -4158 -8747 -4120 -8730
rect -4254 -8764 -4238 -8747
rect -4314 -8780 -4238 -8764
rect -4136 -8764 -4120 -8747
rect -4076 -8747 -4038 -8730
rect -4076 -8764 -4060 -8747
rect -4136 -8780 -4060 -8764
rect 6580 -8810 6656 -8794
rect 6580 -8827 6596 -8810
rect 6558 -8844 6596 -8827
rect 6640 -8827 6656 -8810
rect 6758 -8810 6834 -8794
rect 6758 -8827 6774 -8810
rect 6640 -8844 6678 -8827
rect -5560 -8890 -5484 -8874
rect -5560 -8907 -5544 -8890
rect -5582 -8924 -5544 -8907
rect -5500 -8907 -5484 -8890
rect -5382 -8890 -5306 -8874
rect -5382 -8907 -5366 -8890
rect -5500 -8924 -5462 -8907
rect -5582 -8962 -5462 -8924
rect -5404 -8924 -5366 -8907
rect -5322 -8907 -5306 -8890
rect -5204 -8890 -5128 -8874
rect -5204 -8907 -5188 -8890
rect -5322 -8924 -5284 -8907
rect -5404 -8962 -5284 -8924
rect -5226 -8924 -5188 -8907
rect -5144 -8907 -5128 -8890
rect -5026 -8890 -4950 -8874
rect -5026 -8907 -5010 -8890
rect -5144 -8924 -5106 -8907
rect -5226 -8962 -5106 -8924
rect -5048 -8924 -5010 -8907
rect -4966 -8907 -4950 -8890
rect -4848 -8890 -4772 -8874
rect -4848 -8907 -4832 -8890
rect -4966 -8924 -4928 -8907
rect -5048 -8962 -4928 -8924
rect -4870 -8924 -4832 -8907
rect -4788 -8907 -4772 -8890
rect -4670 -8890 -4594 -8874
rect -4670 -8907 -4654 -8890
rect -4788 -8924 -4750 -8907
rect -4870 -8962 -4750 -8924
rect -4692 -8924 -4654 -8907
rect -4610 -8907 -4594 -8890
rect -4492 -8890 -4416 -8874
rect -4492 -8907 -4476 -8890
rect -4610 -8924 -4572 -8907
rect -4692 -8962 -4572 -8924
rect -4514 -8924 -4476 -8907
rect -4432 -8907 -4416 -8890
rect -4314 -8890 -4238 -8874
rect -4314 -8907 -4298 -8890
rect -4432 -8924 -4394 -8907
rect -4514 -8962 -4394 -8924
rect -4336 -8924 -4298 -8907
rect -4254 -8907 -4238 -8890
rect -4136 -8890 -4060 -8874
rect 6558 -8882 6678 -8844
rect 6736 -8844 6774 -8827
rect 6818 -8827 6834 -8810
rect 6936 -8810 7012 -8794
rect 6936 -8827 6952 -8810
rect 6818 -8844 6856 -8827
rect 6736 -8882 6856 -8844
rect 6914 -8844 6952 -8827
rect 6996 -8827 7012 -8810
rect 7114 -8810 7190 -8794
rect 7114 -8827 7130 -8810
rect 6996 -8844 7034 -8827
rect 6914 -8882 7034 -8844
rect 7092 -8844 7130 -8827
rect 7174 -8827 7190 -8810
rect 7292 -8810 7368 -8794
rect 7292 -8827 7308 -8810
rect 7174 -8844 7212 -8827
rect 7092 -8882 7212 -8844
rect 7270 -8844 7308 -8827
rect 7352 -8827 7368 -8810
rect 7470 -8810 7546 -8794
rect 7470 -8827 7486 -8810
rect 7352 -8844 7390 -8827
rect 7270 -8882 7390 -8844
rect 7448 -8844 7486 -8827
rect 7530 -8827 7546 -8810
rect 7648 -8810 7724 -8794
rect 7648 -8827 7664 -8810
rect 7530 -8844 7568 -8827
rect 7448 -8882 7568 -8844
rect 7626 -8844 7664 -8827
rect 7708 -8827 7724 -8810
rect 7826 -8810 7902 -8794
rect 7826 -8827 7842 -8810
rect 7708 -8844 7746 -8827
rect 7626 -8882 7746 -8844
rect 7804 -8844 7842 -8827
rect 7886 -8827 7902 -8810
rect 8004 -8810 8080 -8794
rect 8004 -8827 8020 -8810
rect 7886 -8844 7924 -8827
rect 7804 -8882 7924 -8844
rect 7982 -8844 8020 -8827
rect 8064 -8827 8080 -8810
rect 8182 -8810 8258 -8794
rect 8182 -8827 8198 -8810
rect 8064 -8844 8102 -8827
rect 7982 -8882 8102 -8844
rect 8160 -8844 8198 -8827
rect 8242 -8827 8258 -8810
rect 8360 -8810 8436 -8794
rect 8360 -8827 8376 -8810
rect 8242 -8844 8280 -8827
rect 8160 -8882 8280 -8844
rect 8338 -8844 8376 -8827
rect 8420 -8827 8436 -8810
rect 8538 -8810 8614 -8794
rect 8538 -8827 8554 -8810
rect 8420 -8844 8458 -8827
rect 8338 -8882 8458 -8844
rect 8516 -8844 8554 -8827
rect 8598 -8827 8614 -8810
rect 8716 -8810 8792 -8794
rect 8716 -8827 8732 -8810
rect 8598 -8844 8636 -8827
rect 8516 -8882 8636 -8844
rect 8694 -8844 8732 -8827
rect 8776 -8827 8792 -8810
rect 8894 -8810 8970 -8794
rect 8894 -8827 8910 -8810
rect 8776 -8844 8814 -8827
rect 8694 -8882 8814 -8844
rect 8872 -8844 8910 -8827
rect 8954 -8827 8970 -8810
rect 9072 -8810 9148 -8794
rect 9072 -8827 9088 -8810
rect 8954 -8844 8992 -8827
rect 8872 -8882 8992 -8844
rect 9050 -8844 9088 -8827
rect 9132 -8827 9148 -8810
rect 9250 -8810 9326 -8794
rect 9250 -8827 9266 -8810
rect 9132 -8844 9170 -8827
rect 9050 -8882 9170 -8844
rect 9228 -8844 9266 -8827
rect 9310 -8827 9326 -8810
rect 9310 -8844 9348 -8827
rect 9228 -8882 9348 -8844
rect 10840 -8840 10916 -8824
rect 10840 -8857 10856 -8840
rect 10818 -8874 10856 -8857
rect 10900 -8857 10916 -8840
rect 11132 -8840 11208 -8824
rect 11132 -8857 11148 -8840
rect 10900 -8874 10938 -8857
rect -4136 -8907 -4120 -8890
rect -4254 -8924 -4216 -8907
rect -4336 -8962 -4216 -8924
rect -4158 -8924 -4120 -8907
rect -4076 -8907 -4060 -8890
rect -4076 -8924 -4038 -8907
rect -4158 -8962 -4038 -8924
rect -2105 -9048 -2029 -9032
rect -2105 -9065 -2089 -9048
rect -2127 -9082 -2089 -9065
rect -2045 -9065 -2029 -9048
rect -1927 -9048 -1851 -9032
rect -1927 -9065 -1911 -9048
rect -2045 -9082 -2007 -9065
rect -2127 -9120 -2007 -9082
rect -1949 -9082 -1911 -9065
rect -1867 -9065 -1851 -9048
rect -1749 -9048 -1673 -9032
rect -1749 -9065 -1733 -9048
rect -1867 -9082 -1829 -9065
rect -1949 -9120 -1829 -9082
rect -1771 -9082 -1733 -9065
rect -1689 -9065 -1673 -9048
rect -1571 -9048 -1495 -9032
rect -1571 -9065 -1555 -9048
rect -1689 -9082 -1651 -9065
rect -1771 -9120 -1651 -9082
rect -1593 -9082 -1555 -9065
rect -1511 -9065 -1495 -9048
rect -1393 -9048 -1317 -9032
rect -1393 -9065 -1377 -9048
rect -1511 -9082 -1473 -9065
rect -1593 -9120 -1473 -9082
rect -1415 -9082 -1377 -9065
rect -1333 -9065 -1317 -9048
rect -1215 -9048 -1139 -9032
rect -1215 -9065 -1199 -9048
rect -1333 -9082 -1295 -9065
rect -1415 -9120 -1295 -9082
rect -1237 -9082 -1199 -9065
rect -1155 -9065 -1139 -9048
rect -1037 -9048 -961 -9032
rect -1037 -9065 -1021 -9048
rect -1155 -9082 -1117 -9065
rect -1237 -9120 -1117 -9082
rect -1059 -9082 -1021 -9065
rect -977 -9065 -961 -9048
rect -859 -9048 -783 -9032
rect -859 -9065 -843 -9048
rect -977 -9082 -939 -9065
rect -1059 -9120 -939 -9082
rect -881 -9082 -843 -9065
rect -799 -9065 -783 -9048
rect -681 -9048 -605 -9032
rect -681 -9065 -665 -9048
rect -799 -9082 -761 -9065
rect -881 -9120 -761 -9082
rect -703 -9082 -665 -9065
rect -621 -9065 -605 -9048
rect -503 -9048 -427 -9032
rect -503 -9065 -487 -9048
rect -621 -9082 -583 -9065
rect -703 -9120 -583 -9082
rect -525 -9082 -487 -9065
rect -443 -9065 -427 -9048
rect -325 -9048 -249 -9032
rect -325 -9065 -309 -9048
rect -443 -9082 -405 -9065
rect -525 -9120 -405 -9082
rect -347 -9082 -309 -9065
rect -265 -9065 -249 -9048
rect -147 -9048 -71 -9032
rect -147 -9065 -131 -9048
rect -265 -9082 -227 -9065
rect -347 -9120 -227 -9082
rect -169 -9082 -131 -9065
rect -87 -9065 -71 -9048
rect 31 -9048 107 -9032
rect 31 -9065 47 -9048
rect -87 -9082 -49 -9065
rect -169 -9120 -49 -9082
rect 9 -9082 47 -9065
rect 91 -9065 107 -9048
rect 209 -9048 285 -9032
rect 209 -9065 225 -9048
rect 91 -9082 129 -9065
rect 9 -9120 129 -9082
rect 187 -9082 225 -9065
rect 269 -9065 285 -9048
rect 387 -9048 463 -9032
rect 387 -9065 403 -9048
rect 269 -9082 307 -9065
rect 187 -9120 307 -9082
rect 365 -9082 403 -9065
rect 447 -9065 463 -9048
rect 565 -9048 641 -9032
rect 565 -9065 581 -9048
rect 447 -9082 485 -9065
rect 365 -9120 485 -9082
rect 543 -9082 581 -9065
rect 625 -9065 641 -9048
rect 743 -9048 819 -9032
rect 743 -9065 759 -9048
rect 625 -9082 663 -9065
rect 543 -9120 663 -9082
rect 721 -9082 759 -9065
rect 803 -9065 819 -9048
rect 921 -9048 997 -9032
rect 921 -9065 937 -9048
rect 803 -9082 841 -9065
rect 721 -9120 841 -9082
rect 899 -9082 937 -9065
rect 981 -9065 997 -9048
rect 1099 -9048 1175 -9032
rect 1099 -9065 1115 -9048
rect 981 -9082 1019 -9065
rect 899 -9120 1019 -9082
rect 1077 -9082 1115 -9065
rect 1159 -9065 1175 -9048
rect 1277 -9048 1353 -9032
rect 1277 -9065 1293 -9048
rect 1159 -9082 1197 -9065
rect 1077 -9120 1197 -9082
rect 1255 -9082 1293 -9065
rect 1337 -9065 1353 -9048
rect 1455 -9048 1531 -9032
rect 1455 -9065 1471 -9048
rect 1337 -9082 1375 -9065
rect 1255 -9120 1375 -9082
rect 1433 -9082 1471 -9065
rect 1515 -9065 1531 -9048
rect 1633 -9048 1709 -9032
rect 1633 -9065 1649 -9048
rect 1515 -9082 1553 -9065
rect 1433 -9120 1553 -9082
rect 1611 -9082 1649 -9065
rect 1693 -9065 1709 -9048
rect 1811 -9048 1887 -9032
rect 1811 -9065 1827 -9048
rect 1693 -9082 1731 -9065
rect 1611 -9120 1731 -9082
rect 1789 -9082 1827 -9065
rect 1871 -9065 1887 -9048
rect 1989 -9048 2065 -9032
rect 1989 -9065 2005 -9048
rect 1871 -9082 1909 -9065
rect 1789 -9120 1909 -9082
rect 1967 -9082 2005 -9065
rect 2049 -9065 2065 -9048
rect 2167 -9048 2243 -9032
rect 2167 -9065 2183 -9048
rect 2049 -9082 2087 -9065
rect 1967 -9120 2087 -9082
rect 2145 -9082 2183 -9065
rect 2227 -9065 2243 -9048
rect 2345 -9048 2421 -9032
rect 2345 -9065 2361 -9048
rect 2227 -9082 2265 -9065
rect 2145 -9120 2265 -9082
rect 2323 -9082 2361 -9065
rect 2405 -9065 2421 -9048
rect 2523 -9048 2599 -9032
rect 2523 -9065 2539 -9048
rect 2405 -9082 2443 -9065
rect 2323 -9120 2443 -9082
rect 2501 -9082 2539 -9065
rect 2583 -9065 2599 -9048
rect 2701 -9048 2777 -9032
rect 2701 -9065 2717 -9048
rect 2583 -9082 2621 -9065
rect 2501 -9120 2621 -9082
rect 2679 -9082 2717 -9065
rect 2761 -9065 2777 -9048
rect 2879 -9048 2955 -9032
rect 2879 -9065 2895 -9048
rect 2761 -9082 2799 -9065
rect 2679 -9120 2799 -9082
rect 2857 -9082 2895 -9065
rect 2939 -9065 2955 -9048
rect 3057 -9048 3133 -9032
rect 3057 -9065 3073 -9048
rect 2939 -9082 2977 -9065
rect 2857 -9120 2977 -9082
rect 3035 -9082 3073 -9065
rect 3117 -9065 3133 -9048
rect 3235 -9048 3311 -9032
rect 3235 -9065 3251 -9048
rect 3117 -9082 3155 -9065
rect 3035 -9120 3155 -9082
rect 3213 -9082 3251 -9065
rect 3295 -9065 3311 -9048
rect 3413 -9048 3489 -9032
rect 3413 -9065 3429 -9048
rect 3295 -9082 3333 -9065
rect 3213 -9120 3333 -9082
rect 3391 -9082 3429 -9065
rect 3473 -9065 3489 -9048
rect 3591 -9048 3667 -9032
rect 3591 -9065 3607 -9048
rect 3473 -9082 3511 -9065
rect 3391 -9120 3511 -9082
rect 3569 -9082 3607 -9065
rect 3651 -9065 3667 -9048
rect 3769 -9048 3845 -9032
rect 3769 -9065 3785 -9048
rect 3651 -9082 3689 -9065
rect 3569 -9120 3689 -9082
rect 3747 -9082 3785 -9065
rect 3829 -9065 3845 -9048
rect 3947 -9048 4023 -9032
rect 3947 -9065 3963 -9048
rect 3829 -9082 3867 -9065
rect 3747 -9120 3867 -9082
rect 3925 -9082 3963 -9065
rect 4007 -9065 4023 -9048
rect 4007 -9082 4045 -9065
rect 3925 -9120 4045 -9082
rect -5582 -9280 -5462 -9242
rect -5582 -9297 -5544 -9280
rect -5560 -9314 -5544 -9297
rect -5500 -9297 -5462 -9280
rect -5404 -9280 -5284 -9242
rect -5404 -9297 -5366 -9280
rect -5500 -9314 -5484 -9297
rect -5560 -9330 -5484 -9314
rect -5382 -9314 -5366 -9297
rect -5322 -9297 -5284 -9280
rect -5226 -9280 -5106 -9242
rect -5226 -9297 -5188 -9280
rect -5322 -9314 -5306 -9297
rect -5382 -9330 -5306 -9314
rect -5204 -9314 -5188 -9297
rect -5144 -9297 -5106 -9280
rect -5048 -9280 -4928 -9242
rect -5048 -9297 -5010 -9280
rect -5144 -9314 -5128 -9297
rect -5204 -9330 -5128 -9314
rect -5026 -9314 -5010 -9297
rect -4966 -9297 -4928 -9280
rect -4870 -9280 -4750 -9242
rect -4870 -9297 -4832 -9280
rect -4966 -9314 -4950 -9297
rect -5026 -9330 -4950 -9314
rect -4848 -9314 -4832 -9297
rect -4788 -9297 -4750 -9280
rect -4692 -9280 -4572 -9242
rect -4692 -9297 -4654 -9280
rect -4788 -9314 -4772 -9297
rect -4848 -9330 -4772 -9314
rect -4670 -9314 -4654 -9297
rect -4610 -9297 -4572 -9280
rect -4514 -9280 -4394 -9242
rect -4514 -9297 -4476 -9280
rect -4610 -9314 -4594 -9297
rect -4670 -9330 -4594 -9314
rect -4492 -9314 -4476 -9297
rect -4432 -9297 -4394 -9280
rect -4336 -9280 -4216 -9242
rect -4336 -9297 -4298 -9280
rect -4432 -9314 -4416 -9297
rect -4492 -9330 -4416 -9314
rect -4314 -9314 -4298 -9297
rect -4254 -9297 -4216 -9280
rect -4158 -9280 -4038 -9242
rect -4158 -9297 -4120 -9280
rect -4254 -9314 -4238 -9297
rect -4314 -9330 -4238 -9314
rect -4136 -9314 -4120 -9297
rect -4076 -9297 -4038 -9280
rect -4076 -9314 -4060 -9297
rect -4136 -9330 -4060 -9314
rect 10818 -8912 10938 -8874
rect 11110 -8874 11148 -8857
rect 11192 -8857 11208 -8840
rect 11424 -8840 11500 -8824
rect 11424 -8857 11440 -8840
rect 11192 -8874 11230 -8857
rect 11110 -8912 11230 -8874
rect 11402 -8874 11440 -8857
rect 11484 -8857 11500 -8840
rect 11716 -8840 11792 -8824
rect 11716 -8857 11732 -8840
rect 11484 -8874 11522 -8857
rect 11402 -8912 11522 -8874
rect 11694 -8874 11732 -8857
rect 11776 -8857 11792 -8840
rect 12008 -8840 12084 -8824
rect 12008 -8857 12024 -8840
rect 11776 -8874 11814 -8857
rect 11694 -8912 11814 -8874
rect 11986 -8874 12024 -8857
rect 12068 -8857 12084 -8840
rect 12300 -8840 12376 -8824
rect 12300 -8857 12316 -8840
rect 12068 -8874 12106 -8857
rect 11986 -8912 12106 -8874
rect 12278 -8874 12316 -8857
rect 12360 -8857 12376 -8840
rect 12592 -8840 12668 -8824
rect 12592 -8857 12608 -8840
rect 12360 -8874 12398 -8857
rect 12278 -8912 12398 -8874
rect 12570 -8874 12608 -8857
rect 12652 -8857 12668 -8840
rect 12652 -8874 12690 -8857
rect 12570 -8912 12690 -8874
rect 6558 -9200 6678 -9162
rect 6558 -9217 6596 -9200
rect 6580 -9234 6596 -9217
rect 6640 -9217 6678 -9200
rect 6736 -9200 6856 -9162
rect 6736 -9217 6774 -9200
rect 6640 -9234 6656 -9217
rect 6580 -9250 6656 -9234
rect 6758 -9234 6774 -9217
rect 6818 -9217 6856 -9200
rect 6914 -9200 7034 -9162
rect 6914 -9217 6952 -9200
rect 6818 -9234 6834 -9217
rect 6758 -9250 6834 -9234
rect 6936 -9234 6952 -9217
rect 6996 -9217 7034 -9200
rect 7092 -9200 7212 -9162
rect 7092 -9217 7130 -9200
rect 6996 -9234 7012 -9217
rect 6936 -9250 7012 -9234
rect 7114 -9234 7130 -9217
rect 7174 -9217 7212 -9200
rect 7270 -9200 7390 -9162
rect 7270 -9217 7308 -9200
rect 7174 -9234 7190 -9217
rect 7114 -9250 7190 -9234
rect 7292 -9234 7308 -9217
rect 7352 -9217 7390 -9200
rect 7448 -9200 7568 -9162
rect 7448 -9217 7486 -9200
rect 7352 -9234 7368 -9217
rect 7292 -9250 7368 -9234
rect 7470 -9234 7486 -9217
rect 7530 -9217 7568 -9200
rect 7626 -9200 7746 -9162
rect 7626 -9217 7664 -9200
rect 7530 -9234 7546 -9217
rect 7470 -9250 7546 -9234
rect 7648 -9234 7664 -9217
rect 7708 -9217 7746 -9200
rect 7804 -9200 7924 -9162
rect 7804 -9217 7842 -9200
rect 7708 -9234 7724 -9217
rect 7648 -9250 7724 -9234
rect 7826 -9234 7842 -9217
rect 7886 -9217 7924 -9200
rect 7982 -9200 8102 -9162
rect 7982 -9217 8020 -9200
rect 7886 -9234 7902 -9217
rect 7826 -9250 7902 -9234
rect 8004 -9234 8020 -9217
rect 8064 -9217 8102 -9200
rect 8160 -9200 8280 -9162
rect 8160 -9217 8198 -9200
rect 8064 -9234 8080 -9217
rect 8004 -9250 8080 -9234
rect 8182 -9234 8198 -9217
rect 8242 -9217 8280 -9200
rect 8338 -9200 8458 -9162
rect 8338 -9217 8376 -9200
rect 8242 -9234 8258 -9217
rect 8182 -9250 8258 -9234
rect 8360 -9234 8376 -9217
rect 8420 -9217 8458 -9200
rect 8516 -9200 8636 -9162
rect 8516 -9217 8554 -9200
rect 8420 -9234 8436 -9217
rect 8360 -9250 8436 -9234
rect 8538 -9234 8554 -9217
rect 8598 -9217 8636 -9200
rect 8694 -9200 8814 -9162
rect 8694 -9217 8732 -9200
rect 8598 -9234 8614 -9217
rect 8538 -9250 8614 -9234
rect 8716 -9234 8732 -9217
rect 8776 -9217 8814 -9200
rect 8872 -9200 8992 -9162
rect 8872 -9217 8910 -9200
rect 8776 -9234 8792 -9217
rect 8716 -9250 8792 -9234
rect 8894 -9234 8910 -9217
rect 8954 -9217 8992 -9200
rect 9050 -9200 9170 -9162
rect 9050 -9217 9088 -9200
rect 8954 -9234 8970 -9217
rect 8894 -9250 8970 -9234
rect 9072 -9234 9088 -9217
rect 9132 -9217 9170 -9200
rect 9228 -9200 9348 -9162
rect 9228 -9217 9266 -9200
rect 9132 -9234 9148 -9217
rect 9072 -9250 9148 -9234
rect 9250 -9234 9266 -9217
rect 9310 -9217 9348 -9200
rect 9310 -9234 9326 -9217
rect 9250 -9250 9326 -9234
rect 10818 -9230 10938 -9192
rect 10818 -9247 10856 -9230
rect 10840 -9264 10856 -9247
rect 10900 -9247 10938 -9230
rect 11110 -9230 11230 -9192
rect 11110 -9247 11148 -9230
rect 10900 -9264 10916 -9247
rect 10840 -9280 10916 -9264
rect 11132 -9264 11148 -9247
rect 11192 -9247 11230 -9230
rect 11402 -9230 11522 -9192
rect 11402 -9247 11440 -9230
rect 11192 -9264 11208 -9247
rect 11132 -9280 11208 -9264
rect 11424 -9264 11440 -9247
rect 11484 -9247 11522 -9230
rect 11694 -9230 11814 -9192
rect 11694 -9247 11732 -9230
rect 11484 -9264 11500 -9247
rect 11424 -9280 11500 -9264
rect 11716 -9264 11732 -9247
rect 11776 -9247 11814 -9230
rect 11986 -9230 12106 -9192
rect 11986 -9247 12024 -9230
rect 11776 -9264 11792 -9247
rect 11716 -9280 11792 -9264
rect 12008 -9264 12024 -9247
rect 12068 -9247 12106 -9230
rect 12278 -9230 12398 -9192
rect 12278 -9247 12316 -9230
rect 12068 -9264 12084 -9247
rect 12008 -9280 12084 -9264
rect 12300 -9264 12316 -9247
rect 12360 -9247 12398 -9230
rect 12570 -9230 12690 -9192
rect 12570 -9247 12608 -9230
rect 12360 -9264 12376 -9247
rect 12300 -9280 12376 -9264
rect 12592 -9264 12608 -9247
rect 12652 -9247 12690 -9230
rect 12652 -9264 12668 -9247
rect 12592 -9280 12668 -9264
rect -5560 -9440 -5484 -9424
rect -5560 -9457 -5544 -9440
rect -5582 -9474 -5544 -9457
rect -5500 -9457 -5484 -9440
rect -5382 -9440 -5306 -9424
rect -5382 -9457 -5366 -9440
rect -5500 -9474 -5462 -9457
rect -5582 -9512 -5462 -9474
rect -5404 -9474 -5366 -9457
rect -5322 -9457 -5306 -9440
rect -5204 -9440 -5128 -9424
rect -5204 -9457 -5188 -9440
rect -5322 -9474 -5284 -9457
rect -5404 -9512 -5284 -9474
rect -5226 -9474 -5188 -9457
rect -5144 -9457 -5128 -9440
rect -5026 -9440 -4950 -9424
rect -5026 -9457 -5010 -9440
rect -5144 -9474 -5106 -9457
rect -5226 -9512 -5106 -9474
rect -5048 -9474 -5010 -9457
rect -4966 -9457 -4950 -9440
rect -4848 -9440 -4772 -9424
rect -4848 -9457 -4832 -9440
rect -4966 -9474 -4928 -9457
rect -5048 -9512 -4928 -9474
rect -4870 -9474 -4832 -9457
rect -4788 -9457 -4772 -9440
rect -4670 -9440 -4594 -9424
rect -4670 -9457 -4654 -9440
rect -4788 -9474 -4750 -9457
rect -4870 -9512 -4750 -9474
rect -4692 -9474 -4654 -9457
rect -4610 -9457 -4594 -9440
rect -4492 -9440 -4416 -9424
rect -4492 -9457 -4476 -9440
rect -4610 -9474 -4572 -9457
rect -4692 -9512 -4572 -9474
rect -4514 -9474 -4476 -9457
rect -4432 -9457 -4416 -9440
rect -4314 -9440 -4238 -9424
rect -4314 -9457 -4298 -9440
rect -4432 -9474 -4394 -9457
rect -4514 -9512 -4394 -9474
rect -4336 -9474 -4298 -9457
rect -4254 -9457 -4238 -9440
rect -4136 -9440 -4060 -9424
rect -4136 -9457 -4120 -9440
rect -4254 -9474 -4216 -9457
rect -4336 -9512 -4216 -9474
rect -4158 -9474 -4120 -9457
rect -4076 -9457 -4060 -9440
rect -2127 -9438 -2007 -9400
rect -2127 -9455 -2089 -9438
rect -4076 -9474 -4038 -9457
rect -4158 -9512 -4038 -9474
rect -2105 -9472 -2089 -9455
rect -2045 -9455 -2007 -9438
rect -1949 -9438 -1829 -9400
rect -1949 -9455 -1911 -9438
rect -2045 -9472 -2029 -9455
rect -2105 -9488 -2029 -9472
rect -1927 -9472 -1911 -9455
rect -1867 -9455 -1829 -9438
rect -1771 -9438 -1651 -9400
rect -1771 -9455 -1733 -9438
rect -1867 -9472 -1851 -9455
rect -1927 -9488 -1851 -9472
rect -1749 -9472 -1733 -9455
rect -1689 -9455 -1651 -9438
rect -1593 -9438 -1473 -9400
rect -1593 -9455 -1555 -9438
rect -1689 -9472 -1673 -9455
rect -1749 -9488 -1673 -9472
rect -1571 -9472 -1555 -9455
rect -1511 -9455 -1473 -9438
rect -1415 -9438 -1295 -9400
rect -1415 -9455 -1377 -9438
rect -1511 -9472 -1495 -9455
rect -1571 -9488 -1495 -9472
rect -1393 -9472 -1377 -9455
rect -1333 -9455 -1295 -9438
rect -1237 -9438 -1117 -9400
rect -1237 -9455 -1199 -9438
rect -1333 -9472 -1317 -9455
rect -1393 -9488 -1317 -9472
rect -1215 -9472 -1199 -9455
rect -1155 -9455 -1117 -9438
rect -1059 -9438 -939 -9400
rect -1059 -9455 -1021 -9438
rect -1155 -9472 -1139 -9455
rect -1215 -9488 -1139 -9472
rect -1037 -9472 -1021 -9455
rect -977 -9455 -939 -9438
rect -881 -9438 -761 -9400
rect -881 -9455 -843 -9438
rect -977 -9472 -961 -9455
rect -1037 -9488 -961 -9472
rect -859 -9472 -843 -9455
rect -799 -9455 -761 -9438
rect -703 -9438 -583 -9400
rect -703 -9455 -665 -9438
rect -799 -9472 -783 -9455
rect -859 -9488 -783 -9472
rect -681 -9472 -665 -9455
rect -621 -9455 -583 -9438
rect -525 -9438 -405 -9400
rect -525 -9455 -487 -9438
rect -621 -9472 -605 -9455
rect -681 -9488 -605 -9472
rect -503 -9472 -487 -9455
rect -443 -9455 -405 -9438
rect -347 -9438 -227 -9400
rect -347 -9455 -309 -9438
rect -443 -9472 -427 -9455
rect -503 -9488 -427 -9472
rect -325 -9472 -309 -9455
rect -265 -9455 -227 -9438
rect -169 -9438 -49 -9400
rect -169 -9455 -131 -9438
rect -265 -9472 -249 -9455
rect -325 -9488 -249 -9472
rect -147 -9472 -131 -9455
rect -87 -9455 -49 -9438
rect 9 -9438 129 -9400
rect 9 -9455 47 -9438
rect -87 -9472 -71 -9455
rect -147 -9488 -71 -9472
rect 31 -9472 47 -9455
rect 91 -9455 129 -9438
rect 187 -9438 307 -9400
rect 187 -9455 225 -9438
rect 91 -9472 107 -9455
rect 31 -9488 107 -9472
rect 209 -9472 225 -9455
rect 269 -9455 307 -9438
rect 365 -9438 485 -9400
rect 365 -9455 403 -9438
rect 269 -9472 285 -9455
rect 209 -9488 285 -9472
rect 387 -9472 403 -9455
rect 447 -9455 485 -9438
rect 543 -9438 663 -9400
rect 543 -9455 581 -9438
rect 447 -9472 463 -9455
rect 387 -9488 463 -9472
rect 565 -9472 581 -9455
rect 625 -9455 663 -9438
rect 721 -9438 841 -9400
rect 721 -9455 759 -9438
rect 625 -9472 641 -9455
rect 565 -9488 641 -9472
rect 743 -9472 759 -9455
rect 803 -9455 841 -9438
rect 899 -9438 1019 -9400
rect 899 -9455 937 -9438
rect 803 -9472 819 -9455
rect 743 -9488 819 -9472
rect 921 -9472 937 -9455
rect 981 -9455 1019 -9438
rect 1077 -9438 1197 -9400
rect 1077 -9455 1115 -9438
rect 981 -9472 997 -9455
rect 921 -9488 997 -9472
rect 1099 -9472 1115 -9455
rect 1159 -9455 1197 -9438
rect 1255 -9438 1375 -9400
rect 1255 -9455 1293 -9438
rect 1159 -9472 1175 -9455
rect 1099 -9488 1175 -9472
rect 1277 -9472 1293 -9455
rect 1337 -9455 1375 -9438
rect 1433 -9438 1553 -9400
rect 1433 -9455 1471 -9438
rect 1337 -9472 1353 -9455
rect 1277 -9488 1353 -9472
rect 1455 -9472 1471 -9455
rect 1515 -9455 1553 -9438
rect 1611 -9438 1731 -9400
rect 1611 -9455 1649 -9438
rect 1515 -9472 1531 -9455
rect 1455 -9488 1531 -9472
rect 1633 -9472 1649 -9455
rect 1693 -9455 1731 -9438
rect 1789 -9438 1909 -9400
rect 1789 -9455 1827 -9438
rect 1693 -9472 1709 -9455
rect 1633 -9488 1709 -9472
rect 1811 -9472 1827 -9455
rect 1871 -9455 1909 -9438
rect 1967 -9438 2087 -9400
rect 1967 -9455 2005 -9438
rect 1871 -9472 1887 -9455
rect 1811 -9488 1887 -9472
rect 1989 -9472 2005 -9455
rect 2049 -9455 2087 -9438
rect 2145 -9438 2265 -9400
rect 2145 -9455 2183 -9438
rect 2049 -9472 2065 -9455
rect 1989 -9488 2065 -9472
rect 2167 -9472 2183 -9455
rect 2227 -9455 2265 -9438
rect 2323 -9438 2443 -9400
rect 2323 -9455 2361 -9438
rect 2227 -9472 2243 -9455
rect 2167 -9488 2243 -9472
rect 2345 -9472 2361 -9455
rect 2405 -9455 2443 -9438
rect 2501 -9438 2621 -9400
rect 2501 -9455 2539 -9438
rect 2405 -9472 2421 -9455
rect 2345 -9488 2421 -9472
rect 2523 -9472 2539 -9455
rect 2583 -9455 2621 -9438
rect 2679 -9438 2799 -9400
rect 2679 -9455 2717 -9438
rect 2583 -9472 2599 -9455
rect 2523 -9488 2599 -9472
rect 2701 -9472 2717 -9455
rect 2761 -9455 2799 -9438
rect 2857 -9438 2977 -9400
rect 2857 -9455 2895 -9438
rect 2761 -9472 2777 -9455
rect 2701 -9488 2777 -9472
rect 2879 -9472 2895 -9455
rect 2939 -9455 2977 -9438
rect 3035 -9438 3155 -9400
rect 3035 -9455 3073 -9438
rect 2939 -9472 2955 -9455
rect 2879 -9488 2955 -9472
rect 3057 -9472 3073 -9455
rect 3117 -9455 3155 -9438
rect 3213 -9438 3333 -9400
rect 3213 -9455 3251 -9438
rect 3117 -9472 3133 -9455
rect 3057 -9488 3133 -9472
rect 3235 -9472 3251 -9455
rect 3295 -9455 3333 -9438
rect 3391 -9438 3511 -9400
rect 3391 -9455 3429 -9438
rect 3295 -9472 3311 -9455
rect 3235 -9488 3311 -9472
rect 3413 -9472 3429 -9455
rect 3473 -9455 3511 -9438
rect 3569 -9438 3689 -9400
rect 3569 -9455 3607 -9438
rect 3473 -9472 3489 -9455
rect 3413 -9488 3489 -9472
rect 3591 -9472 3607 -9455
rect 3651 -9455 3689 -9438
rect 3747 -9438 3867 -9400
rect 3747 -9455 3785 -9438
rect 3651 -9472 3667 -9455
rect 3591 -9488 3667 -9472
rect 3769 -9472 3785 -9455
rect 3829 -9455 3867 -9438
rect 3925 -9438 4045 -9400
rect 3925 -9455 3963 -9438
rect 3829 -9472 3845 -9455
rect 3769 -9488 3845 -9472
rect 3947 -9472 3963 -9455
rect 4007 -9455 4045 -9438
rect 4007 -9472 4023 -9455
rect 3947 -9488 4023 -9472
rect 10840 -9610 10916 -9594
rect 10840 -9627 10856 -9610
rect 10818 -9644 10856 -9627
rect 10900 -9627 10916 -9610
rect 11132 -9610 11208 -9594
rect 11132 -9627 11148 -9610
rect 10900 -9644 10938 -9627
rect 10818 -9682 10938 -9644
rect 11110 -9644 11148 -9627
rect 11192 -9627 11208 -9610
rect 11424 -9610 11500 -9594
rect 11424 -9627 11440 -9610
rect 11192 -9644 11230 -9627
rect 11110 -9682 11230 -9644
rect 11402 -9644 11440 -9627
rect 11484 -9627 11500 -9610
rect 11716 -9610 11792 -9594
rect 11716 -9627 11732 -9610
rect 11484 -9644 11522 -9627
rect 11402 -9682 11522 -9644
rect 11694 -9644 11732 -9627
rect 11776 -9627 11792 -9610
rect 12008 -9610 12084 -9594
rect 12008 -9627 12024 -9610
rect 11776 -9644 11814 -9627
rect 11694 -9682 11814 -9644
rect 11986 -9644 12024 -9627
rect 12068 -9627 12084 -9610
rect 12300 -9610 12376 -9594
rect 12300 -9627 12316 -9610
rect 12068 -9644 12106 -9627
rect 11986 -9682 12106 -9644
rect 12278 -9644 12316 -9627
rect 12360 -9627 12376 -9610
rect 12592 -9610 12668 -9594
rect 12592 -9627 12608 -9610
rect 12360 -9644 12398 -9627
rect 12278 -9682 12398 -9644
rect 12570 -9644 12608 -9627
rect 12652 -9627 12668 -9610
rect 12652 -9644 12690 -9627
rect 12570 -9682 12690 -9644
rect 6580 -9710 6656 -9694
rect 6580 -9727 6596 -9710
rect 6558 -9744 6596 -9727
rect 6640 -9727 6656 -9710
rect 6758 -9710 6834 -9694
rect 6758 -9727 6774 -9710
rect 6640 -9744 6678 -9727
rect 6558 -9782 6678 -9744
rect 6736 -9744 6774 -9727
rect 6818 -9727 6834 -9710
rect 6936 -9710 7012 -9694
rect 6936 -9727 6952 -9710
rect 6818 -9744 6856 -9727
rect 6736 -9782 6856 -9744
rect 6914 -9744 6952 -9727
rect 6996 -9727 7012 -9710
rect 7114 -9710 7190 -9694
rect 7114 -9727 7130 -9710
rect 6996 -9744 7034 -9727
rect 6914 -9782 7034 -9744
rect 7092 -9744 7130 -9727
rect 7174 -9727 7190 -9710
rect 7292 -9710 7368 -9694
rect 7292 -9727 7308 -9710
rect 7174 -9744 7212 -9727
rect 7092 -9782 7212 -9744
rect 7270 -9744 7308 -9727
rect 7352 -9727 7368 -9710
rect 7470 -9710 7546 -9694
rect 7470 -9727 7486 -9710
rect 7352 -9744 7390 -9727
rect 7270 -9782 7390 -9744
rect 7448 -9744 7486 -9727
rect 7530 -9727 7546 -9710
rect 7648 -9710 7724 -9694
rect 7648 -9727 7664 -9710
rect 7530 -9744 7568 -9727
rect 7448 -9782 7568 -9744
rect 7626 -9744 7664 -9727
rect 7708 -9727 7724 -9710
rect 7826 -9710 7902 -9694
rect 7826 -9727 7842 -9710
rect 7708 -9744 7746 -9727
rect 7626 -9782 7746 -9744
rect 7804 -9744 7842 -9727
rect 7886 -9727 7902 -9710
rect 8004 -9710 8080 -9694
rect 8004 -9727 8020 -9710
rect 7886 -9744 7924 -9727
rect 7804 -9782 7924 -9744
rect 7982 -9744 8020 -9727
rect 8064 -9727 8080 -9710
rect 8182 -9710 8258 -9694
rect 8182 -9727 8198 -9710
rect 8064 -9744 8102 -9727
rect 7982 -9782 8102 -9744
rect 8160 -9744 8198 -9727
rect 8242 -9727 8258 -9710
rect 8360 -9710 8436 -9694
rect 8360 -9727 8376 -9710
rect 8242 -9744 8280 -9727
rect 8160 -9782 8280 -9744
rect 8338 -9744 8376 -9727
rect 8420 -9727 8436 -9710
rect 8538 -9710 8614 -9694
rect 8538 -9727 8554 -9710
rect 8420 -9744 8458 -9727
rect 8338 -9782 8458 -9744
rect 8516 -9744 8554 -9727
rect 8598 -9727 8614 -9710
rect 8716 -9710 8792 -9694
rect 8716 -9727 8732 -9710
rect 8598 -9744 8636 -9727
rect 8516 -9782 8636 -9744
rect 8694 -9744 8732 -9727
rect 8776 -9727 8792 -9710
rect 8894 -9710 8970 -9694
rect 8894 -9727 8910 -9710
rect 8776 -9744 8814 -9727
rect 8694 -9782 8814 -9744
rect 8872 -9744 8910 -9727
rect 8954 -9727 8970 -9710
rect 9072 -9710 9148 -9694
rect 9072 -9727 9088 -9710
rect 8954 -9744 8992 -9727
rect 8872 -9782 8992 -9744
rect 9050 -9744 9088 -9727
rect 9132 -9727 9148 -9710
rect 9250 -9710 9326 -9694
rect 9250 -9727 9266 -9710
rect 9132 -9744 9170 -9727
rect 9050 -9782 9170 -9744
rect 9228 -9744 9266 -9727
rect 9310 -9727 9326 -9710
rect 9310 -9744 9348 -9727
rect 9228 -9782 9348 -9744
rect -5582 -9830 -5462 -9792
rect -5582 -9847 -5544 -9830
rect -5560 -9864 -5544 -9847
rect -5500 -9847 -5462 -9830
rect -5404 -9830 -5284 -9792
rect -5404 -9847 -5366 -9830
rect -5500 -9864 -5484 -9847
rect -5560 -9880 -5484 -9864
rect -5382 -9864 -5366 -9847
rect -5322 -9847 -5284 -9830
rect -5226 -9830 -5106 -9792
rect -5226 -9847 -5188 -9830
rect -5322 -9864 -5306 -9847
rect -5382 -9880 -5306 -9864
rect -5204 -9864 -5188 -9847
rect -5144 -9847 -5106 -9830
rect -5048 -9830 -4928 -9792
rect -5048 -9847 -5010 -9830
rect -5144 -9864 -5128 -9847
rect -5204 -9880 -5128 -9864
rect -5026 -9864 -5010 -9847
rect -4966 -9847 -4928 -9830
rect -4870 -9830 -4750 -9792
rect -4870 -9847 -4832 -9830
rect -4966 -9864 -4950 -9847
rect -5026 -9880 -4950 -9864
rect -4848 -9864 -4832 -9847
rect -4788 -9847 -4750 -9830
rect -4692 -9830 -4572 -9792
rect -4692 -9847 -4654 -9830
rect -4788 -9864 -4772 -9847
rect -4848 -9880 -4772 -9864
rect -4670 -9864 -4654 -9847
rect -4610 -9847 -4572 -9830
rect -4514 -9830 -4394 -9792
rect -4514 -9847 -4476 -9830
rect -4610 -9864 -4594 -9847
rect -4670 -9880 -4594 -9864
rect -4492 -9864 -4476 -9847
rect -4432 -9847 -4394 -9830
rect -4336 -9830 -4216 -9792
rect -4336 -9847 -4298 -9830
rect -4432 -9864 -4416 -9847
rect -4492 -9880 -4416 -9864
rect -4314 -9864 -4298 -9847
rect -4254 -9847 -4216 -9830
rect -4158 -9830 -4038 -9792
rect -4158 -9847 -4120 -9830
rect -4254 -9864 -4238 -9847
rect -4314 -9880 -4238 -9864
rect -4136 -9864 -4120 -9847
rect -4076 -9847 -4038 -9830
rect -4076 -9864 -4060 -9847
rect -4136 -9880 -4060 -9864
rect -5560 -9990 -5484 -9974
rect -5560 -10007 -5544 -9990
rect -5582 -10024 -5544 -10007
rect -5500 -10007 -5484 -9990
rect -5382 -9990 -5306 -9974
rect -5382 -10007 -5366 -9990
rect -5500 -10024 -5462 -10007
rect -5582 -10062 -5462 -10024
rect -5404 -10024 -5366 -10007
rect -5322 -10007 -5306 -9990
rect -5204 -9990 -5128 -9974
rect -5204 -10007 -5188 -9990
rect -5322 -10024 -5284 -10007
rect -5404 -10062 -5284 -10024
rect -5226 -10024 -5188 -10007
rect -5144 -10007 -5128 -9990
rect -5026 -9990 -4950 -9974
rect -5026 -10007 -5010 -9990
rect -5144 -10024 -5106 -10007
rect -5226 -10062 -5106 -10024
rect -5048 -10024 -5010 -10007
rect -4966 -10007 -4950 -9990
rect -4848 -9990 -4772 -9974
rect -4848 -10007 -4832 -9990
rect -4966 -10024 -4928 -10007
rect -5048 -10062 -4928 -10024
rect -4870 -10024 -4832 -10007
rect -4788 -10007 -4772 -9990
rect -4670 -9990 -4594 -9974
rect -4670 -10007 -4654 -9990
rect -4788 -10024 -4750 -10007
rect -4870 -10062 -4750 -10024
rect -4692 -10024 -4654 -10007
rect -4610 -10007 -4594 -9990
rect -4492 -9990 -4416 -9974
rect -4492 -10007 -4476 -9990
rect -4610 -10024 -4572 -10007
rect -4692 -10062 -4572 -10024
rect -4514 -10024 -4476 -10007
rect -4432 -10007 -4416 -9990
rect -4314 -9990 -4238 -9974
rect -4314 -10007 -4298 -9990
rect -4432 -10024 -4394 -10007
rect -4514 -10062 -4394 -10024
rect -4336 -10024 -4298 -10007
rect -4254 -10007 -4238 -9990
rect -4136 -9990 -4060 -9974
rect -4136 -10007 -4120 -9990
rect -4254 -10024 -4216 -10007
rect -4336 -10062 -4216 -10024
rect -4158 -10024 -4120 -10007
rect -4076 -10007 -4060 -9990
rect -4076 -10024 -4038 -10007
rect -4158 -10062 -4038 -10024
rect -2105 -10048 -2029 -10032
rect -2105 -10065 -2089 -10048
rect -2127 -10082 -2089 -10065
rect -2045 -10065 -2029 -10048
rect -1927 -10048 -1851 -10032
rect -1927 -10065 -1911 -10048
rect -2045 -10082 -2007 -10065
rect -2127 -10120 -2007 -10082
rect -1949 -10082 -1911 -10065
rect -1867 -10065 -1851 -10048
rect -1749 -10048 -1673 -10032
rect -1749 -10065 -1733 -10048
rect -1867 -10082 -1829 -10065
rect -1949 -10120 -1829 -10082
rect -1771 -10082 -1733 -10065
rect -1689 -10065 -1673 -10048
rect -1571 -10048 -1495 -10032
rect -1571 -10065 -1555 -10048
rect -1689 -10082 -1651 -10065
rect -1771 -10120 -1651 -10082
rect -1593 -10082 -1555 -10065
rect -1511 -10065 -1495 -10048
rect -1393 -10048 -1317 -10032
rect -1393 -10065 -1377 -10048
rect -1511 -10082 -1473 -10065
rect -1593 -10120 -1473 -10082
rect -1415 -10082 -1377 -10065
rect -1333 -10065 -1317 -10048
rect -1215 -10048 -1139 -10032
rect -1215 -10065 -1199 -10048
rect -1333 -10082 -1295 -10065
rect -1415 -10120 -1295 -10082
rect -1237 -10082 -1199 -10065
rect -1155 -10065 -1139 -10048
rect -1037 -10048 -961 -10032
rect -1037 -10065 -1021 -10048
rect -1155 -10082 -1117 -10065
rect -1237 -10120 -1117 -10082
rect -1059 -10082 -1021 -10065
rect -977 -10065 -961 -10048
rect -859 -10048 -783 -10032
rect -859 -10065 -843 -10048
rect -977 -10082 -939 -10065
rect -1059 -10120 -939 -10082
rect -881 -10082 -843 -10065
rect -799 -10065 -783 -10048
rect -681 -10048 -605 -10032
rect -681 -10065 -665 -10048
rect -799 -10082 -761 -10065
rect -881 -10120 -761 -10082
rect -703 -10082 -665 -10065
rect -621 -10065 -605 -10048
rect -503 -10048 -427 -10032
rect -503 -10065 -487 -10048
rect -621 -10082 -583 -10065
rect -703 -10120 -583 -10082
rect -525 -10082 -487 -10065
rect -443 -10065 -427 -10048
rect -325 -10048 -249 -10032
rect -325 -10065 -309 -10048
rect -443 -10082 -405 -10065
rect -525 -10120 -405 -10082
rect -347 -10082 -309 -10065
rect -265 -10065 -249 -10048
rect -147 -10048 -71 -10032
rect -147 -10065 -131 -10048
rect -265 -10082 -227 -10065
rect -347 -10120 -227 -10082
rect -169 -10082 -131 -10065
rect -87 -10065 -71 -10048
rect 31 -10048 107 -10032
rect 31 -10065 47 -10048
rect -87 -10082 -49 -10065
rect -169 -10120 -49 -10082
rect 9 -10082 47 -10065
rect 91 -10065 107 -10048
rect 209 -10048 285 -10032
rect 209 -10065 225 -10048
rect 91 -10082 129 -10065
rect 9 -10120 129 -10082
rect 187 -10082 225 -10065
rect 269 -10065 285 -10048
rect 387 -10048 463 -10032
rect 387 -10065 403 -10048
rect 269 -10082 307 -10065
rect 187 -10120 307 -10082
rect 365 -10082 403 -10065
rect 447 -10065 463 -10048
rect 565 -10048 641 -10032
rect 565 -10065 581 -10048
rect 447 -10082 485 -10065
rect 365 -10120 485 -10082
rect 543 -10082 581 -10065
rect 625 -10065 641 -10048
rect 743 -10048 819 -10032
rect 743 -10065 759 -10048
rect 625 -10082 663 -10065
rect 543 -10120 663 -10082
rect 721 -10082 759 -10065
rect 803 -10065 819 -10048
rect 921 -10048 997 -10032
rect 921 -10065 937 -10048
rect 803 -10082 841 -10065
rect 721 -10120 841 -10082
rect 899 -10082 937 -10065
rect 981 -10065 997 -10048
rect 1099 -10048 1175 -10032
rect 1099 -10065 1115 -10048
rect 981 -10082 1019 -10065
rect 899 -10120 1019 -10082
rect 1077 -10082 1115 -10065
rect 1159 -10065 1175 -10048
rect 1277 -10048 1353 -10032
rect 1277 -10065 1293 -10048
rect 1159 -10082 1197 -10065
rect 1077 -10120 1197 -10082
rect 1255 -10082 1293 -10065
rect 1337 -10065 1353 -10048
rect 1455 -10048 1531 -10032
rect 1455 -10065 1471 -10048
rect 1337 -10082 1375 -10065
rect 1255 -10120 1375 -10082
rect 1433 -10082 1471 -10065
rect 1515 -10065 1531 -10048
rect 1633 -10048 1709 -10032
rect 1633 -10065 1649 -10048
rect 1515 -10082 1553 -10065
rect 1433 -10120 1553 -10082
rect 1611 -10082 1649 -10065
rect 1693 -10065 1709 -10048
rect 1811 -10048 1887 -10032
rect 1811 -10065 1827 -10048
rect 1693 -10082 1731 -10065
rect 1611 -10120 1731 -10082
rect 1789 -10082 1827 -10065
rect 1871 -10065 1887 -10048
rect 1989 -10048 2065 -10032
rect 1989 -10065 2005 -10048
rect 1871 -10082 1909 -10065
rect 1789 -10120 1909 -10082
rect 1967 -10082 2005 -10065
rect 2049 -10065 2065 -10048
rect 2167 -10048 2243 -10032
rect 2167 -10065 2183 -10048
rect 2049 -10082 2087 -10065
rect 1967 -10120 2087 -10082
rect 2145 -10082 2183 -10065
rect 2227 -10065 2243 -10048
rect 2345 -10048 2421 -10032
rect 2345 -10065 2361 -10048
rect 2227 -10082 2265 -10065
rect 2145 -10120 2265 -10082
rect 2323 -10082 2361 -10065
rect 2405 -10065 2421 -10048
rect 2523 -10048 2599 -10032
rect 2523 -10065 2539 -10048
rect 2405 -10082 2443 -10065
rect 2323 -10120 2443 -10082
rect 2501 -10082 2539 -10065
rect 2583 -10065 2599 -10048
rect 2701 -10048 2777 -10032
rect 2701 -10065 2717 -10048
rect 2583 -10082 2621 -10065
rect 2501 -10120 2621 -10082
rect 2679 -10082 2717 -10065
rect 2761 -10065 2777 -10048
rect 2879 -10048 2955 -10032
rect 2879 -10065 2895 -10048
rect 2761 -10082 2799 -10065
rect 2679 -10120 2799 -10082
rect 2857 -10082 2895 -10065
rect 2939 -10065 2955 -10048
rect 3057 -10048 3133 -10032
rect 3057 -10065 3073 -10048
rect 2939 -10082 2977 -10065
rect 2857 -10120 2977 -10082
rect 3035 -10082 3073 -10065
rect 3117 -10065 3133 -10048
rect 3235 -10048 3311 -10032
rect 3235 -10065 3251 -10048
rect 3117 -10082 3155 -10065
rect 3035 -10120 3155 -10082
rect 3213 -10082 3251 -10065
rect 3295 -10065 3311 -10048
rect 3413 -10048 3489 -10032
rect 3413 -10065 3429 -10048
rect 3295 -10082 3333 -10065
rect 3213 -10120 3333 -10082
rect 3391 -10082 3429 -10065
rect 3473 -10065 3489 -10048
rect 3591 -10048 3667 -10032
rect 3591 -10065 3607 -10048
rect 3473 -10082 3511 -10065
rect 3391 -10120 3511 -10082
rect 3569 -10082 3607 -10065
rect 3651 -10065 3667 -10048
rect 3769 -10048 3845 -10032
rect 3769 -10065 3785 -10048
rect 3651 -10082 3689 -10065
rect 3569 -10120 3689 -10082
rect 3747 -10082 3785 -10065
rect 3829 -10065 3845 -10048
rect 3947 -10048 4023 -10032
rect 3947 -10065 3963 -10048
rect 3829 -10082 3867 -10065
rect 3747 -10120 3867 -10082
rect 3925 -10082 3963 -10065
rect 4007 -10065 4023 -10048
rect 10818 -10000 10938 -9962
rect 10818 -10017 10856 -10000
rect 10840 -10034 10856 -10017
rect 10900 -10017 10938 -10000
rect 11110 -10000 11230 -9962
rect 11110 -10017 11148 -10000
rect 10900 -10034 10916 -10017
rect 10840 -10050 10916 -10034
rect 11132 -10034 11148 -10017
rect 11192 -10017 11230 -10000
rect 11402 -10000 11522 -9962
rect 11402 -10017 11440 -10000
rect 11192 -10034 11208 -10017
rect 11132 -10050 11208 -10034
rect 11424 -10034 11440 -10017
rect 11484 -10017 11522 -10000
rect 11694 -10000 11814 -9962
rect 11694 -10017 11732 -10000
rect 11484 -10034 11500 -10017
rect 11424 -10050 11500 -10034
rect 11716 -10034 11732 -10017
rect 11776 -10017 11814 -10000
rect 11986 -10000 12106 -9962
rect 11986 -10017 12024 -10000
rect 11776 -10034 11792 -10017
rect 11716 -10050 11792 -10034
rect 12008 -10034 12024 -10017
rect 12068 -10017 12106 -10000
rect 12278 -10000 12398 -9962
rect 12278 -10017 12316 -10000
rect 12068 -10034 12084 -10017
rect 12008 -10050 12084 -10034
rect 12300 -10034 12316 -10017
rect 12360 -10017 12398 -10000
rect 12570 -10000 12690 -9962
rect 12570 -10017 12608 -10000
rect 12360 -10034 12376 -10017
rect 12300 -10050 12376 -10034
rect 12592 -10034 12608 -10017
rect 12652 -10017 12690 -10000
rect 12652 -10034 12668 -10017
rect 12592 -10050 12668 -10034
rect 4007 -10082 4045 -10065
rect 3925 -10120 4045 -10082
rect 6558 -10100 6678 -10062
rect 6558 -10117 6596 -10100
rect -5582 -10380 -5462 -10342
rect -5582 -10397 -5544 -10380
rect -5560 -10414 -5544 -10397
rect -5500 -10397 -5462 -10380
rect -5404 -10380 -5284 -10342
rect -5404 -10397 -5366 -10380
rect -5500 -10414 -5484 -10397
rect -5560 -10430 -5484 -10414
rect -5382 -10414 -5366 -10397
rect -5322 -10397 -5284 -10380
rect -5226 -10380 -5106 -10342
rect -5226 -10397 -5188 -10380
rect -5322 -10414 -5306 -10397
rect -5382 -10430 -5306 -10414
rect -5204 -10414 -5188 -10397
rect -5144 -10397 -5106 -10380
rect -5048 -10380 -4928 -10342
rect -5048 -10397 -5010 -10380
rect -5144 -10414 -5128 -10397
rect -5204 -10430 -5128 -10414
rect -5026 -10414 -5010 -10397
rect -4966 -10397 -4928 -10380
rect -4870 -10380 -4750 -10342
rect -4870 -10397 -4832 -10380
rect -4966 -10414 -4950 -10397
rect -5026 -10430 -4950 -10414
rect -4848 -10414 -4832 -10397
rect -4788 -10397 -4750 -10380
rect -4692 -10380 -4572 -10342
rect -4692 -10397 -4654 -10380
rect -4788 -10414 -4772 -10397
rect -4848 -10430 -4772 -10414
rect -4670 -10414 -4654 -10397
rect -4610 -10397 -4572 -10380
rect -4514 -10380 -4394 -10342
rect -4514 -10397 -4476 -10380
rect -4610 -10414 -4594 -10397
rect -4670 -10430 -4594 -10414
rect -4492 -10414 -4476 -10397
rect -4432 -10397 -4394 -10380
rect -4336 -10380 -4216 -10342
rect -4336 -10397 -4298 -10380
rect -4432 -10414 -4416 -10397
rect -4492 -10430 -4416 -10414
rect -4314 -10414 -4298 -10397
rect -4254 -10397 -4216 -10380
rect -4158 -10380 -4038 -10342
rect -4158 -10397 -4120 -10380
rect -4254 -10414 -4238 -10397
rect -4314 -10430 -4238 -10414
rect -4136 -10414 -4120 -10397
rect -4076 -10397 -4038 -10380
rect -4076 -10414 -4060 -10397
rect 6580 -10134 6596 -10117
rect 6640 -10117 6678 -10100
rect 6736 -10100 6856 -10062
rect 6736 -10117 6774 -10100
rect 6640 -10134 6656 -10117
rect 6580 -10150 6656 -10134
rect 6758 -10134 6774 -10117
rect 6818 -10117 6856 -10100
rect 6914 -10100 7034 -10062
rect 6914 -10117 6952 -10100
rect 6818 -10134 6834 -10117
rect 6758 -10150 6834 -10134
rect 6936 -10134 6952 -10117
rect 6996 -10117 7034 -10100
rect 7092 -10100 7212 -10062
rect 7092 -10117 7130 -10100
rect 6996 -10134 7012 -10117
rect 6936 -10150 7012 -10134
rect 7114 -10134 7130 -10117
rect 7174 -10117 7212 -10100
rect 7270 -10100 7390 -10062
rect 7270 -10117 7308 -10100
rect 7174 -10134 7190 -10117
rect 7114 -10150 7190 -10134
rect 7292 -10134 7308 -10117
rect 7352 -10117 7390 -10100
rect 7448 -10100 7568 -10062
rect 7448 -10117 7486 -10100
rect 7352 -10134 7368 -10117
rect 7292 -10150 7368 -10134
rect 7470 -10134 7486 -10117
rect 7530 -10117 7568 -10100
rect 7626 -10100 7746 -10062
rect 7626 -10117 7664 -10100
rect 7530 -10134 7546 -10117
rect 7470 -10150 7546 -10134
rect 7648 -10134 7664 -10117
rect 7708 -10117 7746 -10100
rect 7804 -10100 7924 -10062
rect 7804 -10117 7842 -10100
rect 7708 -10134 7724 -10117
rect 7648 -10150 7724 -10134
rect 7826 -10134 7842 -10117
rect 7886 -10117 7924 -10100
rect 7982 -10100 8102 -10062
rect 7982 -10117 8020 -10100
rect 7886 -10134 7902 -10117
rect 7826 -10150 7902 -10134
rect 8004 -10134 8020 -10117
rect 8064 -10117 8102 -10100
rect 8160 -10100 8280 -10062
rect 8160 -10117 8198 -10100
rect 8064 -10134 8080 -10117
rect 8004 -10150 8080 -10134
rect 8182 -10134 8198 -10117
rect 8242 -10117 8280 -10100
rect 8338 -10100 8458 -10062
rect 8338 -10117 8376 -10100
rect 8242 -10134 8258 -10117
rect 8182 -10150 8258 -10134
rect 8360 -10134 8376 -10117
rect 8420 -10117 8458 -10100
rect 8516 -10100 8636 -10062
rect 8516 -10117 8554 -10100
rect 8420 -10134 8436 -10117
rect 8360 -10150 8436 -10134
rect 8538 -10134 8554 -10117
rect 8598 -10117 8636 -10100
rect 8694 -10100 8814 -10062
rect 8694 -10117 8732 -10100
rect 8598 -10134 8614 -10117
rect 8538 -10150 8614 -10134
rect 8716 -10134 8732 -10117
rect 8776 -10117 8814 -10100
rect 8872 -10100 8992 -10062
rect 8872 -10117 8910 -10100
rect 8776 -10134 8792 -10117
rect 8716 -10150 8792 -10134
rect 8894 -10134 8910 -10117
rect 8954 -10117 8992 -10100
rect 9050 -10100 9170 -10062
rect 9050 -10117 9088 -10100
rect 8954 -10134 8970 -10117
rect 8894 -10150 8970 -10134
rect 9072 -10134 9088 -10117
rect 9132 -10117 9170 -10100
rect 9228 -10100 9348 -10062
rect 9228 -10117 9266 -10100
rect 9132 -10134 9148 -10117
rect 9072 -10150 9148 -10134
rect 9250 -10134 9266 -10117
rect 9310 -10117 9348 -10100
rect 9310 -10134 9326 -10117
rect 9250 -10150 9326 -10134
rect 10840 -10380 10916 -10364
rect 10840 -10397 10856 -10380
rect -4136 -10430 -4060 -10414
rect -2127 -10438 -2007 -10400
rect -2127 -10455 -2089 -10438
rect -2105 -10472 -2089 -10455
rect -2045 -10455 -2007 -10438
rect -1949 -10438 -1829 -10400
rect -1949 -10455 -1911 -10438
rect -2045 -10472 -2029 -10455
rect -2105 -10488 -2029 -10472
rect -1927 -10472 -1911 -10455
rect -1867 -10455 -1829 -10438
rect -1771 -10438 -1651 -10400
rect -1771 -10455 -1733 -10438
rect -1867 -10472 -1851 -10455
rect -1927 -10488 -1851 -10472
rect -1749 -10472 -1733 -10455
rect -1689 -10455 -1651 -10438
rect -1593 -10438 -1473 -10400
rect -1593 -10455 -1555 -10438
rect -1689 -10472 -1673 -10455
rect -1749 -10488 -1673 -10472
rect -1571 -10472 -1555 -10455
rect -1511 -10455 -1473 -10438
rect -1415 -10438 -1295 -10400
rect -1415 -10455 -1377 -10438
rect -1511 -10472 -1495 -10455
rect -1571 -10488 -1495 -10472
rect -1393 -10472 -1377 -10455
rect -1333 -10455 -1295 -10438
rect -1237 -10438 -1117 -10400
rect -1237 -10455 -1199 -10438
rect -1333 -10472 -1317 -10455
rect -1393 -10488 -1317 -10472
rect -1215 -10472 -1199 -10455
rect -1155 -10455 -1117 -10438
rect -1059 -10438 -939 -10400
rect -1059 -10455 -1021 -10438
rect -1155 -10472 -1139 -10455
rect -1215 -10488 -1139 -10472
rect -1037 -10472 -1021 -10455
rect -977 -10455 -939 -10438
rect -881 -10438 -761 -10400
rect -881 -10455 -843 -10438
rect -977 -10472 -961 -10455
rect -1037 -10488 -961 -10472
rect -859 -10472 -843 -10455
rect -799 -10455 -761 -10438
rect -703 -10438 -583 -10400
rect -703 -10455 -665 -10438
rect -799 -10472 -783 -10455
rect -859 -10488 -783 -10472
rect -681 -10472 -665 -10455
rect -621 -10455 -583 -10438
rect -525 -10438 -405 -10400
rect -525 -10455 -487 -10438
rect -621 -10472 -605 -10455
rect -681 -10488 -605 -10472
rect -503 -10472 -487 -10455
rect -443 -10455 -405 -10438
rect -347 -10438 -227 -10400
rect -347 -10455 -309 -10438
rect -443 -10472 -427 -10455
rect -503 -10488 -427 -10472
rect -325 -10472 -309 -10455
rect -265 -10455 -227 -10438
rect -169 -10438 -49 -10400
rect -169 -10455 -131 -10438
rect -265 -10472 -249 -10455
rect -325 -10488 -249 -10472
rect -147 -10472 -131 -10455
rect -87 -10455 -49 -10438
rect 9 -10438 129 -10400
rect 9 -10455 47 -10438
rect -87 -10472 -71 -10455
rect -147 -10488 -71 -10472
rect 31 -10472 47 -10455
rect 91 -10455 129 -10438
rect 187 -10438 307 -10400
rect 187 -10455 225 -10438
rect 91 -10472 107 -10455
rect 31 -10488 107 -10472
rect 209 -10472 225 -10455
rect 269 -10455 307 -10438
rect 365 -10438 485 -10400
rect 365 -10455 403 -10438
rect 269 -10472 285 -10455
rect 209 -10488 285 -10472
rect 387 -10472 403 -10455
rect 447 -10455 485 -10438
rect 543 -10438 663 -10400
rect 543 -10455 581 -10438
rect 447 -10472 463 -10455
rect 387 -10488 463 -10472
rect 565 -10472 581 -10455
rect 625 -10455 663 -10438
rect 721 -10438 841 -10400
rect 721 -10455 759 -10438
rect 625 -10472 641 -10455
rect 565 -10488 641 -10472
rect 743 -10472 759 -10455
rect 803 -10455 841 -10438
rect 899 -10438 1019 -10400
rect 899 -10455 937 -10438
rect 803 -10472 819 -10455
rect 743 -10488 819 -10472
rect 921 -10472 937 -10455
rect 981 -10455 1019 -10438
rect 1077 -10438 1197 -10400
rect 1077 -10455 1115 -10438
rect 981 -10472 997 -10455
rect 921 -10488 997 -10472
rect 1099 -10472 1115 -10455
rect 1159 -10455 1197 -10438
rect 1255 -10438 1375 -10400
rect 1255 -10455 1293 -10438
rect 1159 -10472 1175 -10455
rect 1099 -10488 1175 -10472
rect 1277 -10472 1293 -10455
rect 1337 -10455 1375 -10438
rect 1433 -10438 1553 -10400
rect 1433 -10455 1471 -10438
rect 1337 -10472 1353 -10455
rect 1277 -10488 1353 -10472
rect 1455 -10472 1471 -10455
rect 1515 -10455 1553 -10438
rect 1611 -10438 1731 -10400
rect 1611 -10455 1649 -10438
rect 1515 -10472 1531 -10455
rect 1455 -10488 1531 -10472
rect 1633 -10472 1649 -10455
rect 1693 -10455 1731 -10438
rect 1789 -10438 1909 -10400
rect 1789 -10455 1827 -10438
rect 1693 -10472 1709 -10455
rect 1633 -10488 1709 -10472
rect 1811 -10472 1827 -10455
rect 1871 -10455 1909 -10438
rect 1967 -10438 2087 -10400
rect 1967 -10455 2005 -10438
rect 1871 -10472 1887 -10455
rect 1811 -10488 1887 -10472
rect 1989 -10472 2005 -10455
rect 2049 -10455 2087 -10438
rect 2145 -10438 2265 -10400
rect 2145 -10455 2183 -10438
rect 2049 -10472 2065 -10455
rect 1989 -10488 2065 -10472
rect 2167 -10472 2183 -10455
rect 2227 -10455 2265 -10438
rect 2323 -10438 2443 -10400
rect 2323 -10455 2361 -10438
rect 2227 -10472 2243 -10455
rect 2167 -10488 2243 -10472
rect 2345 -10472 2361 -10455
rect 2405 -10455 2443 -10438
rect 2501 -10438 2621 -10400
rect 2501 -10455 2539 -10438
rect 2405 -10472 2421 -10455
rect 2345 -10488 2421 -10472
rect 2523 -10472 2539 -10455
rect 2583 -10455 2621 -10438
rect 2679 -10438 2799 -10400
rect 2679 -10455 2717 -10438
rect 2583 -10472 2599 -10455
rect 2523 -10488 2599 -10472
rect 2701 -10472 2717 -10455
rect 2761 -10455 2799 -10438
rect 2857 -10438 2977 -10400
rect 2857 -10455 2895 -10438
rect 2761 -10472 2777 -10455
rect 2701 -10488 2777 -10472
rect 2879 -10472 2895 -10455
rect 2939 -10455 2977 -10438
rect 3035 -10438 3155 -10400
rect 3035 -10455 3073 -10438
rect 2939 -10472 2955 -10455
rect 2879 -10488 2955 -10472
rect 3057 -10472 3073 -10455
rect 3117 -10455 3155 -10438
rect 3213 -10438 3333 -10400
rect 3213 -10455 3251 -10438
rect 3117 -10472 3133 -10455
rect 3057 -10488 3133 -10472
rect 3235 -10472 3251 -10455
rect 3295 -10455 3333 -10438
rect 3391 -10438 3511 -10400
rect 3391 -10455 3429 -10438
rect 3295 -10472 3311 -10455
rect 3235 -10488 3311 -10472
rect 3413 -10472 3429 -10455
rect 3473 -10455 3511 -10438
rect 3569 -10438 3689 -10400
rect 3569 -10455 3607 -10438
rect 3473 -10472 3489 -10455
rect 3413 -10488 3489 -10472
rect 3591 -10472 3607 -10455
rect 3651 -10455 3689 -10438
rect 3747 -10438 3867 -10400
rect 3747 -10455 3785 -10438
rect 3651 -10472 3667 -10455
rect 3591 -10488 3667 -10472
rect 3769 -10472 3785 -10455
rect 3829 -10455 3867 -10438
rect 3925 -10438 4045 -10400
rect 3925 -10455 3963 -10438
rect 3829 -10472 3845 -10455
rect 3769 -10488 3845 -10472
rect 3947 -10472 3963 -10455
rect 4007 -10455 4045 -10438
rect 10818 -10414 10856 -10397
rect 10900 -10397 10916 -10380
rect 11132 -10380 11208 -10364
rect 11132 -10397 11148 -10380
rect 10900 -10414 10938 -10397
rect 10818 -10452 10938 -10414
rect 11110 -10414 11148 -10397
rect 11192 -10397 11208 -10380
rect 11424 -10380 11500 -10364
rect 11424 -10397 11440 -10380
rect 11192 -10414 11230 -10397
rect 11110 -10452 11230 -10414
rect 11402 -10414 11440 -10397
rect 11484 -10397 11500 -10380
rect 11716 -10380 11792 -10364
rect 11716 -10397 11732 -10380
rect 11484 -10414 11522 -10397
rect 11402 -10452 11522 -10414
rect 11694 -10414 11732 -10397
rect 11776 -10397 11792 -10380
rect 12008 -10380 12084 -10364
rect 12008 -10397 12024 -10380
rect 11776 -10414 11814 -10397
rect 11694 -10452 11814 -10414
rect 11986 -10414 12024 -10397
rect 12068 -10397 12084 -10380
rect 12300 -10380 12376 -10364
rect 12300 -10397 12316 -10380
rect 12068 -10414 12106 -10397
rect 11986 -10452 12106 -10414
rect 12278 -10414 12316 -10397
rect 12360 -10397 12376 -10380
rect 12592 -10380 12668 -10364
rect 12592 -10397 12608 -10380
rect 12360 -10414 12398 -10397
rect 12278 -10452 12398 -10414
rect 12570 -10414 12608 -10397
rect 12652 -10397 12668 -10380
rect 12652 -10414 12690 -10397
rect 12570 -10452 12690 -10414
rect 4007 -10472 4023 -10455
rect 3947 -10488 4023 -10472
rect -5560 -10540 -5484 -10524
rect -5560 -10557 -5544 -10540
rect -5582 -10574 -5544 -10557
rect -5500 -10557 -5484 -10540
rect -5382 -10540 -5306 -10524
rect -5382 -10557 -5366 -10540
rect -5500 -10574 -5462 -10557
rect -5582 -10612 -5462 -10574
rect -5404 -10574 -5366 -10557
rect -5322 -10557 -5306 -10540
rect -5204 -10540 -5128 -10524
rect -5204 -10557 -5188 -10540
rect -5322 -10574 -5284 -10557
rect -5404 -10612 -5284 -10574
rect -5226 -10574 -5188 -10557
rect -5144 -10557 -5128 -10540
rect -5026 -10540 -4950 -10524
rect -5026 -10557 -5010 -10540
rect -5144 -10574 -5106 -10557
rect -5226 -10612 -5106 -10574
rect -5048 -10574 -5010 -10557
rect -4966 -10557 -4950 -10540
rect -4848 -10540 -4772 -10524
rect -4848 -10557 -4832 -10540
rect -4966 -10574 -4928 -10557
rect -5048 -10612 -4928 -10574
rect -4870 -10574 -4832 -10557
rect -4788 -10557 -4772 -10540
rect -4670 -10540 -4594 -10524
rect -4670 -10557 -4654 -10540
rect -4788 -10574 -4750 -10557
rect -4870 -10612 -4750 -10574
rect -4692 -10574 -4654 -10557
rect -4610 -10557 -4594 -10540
rect -4492 -10540 -4416 -10524
rect -4492 -10557 -4476 -10540
rect -4610 -10574 -4572 -10557
rect -4692 -10612 -4572 -10574
rect -4514 -10574 -4476 -10557
rect -4432 -10557 -4416 -10540
rect -4314 -10540 -4238 -10524
rect -4314 -10557 -4298 -10540
rect -4432 -10574 -4394 -10557
rect -4514 -10612 -4394 -10574
rect -4336 -10574 -4298 -10557
rect -4254 -10557 -4238 -10540
rect -4136 -10540 -4060 -10524
rect -4136 -10557 -4120 -10540
rect -4254 -10574 -4216 -10557
rect -4336 -10612 -4216 -10574
rect -4158 -10574 -4120 -10557
rect -4076 -10557 -4060 -10540
rect -4076 -10574 -4038 -10557
rect -4158 -10612 -4038 -10574
rect 6580 -10610 6656 -10594
rect 6580 -10627 6596 -10610
rect 6558 -10644 6596 -10627
rect 6640 -10627 6656 -10610
rect 6758 -10610 6834 -10594
rect 6758 -10627 6774 -10610
rect 6640 -10644 6678 -10627
rect 6558 -10682 6678 -10644
rect 6736 -10644 6774 -10627
rect 6818 -10627 6834 -10610
rect 6936 -10610 7012 -10594
rect 6936 -10627 6952 -10610
rect 6818 -10644 6856 -10627
rect 6736 -10682 6856 -10644
rect 6914 -10644 6952 -10627
rect 6996 -10627 7012 -10610
rect 7114 -10610 7190 -10594
rect 7114 -10627 7130 -10610
rect 6996 -10644 7034 -10627
rect 6914 -10682 7034 -10644
rect 7092 -10644 7130 -10627
rect 7174 -10627 7190 -10610
rect 7292 -10610 7368 -10594
rect 7292 -10627 7308 -10610
rect 7174 -10644 7212 -10627
rect 7092 -10682 7212 -10644
rect 7270 -10644 7308 -10627
rect 7352 -10627 7368 -10610
rect 7470 -10610 7546 -10594
rect 7470 -10627 7486 -10610
rect 7352 -10644 7390 -10627
rect 7270 -10682 7390 -10644
rect 7448 -10644 7486 -10627
rect 7530 -10627 7546 -10610
rect 7648 -10610 7724 -10594
rect 7648 -10627 7664 -10610
rect 7530 -10644 7568 -10627
rect 7448 -10682 7568 -10644
rect 7626 -10644 7664 -10627
rect 7708 -10627 7724 -10610
rect 7826 -10610 7902 -10594
rect 7826 -10627 7842 -10610
rect 7708 -10644 7746 -10627
rect 7626 -10682 7746 -10644
rect 7804 -10644 7842 -10627
rect 7886 -10627 7902 -10610
rect 8004 -10610 8080 -10594
rect 8004 -10627 8020 -10610
rect 7886 -10644 7924 -10627
rect 7804 -10682 7924 -10644
rect 7982 -10644 8020 -10627
rect 8064 -10627 8080 -10610
rect 8182 -10610 8258 -10594
rect 8182 -10627 8198 -10610
rect 8064 -10644 8102 -10627
rect 7982 -10682 8102 -10644
rect 8160 -10644 8198 -10627
rect 8242 -10627 8258 -10610
rect 8360 -10610 8436 -10594
rect 8360 -10627 8376 -10610
rect 8242 -10644 8280 -10627
rect 8160 -10682 8280 -10644
rect 8338 -10644 8376 -10627
rect 8420 -10627 8436 -10610
rect 8538 -10610 8614 -10594
rect 8538 -10627 8554 -10610
rect 8420 -10644 8458 -10627
rect 8338 -10682 8458 -10644
rect 8516 -10644 8554 -10627
rect 8598 -10627 8614 -10610
rect 8716 -10610 8792 -10594
rect 8716 -10627 8732 -10610
rect 8598 -10644 8636 -10627
rect 8516 -10682 8636 -10644
rect 8694 -10644 8732 -10627
rect 8776 -10627 8792 -10610
rect 8894 -10610 8970 -10594
rect 8894 -10627 8910 -10610
rect 8776 -10644 8814 -10627
rect 8694 -10682 8814 -10644
rect 8872 -10644 8910 -10627
rect 8954 -10627 8970 -10610
rect 9072 -10610 9148 -10594
rect 9072 -10627 9088 -10610
rect 8954 -10644 8992 -10627
rect 8872 -10682 8992 -10644
rect 9050 -10644 9088 -10627
rect 9132 -10627 9148 -10610
rect 9250 -10610 9326 -10594
rect 9250 -10627 9266 -10610
rect 9132 -10644 9170 -10627
rect 9050 -10682 9170 -10644
rect 9228 -10644 9266 -10627
rect 9310 -10627 9326 -10610
rect 9310 -10644 9348 -10627
rect 9228 -10682 9348 -10644
rect -5582 -10930 -5462 -10892
rect -5582 -10947 -5544 -10930
rect -5560 -10964 -5544 -10947
rect -5500 -10947 -5462 -10930
rect -5404 -10930 -5284 -10892
rect -5404 -10947 -5366 -10930
rect -5500 -10964 -5484 -10947
rect -5560 -10980 -5484 -10964
rect -5382 -10964 -5366 -10947
rect -5322 -10947 -5284 -10930
rect -5226 -10930 -5106 -10892
rect -5226 -10947 -5188 -10930
rect -5322 -10964 -5306 -10947
rect -5382 -10980 -5306 -10964
rect -5204 -10964 -5188 -10947
rect -5144 -10947 -5106 -10930
rect -5048 -10930 -4928 -10892
rect -5048 -10947 -5010 -10930
rect -5144 -10964 -5128 -10947
rect -5204 -10980 -5128 -10964
rect -5026 -10964 -5010 -10947
rect -4966 -10947 -4928 -10930
rect -4870 -10930 -4750 -10892
rect -4870 -10947 -4832 -10930
rect -4966 -10964 -4950 -10947
rect -5026 -10980 -4950 -10964
rect -4848 -10964 -4832 -10947
rect -4788 -10947 -4750 -10930
rect -4692 -10930 -4572 -10892
rect -4692 -10947 -4654 -10930
rect -4788 -10964 -4772 -10947
rect -4848 -10980 -4772 -10964
rect -4670 -10964 -4654 -10947
rect -4610 -10947 -4572 -10930
rect -4514 -10930 -4394 -10892
rect -4514 -10947 -4476 -10930
rect -4610 -10964 -4594 -10947
rect -4670 -10980 -4594 -10964
rect -4492 -10964 -4476 -10947
rect -4432 -10947 -4394 -10930
rect -4336 -10930 -4216 -10892
rect -4336 -10947 -4298 -10930
rect -4432 -10964 -4416 -10947
rect -4492 -10980 -4416 -10964
rect -4314 -10964 -4298 -10947
rect -4254 -10947 -4216 -10930
rect -4158 -10930 -4038 -10892
rect -4158 -10947 -4120 -10930
rect -4254 -10964 -4238 -10947
rect -4314 -10980 -4238 -10964
rect -4136 -10964 -4120 -10947
rect -4076 -10947 -4038 -10930
rect -4076 -10964 -4060 -10947
rect 10818 -10770 10938 -10732
rect 10818 -10787 10856 -10770
rect 10840 -10804 10856 -10787
rect 10900 -10787 10938 -10770
rect 11110 -10770 11230 -10732
rect 11110 -10787 11148 -10770
rect 10900 -10804 10916 -10787
rect 10840 -10820 10916 -10804
rect 11132 -10804 11148 -10787
rect 11192 -10787 11230 -10770
rect 11402 -10770 11522 -10732
rect 11402 -10787 11440 -10770
rect 11192 -10804 11208 -10787
rect 11132 -10820 11208 -10804
rect 11424 -10804 11440 -10787
rect 11484 -10787 11522 -10770
rect 11694 -10770 11814 -10732
rect 11694 -10787 11732 -10770
rect 11484 -10804 11500 -10787
rect 11424 -10820 11500 -10804
rect 11716 -10804 11732 -10787
rect 11776 -10787 11814 -10770
rect 11986 -10770 12106 -10732
rect 11986 -10787 12024 -10770
rect 11776 -10804 11792 -10787
rect 11716 -10820 11792 -10804
rect 12008 -10804 12024 -10787
rect 12068 -10787 12106 -10770
rect 12278 -10770 12398 -10732
rect 12278 -10787 12316 -10770
rect 12068 -10804 12084 -10787
rect 12008 -10820 12084 -10804
rect 12300 -10804 12316 -10787
rect 12360 -10787 12398 -10770
rect 12570 -10770 12690 -10732
rect 12570 -10787 12608 -10770
rect 12360 -10804 12376 -10787
rect 12300 -10820 12376 -10804
rect 12592 -10804 12608 -10787
rect 12652 -10787 12690 -10770
rect 12652 -10804 12668 -10787
rect 12592 -10820 12668 -10804
rect -4136 -10980 -4060 -10964
rect 6558 -11000 6678 -10962
rect 6558 -11017 6596 -11000
rect -2105 -11048 -2029 -11032
rect -2105 -11065 -2089 -11048
rect -5560 -11090 -5484 -11074
rect -5560 -11107 -5544 -11090
rect -5582 -11124 -5544 -11107
rect -5500 -11107 -5484 -11090
rect -5382 -11090 -5306 -11074
rect -5382 -11107 -5366 -11090
rect -5500 -11124 -5462 -11107
rect -5582 -11162 -5462 -11124
rect -5404 -11124 -5366 -11107
rect -5322 -11107 -5306 -11090
rect -5204 -11090 -5128 -11074
rect -5204 -11107 -5188 -11090
rect -5322 -11124 -5284 -11107
rect -5404 -11162 -5284 -11124
rect -5226 -11124 -5188 -11107
rect -5144 -11107 -5128 -11090
rect -5026 -11090 -4950 -11074
rect -5026 -11107 -5010 -11090
rect -5144 -11124 -5106 -11107
rect -5226 -11162 -5106 -11124
rect -5048 -11124 -5010 -11107
rect -4966 -11107 -4950 -11090
rect -4848 -11090 -4772 -11074
rect -4848 -11107 -4832 -11090
rect -4966 -11124 -4928 -11107
rect -5048 -11162 -4928 -11124
rect -4870 -11124 -4832 -11107
rect -4788 -11107 -4772 -11090
rect -4670 -11090 -4594 -11074
rect -4670 -11107 -4654 -11090
rect -4788 -11124 -4750 -11107
rect -4870 -11162 -4750 -11124
rect -4692 -11124 -4654 -11107
rect -4610 -11107 -4594 -11090
rect -4492 -11090 -4416 -11074
rect -4492 -11107 -4476 -11090
rect -4610 -11124 -4572 -11107
rect -4692 -11162 -4572 -11124
rect -4514 -11124 -4476 -11107
rect -4432 -11107 -4416 -11090
rect -4314 -11090 -4238 -11074
rect -4314 -11107 -4298 -11090
rect -4432 -11124 -4394 -11107
rect -4514 -11162 -4394 -11124
rect -4336 -11124 -4298 -11107
rect -4254 -11107 -4238 -11090
rect -4136 -11090 -4060 -11074
rect -4136 -11107 -4120 -11090
rect -4254 -11124 -4216 -11107
rect -4336 -11162 -4216 -11124
rect -4158 -11124 -4120 -11107
rect -4076 -11107 -4060 -11090
rect -2127 -11082 -2089 -11065
rect -2045 -11065 -2029 -11048
rect -1927 -11048 -1851 -11032
rect -1927 -11065 -1911 -11048
rect -2045 -11082 -2007 -11065
rect -4076 -11124 -4038 -11107
rect -2127 -11120 -2007 -11082
rect -1949 -11082 -1911 -11065
rect -1867 -11065 -1851 -11048
rect -1749 -11048 -1673 -11032
rect -1749 -11065 -1733 -11048
rect -1867 -11082 -1829 -11065
rect -1949 -11120 -1829 -11082
rect -1771 -11082 -1733 -11065
rect -1689 -11065 -1673 -11048
rect -1571 -11048 -1495 -11032
rect -1571 -11065 -1555 -11048
rect -1689 -11082 -1651 -11065
rect -1771 -11120 -1651 -11082
rect -1593 -11082 -1555 -11065
rect -1511 -11065 -1495 -11048
rect -1393 -11048 -1317 -11032
rect -1393 -11065 -1377 -11048
rect -1511 -11082 -1473 -11065
rect -1593 -11120 -1473 -11082
rect -1415 -11082 -1377 -11065
rect -1333 -11065 -1317 -11048
rect -1215 -11048 -1139 -11032
rect -1215 -11065 -1199 -11048
rect -1333 -11082 -1295 -11065
rect -1415 -11120 -1295 -11082
rect -1237 -11082 -1199 -11065
rect -1155 -11065 -1139 -11048
rect -1037 -11048 -961 -11032
rect -1037 -11065 -1021 -11048
rect -1155 -11082 -1117 -11065
rect -1237 -11120 -1117 -11082
rect -1059 -11082 -1021 -11065
rect -977 -11065 -961 -11048
rect -859 -11048 -783 -11032
rect -859 -11065 -843 -11048
rect -977 -11082 -939 -11065
rect -1059 -11120 -939 -11082
rect -881 -11082 -843 -11065
rect -799 -11065 -783 -11048
rect -681 -11048 -605 -11032
rect -681 -11065 -665 -11048
rect -799 -11082 -761 -11065
rect -881 -11120 -761 -11082
rect -703 -11082 -665 -11065
rect -621 -11065 -605 -11048
rect -503 -11048 -427 -11032
rect -503 -11065 -487 -11048
rect -621 -11082 -583 -11065
rect -703 -11120 -583 -11082
rect -525 -11082 -487 -11065
rect -443 -11065 -427 -11048
rect -325 -11048 -249 -11032
rect -325 -11065 -309 -11048
rect -443 -11082 -405 -11065
rect -525 -11120 -405 -11082
rect -347 -11082 -309 -11065
rect -265 -11065 -249 -11048
rect -147 -11048 -71 -11032
rect -147 -11065 -131 -11048
rect -265 -11082 -227 -11065
rect -347 -11120 -227 -11082
rect -169 -11082 -131 -11065
rect -87 -11065 -71 -11048
rect 31 -11048 107 -11032
rect 31 -11065 47 -11048
rect -87 -11082 -49 -11065
rect -169 -11120 -49 -11082
rect 9 -11082 47 -11065
rect 91 -11065 107 -11048
rect 209 -11048 285 -11032
rect 209 -11065 225 -11048
rect 91 -11082 129 -11065
rect 9 -11120 129 -11082
rect 187 -11082 225 -11065
rect 269 -11065 285 -11048
rect 387 -11048 463 -11032
rect 387 -11065 403 -11048
rect 269 -11082 307 -11065
rect 187 -11120 307 -11082
rect 365 -11082 403 -11065
rect 447 -11065 463 -11048
rect 565 -11048 641 -11032
rect 565 -11065 581 -11048
rect 447 -11082 485 -11065
rect 365 -11120 485 -11082
rect 543 -11082 581 -11065
rect 625 -11065 641 -11048
rect 743 -11048 819 -11032
rect 743 -11065 759 -11048
rect 625 -11082 663 -11065
rect 543 -11120 663 -11082
rect 721 -11082 759 -11065
rect 803 -11065 819 -11048
rect 921 -11048 997 -11032
rect 921 -11065 937 -11048
rect 803 -11082 841 -11065
rect 721 -11120 841 -11082
rect 899 -11082 937 -11065
rect 981 -11065 997 -11048
rect 1099 -11048 1175 -11032
rect 1099 -11065 1115 -11048
rect 981 -11082 1019 -11065
rect 899 -11120 1019 -11082
rect 1077 -11082 1115 -11065
rect 1159 -11065 1175 -11048
rect 1277 -11048 1353 -11032
rect 1277 -11065 1293 -11048
rect 1159 -11082 1197 -11065
rect 1077 -11120 1197 -11082
rect 1255 -11082 1293 -11065
rect 1337 -11065 1353 -11048
rect 1455 -11048 1531 -11032
rect 1455 -11065 1471 -11048
rect 1337 -11082 1375 -11065
rect 1255 -11120 1375 -11082
rect 1433 -11082 1471 -11065
rect 1515 -11065 1531 -11048
rect 1633 -11048 1709 -11032
rect 1633 -11065 1649 -11048
rect 1515 -11082 1553 -11065
rect 1433 -11120 1553 -11082
rect 1611 -11082 1649 -11065
rect 1693 -11065 1709 -11048
rect 1811 -11048 1887 -11032
rect 1811 -11065 1827 -11048
rect 1693 -11082 1731 -11065
rect 1611 -11120 1731 -11082
rect 1789 -11082 1827 -11065
rect 1871 -11065 1887 -11048
rect 1989 -11048 2065 -11032
rect 1989 -11065 2005 -11048
rect 1871 -11082 1909 -11065
rect 1789 -11120 1909 -11082
rect 1967 -11082 2005 -11065
rect 2049 -11065 2065 -11048
rect 2167 -11048 2243 -11032
rect 2167 -11065 2183 -11048
rect 2049 -11082 2087 -11065
rect 1967 -11120 2087 -11082
rect 2145 -11082 2183 -11065
rect 2227 -11065 2243 -11048
rect 2345 -11048 2421 -11032
rect 2345 -11065 2361 -11048
rect 2227 -11082 2265 -11065
rect 2145 -11120 2265 -11082
rect 2323 -11082 2361 -11065
rect 2405 -11065 2421 -11048
rect 2523 -11048 2599 -11032
rect 2523 -11065 2539 -11048
rect 2405 -11082 2443 -11065
rect 2323 -11120 2443 -11082
rect 2501 -11082 2539 -11065
rect 2583 -11065 2599 -11048
rect 2701 -11048 2777 -11032
rect 2701 -11065 2717 -11048
rect 2583 -11082 2621 -11065
rect 2501 -11120 2621 -11082
rect 2679 -11082 2717 -11065
rect 2761 -11065 2777 -11048
rect 2879 -11048 2955 -11032
rect 2879 -11065 2895 -11048
rect 2761 -11082 2799 -11065
rect 2679 -11120 2799 -11082
rect 2857 -11082 2895 -11065
rect 2939 -11065 2955 -11048
rect 3057 -11048 3133 -11032
rect 3057 -11065 3073 -11048
rect 2939 -11082 2977 -11065
rect 2857 -11120 2977 -11082
rect 3035 -11082 3073 -11065
rect 3117 -11065 3133 -11048
rect 3235 -11048 3311 -11032
rect 3235 -11065 3251 -11048
rect 3117 -11082 3155 -11065
rect 3035 -11120 3155 -11082
rect 3213 -11082 3251 -11065
rect 3295 -11065 3311 -11048
rect 3413 -11048 3489 -11032
rect 3413 -11065 3429 -11048
rect 3295 -11082 3333 -11065
rect 3213 -11120 3333 -11082
rect 3391 -11082 3429 -11065
rect 3473 -11065 3489 -11048
rect 3591 -11048 3667 -11032
rect 3591 -11065 3607 -11048
rect 3473 -11082 3511 -11065
rect 3391 -11120 3511 -11082
rect 3569 -11082 3607 -11065
rect 3651 -11065 3667 -11048
rect 3769 -11048 3845 -11032
rect 3769 -11065 3785 -11048
rect 3651 -11082 3689 -11065
rect 3569 -11120 3689 -11082
rect 3747 -11082 3785 -11065
rect 3829 -11065 3845 -11048
rect 3947 -11048 4023 -11032
rect 3947 -11065 3963 -11048
rect 3829 -11082 3867 -11065
rect 3747 -11120 3867 -11082
rect 3925 -11082 3963 -11065
rect 4007 -11065 4023 -11048
rect 6580 -11034 6596 -11017
rect 6640 -11017 6678 -11000
rect 6736 -11000 6856 -10962
rect 6736 -11017 6774 -11000
rect 6640 -11034 6656 -11017
rect 6580 -11050 6656 -11034
rect 6758 -11034 6774 -11017
rect 6818 -11017 6856 -11000
rect 6914 -11000 7034 -10962
rect 6914 -11017 6952 -11000
rect 6818 -11034 6834 -11017
rect 6758 -11050 6834 -11034
rect 6936 -11034 6952 -11017
rect 6996 -11017 7034 -11000
rect 7092 -11000 7212 -10962
rect 7092 -11017 7130 -11000
rect 6996 -11034 7012 -11017
rect 6936 -11050 7012 -11034
rect 7114 -11034 7130 -11017
rect 7174 -11017 7212 -11000
rect 7270 -11000 7390 -10962
rect 7270 -11017 7308 -11000
rect 7174 -11034 7190 -11017
rect 7114 -11050 7190 -11034
rect 7292 -11034 7308 -11017
rect 7352 -11017 7390 -11000
rect 7448 -11000 7568 -10962
rect 7448 -11017 7486 -11000
rect 7352 -11034 7368 -11017
rect 7292 -11050 7368 -11034
rect 7470 -11034 7486 -11017
rect 7530 -11017 7568 -11000
rect 7626 -11000 7746 -10962
rect 7626 -11017 7664 -11000
rect 7530 -11034 7546 -11017
rect 7470 -11050 7546 -11034
rect 7648 -11034 7664 -11017
rect 7708 -11017 7746 -11000
rect 7804 -11000 7924 -10962
rect 7804 -11017 7842 -11000
rect 7708 -11034 7724 -11017
rect 7648 -11050 7724 -11034
rect 7826 -11034 7842 -11017
rect 7886 -11017 7924 -11000
rect 7982 -11000 8102 -10962
rect 7982 -11017 8020 -11000
rect 7886 -11034 7902 -11017
rect 7826 -11050 7902 -11034
rect 8004 -11034 8020 -11017
rect 8064 -11017 8102 -11000
rect 8160 -11000 8280 -10962
rect 8160 -11017 8198 -11000
rect 8064 -11034 8080 -11017
rect 8004 -11050 8080 -11034
rect 8182 -11034 8198 -11017
rect 8242 -11017 8280 -11000
rect 8338 -11000 8458 -10962
rect 8338 -11017 8376 -11000
rect 8242 -11034 8258 -11017
rect 8182 -11050 8258 -11034
rect 8360 -11034 8376 -11017
rect 8420 -11017 8458 -11000
rect 8516 -11000 8636 -10962
rect 8516 -11017 8554 -11000
rect 8420 -11034 8436 -11017
rect 8360 -11050 8436 -11034
rect 8538 -11034 8554 -11017
rect 8598 -11017 8636 -11000
rect 8694 -11000 8814 -10962
rect 8694 -11017 8732 -11000
rect 8598 -11034 8614 -11017
rect 8538 -11050 8614 -11034
rect 8716 -11034 8732 -11017
rect 8776 -11017 8814 -11000
rect 8872 -11000 8992 -10962
rect 8872 -11017 8910 -11000
rect 8776 -11034 8792 -11017
rect 8716 -11050 8792 -11034
rect 8894 -11034 8910 -11017
rect 8954 -11017 8992 -11000
rect 9050 -11000 9170 -10962
rect 9050 -11017 9088 -11000
rect 8954 -11034 8970 -11017
rect 8894 -11050 8970 -11034
rect 9072 -11034 9088 -11017
rect 9132 -11017 9170 -11000
rect 9228 -11000 9348 -10962
rect 9228 -11017 9266 -11000
rect 9132 -11034 9148 -11017
rect 9072 -11050 9148 -11034
rect 9250 -11034 9266 -11017
rect 9310 -11017 9348 -11000
rect 9310 -11034 9326 -11017
rect 9250 -11050 9326 -11034
rect 4007 -11082 4045 -11065
rect 3925 -11120 4045 -11082
rect -4158 -11162 -4038 -11124
rect 10840 -11150 10916 -11134
rect 10840 -11167 10856 -11150
rect 10818 -11184 10856 -11167
rect 10900 -11167 10916 -11150
rect 11132 -11150 11208 -11134
rect 11132 -11167 11148 -11150
rect 10900 -11184 10938 -11167
rect 10818 -11222 10938 -11184
rect 11110 -11184 11148 -11167
rect 11192 -11167 11208 -11150
rect 11424 -11150 11500 -11134
rect 11424 -11167 11440 -11150
rect 11192 -11184 11230 -11167
rect 11110 -11222 11230 -11184
rect 11402 -11184 11440 -11167
rect 11484 -11167 11500 -11150
rect 11716 -11150 11792 -11134
rect 11716 -11167 11732 -11150
rect 11484 -11184 11522 -11167
rect 11402 -11222 11522 -11184
rect 11694 -11184 11732 -11167
rect 11776 -11167 11792 -11150
rect 12008 -11150 12084 -11134
rect 12008 -11167 12024 -11150
rect 11776 -11184 11814 -11167
rect 11694 -11222 11814 -11184
rect 11986 -11184 12024 -11167
rect 12068 -11167 12084 -11150
rect 12300 -11150 12376 -11134
rect 12300 -11167 12316 -11150
rect 12068 -11184 12106 -11167
rect 11986 -11222 12106 -11184
rect 12278 -11184 12316 -11167
rect 12360 -11167 12376 -11150
rect 12592 -11150 12668 -11134
rect 12592 -11167 12608 -11150
rect 12360 -11184 12398 -11167
rect 12278 -11222 12398 -11184
rect 12570 -11184 12608 -11167
rect 12652 -11167 12668 -11150
rect 12652 -11184 12690 -11167
rect 12570 -11222 12690 -11184
rect -2127 -11438 -2007 -11400
rect -5582 -11480 -5462 -11442
rect -5582 -11497 -5544 -11480
rect -5560 -11514 -5544 -11497
rect -5500 -11497 -5462 -11480
rect -5404 -11480 -5284 -11442
rect -5404 -11497 -5366 -11480
rect -5500 -11514 -5484 -11497
rect -5560 -11530 -5484 -11514
rect -5382 -11514 -5366 -11497
rect -5322 -11497 -5284 -11480
rect -5226 -11480 -5106 -11442
rect -5226 -11497 -5188 -11480
rect -5322 -11514 -5306 -11497
rect -5382 -11530 -5306 -11514
rect -5204 -11514 -5188 -11497
rect -5144 -11497 -5106 -11480
rect -5048 -11480 -4928 -11442
rect -5048 -11497 -5010 -11480
rect -5144 -11514 -5128 -11497
rect -5204 -11530 -5128 -11514
rect -5026 -11514 -5010 -11497
rect -4966 -11497 -4928 -11480
rect -4870 -11480 -4750 -11442
rect -4870 -11497 -4832 -11480
rect -4966 -11514 -4950 -11497
rect -5026 -11530 -4950 -11514
rect -4848 -11514 -4832 -11497
rect -4788 -11497 -4750 -11480
rect -4692 -11480 -4572 -11442
rect -4692 -11497 -4654 -11480
rect -4788 -11514 -4772 -11497
rect -4848 -11530 -4772 -11514
rect -4670 -11514 -4654 -11497
rect -4610 -11497 -4572 -11480
rect -4514 -11480 -4394 -11442
rect -4514 -11497 -4476 -11480
rect -4610 -11514 -4594 -11497
rect -4670 -11530 -4594 -11514
rect -4492 -11514 -4476 -11497
rect -4432 -11497 -4394 -11480
rect -4336 -11480 -4216 -11442
rect -4336 -11497 -4298 -11480
rect -4432 -11514 -4416 -11497
rect -4492 -11530 -4416 -11514
rect -4314 -11514 -4298 -11497
rect -4254 -11497 -4216 -11480
rect -4158 -11480 -4038 -11442
rect -2127 -11455 -2089 -11438
rect -4158 -11497 -4120 -11480
rect -4254 -11514 -4238 -11497
rect -4314 -11530 -4238 -11514
rect -4136 -11514 -4120 -11497
rect -4076 -11497 -4038 -11480
rect -2105 -11472 -2089 -11455
rect -2045 -11455 -2007 -11438
rect -1949 -11438 -1829 -11400
rect -1949 -11455 -1911 -11438
rect -2045 -11472 -2029 -11455
rect -2105 -11488 -2029 -11472
rect -1927 -11472 -1911 -11455
rect -1867 -11455 -1829 -11438
rect -1771 -11438 -1651 -11400
rect -1771 -11455 -1733 -11438
rect -1867 -11472 -1851 -11455
rect -1927 -11488 -1851 -11472
rect -1749 -11472 -1733 -11455
rect -1689 -11455 -1651 -11438
rect -1593 -11438 -1473 -11400
rect -1593 -11455 -1555 -11438
rect -1689 -11472 -1673 -11455
rect -1749 -11488 -1673 -11472
rect -1571 -11472 -1555 -11455
rect -1511 -11455 -1473 -11438
rect -1415 -11438 -1295 -11400
rect -1415 -11455 -1377 -11438
rect -1511 -11472 -1495 -11455
rect -1571 -11488 -1495 -11472
rect -1393 -11472 -1377 -11455
rect -1333 -11455 -1295 -11438
rect -1237 -11438 -1117 -11400
rect -1237 -11455 -1199 -11438
rect -1333 -11472 -1317 -11455
rect -1393 -11488 -1317 -11472
rect -1215 -11472 -1199 -11455
rect -1155 -11455 -1117 -11438
rect -1059 -11438 -939 -11400
rect -1059 -11455 -1021 -11438
rect -1155 -11472 -1139 -11455
rect -1215 -11488 -1139 -11472
rect -1037 -11472 -1021 -11455
rect -977 -11455 -939 -11438
rect -881 -11438 -761 -11400
rect -881 -11455 -843 -11438
rect -977 -11472 -961 -11455
rect -1037 -11488 -961 -11472
rect -859 -11472 -843 -11455
rect -799 -11455 -761 -11438
rect -703 -11438 -583 -11400
rect -703 -11455 -665 -11438
rect -799 -11472 -783 -11455
rect -859 -11488 -783 -11472
rect -681 -11472 -665 -11455
rect -621 -11455 -583 -11438
rect -525 -11438 -405 -11400
rect -525 -11455 -487 -11438
rect -621 -11472 -605 -11455
rect -681 -11488 -605 -11472
rect -503 -11472 -487 -11455
rect -443 -11455 -405 -11438
rect -347 -11438 -227 -11400
rect -347 -11455 -309 -11438
rect -443 -11472 -427 -11455
rect -503 -11488 -427 -11472
rect -325 -11472 -309 -11455
rect -265 -11455 -227 -11438
rect -169 -11438 -49 -11400
rect -169 -11455 -131 -11438
rect -265 -11472 -249 -11455
rect -325 -11488 -249 -11472
rect -147 -11472 -131 -11455
rect -87 -11455 -49 -11438
rect 9 -11438 129 -11400
rect 9 -11455 47 -11438
rect -87 -11472 -71 -11455
rect -147 -11488 -71 -11472
rect 31 -11472 47 -11455
rect 91 -11455 129 -11438
rect 187 -11438 307 -11400
rect 187 -11455 225 -11438
rect 91 -11472 107 -11455
rect 31 -11488 107 -11472
rect 209 -11472 225 -11455
rect 269 -11455 307 -11438
rect 365 -11438 485 -11400
rect 365 -11455 403 -11438
rect 269 -11472 285 -11455
rect 209 -11488 285 -11472
rect 387 -11472 403 -11455
rect 447 -11455 485 -11438
rect 543 -11438 663 -11400
rect 543 -11455 581 -11438
rect 447 -11472 463 -11455
rect 387 -11488 463 -11472
rect 565 -11472 581 -11455
rect 625 -11455 663 -11438
rect 721 -11438 841 -11400
rect 721 -11455 759 -11438
rect 625 -11472 641 -11455
rect 565 -11488 641 -11472
rect 743 -11472 759 -11455
rect 803 -11455 841 -11438
rect 899 -11438 1019 -11400
rect 899 -11455 937 -11438
rect 803 -11472 819 -11455
rect 743 -11488 819 -11472
rect 921 -11472 937 -11455
rect 981 -11455 1019 -11438
rect 1077 -11438 1197 -11400
rect 1077 -11455 1115 -11438
rect 981 -11472 997 -11455
rect 921 -11488 997 -11472
rect 1099 -11472 1115 -11455
rect 1159 -11455 1197 -11438
rect 1255 -11438 1375 -11400
rect 1255 -11455 1293 -11438
rect 1159 -11472 1175 -11455
rect 1099 -11488 1175 -11472
rect 1277 -11472 1293 -11455
rect 1337 -11455 1375 -11438
rect 1433 -11438 1553 -11400
rect 1433 -11455 1471 -11438
rect 1337 -11472 1353 -11455
rect 1277 -11488 1353 -11472
rect 1455 -11472 1471 -11455
rect 1515 -11455 1553 -11438
rect 1611 -11438 1731 -11400
rect 1611 -11455 1649 -11438
rect 1515 -11472 1531 -11455
rect 1455 -11488 1531 -11472
rect 1633 -11472 1649 -11455
rect 1693 -11455 1731 -11438
rect 1789 -11438 1909 -11400
rect 1789 -11455 1827 -11438
rect 1693 -11472 1709 -11455
rect 1633 -11488 1709 -11472
rect 1811 -11472 1827 -11455
rect 1871 -11455 1909 -11438
rect 1967 -11438 2087 -11400
rect 1967 -11455 2005 -11438
rect 1871 -11472 1887 -11455
rect 1811 -11488 1887 -11472
rect 1989 -11472 2005 -11455
rect 2049 -11455 2087 -11438
rect 2145 -11438 2265 -11400
rect 2145 -11455 2183 -11438
rect 2049 -11472 2065 -11455
rect 1989 -11488 2065 -11472
rect 2167 -11472 2183 -11455
rect 2227 -11455 2265 -11438
rect 2323 -11438 2443 -11400
rect 2323 -11455 2361 -11438
rect 2227 -11472 2243 -11455
rect 2167 -11488 2243 -11472
rect 2345 -11472 2361 -11455
rect 2405 -11455 2443 -11438
rect 2501 -11438 2621 -11400
rect 2501 -11455 2539 -11438
rect 2405 -11472 2421 -11455
rect 2345 -11488 2421 -11472
rect 2523 -11472 2539 -11455
rect 2583 -11455 2621 -11438
rect 2679 -11438 2799 -11400
rect 2679 -11455 2717 -11438
rect 2583 -11472 2599 -11455
rect 2523 -11488 2599 -11472
rect 2701 -11472 2717 -11455
rect 2761 -11455 2799 -11438
rect 2857 -11438 2977 -11400
rect 2857 -11455 2895 -11438
rect 2761 -11472 2777 -11455
rect 2701 -11488 2777 -11472
rect 2879 -11472 2895 -11455
rect 2939 -11455 2977 -11438
rect 3035 -11438 3155 -11400
rect 3035 -11455 3073 -11438
rect 2939 -11472 2955 -11455
rect 2879 -11488 2955 -11472
rect 3057 -11472 3073 -11455
rect 3117 -11455 3155 -11438
rect 3213 -11438 3333 -11400
rect 3213 -11455 3251 -11438
rect 3117 -11472 3133 -11455
rect 3057 -11488 3133 -11472
rect 3235 -11472 3251 -11455
rect 3295 -11455 3333 -11438
rect 3391 -11438 3511 -11400
rect 3391 -11455 3429 -11438
rect 3295 -11472 3311 -11455
rect 3235 -11488 3311 -11472
rect 3413 -11472 3429 -11455
rect 3473 -11455 3511 -11438
rect 3569 -11438 3689 -11400
rect 3569 -11455 3607 -11438
rect 3473 -11472 3489 -11455
rect 3413 -11488 3489 -11472
rect 3591 -11472 3607 -11455
rect 3651 -11455 3689 -11438
rect 3747 -11438 3867 -11400
rect 3747 -11455 3785 -11438
rect 3651 -11472 3667 -11455
rect 3591 -11488 3667 -11472
rect 3769 -11472 3785 -11455
rect 3829 -11455 3867 -11438
rect 3925 -11438 4045 -11400
rect 3925 -11455 3963 -11438
rect 3829 -11472 3845 -11455
rect 3769 -11488 3845 -11472
rect 3947 -11472 3963 -11455
rect 4007 -11455 4045 -11438
rect 4007 -11472 4023 -11455
rect 3947 -11488 4023 -11472
rect -4076 -11514 -4060 -11497
rect -4136 -11530 -4060 -11514
rect 6580 -11510 6656 -11494
rect 6580 -11527 6596 -11510
rect 6558 -11544 6596 -11527
rect 6640 -11527 6656 -11510
rect 6758 -11510 6834 -11494
rect 6758 -11527 6774 -11510
rect 6640 -11544 6678 -11527
rect 6558 -11582 6678 -11544
rect 6736 -11544 6774 -11527
rect 6818 -11527 6834 -11510
rect 6936 -11510 7012 -11494
rect 6936 -11527 6952 -11510
rect 6818 -11544 6856 -11527
rect 6736 -11582 6856 -11544
rect 6914 -11544 6952 -11527
rect 6996 -11527 7012 -11510
rect 7114 -11510 7190 -11494
rect 7114 -11527 7130 -11510
rect 6996 -11544 7034 -11527
rect 6914 -11582 7034 -11544
rect 7092 -11544 7130 -11527
rect 7174 -11527 7190 -11510
rect 7292 -11510 7368 -11494
rect 7292 -11527 7308 -11510
rect 7174 -11544 7212 -11527
rect 7092 -11582 7212 -11544
rect 7270 -11544 7308 -11527
rect 7352 -11527 7368 -11510
rect 7470 -11510 7546 -11494
rect 7470 -11527 7486 -11510
rect 7352 -11544 7390 -11527
rect 7270 -11582 7390 -11544
rect 7448 -11544 7486 -11527
rect 7530 -11527 7546 -11510
rect 7648 -11510 7724 -11494
rect 7648 -11527 7664 -11510
rect 7530 -11544 7568 -11527
rect 7448 -11582 7568 -11544
rect 7626 -11544 7664 -11527
rect 7708 -11527 7724 -11510
rect 7826 -11510 7902 -11494
rect 7826 -11527 7842 -11510
rect 7708 -11544 7746 -11527
rect 7626 -11582 7746 -11544
rect 7804 -11544 7842 -11527
rect 7886 -11527 7902 -11510
rect 8004 -11510 8080 -11494
rect 8004 -11527 8020 -11510
rect 7886 -11544 7924 -11527
rect 7804 -11582 7924 -11544
rect 7982 -11544 8020 -11527
rect 8064 -11527 8080 -11510
rect 8182 -11510 8258 -11494
rect 8182 -11527 8198 -11510
rect 8064 -11544 8102 -11527
rect 7982 -11582 8102 -11544
rect 8160 -11544 8198 -11527
rect 8242 -11527 8258 -11510
rect 8360 -11510 8436 -11494
rect 8360 -11527 8376 -11510
rect 8242 -11544 8280 -11527
rect 8160 -11582 8280 -11544
rect 8338 -11544 8376 -11527
rect 8420 -11527 8436 -11510
rect 8538 -11510 8614 -11494
rect 8538 -11527 8554 -11510
rect 8420 -11544 8458 -11527
rect 8338 -11582 8458 -11544
rect 8516 -11544 8554 -11527
rect 8598 -11527 8614 -11510
rect 8716 -11510 8792 -11494
rect 8716 -11527 8732 -11510
rect 8598 -11544 8636 -11527
rect 8516 -11582 8636 -11544
rect 8694 -11544 8732 -11527
rect 8776 -11527 8792 -11510
rect 8894 -11510 8970 -11494
rect 8894 -11527 8910 -11510
rect 8776 -11544 8814 -11527
rect 8694 -11582 8814 -11544
rect 8872 -11544 8910 -11527
rect 8954 -11527 8970 -11510
rect 9072 -11510 9148 -11494
rect 9072 -11527 9088 -11510
rect 8954 -11544 8992 -11527
rect 8872 -11582 8992 -11544
rect 9050 -11544 9088 -11527
rect 9132 -11527 9148 -11510
rect 9250 -11510 9326 -11494
rect 9250 -11527 9266 -11510
rect 9132 -11544 9170 -11527
rect 9050 -11582 9170 -11544
rect 9228 -11544 9266 -11527
rect 9310 -11527 9326 -11510
rect 9310 -11544 9348 -11527
rect 9228 -11582 9348 -11544
rect 10818 -11540 10938 -11502
rect 10818 -11557 10856 -11540
rect 10840 -11574 10856 -11557
rect 10900 -11557 10938 -11540
rect 11110 -11540 11230 -11502
rect 11110 -11557 11148 -11540
rect 10900 -11574 10916 -11557
rect -5560 -11640 -5484 -11624
rect -5560 -11657 -5544 -11640
rect -5582 -11674 -5544 -11657
rect -5500 -11657 -5484 -11640
rect -5382 -11640 -5306 -11624
rect -5382 -11657 -5366 -11640
rect -5500 -11674 -5462 -11657
rect -5582 -11712 -5462 -11674
rect -5404 -11674 -5366 -11657
rect -5322 -11657 -5306 -11640
rect -5204 -11640 -5128 -11624
rect -5204 -11657 -5188 -11640
rect -5322 -11674 -5284 -11657
rect -5404 -11712 -5284 -11674
rect -5226 -11674 -5188 -11657
rect -5144 -11657 -5128 -11640
rect -5026 -11640 -4950 -11624
rect -5026 -11657 -5010 -11640
rect -5144 -11674 -5106 -11657
rect -5226 -11712 -5106 -11674
rect -5048 -11674 -5010 -11657
rect -4966 -11657 -4950 -11640
rect -4848 -11640 -4772 -11624
rect -4848 -11657 -4832 -11640
rect -4966 -11674 -4928 -11657
rect -5048 -11712 -4928 -11674
rect -4870 -11674 -4832 -11657
rect -4788 -11657 -4772 -11640
rect -4670 -11640 -4594 -11624
rect -4670 -11657 -4654 -11640
rect -4788 -11674 -4750 -11657
rect -4870 -11712 -4750 -11674
rect -4692 -11674 -4654 -11657
rect -4610 -11657 -4594 -11640
rect -4492 -11640 -4416 -11624
rect -4492 -11657 -4476 -11640
rect -4610 -11674 -4572 -11657
rect -4692 -11712 -4572 -11674
rect -4514 -11674 -4476 -11657
rect -4432 -11657 -4416 -11640
rect -4314 -11640 -4238 -11624
rect -4314 -11657 -4298 -11640
rect -4432 -11674 -4394 -11657
rect -4514 -11712 -4394 -11674
rect -4336 -11674 -4298 -11657
rect -4254 -11657 -4238 -11640
rect -4136 -11640 -4060 -11624
rect -4136 -11657 -4120 -11640
rect -4254 -11674 -4216 -11657
rect -4336 -11712 -4216 -11674
rect -4158 -11674 -4120 -11657
rect -4076 -11657 -4060 -11640
rect -4076 -11674 -4038 -11657
rect -4158 -11712 -4038 -11674
rect 10840 -11590 10916 -11574
rect 11132 -11574 11148 -11557
rect 11192 -11557 11230 -11540
rect 11402 -11540 11522 -11502
rect 11402 -11557 11440 -11540
rect 11192 -11574 11208 -11557
rect 11132 -11590 11208 -11574
rect 11424 -11574 11440 -11557
rect 11484 -11557 11522 -11540
rect 11694 -11540 11814 -11502
rect 11694 -11557 11732 -11540
rect 11484 -11574 11500 -11557
rect 11424 -11590 11500 -11574
rect 11716 -11574 11732 -11557
rect 11776 -11557 11814 -11540
rect 11986 -11540 12106 -11502
rect 11986 -11557 12024 -11540
rect 11776 -11574 11792 -11557
rect 11716 -11590 11792 -11574
rect 12008 -11574 12024 -11557
rect 12068 -11557 12106 -11540
rect 12278 -11540 12398 -11502
rect 12278 -11557 12316 -11540
rect 12068 -11574 12084 -11557
rect 12008 -11590 12084 -11574
rect 12300 -11574 12316 -11557
rect 12360 -11557 12398 -11540
rect 12570 -11540 12690 -11502
rect 12570 -11557 12608 -11540
rect 12360 -11574 12376 -11557
rect 12300 -11590 12376 -11574
rect 12592 -11574 12608 -11557
rect 12652 -11557 12690 -11540
rect 12652 -11574 12668 -11557
rect 12592 -11590 12668 -11574
rect 6558 -11900 6678 -11862
rect 6558 -11917 6596 -11900
rect 6580 -11934 6596 -11917
rect 6640 -11917 6678 -11900
rect 6736 -11900 6856 -11862
rect 6736 -11917 6774 -11900
rect 6640 -11934 6656 -11917
rect 6580 -11950 6656 -11934
rect 6758 -11934 6774 -11917
rect 6818 -11917 6856 -11900
rect 6914 -11900 7034 -11862
rect 6914 -11917 6952 -11900
rect 6818 -11934 6834 -11917
rect 6758 -11950 6834 -11934
rect 6936 -11934 6952 -11917
rect 6996 -11917 7034 -11900
rect 7092 -11900 7212 -11862
rect 7092 -11917 7130 -11900
rect 6996 -11934 7012 -11917
rect 6936 -11950 7012 -11934
rect 7114 -11934 7130 -11917
rect 7174 -11917 7212 -11900
rect 7270 -11900 7390 -11862
rect 7270 -11917 7308 -11900
rect 7174 -11934 7190 -11917
rect 7114 -11950 7190 -11934
rect 7292 -11934 7308 -11917
rect 7352 -11917 7390 -11900
rect 7448 -11900 7568 -11862
rect 7448 -11917 7486 -11900
rect 7352 -11934 7368 -11917
rect 7292 -11950 7368 -11934
rect 7470 -11934 7486 -11917
rect 7530 -11917 7568 -11900
rect 7626 -11900 7746 -11862
rect 7626 -11917 7664 -11900
rect 7530 -11934 7546 -11917
rect 7470 -11950 7546 -11934
rect 7648 -11934 7664 -11917
rect 7708 -11917 7746 -11900
rect 7804 -11900 7924 -11862
rect 7804 -11917 7842 -11900
rect 7708 -11934 7724 -11917
rect 7648 -11950 7724 -11934
rect 7826 -11934 7842 -11917
rect 7886 -11917 7924 -11900
rect 7982 -11900 8102 -11862
rect 7982 -11917 8020 -11900
rect 7886 -11934 7902 -11917
rect 7826 -11950 7902 -11934
rect 8004 -11934 8020 -11917
rect 8064 -11917 8102 -11900
rect 8160 -11900 8280 -11862
rect 8160 -11917 8198 -11900
rect 8064 -11934 8080 -11917
rect 8004 -11950 8080 -11934
rect 8182 -11934 8198 -11917
rect 8242 -11917 8280 -11900
rect 8338 -11900 8458 -11862
rect 8338 -11917 8376 -11900
rect 8242 -11934 8258 -11917
rect 8182 -11950 8258 -11934
rect 8360 -11934 8376 -11917
rect 8420 -11917 8458 -11900
rect 8516 -11900 8636 -11862
rect 8516 -11917 8554 -11900
rect 8420 -11934 8436 -11917
rect 8360 -11950 8436 -11934
rect 8538 -11934 8554 -11917
rect 8598 -11917 8636 -11900
rect 8694 -11900 8814 -11862
rect 8694 -11917 8732 -11900
rect 8598 -11934 8614 -11917
rect 8538 -11950 8614 -11934
rect 8716 -11934 8732 -11917
rect 8776 -11917 8814 -11900
rect 8872 -11900 8992 -11862
rect 8872 -11917 8910 -11900
rect 8776 -11934 8792 -11917
rect 8716 -11950 8792 -11934
rect 8894 -11934 8910 -11917
rect 8954 -11917 8992 -11900
rect 9050 -11900 9170 -11862
rect 9050 -11917 9088 -11900
rect 8954 -11934 8970 -11917
rect 8894 -11950 8970 -11934
rect 9072 -11934 9088 -11917
rect 9132 -11917 9170 -11900
rect 9228 -11900 9348 -11862
rect 9228 -11917 9266 -11900
rect 9132 -11934 9148 -11917
rect 9072 -11950 9148 -11934
rect 9250 -11934 9266 -11917
rect 9310 -11917 9348 -11900
rect 9310 -11934 9326 -11917
rect 9250 -11950 9326 -11934
rect -5582 -12030 -5462 -11992
rect -5582 -12047 -5544 -12030
rect -5560 -12064 -5544 -12047
rect -5500 -12047 -5462 -12030
rect -5404 -12030 -5284 -11992
rect -5404 -12047 -5366 -12030
rect -5500 -12064 -5484 -12047
rect -5560 -12080 -5484 -12064
rect -5382 -12064 -5366 -12047
rect -5322 -12047 -5284 -12030
rect -5226 -12030 -5106 -11992
rect -5226 -12047 -5188 -12030
rect -5322 -12064 -5306 -12047
rect -5382 -12080 -5306 -12064
rect -5204 -12064 -5188 -12047
rect -5144 -12047 -5106 -12030
rect -5048 -12030 -4928 -11992
rect -5048 -12047 -5010 -12030
rect -5144 -12064 -5128 -12047
rect -5204 -12080 -5128 -12064
rect -5026 -12064 -5010 -12047
rect -4966 -12047 -4928 -12030
rect -4870 -12030 -4750 -11992
rect -4870 -12047 -4832 -12030
rect -4966 -12064 -4950 -12047
rect -5026 -12080 -4950 -12064
rect -4848 -12064 -4832 -12047
rect -4788 -12047 -4750 -12030
rect -4692 -12030 -4572 -11992
rect -4692 -12047 -4654 -12030
rect -4788 -12064 -4772 -12047
rect -4848 -12080 -4772 -12064
rect -4670 -12064 -4654 -12047
rect -4610 -12047 -4572 -12030
rect -4514 -12030 -4394 -11992
rect -4514 -12047 -4476 -12030
rect -4610 -12064 -4594 -12047
rect -4670 -12080 -4594 -12064
rect -4492 -12064 -4476 -12047
rect -4432 -12047 -4394 -12030
rect -4336 -12030 -4216 -11992
rect -4336 -12047 -4298 -12030
rect -4432 -12064 -4416 -12047
rect -4492 -12080 -4416 -12064
rect -4314 -12064 -4298 -12047
rect -4254 -12047 -4216 -12030
rect -4158 -12030 -4038 -11992
rect -4158 -12047 -4120 -12030
rect -4254 -12064 -4238 -12047
rect -4314 -12080 -4238 -12064
rect -4136 -12064 -4120 -12047
rect -4076 -12047 -4038 -12030
rect -4076 -12064 -4060 -12047
rect -4136 -12080 -4060 -12064
rect -2105 -12048 -2029 -12032
rect -2105 -12065 -2089 -12048
rect -2127 -12082 -2089 -12065
rect -2045 -12065 -2029 -12048
rect -1927 -12048 -1851 -12032
rect -1927 -12065 -1911 -12048
rect -2045 -12082 -2007 -12065
rect -2127 -12120 -2007 -12082
rect -1949 -12082 -1911 -12065
rect -1867 -12065 -1851 -12048
rect -1749 -12048 -1673 -12032
rect -1749 -12065 -1733 -12048
rect -1867 -12082 -1829 -12065
rect -1949 -12120 -1829 -12082
rect -1771 -12082 -1733 -12065
rect -1689 -12065 -1673 -12048
rect -1571 -12048 -1495 -12032
rect -1571 -12065 -1555 -12048
rect -1689 -12082 -1651 -12065
rect -1771 -12120 -1651 -12082
rect -1593 -12082 -1555 -12065
rect -1511 -12065 -1495 -12048
rect -1393 -12048 -1317 -12032
rect -1393 -12065 -1377 -12048
rect -1511 -12082 -1473 -12065
rect -1593 -12120 -1473 -12082
rect -1415 -12082 -1377 -12065
rect -1333 -12065 -1317 -12048
rect -1215 -12048 -1139 -12032
rect -1215 -12065 -1199 -12048
rect -1333 -12082 -1295 -12065
rect -1415 -12120 -1295 -12082
rect -1237 -12082 -1199 -12065
rect -1155 -12065 -1139 -12048
rect -1037 -12048 -961 -12032
rect -1037 -12065 -1021 -12048
rect -1155 -12082 -1117 -12065
rect -1237 -12120 -1117 -12082
rect -1059 -12082 -1021 -12065
rect -977 -12065 -961 -12048
rect -859 -12048 -783 -12032
rect -859 -12065 -843 -12048
rect -977 -12082 -939 -12065
rect -1059 -12120 -939 -12082
rect -881 -12082 -843 -12065
rect -799 -12065 -783 -12048
rect -681 -12048 -605 -12032
rect -681 -12065 -665 -12048
rect -799 -12082 -761 -12065
rect -881 -12120 -761 -12082
rect -703 -12082 -665 -12065
rect -621 -12065 -605 -12048
rect -503 -12048 -427 -12032
rect -503 -12065 -487 -12048
rect -621 -12082 -583 -12065
rect -703 -12120 -583 -12082
rect -525 -12082 -487 -12065
rect -443 -12065 -427 -12048
rect -325 -12048 -249 -12032
rect -325 -12065 -309 -12048
rect -443 -12082 -405 -12065
rect -525 -12120 -405 -12082
rect -347 -12082 -309 -12065
rect -265 -12065 -249 -12048
rect -147 -12048 -71 -12032
rect -147 -12065 -131 -12048
rect -265 -12082 -227 -12065
rect -347 -12120 -227 -12082
rect -169 -12082 -131 -12065
rect -87 -12065 -71 -12048
rect 31 -12048 107 -12032
rect 31 -12065 47 -12048
rect -87 -12082 -49 -12065
rect -169 -12120 -49 -12082
rect 9 -12082 47 -12065
rect 91 -12065 107 -12048
rect 209 -12048 285 -12032
rect 209 -12065 225 -12048
rect 91 -12082 129 -12065
rect 9 -12120 129 -12082
rect 187 -12082 225 -12065
rect 269 -12065 285 -12048
rect 387 -12048 463 -12032
rect 387 -12065 403 -12048
rect 269 -12082 307 -12065
rect 187 -12120 307 -12082
rect 365 -12082 403 -12065
rect 447 -12065 463 -12048
rect 565 -12048 641 -12032
rect 565 -12065 581 -12048
rect 447 -12082 485 -12065
rect 365 -12120 485 -12082
rect 543 -12082 581 -12065
rect 625 -12065 641 -12048
rect 743 -12048 819 -12032
rect 743 -12065 759 -12048
rect 625 -12082 663 -12065
rect 543 -12120 663 -12082
rect 721 -12082 759 -12065
rect 803 -12065 819 -12048
rect 921 -12048 997 -12032
rect 921 -12065 937 -12048
rect 803 -12082 841 -12065
rect 721 -12120 841 -12082
rect 899 -12082 937 -12065
rect 981 -12065 997 -12048
rect 1099 -12048 1175 -12032
rect 1099 -12065 1115 -12048
rect 981 -12082 1019 -12065
rect 899 -12120 1019 -12082
rect 1077 -12082 1115 -12065
rect 1159 -12065 1175 -12048
rect 1277 -12048 1353 -12032
rect 1277 -12065 1293 -12048
rect 1159 -12082 1197 -12065
rect 1077 -12120 1197 -12082
rect 1255 -12082 1293 -12065
rect 1337 -12065 1353 -12048
rect 1455 -12048 1531 -12032
rect 1455 -12065 1471 -12048
rect 1337 -12082 1375 -12065
rect 1255 -12120 1375 -12082
rect 1433 -12082 1471 -12065
rect 1515 -12065 1531 -12048
rect 1633 -12048 1709 -12032
rect 1633 -12065 1649 -12048
rect 1515 -12082 1553 -12065
rect 1433 -12120 1553 -12082
rect 1611 -12082 1649 -12065
rect 1693 -12065 1709 -12048
rect 1811 -12048 1887 -12032
rect 1811 -12065 1827 -12048
rect 1693 -12082 1731 -12065
rect 1611 -12120 1731 -12082
rect 1789 -12082 1827 -12065
rect 1871 -12065 1887 -12048
rect 1989 -12048 2065 -12032
rect 1989 -12065 2005 -12048
rect 1871 -12082 1909 -12065
rect 1789 -12120 1909 -12082
rect 1967 -12082 2005 -12065
rect 2049 -12065 2065 -12048
rect 2167 -12048 2243 -12032
rect 2167 -12065 2183 -12048
rect 2049 -12082 2087 -12065
rect 1967 -12120 2087 -12082
rect 2145 -12082 2183 -12065
rect 2227 -12065 2243 -12048
rect 2345 -12048 2421 -12032
rect 2345 -12065 2361 -12048
rect 2227 -12082 2265 -12065
rect 2145 -12120 2265 -12082
rect 2323 -12082 2361 -12065
rect 2405 -12065 2421 -12048
rect 2523 -12048 2599 -12032
rect 2523 -12065 2539 -12048
rect 2405 -12082 2443 -12065
rect 2323 -12120 2443 -12082
rect 2501 -12082 2539 -12065
rect 2583 -12065 2599 -12048
rect 2701 -12048 2777 -12032
rect 2701 -12065 2717 -12048
rect 2583 -12082 2621 -12065
rect 2501 -12120 2621 -12082
rect 2679 -12082 2717 -12065
rect 2761 -12065 2777 -12048
rect 2879 -12048 2955 -12032
rect 2879 -12065 2895 -12048
rect 2761 -12082 2799 -12065
rect 2679 -12120 2799 -12082
rect 2857 -12082 2895 -12065
rect 2939 -12065 2955 -12048
rect 3057 -12048 3133 -12032
rect 3057 -12065 3073 -12048
rect 2939 -12082 2977 -12065
rect 2857 -12120 2977 -12082
rect 3035 -12082 3073 -12065
rect 3117 -12065 3133 -12048
rect 3235 -12048 3311 -12032
rect 3235 -12065 3251 -12048
rect 3117 -12082 3155 -12065
rect 3035 -12120 3155 -12082
rect 3213 -12082 3251 -12065
rect 3295 -12065 3311 -12048
rect 3413 -12048 3489 -12032
rect 3413 -12065 3429 -12048
rect 3295 -12082 3333 -12065
rect 3213 -12120 3333 -12082
rect 3391 -12082 3429 -12065
rect 3473 -12065 3489 -12048
rect 3591 -12048 3667 -12032
rect 3591 -12065 3607 -12048
rect 3473 -12082 3511 -12065
rect 3391 -12120 3511 -12082
rect 3569 -12082 3607 -12065
rect 3651 -12065 3667 -12048
rect 3769 -12048 3845 -12032
rect 3769 -12065 3785 -12048
rect 3651 -12082 3689 -12065
rect 3569 -12120 3689 -12082
rect 3747 -12082 3785 -12065
rect 3829 -12065 3845 -12048
rect 3947 -12048 4023 -12032
rect 3947 -12065 3963 -12048
rect 3829 -12082 3867 -12065
rect 3747 -12120 3867 -12082
rect 3925 -12082 3963 -12065
rect 4007 -12065 4023 -12048
rect 4007 -12082 4045 -12065
rect 3925 -12120 4045 -12082
rect -2127 -12438 -2007 -12400
rect -2127 -12455 -2089 -12438
rect -2105 -12472 -2089 -12455
rect -2045 -12455 -2007 -12438
rect -1949 -12438 -1829 -12400
rect -1949 -12455 -1911 -12438
rect -2045 -12472 -2029 -12455
rect -2105 -12488 -2029 -12472
rect -1927 -12472 -1911 -12455
rect -1867 -12455 -1829 -12438
rect -1771 -12438 -1651 -12400
rect -1771 -12455 -1733 -12438
rect -1867 -12472 -1851 -12455
rect -1927 -12488 -1851 -12472
rect -1749 -12472 -1733 -12455
rect -1689 -12455 -1651 -12438
rect -1593 -12438 -1473 -12400
rect -1593 -12455 -1555 -12438
rect -1689 -12472 -1673 -12455
rect -1749 -12488 -1673 -12472
rect -1571 -12472 -1555 -12455
rect -1511 -12455 -1473 -12438
rect -1415 -12438 -1295 -12400
rect -1415 -12455 -1377 -12438
rect -1511 -12472 -1495 -12455
rect -1571 -12488 -1495 -12472
rect -1393 -12472 -1377 -12455
rect -1333 -12455 -1295 -12438
rect -1237 -12438 -1117 -12400
rect -1237 -12455 -1199 -12438
rect -1333 -12472 -1317 -12455
rect -1393 -12488 -1317 -12472
rect -1215 -12472 -1199 -12455
rect -1155 -12455 -1117 -12438
rect -1059 -12438 -939 -12400
rect -1059 -12455 -1021 -12438
rect -1155 -12472 -1139 -12455
rect -1215 -12488 -1139 -12472
rect -1037 -12472 -1021 -12455
rect -977 -12455 -939 -12438
rect -881 -12438 -761 -12400
rect -881 -12455 -843 -12438
rect -977 -12472 -961 -12455
rect -1037 -12488 -961 -12472
rect -859 -12472 -843 -12455
rect -799 -12455 -761 -12438
rect -703 -12438 -583 -12400
rect -703 -12455 -665 -12438
rect -799 -12472 -783 -12455
rect -859 -12488 -783 -12472
rect -681 -12472 -665 -12455
rect -621 -12455 -583 -12438
rect -525 -12438 -405 -12400
rect -525 -12455 -487 -12438
rect -621 -12472 -605 -12455
rect -681 -12488 -605 -12472
rect -503 -12472 -487 -12455
rect -443 -12455 -405 -12438
rect -347 -12438 -227 -12400
rect -347 -12455 -309 -12438
rect -443 -12472 -427 -12455
rect -503 -12488 -427 -12472
rect -325 -12472 -309 -12455
rect -265 -12455 -227 -12438
rect -169 -12438 -49 -12400
rect -169 -12455 -131 -12438
rect -265 -12472 -249 -12455
rect -325 -12488 -249 -12472
rect -147 -12472 -131 -12455
rect -87 -12455 -49 -12438
rect 9 -12438 129 -12400
rect 9 -12455 47 -12438
rect -87 -12472 -71 -12455
rect -147 -12488 -71 -12472
rect 31 -12472 47 -12455
rect 91 -12455 129 -12438
rect 187 -12438 307 -12400
rect 187 -12455 225 -12438
rect 91 -12472 107 -12455
rect 31 -12488 107 -12472
rect 209 -12472 225 -12455
rect 269 -12455 307 -12438
rect 365 -12438 485 -12400
rect 365 -12455 403 -12438
rect 269 -12472 285 -12455
rect 209 -12488 285 -12472
rect 387 -12472 403 -12455
rect 447 -12455 485 -12438
rect 543 -12438 663 -12400
rect 543 -12455 581 -12438
rect 447 -12472 463 -12455
rect 387 -12488 463 -12472
rect 565 -12472 581 -12455
rect 625 -12455 663 -12438
rect 721 -12438 841 -12400
rect 721 -12455 759 -12438
rect 625 -12472 641 -12455
rect 565 -12488 641 -12472
rect 743 -12472 759 -12455
rect 803 -12455 841 -12438
rect 899 -12438 1019 -12400
rect 899 -12455 937 -12438
rect 803 -12472 819 -12455
rect 743 -12488 819 -12472
rect 921 -12472 937 -12455
rect 981 -12455 1019 -12438
rect 1077 -12438 1197 -12400
rect 1077 -12455 1115 -12438
rect 981 -12472 997 -12455
rect 921 -12488 997 -12472
rect 1099 -12472 1115 -12455
rect 1159 -12455 1197 -12438
rect 1255 -12438 1375 -12400
rect 1255 -12455 1293 -12438
rect 1159 -12472 1175 -12455
rect 1099 -12488 1175 -12472
rect 1277 -12472 1293 -12455
rect 1337 -12455 1375 -12438
rect 1433 -12438 1553 -12400
rect 1433 -12455 1471 -12438
rect 1337 -12472 1353 -12455
rect 1277 -12488 1353 -12472
rect 1455 -12472 1471 -12455
rect 1515 -12455 1553 -12438
rect 1611 -12438 1731 -12400
rect 1611 -12455 1649 -12438
rect 1515 -12472 1531 -12455
rect 1455 -12488 1531 -12472
rect 1633 -12472 1649 -12455
rect 1693 -12455 1731 -12438
rect 1789 -12438 1909 -12400
rect 1789 -12455 1827 -12438
rect 1693 -12472 1709 -12455
rect 1633 -12488 1709 -12472
rect 1811 -12472 1827 -12455
rect 1871 -12455 1909 -12438
rect 1967 -12438 2087 -12400
rect 1967 -12455 2005 -12438
rect 1871 -12472 1887 -12455
rect 1811 -12488 1887 -12472
rect 1989 -12472 2005 -12455
rect 2049 -12455 2087 -12438
rect 2145 -12438 2265 -12400
rect 2145 -12455 2183 -12438
rect 2049 -12472 2065 -12455
rect 1989 -12488 2065 -12472
rect 2167 -12472 2183 -12455
rect 2227 -12455 2265 -12438
rect 2323 -12438 2443 -12400
rect 2323 -12455 2361 -12438
rect 2227 -12472 2243 -12455
rect 2167 -12488 2243 -12472
rect 2345 -12472 2361 -12455
rect 2405 -12455 2443 -12438
rect 2501 -12438 2621 -12400
rect 2501 -12455 2539 -12438
rect 2405 -12472 2421 -12455
rect 2345 -12488 2421 -12472
rect 2523 -12472 2539 -12455
rect 2583 -12455 2621 -12438
rect 2679 -12438 2799 -12400
rect 2679 -12455 2717 -12438
rect 2583 -12472 2599 -12455
rect 2523 -12488 2599 -12472
rect 2701 -12472 2717 -12455
rect 2761 -12455 2799 -12438
rect 2857 -12438 2977 -12400
rect 2857 -12455 2895 -12438
rect 2761 -12472 2777 -12455
rect 2701 -12488 2777 -12472
rect 2879 -12472 2895 -12455
rect 2939 -12455 2977 -12438
rect 3035 -12438 3155 -12400
rect 3035 -12455 3073 -12438
rect 2939 -12472 2955 -12455
rect 2879 -12488 2955 -12472
rect 3057 -12472 3073 -12455
rect 3117 -12455 3155 -12438
rect 3213 -12438 3333 -12400
rect 3213 -12455 3251 -12438
rect 3117 -12472 3133 -12455
rect 3057 -12488 3133 -12472
rect 3235 -12472 3251 -12455
rect 3295 -12455 3333 -12438
rect 3391 -12438 3511 -12400
rect 3391 -12455 3429 -12438
rect 3295 -12472 3311 -12455
rect 3235 -12488 3311 -12472
rect 3413 -12472 3429 -12455
rect 3473 -12455 3511 -12438
rect 3569 -12438 3689 -12400
rect 3569 -12455 3607 -12438
rect 3473 -12472 3489 -12455
rect 3413 -12488 3489 -12472
rect 3591 -12472 3607 -12455
rect 3651 -12455 3689 -12438
rect 3747 -12438 3867 -12400
rect 3747 -12455 3785 -12438
rect 3651 -12472 3667 -12455
rect 3591 -12488 3667 -12472
rect 3769 -12472 3785 -12455
rect 3829 -12455 3867 -12438
rect 3925 -12438 4045 -12400
rect 3925 -12455 3963 -12438
rect 3829 -12472 3845 -12455
rect 3769 -12488 3845 -12472
rect 3947 -12472 3963 -12455
rect 4007 -12455 4045 -12438
rect 4007 -12472 4023 -12455
rect 3947 -12488 4023 -12472
rect -5883 -12628 -5817 -12612
rect -5883 -12662 -5867 -12628
rect -5833 -12662 -5817 -12628
rect -5883 -12678 -5817 -12662
rect -5633 -12628 -5567 -12612
rect -5633 -12662 -5617 -12628
rect -5583 -12662 -5567 -12628
rect -5633 -12678 -5567 -12662
rect -5383 -12628 -5317 -12612
rect -5383 -12662 -5367 -12628
rect -5333 -12662 -5317 -12628
rect -5383 -12678 -5317 -12662
rect -5133 -12628 -5067 -12612
rect -5133 -12662 -5117 -12628
rect -5083 -12662 -5067 -12628
rect -5133 -12678 -5067 -12662
rect -4883 -12628 -4817 -12612
rect -4883 -12662 -4867 -12628
rect -4833 -12662 -4817 -12628
rect -4883 -12678 -4817 -12662
rect -4633 -12628 -4567 -12612
rect -4633 -12662 -4617 -12628
rect -4583 -12662 -4567 -12628
rect -4633 -12678 -4567 -12662
rect -4383 -12628 -4317 -12612
rect -4383 -12662 -4367 -12628
rect -4333 -12662 -4317 -12628
rect -4383 -12678 -4317 -12662
rect -4133 -12628 -4067 -12612
rect -4133 -12662 -4117 -12628
rect -4083 -12662 -4067 -12628
rect -4133 -12678 -4067 -12662
rect -5870 -12700 -5830 -12678
rect -5620 -12700 -5580 -12678
rect -5370 -12700 -5330 -12678
rect -5120 -12700 -5080 -12678
rect -4870 -12700 -4830 -12678
rect -4620 -12700 -4580 -12678
rect -4370 -12700 -4330 -12678
rect -4120 -12700 -4080 -12678
rect -5870 -12962 -5830 -12940
rect -5620 -12962 -5580 -12940
rect -5370 -12962 -5330 -12940
rect -5120 -12962 -5080 -12940
rect -4870 -12962 -4830 -12940
rect -4620 -12962 -4580 -12940
rect -4370 -12962 -4330 -12940
rect -4120 -12962 -4080 -12940
rect -5883 -12978 -5817 -12962
rect -5883 -13012 -5867 -12978
rect -5833 -13012 -5817 -12978
rect -5883 -13028 -5817 -13012
rect -5633 -12978 -5567 -12962
rect -5633 -13012 -5617 -12978
rect -5583 -13012 -5567 -12978
rect -5633 -13028 -5567 -13012
rect -5383 -12978 -5317 -12962
rect -5383 -13012 -5367 -12978
rect -5333 -13012 -5317 -12978
rect -5383 -13028 -5317 -13012
rect -5133 -12978 -5067 -12962
rect -5133 -13012 -5117 -12978
rect -5083 -13012 -5067 -12978
rect -5133 -13028 -5067 -13012
rect -4883 -12978 -4817 -12962
rect -4883 -13012 -4867 -12978
rect -4833 -13012 -4817 -12978
rect -4883 -13028 -4817 -13012
rect -4633 -12978 -4567 -12962
rect -4633 -13012 -4617 -12978
rect -4583 -13012 -4567 -12978
rect -4633 -13028 -4567 -13012
rect -4383 -12978 -4317 -12962
rect -4383 -13012 -4367 -12978
rect -4333 -13012 -4317 -12978
rect -4383 -13028 -4317 -13012
rect -4133 -12978 -4067 -12962
rect -4133 -13012 -4117 -12978
rect -4083 -13012 -4067 -12978
rect -4133 -13028 -4067 -13012
rect -2105 -13048 -2029 -13032
rect -2105 -13065 -2089 -13048
rect -2127 -13082 -2089 -13065
rect -2045 -13065 -2029 -13048
rect -1927 -13048 -1851 -13032
rect -1927 -13065 -1911 -13048
rect -2045 -13082 -2007 -13065
rect -2127 -13120 -2007 -13082
rect -1949 -13082 -1911 -13065
rect -1867 -13065 -1851 -13048
rect -1749 -13048 -1673 -13032
rect -1749 -13065 -1733 -13048
rect -1867 -13082 -1829 -13065
rect -1949 -13120 -1829 -13082
rect -1771 -13082 -1733 -13065
rect -1689 -13065 -1673 -13048
rect -1571 -13048 -1495 -13032
rect -1571 -13065 -1555 -13048
rect -1689 -13082 -1651 -13065
rect -1771 -13120 -1651 -13082
rect -1593 -13082 -1555 -13065
rect -1511 -13065 -1495 -13048
rect -1393 -13048 -1317 -13032
rect -1393 -13065 -1377 -13048
rect -1511 -13082 -1473 -13065
rect -1593 -13120 -1473 -13082
rect -1415 -13082 -1377 -13065
rect -1333 -13065 -1317 -13048
rect -1215 -13048 -1139 -13032
rect -1215 -13065 -1199 -13048
rect -1333 -13082 -1295 -13065
rect -1415 -13120 -1295 -13082
rect -1237 -13082 -1199 -13065
rect -1155 -13065 -1139 -13048
rect -1037 -13048 -961 -13032
rect -1037 -13065 -1021 -13048
rect -1155 -13082 -1117 -13065
rect -1237 -13120 -1117 -13082
rect -1059 -13082 -1021 -13065
rect -977 -13065 -961 -13048
rect -859 -13048 -783 -13032
rect -859 -13065 -843 -13048
rect -977 -13082 -939 -13065
rect -1059 -13120 -939 -13082
rect -881 -13082 -843 -13065
rect -799 -13065 -783 -13048
rect -681 -13048 -605 -13032
rect -681 -13065 -665 -13048
rect -799 -13082 -761 -13065
rect -881 -13120 -761 -13082
rect -703 -13082 -665 -13065
rect -621 -13065 -605 -13048
rect -503 -13048 -427 -13032
rect -503 -13065 -487 -13048
rect -621 -13082 -583 -13065
rect -703 -13120 -583 -13082
rect -525 -13082 -487 -13065
rect -443 -13065 -427 -13048
rect -325 -13048 -249 -13032
rect -325 -13065 -309 -13048
rect -443 -13082 -405 -13065
rect -525 -13120 -405 -13082
rect -347 -13082 -309 -13065
rect -265 -13065 -249 -13048
rect -147 -13048 -71 -13032
rect -147 -13065 -131 -13048
rect -265 -13082 -227 -13065
rect -347 -13120 -227 -13082
rect -169 -13082 -131 -13065
rect -87 -13065 -71 -13048
rect 31 -13048 107 -13032
rect 31 -13065 47 -13048
rect -87 -13082 -49 -13065
rect -169 -13120 -49 -13082
rect 9 -13082 47 -13065
rect 91 -13065 107 -13048
rect 209 -13048 285 -13032
rect 209 -13065 225 -13048
rect 91 -13082 129 -13065
rect 9 -13120 129 -13082
rect 187 -13082 225 -13065
rect 269 -13065 285 -13048
rect 387 -13048 463 -13032
rect 387 -13065 403 -13048
rect 269 -13082 307 -13065
rect 187 -13120 307 -13082
rect 365 -13082 403 -13065
rect 447 -13065 463 -13048
rect 565 -13048 641 -13032
rect 565 -13065 581 -13048
rect 447 -13082 485 -13065
rect 365 -13120 485 -13082
rect 543 -13082 581 -13065
rect 625 -13065 641 -13048
rect 743 -13048 819 -13032
rect 743 -13065 759 -13048
rect 625 -13082 663 -13065
rect 543 -13120 663 -13082
rect 721 -13082 759 -13065
rect 803 -13065 819 -13048
rect 921 -13048 997 -13032
rect 921 -13065 937 -13048
rect 803 -13082 841 -13065
rect 721 -13120 841 -13082
rect 899 -13082 937 -13065
rect 981 -13065 997 -13048
rect 1099 -13048 1175 -13032
rect 1099 -13065 1115 -13048
rect 981 -13082 1019 -13065
rect 899 -13120 1019 -13082
rect 1077 -13082 1115 -13065
rect 1159 -13065 1175 -13048
rect 1277 -13048 1353 -13032
rect 1277 -13065 1293 -13048
rect 1159 -13082 1197 -13065
rect 1077 -13120 1197 -13082
rect 1255 -13082 1293 -13065
rect 1337 -13065 1353 -13048
rect 1455 -13048 1531 -13032
rect 1455 -13065 1471 -13048
rect 1337 -13082 1375 -13065
rect 1255 -13120 1375 -13082
rect 1433 -13082 1471 -13065
rect 1515 -13065 1531 -13048
rect 1633 -13048 1709 -13032
rect 1633 -13065 1649 -13048
rect 1515 -13082 1553 -13065
rect 1433 -13120 1553 -13082
rect 1611 -13082 1649 -13065
rect 1693 -13065 1709 -13048
rect 1811 -13048 1887 -13032
rect 1811 -13065 1827 -13048
rect 1693 -13082 1731 -13065
rect 1611 -13120 1731 -13082
rect 1789 -13082 1827 -13065
rect 1871 -13065 1887 -13048
rect 1989 -13048 2065 -13032
rect 1989 -13065 2005 -13048
rect 1871 -13082 1909 -13065
rect 1789 -13120 1909 -13082
rect 1967 -13082 2005 -13065
rect 2049 -13065 2065 -13048
rect 2167 -13048 2243 -13032
rect 2167 -13065 2183 -13048
rect 2049 -13082 2087 -13065
rect 1967 -13120 2087 -13082
rect 2145 -13082 2183 -13065
rect 2227 -13065 2243 -13048
rect 2345 -13048 2421 -13032
rect 2345 -13065 2361 -13048
rect 2227 -13082 2265 -13065
rect 2145 -13120 2265 -13082
rect 2323 -13082 2361 -13065
rect 2405 -13065 2421 -13048
rect 2523 -13048 2599 -13032
rect 2523 -13065 2539 -13048
rect 2405 -13082 2443 -13065
rect 2323 -13120 2443 -13082
rect 2501 -13082 2539 -13065
rect 2583 -13065 2599 -13048
rect 2701 -13048 2777 -13032
rect 2701 -13065 2717 -13048
rect 2583 -13082 2621 -13065
rect 2501 -13120 2621 -13082
rect 2679 -13082 2717 -13065
rect 2761 -13065 2777 -13048
rect 2879 -13048 2955 -13032
rect 2879 -13065 2895 -13048
rect 2761 -13082 2799 -13065
rect 2679 -13120 2799 -13082
rect 2857 -13082 2895 -13065
rect 2939 -13065 2955 -13048
rect 3057 -13048 3133 -13032
rect 3057 -13065 3073 -13048
rect 2939 -13082 2977 -13065
rect 2857 -13120 2977 -13082
rect 3035 -13082 3073 -13065
rect 3117 -13065 3133 -13048
rect 3235 -13048 3311 -13032
rect 3235 -13065 3251 -13048
rect 3117 -13082 3155 -13065
rect 3035 -13120 3155 -13082
rect 3213 -13082 3251 -13065
rect 3295 -13065 3311 -13048
rect 3413 -13048 3489 -13032
rect 3413 -13065 3429 -13048
rect 3295 -13082 3333 -13065
rect 3213 -13120 3333 -13082
rect 3391 -13082 3429 -13065
rect 3473 -13065 3489 -13048
rect 3591 -13048 3667 -13032
rect 3591 -13065 3607 -13048
rect 3473 -13082 3511 -13065
rect 3391 -13120 3511 -13082
rect 3569 -13082 3607 -13065
rect 3651 -13065 3667 -13048
rect 3769 -13048 3845 -13032
rect 3769 -13065 3785 -13048
rect 3651 -13082 3689 -13065
rect 3569 -13120 3689 -13082
rect 3747 -13082 3785 -13065
rect 3829 -13065 3845 -13048
rect 3947 -13048 4023 -13032
rect 3947 -13065 3963 -13048
rect 3829 -13082 3867 -13065
rect 3747 -13120 3867 -13082
rect 3925 -13082 3963 -13065
rect 4007 -13065 4023 -13048
rect 4007 -13082 4045 -13065
rect 3925 -13120 4045 -13082
rect -5883 -13308 -5817 -13292
rect -5883 -13342 -5867 -13308
rect -5833 -13342 -5817 -13308
rect -5883 -13358 -5817 -13342
rect -5633 -13308 -5567 -13292
rect -5633 -13342 -5617 -13308
rect -5583 -13342 -5567 -13308
rect -5633 -13358 -5567 -13342
rect -5383 -13308 -5317 -13292
rect -5383 -13342 -5367 -13308
rect -5333 -13342 -5317 -13308
rect -5383 -13358 -5317 -13342
rect -5133 -13308 -5067 -13292
rect -5133 -13342 -5117 -13308
rect -5083 -13342 -5067 -13308
rect -5133 -13358 -5067 -13342
rect -4883 -13308 -4817 -13292
rect -4883 -13342 -4867 -13308
rect -4833 -13342 -4817 -13308
rect -4883 -13358 -4817 -13342
rect -4633 -13308 -4567 -13292
rect -4633 -13342 -4617 -13308
rect -4583 -13342 -4567 -13308
rect -4633 -13358 -4567 -13342
rect -4383 -13308 -4317 -13292
rect -4383 -13342 -4367 -13308
rect -4333 -13342 -4317 -13308
rect -4383 -13358 -4317 -13342
rect -4133 -13308 -4067 -13292
rect -4133 -13342 -4117 -13308
rect -4083 -13342 -4067 -13308
rect -4133 -13358 -4067 -13342
rect -5870 -13380 -5830 -13358
rect -5620 -13380 -5580 -13358
rect -5370 -13380 -5330 -13358
rect -5120 -13380 -5080 -13358
rect -4870 -13380 -4830 -13358
rect -4620 -13380 -4580 -13358
rect -4370 -13380 -4330 -13358
rect -4120 -13380 -4080 -13358
rect -2127 -13438 -2007 -13400
rect -2127 -13455 -2089 -13438
rect -2105 -13472 -2089 -13455
rect -2045 -13455 -2007 -13438
rect -1949 -13438 -1829 -13400
rect -1949 -13455 -1911 -13438
rect -2045 -13472 -2029 -13455
rect -2105 -13488 -2029 -13472
rect -1927 -13472 -1911 -13455
rect -1867 -13455 -1829 -13438
rect -1771 -13438 -1651 -13400
rect -1771 -13455 -1733 -13438
rect -1867 -13472 -1851 -13455
rect -1927 -13488 -1851 -13472
rect -1749 -13472 -1733 -13455
rect -1689 -13455 -1651 -13438
rect -1593 -13438 -1473 -13400
rect -1593 -13455 -1555 -13438
rect -1689 -13472 -1673 -13455
rect -1749 -13488 -1673 -13472
rect -1571 -13472 -1555 -13455
rect -1511 -13455 -1473 -13438
rect -1415 -13438 -1295 -13400
rect -1415 -13455 -1377 -13438
rect -1511 -13472 -1495 -13455
rect -1571 -13488 -1495 -13472
rect -1393 -13472 -1377 -13455
rect -1333 -13455 -1295 -13438
rect -1237 -13438 -1117 -13400
rect -1237 -13455 -1199 -13438
rect -1333 -13472 -1317 -13455
rect -1393 -13488 -1317 -13472
rect -1215 -13472 -1199 -13455
rect -1155 -13455 -1117 -13438
rect -1059 -13438 -939 -13400
rect -1059 -13455 -1021 -13438
rect -1155 -13472 -1139 -13455
rect -1215 -13488 -1139 -13472
rect -1037 -13472 -1021 -13455
rect -977 -13455 -939 -13438
rect -881 -13438 -761 -13400
rect -881 -13455 -843 -13438
rect -977 -13472 -961 -13455
rect -1037 -13488 -961 -13472
rect -859 -13472 -843 -13455
rect -799 -13455 -761 -13438
rect -703 -13438 -583 -13400
rect -703 -13455 -665 -13438
rect -799 -13472 -783 -13455
rect -859 -13488 -783 -13472
rect -681 -13472 -665 -13455
rect -621 -13455 -583 -13438
rect -525 -13438 -405 -13400
rect -525 -13455 -487 -13438
rect -621 -13472 -605 -13455
rect -681 -13488 -605 -13472
rect -503 -13472 -487 -13455
rect -443 -13455 -405 -13438
rect -347 -13438 -227 -13400
rect -347 -13455 -309 -13438
rect -443 -13472 -427 -13455
rect -503 -13488 -427 -13472
rect -325 -13472 -309 -13455
rect -265 -13455 -227 -13438
rect -169 -13438 -49 -13400
rect -169 -13455 -131 -13438
rect -265 -13472 -249 -13455
rect -325 -13488 -249 -13472
rect -147 -13472 -131 -13455
rect -87 -13455 -49 -13438
rect 9 -13438 129 -13400
rect 9 -13455 47 -13438
rect -87 -13472 -71 -13455
rect -147 -13488 -71 -13472
rect 31 -13472 47 -13455
rect 91 -13455 129 -13438
rect 187 -13438 307 -13400
rect 187 -13455 225 -13438
rect 91 -13472 107 -13455
rect 31 -13488 107 -13472
rect 209 -13472 225 -13455
rect 269 -13455 307 -13438
rect 365 -13438 485 -13400
rect 365 -13455 403 -13438
rect 269 -13472 285 -13455
rect 209 -13488 285 -13472
rect 387 -13472 403 -13455
rect 447 -13455 485 -13438
rect 543 -13438 663 -13400
rect 543 -13455 581 -13438
rect 447 -13472 463 -13455
rect 387 -13488 463 -13472
rect 565 -13472 581 -13455
rect 625 -13455 663 -13438
rect 721 -13438 841 -13400
rect 721 -13455 759 -13438
rect 625 -13472 641 -13455
rect 565 -13488 641 -13472
rect 743 -13472 759 -13455
rect 803 -13455 841 -13438
rect 899 -13438 1019 -13400
rect 899 -13455 937 -13438
rect 803 -13472 819 -13455
rect 743 -13488 819 -13472
rect 921 -13472 937 -13455
rect 981 -13455 1019 -13438
rect 1077 -13438 1197 -13400
rect 1077 -13455 1115 -13438
rect 981 -13472 997 -13455
rect 921 -13488 997 -13472
rect 1099 -13472 1115 -13455
rect 1159 -13455 1197 -13438
rect 1255 -13438 1375 -13400
rect 1255 -13455 1293 -13438
rect 1159 -13472 1175 -13455
rect 1099 -13488 1175 -13472
rect 1277 -13472 1293 -13455
rect 1337 -13455 1375 -13438
rect 1433 -13438 1553 -13400
rect 1433 -13455 1471 -13438
rect 1337 -13472 1353 -13455
rect 1277 -13488 1353 -13472
rect 1455 -13472 1471 -13455
rect 1515 -13455 1553 -13438
rect 1611 -13438 1731 -13400
rect 1611 -13455 1649 -13438
rect 1515 -13472 1531 -13455
rect 1455 -13488 1531 -13472
rect 1633 -13472 1649 -13455
rect 1693 -13455 1731 -13438
rect 1789 -13438 1909 -13400
rect 1789 -13455 1827 -13438
rect 1693 -13472 1709 -13455
rect 1633 -13488 1709 -13472
rect 1811 -13472 1827 -13455
rect 1871 -13455 1909 -13438
rect 1967 -13438 2087 -13400
rect 1967 -13455 2005 -13438
rect 1871 -13472 1887 -13455
rect 1811 -13488 1887 -13472
rect 1989 -13472 2005 -13455
rect 2049 -13455 2087 -13438
rect 2145 -13438 2265 -13400
rect 2145 -13455 2183 -13438
rect 2049 -13472 2065 -13455
rect 1989 -13488 2065 -13472
rect 2167 -13472 2183 -13455
rect 2227 -13455 2265 -13438
rect 2323 -13438 2443 -13400
rect 2323 -13455 2361 -13438
rect 2227 -13472 2243 -13455
rect 2167 -13488 2243 -13472
rect 2345 -13472 2361 -13455
rect 2405 -13455 2443 -13438
rect 2501 -13438 2621 -13400
rect 2501 -13455 2539 -13438
rect 2405 -13472 2421 -13455
rect 2345 -13488 2421 -13472
rect 2523 -13472 2539 -13455
rect 2583 -13455 2621 -13438
rect 2679 -13438 2799 -13400
rect 2679 -13455 2717 -13438
rect 2583 -13472 2599 -13455
rect 2523 -13488 2599 -13472
rect 2701 -13472 2717 -13455
rect 2761 -13455 2799 -13438
rect 2857 -13438 2977 -13400
rect 2857 -13455 2895 -13438
rect 2761 -13472 2777 -13455
rect 2701 -13488 2777 -13472
rect 2879 -13472 2895 -13455
rect 2939 -13455 2977 -13438
rect 3035 -13438 3155 -13400
rect 3035 -13455 3073 -13438
rect 2939 -13472 2955 -13455
rect 2879 -13488 2955 -13472
rect 3057 -13472 3073 -13455
rect 3117 -13455 3155 -13438
rect 3213 -13438 3333 -13400
rect 3213 -13455 3251 -13438
rect 3117 -13472 3133 -13455
rect 3057 -13488 3133 -13472
rect 3235 -13472 3251 -13455
rect 3295 -13455 3333 -13438
rect 3391 -13438 3511 -13400
rect 3391 -13455 3429 -13438
rect 3295 -13472 3311 -13455
rect 3235 -13488 3311 -13472
rect 3413 -13472 3429 -13455
rect 3473 -13455 3511 -13438
rect 3569 -13438 3689 -13400
rect 3569 -13455 3607 -13438
rect 3473 -13472 3489 -13455
rect 3413 -13488 3489 -13472
rect 3591 -13472 3607 -13455
rect 3651 -13455 3689 -13438
rect 3747 -13438 3867 -13400
rect 3747 -13455 3785 -13438
rect 3651 -13472 3667 -13455
rect 3591 -13488 3667 -13472
rect 3769 -13472 3785 -13455
rect 3829 -13455 3867 -13438
rect 3925 -13438 4045 -13400
rect 3925 -13455 3963 -13438
rect 3829 -13472 3845 -13455
rect 3769 -13488 3845 -13472
rect 3947 -13472 3963 -13455
rect 4007 -13455 4045 -13438
rect 4007 -13472 4023 -13455
rect 3947 -13488 4023 -13472
rect -5870 -13642 -5830 -13620
rect -5620 -13642 -5580 -13620
rect -5370 -13642 -5330 -13620
rect -5120 -13642 -5080 -13620
rect -4870 -13642 -4830 -13620
rect -4620 -13642 -4580 -13620
rect -4370 -13642 -4330 -13620
rect -4120 -13642 -4080 -13620
rect -5883 -13658 -5817 -13642
rect -5883 -13692 -5867 -13658
rect -5833 -13692 -5817 -13658
rect -5883 -13708 -5817 -13692
rect -5633 -13658 -5567 -13642
rect -5633 -13692 -5617 -13658
rect -5583 -13692 -5567 -13658
rect -5633 -13708 -5567 -13692
rect -5383 -13658 -5317 -13642
rect -5383 -13692 -5367 -13658
rect -5333 -13692 -5317 -13658
rect -5383 -13708 -5317 -13692
rect -5133 -13658 -5067 -13642
rect -5133 -13692 -5117 -13658
rect -5083 -13692 -5067 -13658
rect -5133 -13708 -5067 -13692
rect -4883 -13658 -4817 -13642
rect -4883 -13692 -4867 -13658
rect -4833 -13692 -4817 -13658
rect -4883 -13708 -4817 -13692
rect -4633 -13658 -4567 -13642
rect -4633 -13692 -4617 -13658
rect -4583 -13692 -4567 -13658
rect -4633 -13708 -4567 -13692
rect -4383 -13658 -4317 -13642
rect -4383 -13692 -4367 -13658
rect -4333 -13692 -4317 -13658
rect -4383 -13708 -4317 -13692
rect -4133 -13658 -4067 -13642
rect -4133 -13692 -4117 -13658
rect -4083 -13692 -4067 -13658
rect -4133 -13708 -4067 -13692
rect -2105 -14048 -2029 -14032
rect -2105 -14065 -2089 -14048
rect -2127 -14082 -2089 -14065
rect -2045 -14065 -2029 -14048
rect -1927 -14048 -1851 -14032
rect -1927 -14065 -1911 -14048
rect -2045 -14082 -2007 -14065
rect -2127 -14120 -2007 -14082
rect -1949 -14082 -1911 -14065
rect -1867 -14065 -1851 -14048
rect -1749 -14048 -1673 -14032
rect -1749 -14065 -1733 -14048
rect -1867 -14082 -1829 -14065
rect -1949 -14120 -1829 -14082
rect -1771 -14082 -1733 -14065
rect -1689 -14065 -1673 -14048
rect -1571 -14048 -1495 -14032
rect -1571 -14065 -1555 -14048
rect -1689 -14082 -1651 -14065
rect -1771 -14120 -1651 -14082
rect -1593 -14082 -1555 -14065
rect -1511 -14065 -1495 -14048
rect -1393 -14048 -1317 -14032
rect -1393 -14065 -1377 -14048
rect -1511 -14082 -1473 -14065
rect -1593 -14120 -1473 -14082
rect -1415 -14082 -1377 -14065
rect -1333 -14065 -1317 -14048
rect -1215 -14048 -1139 -14032
rect -1215 -14065 -1199 -14048
rect -1333 -14082 -1295 -14065
rect -1415 -14120 -1295 -14082
rect -1237 -14082 -1199 -14065
rect -1155 -14065 -1139 -14048
rect -1037 -14048 -961 -14032
rect -1037 -14065 -1021 -14048
rect -1155 -14082 -1117 -14065
rect -1237 -14120 -1117 -14082
rect -1059 -14082 -1021 -14065
rect -977 -14065 -961 -14048
rect -859 -14048 -783 -14032
rect -859 -14065 -843 -14048
rect -977 -14082 -939 -14065
rect -1059 -14120 -939 -14082
rect -881 -14082 -843 -14065
rect -799 -14065 -783 -14048
rect -681 -14048 -605 -14032
rect -681 -14065 -665 -14048
rect -799 -14082 -761 -14065
rect -881 -14120 -761 -14082
rect -703 -14082 -665 -14065
rect -621 -14065 -605 -14048
rect -503 -14048 -427 -14032
rect -503 -14065 -487 -14048
rect -621 -14082 -583 -14065
rect -703 -14120 -583 -14082
rect -525 -14082 -487 -14065
rect -443 -14065 -427 -14048
rect -325 -14048 -249 -14032
rect -325 -14065 -309 -14048
rect -443 -14082 -405 -14065
rect -525 -14120 -405 -14082
rect -347 -14082 -309 -14065
rect -265 -14065 -249 -14048
rect -147 -14048 -71 -14032
rect -147 -14065 -131 -14048
rect -265 -14082 -227 -14065
rect -347 -14120 -227 -14082
rect -169 -14082 -131 -14065
rect -87 -14065 -71 -14048
rect 31 -14048 107 -14032
rect 31 -14065 47 -14048
rect -87 -14082 -49 -14065
rect -169 -14120 -49 -14082
rect 9 -14082 47 -14065
rect 91 -14065 107 -14048
rect 209 -14048 285 -14032
rect 209 -14065 225 -14048
rect 91 -14082 129 -14065
rect 9 -14120 129 -14082
rect 187 -14082 225 -14065
rect 269 -14065 285 -14048
rect 387 -14048 463 -14032
rect 387 -14065 403 -14048
rect 269 -14082 307 -14065
rect 187 -14120 307 -14082
rect 365 -14082 403 -14065
rect 447 -14065 463 -14048
rect 565 -14048 641 -14032
rect 565 -14065 581 -14048
rect 447 -14082 485 -14065
rect 365 -14120 485 -14082
rect 543 -14082 581 -14065
rect 625 -14065 641 -14048
rect 743 -14048 819 -14032
rect 743 -14065 759 -14048
rect 625 -14082 663 -14065
rect 543 -14120 663 -14082
rect 721 -14082 759 -14065
rect 803 -14065 819 -14048
rect 921 -14048 997 -14032
rect 921 -14065 937 -14048
rect 803 -14082 841 -14065
rect 721 -14120 841 -14082
rect 899 -14082 937 -14065
rect 981 -14065 997 -14048
rect 1099 -14048 1175 -14032
rect 1099 -14065 1115 -14048
rect 981 -14082 1019 -14065
rect 899 -14120 1019 -14082
rect 1077 -14082 1115 -14065
rect 1159 -14065 1175 -14048
rect 1277 -14048 1353 -14032
rect 1277 -14065 1293 -14048
rect 1159 -14082 1197 -14065
rect 1077 -14120 1197 -14082
rect 1255 -14082 1293 -14065
rect 1337 -14065 1353 -14048
rect 1455 -14048 1531 -14032
rect 1455 -14065 1471 -14048
rect 1337 -14082 1375 -14065
rect 1255 -14120 1375 -14082
rect 1433 -14082 1471 -14065
rect 1515 -14065 1531 -14048
rect 1633 -14048 1709 -14032
rect 1633 -14065 1649 -14048
rect 1515 -14082 1553 -14065
rect 1433 -14120 1553 -14082
rect 1611 -14082 1649 -14065
rect 1693 -14065 1709 -14048
rect 1811 -14048 1887 -14032
rect 1811 -14065 1827 -14048
rect 1693 -14082 1731 -14065
rect 1611 -14120 1731 -14082
rect 1789 -14082 1827 -14065
rect 1871 -14065 1887 -14048
rect 1989 -14048 2065 -14032
rect 1989 -14065 2005 -14048
rect 1871 -14082 1909 -14065
rect 1789 -14120 1909 -14082
rect 1967 -14082 2005 -14065
rect 2049 -14065 2065 -14048
rect 2167 -14048 2243 -14032
rect 2167 -14065 2183 -14048
rect 2049 -14082 2087 -14065
rect 1967 -14120 2087 -14082
rect 2145 -14082 2183 -14065
rect 2227 -14065 2243 -14048
rect 2345 -14048 2421 -14032
rect 2345 -14065 2361 -14048
rect 2227 -14082 2265 -14065
rect 2145 -14120 2265 -14082
rect 2323 -14082 2361 -14065
rect 2405 -14065 2421 -14048
rect 2523 -14048 2599 -14032
rect 2523 -14065 2539 -14048
rect 2405 -14082 2443 -14065
rect 2323 -14120 2443 -14082
rect 2501 -14082 2539 -14065
rect 2583 -14065 2599 -14048
rect 2701 -14048 2777 -14032
rect 2701 -14065 2717 -14048
rect 2583 -14082 2621 -14065
rect 2501 -14120 2621 -14082
rect 2679 -14082 2717 -14065
rect 2761 -14065 2777 -14048
rect 2879 -14048 2955 -14032
rect 2879 -14065 2895 -14048
rect 2761 -14082 2799 -14065
rect 2679 -14120 2799 -14082
rect 2857 -14082 2895 -14065
rect 2939 -14065 2955 -14048
rect 3057 -14048 3133 -14032
rect 3057 -14065 3073 -14048
rect 2939 -14082 2977 -14065
rect 2857 -14120 2977 -14082
rect 3035 -14082 3073 -14065
rect 3117 -14065 3133 -14048
rect 3235 -14048 3311 -14032
rect 3235 -14065 3251 -14048
rect 3117 -14082 3155 -14065
rect 3035 -14120 3155 -14082
rect 3213 -14082 3251 -14065
rect 3295 -14065 3311 -14048
rect 3413 -14048 3489 -14032
rect 3413 -14065 3429 -14048
rect 3295 -14082 3333 -14065
rect 3213 -14120 3333 -14082
rect 3391 -14082 3429 -14065
rect 3473 -14065 3489 -14048
rect 3591 -14048 3667 -14032
rect 3591 -14065 3607 -14048
rect 3473 -14082 3511 -14065
rect 3391 -14120 3511 -14082
rect 3569 -14082 3607 -14065
rect 3651 -14065 3667 -14048
rect 3769 -14048 3845 -14032
rect 3769 -14065 3785 -14048
rect 3651 -14082 3689 -14065
rect 3569 -14120 3689 -14082
rect 3747 -14082 3785 -14065
rect 3829 -14065 3845 -14048
rect 3947 -14048 4023 -14032
rect 3947 -14065 3963 -14048
rect 3829 -14082 3867 -14065
rect 3747 -14120 3867 -14082
rect 3925 -14082 3963 -14065
rect 4007 -14065 4023 -14048
rect 5645 -14048 5721 -14032
rect 5645 -14065 5661 -14048
rect 4007 -14082 4045 -14065
rect 3925 -14120 4045 -14082
rect 5623 -14082 5661 -14065
rect 5705 -14065 5721 -14048
rect 5823 -14048 5899 -14032
rect 5823 -14065 5839 -14048
rect 5705 -14082 5743 -14065
rect 5623 -14120 5743 -14082
rect 5801 -14082 5839 -14065
rect 5883 -14065 5899 -14048
rect 6001 -14048 6077 -14032
rect 6001 -14065 6017 -14048
rect 5883 -14082 5921 -14065
rect 5801 -14120 5921 -14082
rect 5979 -14082 6017 -14065
rect 6061 -14065 6077 -14048
rect 6179 -14048 6255 -14032
rect 6179 -14065 6195 -14048
rect 6061 -14082 6099 -14065
rect 5979 -14120 6099 -14082
rect 6157 -14082 6195 -14065
rect 6239 -14065 6255 -14048
rect 6357 -14048 6433 -14032
rect 6357 -14065 6373 -14048
rect 6239 -14082 6277 -14065
rect 6157 -14120 6277 -14082
rect 6335 -14082 6373 -14065
rect 6417 -14065 6433 -14048
rect 6535 -14048 6611 -14032
rect 6535 -14065 6551 -14048
rect 6417 -14082 6455 -14065
rect 6335 -14120 6455 -14082
rect 6513 -14082 6551 -14065
rect 6595 -14065 6611 -14048
rect 6713 -14048 6789 -14032
rect 6713 -14065 6729 -14048
rect 6595 -14082 6633 -14065
rect 6513 -14120 6633 -14082
rect 6691 -14082 6729 -14065
rect 6773 -14065 6789 -14048
rect 6891 -14048 6967 -14032
rect 6891 -14065 6907 -14048
rect 6773 -14082 6811 -14065
rect 6691 -14120 6811 -14082
rect 6869 -14082 6907 -14065
rect 6951 -14065 6967 -14048
rect 7069 -14048 7145 -14032
rect 7069 -14065 7085 -14048
rect 6951 -14082 6989 -14065
rect 6869 -14120 6989 -14082
rect 7047 -14082 7085 -14065
rect 7129 -14065 7145 -14048
rect 7247 -14048 7323 -14032
rect 7247 -14065 7263 -14048
rect 7129 -14082 7167 -14065
rect 7047 -14120 7167 -14082
rect 7225 -14082 7263 -14065
rect 7307 -14065 7323 -14048
rect 7425 -14048 7501 -14032
rect 7425 -14065 7441 -14048
rect 7307 -14082 7345 -14065
rect 7225 -14120 7345 -14082
rect 7403 -14082 7441 -14065
rect 7485 -14065 7501 -14048
rect 7603 -14048 7679 -14032
rect 7603 -14065 7619 -14048
rect 7485 -14082 7523 -14065
rect 7403 -14120 7523 -14082
rect 7581 -14082 7619 -14065
rect 7663 -14065 7679 -14048
rect 7781 -14048 7857 -14032
rect 7781 -14065 7797 -14048
rect 7663 -14082 7701 -14065
rect 7581 -14120 7701 -14082
rect 7759 -14082 7797 -14065
rect 7841 -14065 7857 -14048
rect 7959 -14048 8035 -14032
rect 7959 -14065 7975 -14048
rect 7841 -14082 7879 -14065
rect 7759 -14120 7879 -14082
rect 7937 -14082 7975 -14065
rect 8019 -14065 8035 -14048
rect 8137 -14048 8213 -14032
rect 8137 -14065 8153 -14048
rect 8019 -14082 8057 -14065
rect 7937 -14120 8057 -14082
rect 8115 -14082 8153 -14065
rect 8197 -14065 8213 -14048
rect 8315 -14048 8391 -14032
rect 8315 -14065 8331 -14048
rect 8197 -14082 8235 -14065
rect 8115 -14120 8235 -14082
rect 8293 -14082 8331 -14065
rect 8375 -14065 8391 -14048
rect 8493 -14048 8569 -14032
rect 8493 -14065 8509 -14048
rect 8375 -14082 8413 -14065
rect 8293 -14120 8413 -14082
rect 8471 -14082 8509 -14065
rect 8553 -14065 8569 -14048
rect 8671 -14048 8747 -14032
rect 8671 -14065 8687 -14048
rect 8553 -14082 8591 -14065
rect 8471 -14120 8591 -14082
rect 8649 -14082 8687 -14065
rect 8731 -14065 8747 -14048
rect 8849 -14048 8925 -14032
rect 8849 -14065 8865 -14048
rect 8731 -14082 8769 -14065
rect 8649 -14120 8769 -14082
rect 8827 -14082 8865 -14065
rect 8909 -14065 8925 -14048
rect 9027 -14048 9103 -14032
rect 9027 -14065 9043 -14048
rect 8909 -14082 8947 -14065
rect 8827 -14120 8947 -14082
rect 9005 -14082 9043 -14065
rect 9087 -14065 9103 -14048
rect 9205 -14048 9281 -14032
rect 9205 -14065 9221 -14048
rect 9087 -14082 9125 -14065
rect 9005 -14120 9125 -14082
rect 9183 -14082 9221 -14065
rect 9265 -14065 9281 -14048
rect 9383 -14048 9459 -14032
rect 9383 -14065 9399 -14048
rect 9265 -14082 9303 -14065
rect 9183 -14120 9303 -14082
rect 9361 -14082 9399 -14065
rect 9443 -14065 9459 -14048
rect 9561 -14048 9637 -14032
rect 9561 -14065 9577 -14048
rect 9443 -14082 9481 -14065
rect 9361 -14120 9481 -14082
rect 9539 -14082 9577 -14065
rect 9621 -14065 9637 -14048
rect 9739 -14048 9815 -14032
rect 9739 -14065 9755 -14048
rect 9621 -14082 9659 -14065
rect 9539 -14120 9659 -14082
rect 9717 -14082 9755 -14065
rect 9799 -14065 9815 -14048
rect 9917 -14048 9993 -14032
rect 9917 -14065 9933 -14048
rect 9799 -14082 9837 -14065
rect 9717 -14120 9837 -14082
rect 9895 -14082 9933 -14065
rect 9977 -14065 9993 -14048
rect 10095 -14048 10171 -14032
rect 10095 -14065 10111 -14048
rect 9977 -14082 10015 -14065
rect 9895 -14120 10015 -14082
rect 10073 -14082 10111 -14065
rect 10155 -14065 10171 -14048
rect 10273 -14048 10349 -14032
rect 10273 -14065 10289 -14048
rect 10155 -14082 10193 -14065
rect 10073 -14120 10193 -14082
rect 10251 -14082 10289 -14065
rect 10333 -14065 10349 -14048
rect 10451 -14048 10527 -14032
rect 10451 -14065 10467 -14048
rect 10333 -14082 10371 -14065
rect 10251 -14120 10371 -14082
rect 10429 -14082 10467 -14065
rect 10511 -14065 10527 -14048
rect 10629 -14048 10705 -14032
rect 10629 -14065 10645 -14048
rect 10511 -14082 10549 -14065
rect 10429 -14120 10549 -14082
rect 10607 -14082 10645 -14065
rect 10689 -14065 10705 -14048
rect 10807 -14048 10883 -14032
rect 10807 -14065 10823 -14048
rect 10689 -14082 10727 -14065
rect 10607 -14120 10727 -14082
rect 10785 -14082 10823 -14065
rect 10867 -14065 10883 -14048
rect 10985 -14048 11061 -14032
rect 10985 -14065 11001 -14048
rect 10867 -14082 10905 -14065
rect 10785 -14120 10905 -14082
rect 10963 -14082 11001 -14065
rect 11045 -14065 11061 -14048
rect 11163 -14048 11239 -14032
rect 11163 -14065 11179 -14048
rect 11045 -14082 11083 -14065
rect 10963 -14120 11083 -14082
rect 11141 -14082 11179 -14065
rect 11223 -14065 11239 -14048
rect 11341 -14048 11417 -14032
rect 11341 -14065 11357 -14048
rect 11223 -14082 11261 -14065
rect 11141 -14120 11261 -14082
rect 11319 -14082 11357 -14065
rect 11401 -14065 11417 -14048
rect 11519 -14048 11595 -14032
rect 11519 -14065 11535 -14048
rect 11401 -14082 11439 -14065
rect 11319 -14120 11439 -14082
rect 11497 -14082 11535 -14065
rect 11579 -14065 11595 -14048
rect 11697 -14048 11773 -14032
rect 11697 -14065 11713 -14048
rect 11579 -14082 11617 -14065
rect 11497 -14120 11617 -14082
rect 11675 -14082 11713 -14065
rect 11757 -14065 11773 -14048
rect 11875 -14048 11951 -14032
rect 11875 -14065 11891 -14048
rect 11757 -14082 11795 -14065
rect 11675 -14120 11795 -14082
rect 11853 -14082 11891 -14065
rect 11935 -14065 11951 -14048
rect 12053 -14048 12129 -14032
rect 12053 -14065 12069 -14048
rect 11935 -14082 11973 -14065
rect 11853 -14120 11973 -14082
rect 12031 -14082 12069 -14065
rect 12113 -14065 12129 -14048
rect 12231 -14048 12307 -14032
rect 12231 -14065 12247 -14048
rect 12113 -14082 12151 -14065
rect 12031 -14120 12151 -14082
rect 12209 -14082 12247 -14065
rect 12291 -14065 12307 -14048
rect 12409 -14048 12485 -14032
rect 12409 -14065 12425 -14048
rect 12291 -14082 12329 -14065
rect 12209 -14120 12329 -14082
rect 12387 -14082 12425 -14065
rect 12469 -14065 12485 -14048
rect 12587 -14048 12663 -14032
rect 12587 -14065 12603 -14048
rect 12469 -14082 12507 -14065
rect 12387 -14120 12507 -14082
rect 12565 -14082 12603 -14065
rect 12647 -14065 12663 -14048
rect 12647 -14082 12685 -14065
rect 12565 -14120 12685 -14082
rect -5960 -14310 -5884 -14294
rect -5960 -14327 -5944 -14310
rect -5982 -14344 -5944 -14327
rect -5900 -14327 -5884 -14310
rect -5782 -14310 -5706 -14294
rect -5782 -14327 -5766 -14310
rect -5900 -14344 -5862 -14327
rect -5982 -14382 -5862 -14344
rect -5804 -14344 -5766 -14327
rect -5722 -14327 -5706 -14310
rect -5604 -14310 -5528 -14294
rect -5604 -14327 -5588 -14310
rect -5722 -14344 -5684 -14327
rect -5804 -14382 -5684 -14344
rect -5626 -14344 -5588 -14327
rect -5544 -14327 -5528 -14310
rect -5426 -14310 -5350 -14294
rect -5426 -14327 -5410 -14310
rect -5544 -14344 -5506 -14327
rect -5626 -14382 -5506 -14344
rect -5448 -14344 -5410 -14327
rect -5366 -14327 -5350 -14310
rect -5248 -14310 -5172 -14294
rect -5248 -14327 -5232 -14310
rect -5366 -14344 -5328 -14327
rect -5448 -14382 -5328 -14344
rect -5270 -14344 -5232 -14327
rect -5188 -14327 -5172 -14310
rect -5070 -14310 -4994 -14294
rect -5070 -14327 -5054 -14310
rect -5188 -14344 -5150 -14327
rect -5270 -14382 -5150 -14344
rect -5092 -14344 -5054 -14327
rect -5010 -14327 -4994 -14310
rect -4892 -14310 -4816 -14294
rect -4892 -14327 -4876 -14310
rect -5010 -14344 -4972 -14327
rect -5092 -14382 -4972 -14344
rect -4914 -14344 -4876 -14327
rect -4832 -14327 -4816 -14310
rect -4714 -14310 -4638 -14294
rect -4714 -14327 -4698 -14310
rect -4832 -14344 -4794 -14327
rect -4914 -14382 -4794 -14344
rect -4736 -14344 -4698 -14327
rect -4654 -14327 -4638 -14310
rect -4536 -14310 -4460 -14294
rect -4536 -14327 -4520 -14310
rect -4654 -14344 -4616 -14327
rect -4736 -14382 -4616 -14344
rect -4558 -14344 -4520 -14327
rect -4476 -14327 -4460 -14310
rect -4358 -14310 -4282 -14294
rect -4358 -14327 -4342 -14310
rect -4476 -14344 -4438 -14327
rect -4558 -14382 -4438 -14344
rect -4380 -14344 -4342 -14327
rect -4298 -14327 -4282 -14310
rect -4180 -14310 -4104 -14294
rect -4180 -14327 -4164 -14310
rect -4298 -14344 -4260 -14327
rect -4380 -14382 -4260 -14344
rect -4202 -14344 -4164 -14327
rect -4120 -14327 -4104 -14310
rect -4120 -14344 -4082 -14327
rect -4202 -14382 -4082 -14344
rect -2127 -14438 -2007 -14400
rect -2127 -14455 -2089 -14438
rect -2105 -14472 -2089 -14455
rect -2045 -14455 -2007 -14438
rect -1949 -14438 -1829 -14400
rect -1949 -14455 -1911 -14438
rect -2045 -14472 -2029 -14455
rect -2105 -14488 -2029 -14472
rect -1927 -14472 -1911 -14455
rect -1867 -14455 -1829 -14438
rect -1771 -14438 -1651 -14400
rect -1771 -14455 -1733 -14438
rect -1867 -14472 -1851 -14455
rect -1927 -14488 -1851 -14472
rect -1749 -14472 -1733 -14455
rect -1689 -14455 -1651 -14438
rect -1593 -14438 -1473 -14400
rect -1593 -14455 -1555 -14438
rect -1689 -14472 -1673 -14455
rect -1749 -14488 -1673 -14472
rect -1571 -14472 -1555 -14455
rect -1511 -14455 -1473 -14438
rect -1415 -14438 -1295 -14400
rect -1415 -14455 -1377 -14438
rect -1511 -14472 -1495 -14455
rect -1571 -14488 -1495 -14472
rect -1393 -14472 -1377 -14455
rect -1333 -14455 -1295 -14438
rect -1237 -14438 -1117 -14400
rect -1237 -14455 -1199 -14438
rect -1333 -14472 -1317 -14455
rect -1393 -14488 -1317 -14472
rect -1215 -14472 -1199 -14455
rect -1155 -14455 -1117 -14438
rect -1059 -14438 -939 -14400
rect -1059 -14455 -1021 -14438
rect -1155 -14472 -1139 -14455
rect -1215 -14488 -1139 -14472
rect -1037 -14472 -1021 -14455
rect -977 -14455 -939 -14438
rect -881 -14438 -761 -14400
rect -881 -14455 -843 -14438
rect -977 -14472 -961 -14455
rect -1037 -14488 -961 -14472
rect -859 -14472 -843 -14455
rect -799 -14455 -761 -14438
rect -703 -14438 -583 -14400
rect -703 -14455 -665 -14438
rect -799 -14472 -783 -14455
rect -859 -14488 -783 -14472
rect -681 -14472 -665 -14455
rect -621 -14455 -583 -14438
rect -525 -14438 -405 -14400
rect -525 -14455 -487 -14438
rect -621 -14472 -605 -14455
rect -681 -14488 -605 -14472
rect -503 -14472 -487 -14455
rect -443 -14455 -405 -14438
rect -347 -14438 -227 -14400
rect -347 -14455 -309 -14438
rect -443 -14472 -427 -14455
rect -503 -14488 -427 -14472
rect -325 -14472 -309 -14455
rect -265 -14455 -227 -14438
rect -169 -14438 -49 -14400
rect -169 -14455 -131 -14438
rect -265 -14472 -249 -14455
rect -325 -14488 -249 -14472
rect -147 -14472 -131 -14455
rect -87 -14455 -49 -14438
rect 9 -14438 129 -14400
rect 9 -14455 47 -14438
rect -87 -14472 -71 -14455
rect -147 -14488 -71 -14472
rect 31 -14472 47 -14455
rect 91 -14455 129 -14438
rect 187 -14438 307 -14400
rect 187 -14455 225 -14438
rect 91 -14472 107 -14455
rect 31 -14488 107 -14472
rect 209 -14472 225 -14455
rect 269 -14455 307 -14438
rect 365 -14438 485 -14400
rect 365 -14455 403 -14438
rect 269 -14472 285 -14455
rect 209 -14488 285 -14472
rect 387 -14472 403 -14455
rect 447 -14455 485 -14438
rect 543 -14438 663 -14400
rect 543 -14455 581 -14438
rect 447 -14472 463 -14455
rect 387 -14488 463 -14472
rect 565 -14472 581 -14455
rect 625 -14455 663 -14438
rect 721 -14438 841 -14400
rect 721 -14455 759 -14438
rect 625 -14472 641 -14455
rect 565 -14488 641 -14472
rect 743 -14472 759 -14455
rect 803 -14455 841 -14438
rect 899 -14438 1019 -14400
rect 899 -14455 937 -14438
rect 803 -14472 819 -14455
rect 743 -14488 819 -14472
rect 921 -14472 937 -14455
rect 981 -14455 1019 -14438
rect 1077 -14438 1197 -14400
rect 1077 -14455 1115 -14438
rect 981 -14472 997 -14455
rect 921 -14488 997 -14472
rect 1099 -14472 1115 -14455
rect 1159 -14455 1197 -14438
rect 1255 -14438 1375 -14400
rect 1255 -14455 1293 -14438
rect 1159 -14472 1175 -14455
rect 1099 -14488 1175 -14472
rect 1277 -14472 1293 -14455
rect 1337 -14455 1375 -14438
rect 1433 -14438 1553 -14400
rect 1433 -14455 1471 -14438
rect 1337 -14472 1353 -14455
rect 1277 -14488 1353 -14472
rect 1455 -14472 1471 -14455
rect 1515 -14455 1553 -14438
rect 1611 -14438 1731 -14400
rect 1611 -14455 1649 -14438
rect 1515 -14472 1531 -14455
rect 1455 -14488 1531 -14472
rect 1633 -14472 1649 -14455
rect 1693 -14455 1731 -14438
rect 1789 -14438 1909 -14400
rect 1789 -14455 1827 -14438
rect 1693 -14472 1709 -14455
rect 1633 -14488 1709 -14472
rect 1811 -14472 1827 -14455
rect 1871 -14455 1909 -14438
rect 1967 -14438 2087 -14400
rect 1967 -14455 2005 -14438
rect 1871 -14472 1887 -14455
rect 1811 -14488 1887 -14472
rect 1989 -14472 2005 -14455
rect 2049 -14455 2087 -14438
rect 2145 -14438 2265 -14400
rect 2145 -14455 2183 -14438
rect 2049 -14472 2065 -14455
rect 1989 -14488 2065 -14472
rect 2167 -14472 2183 -14455
rect 2227 -14455 2265 -14438
rect 2323 -14438 2443 -14400
rect 2323 -14455 2361 -14438
rect 2227 -14472 2243 -14455
rect 2167 -14488 2243 -14472
rect 2345 -14472 2361 -14455
rect 2405 -14455 2443 -14438
rect 2501 -14438 2621 -14400
rect 2501 -14455 2539 -14438
rect 2405 -14472 2421 -14455
rect 2345 -14488 2421 -14472
rect 2523 -14472 2539 -14455
rect 2583 -14455 2621 -14438
rect 2679 -14438 2799 -14400
rect 2679 -14455 2717 -14438
rect 2583 -14472 2599 -14455
rect 2523 -14488 2599 -14472
rect 2701 -14472 2717 -14455
rect 2761 -14455 2799 -14438
rect 2857 -14438 2977 -14400
rect 2857 -14455 2895 -14438
rect 2761 -14472 2777 -14455
rect 2701 -14488 2777 -14472
rect 2879 -14472 2895 -14455
rect 2939 -14455 2977 -14438
rect 3035 -14438 3155 -14400
rect 3035 -14455 3073 -14438
rect 2939 -14472 2955 -14455
rect 2879 -14488 2955 -14472
rect 3057 -14472 3073 -14455
rect 3117 -14455 3155 -14438
rect 3213 -14438 3333 -14400
rect 3213 -14455 3251 -14438
rect 3117 -14472 3133 -14455
rect 3057 -14488 3133 -14472
rect 3235 -14472 3251 -14455
rect 3295 -14455 3333 -14438
rect 3391 -14438 3511 -14400
rect 3391 -14455 3429 -14438
rect 3295 -14472 3311 -14455
rect 3235 -14488 3311 -14472
rect 3413 -14472 3429 -14455
rect 3473 -14455 3511 -14438
rect 3569 -14438 3689 -14400
rect 3569 -14455 3607 -14438
rect 3473 -14472 3489 -14455
rect 3413 -14488 3489 -14472
rect 3591 -14472 3607 -14455
rect 3651 -14455 3689 -14438
rect 3747 -14438 3867 -14400
rect 3747 -14455 3785 -14438
rect 3651 -14472 3667 -14455
rect 3591 -14488 3667 -14472
rect 3769 -14472 3785 -14455
rect 3829 -14455 3867 -14438
rect 3925 -14438 4045 -14400
rect 3925 -14455 3963 -14438
rect 3829 -14472 3845 -14455
rect 3769 -14488 3845 -14472
rect 3947 -14472 3963 -14455
rect 4007 -14455 4045 -14438
rect 5623 -14438 5743 -14400
rect 5623 -14455 5661 -14438
rect 4007 -14472 4023 -14455
rect 3947 -14488 4023 -14472
rect 5645 -14472 5661 -14455
rect 5705 -14455 5743 -14438
rect 5801 -14438 5921 -14400
rect 5801 -14455 5839 -14438
rect 5705 -14472 5721 -14455
rect 5645 -14488 5721 -14472
rect 5823 -14472 5839 -14455
rect 5883 -14455 5921 -14438
rect 5979 -14438 6099 -14400
rect 5979 -14455 6017 -14438
rect 5883 -14472 5899 -14455
rect 5823 -14488 5899 -14472
rect 6001 -14472 6017 -14455
rect 6061 -14455 6099 -14438
rect 6157 -14438 6277 -14400
rect 6157 -14455 6195 -14438
rect 6061 -14472 6077 -14455
rect 6001 -14488 6077 -14472
rect 6179 -14472 6195 -14455
rect 6239 -14455 6277 -14438
rect 6335 -14438 6455 -14400
rect 6335 -14455 6373 -14438
rect 6239 -14472 6255 -14455
rect 6179 -14488 6255 -14472
rect 6357 -14472 6373 -14455
rect 6417 -14455 6455 -14438
rect 6513 -14438 6633 -14400
rect 6513 -14455 6551 -14438
rect 6417 -14472 6433 -14455
rect 6357 -14488 6433 -14472
rect 6535 -14472 6551 -14455
rect 6595 -14455 6633 -14438
rect 6691 -14438 6811 -14400
rect 6691 -14455 6729 -14438
rect 6595 -14472 6611 -14455
rect 6535 -14488 6611 -14472
rect 6713 -14472 6729 -14455
rect 6773 -14455 6811 -14438
rect 6869 -14438 6989 -14400
rect 6869 -14455 6907 -14438
rect 6773 -14472 6789 -14455
rect 6713 -14488 6789 -14472
rect 6891 -14472 6907 -14455
rect 6951 -14455 6989 -14438
rect 7047 -14438 7167 -14400
rect 7047 -14455 7085 -14438
rect 6951 -14472 6967 -14455
rect 6891 -14488 6967 -14472
rect 7069 -14472 7085 -14455
rect 7129 -14455 7167 -14438
rect 7225 -14438 7345 -14400
rect 7225 -14455 7263 -14438
rect 7129 -14472 7145 -14455
rect 7069 -14488 7145 -14472
rect 7247 -14472 7263 -14455
rect 7307 -14455 7345 -14438
rect 7403 -14438 7523 -14400
rect 7403 -14455 7441 -14438
rect 7307 -14472 7323 -14455
rect 7247 -14488 7323 -14472
rect 7425 -14472 7441 -14455
rect 7485 -14455 7523 -14438
rect 7581 -14438 7701 -14400
rect 7581 -14455 7619 -14438
rect 7485 -14472 7501 -14455
rect 7425 -14488 7501 -14472
rect 7603 -14472 7619 -14455
rect 7663 -14455 7701 -14438
rect 7759 -14438 7879 -14400
rect 7759 -14455 7797 -14438
rect 7663 -14472 7679 -14455
rect 7603 -14488 7679 -14472
rect 7781 -14472 7797 -14455
rect 7841 -14455 7879 -14438
rect 7937 -14438 8057 -14400
rect 7937 -14455 7975 -14438
rect 7841 -14472 7857 -14455
rect 7781 -14488 7857 -14472
rect 7959 -14472 7975 -14455
rect 8019 -14455 8057 -14438
rect 8115 -14438 8235 -14400
rect 8115 -14455 8153 -14438
rect 8019 -14472 8035 -14455
rect 7959 -14488 8035 -14472
rect 8137 -14472 8153 -14455
rect 8197 -14455 8235 -14438
rect 8293 -14438 8413 -14400
rect 8293 -14455 8331 -14438
rect 8197 -14472 8213 -14455
rect 8137 -14488 8213 -14472
rect 8315 -14472 8331 -14455
rect 8375 -14455 8413 -14438
rect 8471 -14438 8591 -14400
rect 8471 -14455 8509 -14438
rect 8375 -14472 8391 -14455
rect 8315 -14488 8391 -14472
rect 8493 -14472 8509 -14455
rect 8553 -14455 8591 -14438
rect 8649 -14438 8769 -14400
rect 8649 -14455 8687 -14438
rect 8553 -14472 8569 -14455
rect 8493 -14488 8569 -14472
rect 8671 -14472 8687 -14455
rect 8731 -14455 8769 -14438
rect 8827 -14438 8947 -14400
rect 8827 -14455 8865 -14438
rect 8731 -14472 8747 -14455
rect 8671 -14488 8747 -14472
rect 8849 -14472 8865 -14455
rect 8909 -14455 8947 -14438
rect 9005 -14438 9125 -14400
rect 9005 -14455 9043 -14438
rect 8909 -14472 8925 -14455
rect 8849 -14488 8925 -14472
rect 9027 -14472 9043 -14455
rect 9087 -14455 9125 -14438
rect 9183 -14438 9303 -14400
rect 9183 -14455 9221 -14438
rect 9087 -14472 9103 -14455
rect 9027 -14488 9103 -14472
rect 9205 -14472 9221 -14455
rect 9265 -14455 9303 -14438
rect 9361 -14438 9481 -14400
rect 9361 -14455 9399 -14438
rect 9265 -14472 9281 -14455
rect 9205 -14488 9281 -14472
rect 9383 -14472 9399 -14455
rect 9443 -14455 9481 -14438
rect 9539 -14438 9659 -14400
rect 9539 -14455 9577 -14438
rect 9443 -14472 9459 -14455
rect 9383 -14488 9459 -14472
rect 9561 -14472 9577 -14455
rect 9621 -14455 9659 -14438
rect 9717 -14438 9837 -14400
rect 9717 -14455 9755 -14438
rect 9621 -14472 9637 -14455
rect 9561 -14488 9637 -14472
rect 9739 -14472 9755 -14455
rect 9799 -14455 9837 -14438
rect 9895 -14438 10015 -14400
rect 9895 -14455 9933 -14438
rect 9799 -14472 9815 -14455
rect 9739 -14488 9815 -14472
rect 9917 -14472 9933 -14455
rect 9977 -14455 10015 -14438
rect 10073 -14438 10193 -14400
rect 10073 -14455 10111 -14438
rect 9977 -14472 9993 -14455
rect 9917 -14488 9993 -14472
rect 10095 -14472 10111 -14455
rect 10155 -14455 10193 -14438
rect 10251 -14438 10371 -14400
rect 10251 -14455 10289 -14438
rect 10155 -14472 10171 -14455
rect 10095 -14488 10171 -14472
rect 10273 -14472 10289 -14455
rect 10333 -14455 10371 -14438
rect 10429 -14438 10549 -14400
rect 10429 -14455 10467 -14438
rect 10333 -14472 10349 -14455
rect 10273 -14488 10349 -14472
rect 10451 -14472 10467 -14455
rect 10511 -14455 10549 -14438
rect 10607 -14438 10727 -14400
rect 10607 -14455 10645 -14438
rect 10511 -14472 10527 -14455
rect 10451 -14488 10527 -14472
rect 10629 -14472 10645 -14455
rect 10689 -14455 10727 -14438
rect 10785 -14438 10905 -14400
rect 10785 -14455 10823 -14438
rect 10689 -14472 10705 -14455
rect 10629 -14488 10705 -14472
rect 10807 -14472 10823 -14455
rect 10867 -14455 10905 -14438
rect 10963 -14438 11083 -14400
rect 10963 -14455 11001 -14438
rect 10867 -14472 10883 -14455
rect 10807 -14488 10883 -14472
rect 10985 -14472 11001 -14455
rect 11045 -14455 11083 -14438
rect 11141 -14438 11261 -14400
rect 11141 -14455 11179 -14438
rect 11045 -14472 11061 -14455
rect 10985 -14488 11061 -14472
rect 11163 -14472 11179 -14455
rect 11223 -14455 11261 -14438
rect 11319 -14438 11439 -14400
rect 11319 -14455 11357 -14438
rect 11223 -14472 11239 -14455
rect 11163 -14488 11239 -14472
rect 11341 -14472 11357 -14455
rect 11401 -14455 11439 -14438
rect 11497 -14438 11617 -14400
rect 11497 -14455 11535 -14438
rect 11401 -14472 11417 -14455
rect 11341 -14488 11417 -14472
rect 11519 -14472 11535 -14455
rect 11579 -14455 11617 -14438
rect 11675 -14438 11795 -14400
rect 11675 -14455 11713 -14438
rect 11579 -14472 11595 -14455
rect 11519 -14488 11595 -14472
rect 11697 -14472 11713 -14455
rect 11757 -14455 11795 -14438
rect 11853 -14438 11973 -14400
rect 11853 -14455 11891 -14438
rect 11757 -14472 11773 -14455
rect 11697 -14488 11773 -14472
rect 11875 -14472 11891 -14455
rect 11935 -14455 11973 -14438
rect 12031 -14438 12151 -14400
rect 12031 -14455 12069 -14438
rect 11935 -14472 11951 -14455
rect 11875 -14488 11951 -14472
rect 12053 -14472 12069 -14455
rect 12113 -14455 12151 -14438
rect 12209 -14438 12329 -14400
rect 12209 -14455 12247 -14438
rect 12113 -14472 12129 -14455
rect 12053 -14488 12129 -14472
rect 12231 -14472 12247 -14455
rect 12291 -14455 12329 -14438
rect 12387 -14438 12507 -14400
rect 12387 -14455 12425 -14438
rect 12291 -14472 12307 -14455
rect 12231 -14488 12307 -14472
rect 12409 -14472 12425 -14455
rect 12469 -14455 12507 -14438
rect 12565 -14438 12685 -14400
rect 12565 -14455 12603 -14438
rect 12469 -14472 12485 -14455
rect 12409 -14488 12485 -14472
rect 12587 -14472 12603 -14455
rect 12647 -14455 12685 -14438
rect 12647 -14472 12663 -14455
rect 12587 -14488 12663 -14472
rect -5982 -14700 -5862 -14662
rect -5982 -14717 -5944 -14700
rect -5960 -14734 -5944 -14717
rect -5900 -14717 -5862 -14700
rect -5804 -14700 -5684 -14662
rect -5804 -14717 -5766 -14700
rect -5900 -14734 -5884 -14717
rect -5960 -14750 -5884 -14734
rect -5782 -14734 -5766 -14717
rect -5722 -14717 -5684 -14700
rect -5626 -14700 -5506 -14662
rect -5626 -14717 -5588 -14700
rect -5722 -14734 -5706 -14717
rect -5782 -14750 -5706 -14734
rect -5604 -14734 -5588 -14717
rect -5544 -14717 -5506 -14700
rect -5448 -14700 -5328 -14662
rect -5448 -14717 -5410 -14700
rect -5544 -14734 -5528 -14717
rect -5604 -14750 -5528 -14734
rect -5426 -14734 -5410 -14717
rect -5366 -14717 -5328 -14700
rect -5270 -14700 -5150 -14662
rect -5270 -14717 -5232 -14700
rect -5366 -14734 -5350 -14717
rect -5426 -14750 -5350 -14734
rect -5248 -14734 -5232 -14717
rect -5188 -14717 -5150 -14700
rect -5092 -14700 -4972 -14662
rect -5092 -14717 -5054 -14700
rect -5188 -14734 -5172 -14717
rect -5248 -14750 -5172 -14734
rect -5070 -14734 -5054 -14717
rect -5010 -14717 -4972 -14700
rect -4914 -14700 -4794 -14662
rect -4914 -14717 -4876 -14700
rect -5010 -14734 -4994 -14717
rect -5070 -14750 -4994 -14734
rect -4892 -14734 -4876 -14717
rect -4832 -14717 -4794 -14700
rect -4736 -14700 -4616 -14662
rect -4736 -14717 -4698 -14700
rect -4832 -14734 -4816 -14717
rect -4892 -14750 -4816 -14734
rect -4714 -14734 -4698 -14717
rect -4654 -14717 -4616 -14700
rect -4558 -14700 -4438 -14662
rect -4558 -14717 -4520 -14700
rect -4654 -14734 -4638 -14717
rect -4714 -14750 -4638 -14734
rect -4536 -14734 -4520 -14717
rect -4476 -14717 -4438 -14700
rect -4380 -14700 -4260 -14662
rect -4380 -14717 -4342 -14700
rect -4476 -14734 -4460 -14717
rect -4536 -14750 -4460 -14734
rect -4358 -14734 -4342 -14717
rect -4298 -14717 -4260 -14700
rect -4202 -14700 -4082 -14662
rect -4202 -14717 -4164 -14700
rect -4298 -14734 -4282 -14717
rect -4358 -14750 -4282 -14734
rect -4180 -14734 -4164 -14717
rect -4120 -14717 -4082 -14700
rect -4120 -14734 -4104 -14717
rect -4180 -14750 -4104 -14734
rect -5960 -15010 -5884 -14994
rect -5960 -15027 -5944 -15010
rect -5982 -15044 -5944 -15027
rect -5900 -15027 -5884 -15010
rect -5782 -15010 -5706 -14994
rect -5782 -15027 -5766 -15010
rect -5900 -15044 -5862 -15027
rect -5982 -15082 -5862 -15044
rect -5804 -15044 -5766 -15027
rect -5722 -15027 -5706 -15010
rect -5604 -15010 -5528 -14994
rect -5604 -15027 -5588 -15010
rect -5722 -15044 -5684 -15027
rect -5804 -15082 -5684 -15044
rect -5626 -15044 -5588 -15027
rect -5544 -15027 -5528 -15010
rect -5426 -15010 -5350 -14994
rect -5426 -15027 -5410 -15010
rect -5544 -15044 -5506 -15027
rect -5626 -15082 -5506 -15044
rect -5448 -15044 -5410 -15027
rect -5366 -15027 -5350 -15010
rect -5248 -15010 -5172 -14994
rect -5248 -15027 -5232 -15010
rect -5366 -15044 -5328 -15027
rect -5448 -15082 -5328 -15044
rect -5270 -15044 -5232 -15027
rect -5188 -15027 -5172 -15010
rect -5070 -15010 -4994 -14994
rect -5070 -15027 -5054 -15010
rect -5188 -15044 -5150 -15027
rect -5270 -15082 -5150 -15044
rect -5092 -15044 -5054 -15027
rect -5010 -15027 -4994 -15010
rect -4892 -15010 -4816 -14994
rect -4892 -15027 -4876 -15010
rect -5010 -15044 -4972 -15027
rect -5092 -15082 -4972 -15044
rect -4914 -15044 -4876 -15027
rect -4832 -15027 -4816 -15010
rect -4714 -15010 -4638 -14994
rect -4714 -15027 -4698 -15010
rect -4832 -15044 -4794 -15027
rect -4914 -15082 -4794 -15044
rect -4736 -15044 -4698 -15027
rect -4654 -15027 -4638 -15010
rect -4536 -15010 -4460 -14994
rect -4536 -15027 -4520 -15010
rect -4654 -15044 -4616 -15027
rect -4736 -15082 -4616 -15044
rect -4558 -15044 -4520 -15027
rect -4476 -15027 -4460 -15010
rect -4358 -15010 -4282 -14994
rect -4358 -15027 -4342 -15010
rect -4476 -15044 -4438 -15027
rect -4558 -15082 -4438 -15044
rect -4380 -15044 -4342 -15027
rect -4298 -15027 -4282 -15010
rect -4180 -15010 -4104 -14994
rect -4180 -15027 -4164 -15010
rect -4298 -15044 -4260 -15027
rect -4380 -15082 -4260 -15044
rect -4202 -15044 -4164 -15027
rect -4120 -15027 -4104 -15010
rect -4120 -15044 -4082 -15027
rect -4202 -15082 -4082 -15044
rect -2105 -15048 -2029 -15032
rect -2105 -15065 -2089 -15048
rect -2127 -15082 -2089 -15065
rect -2045 -15065 -2029 -15048
rect -1927 -15048 -1851 -15032
rect -1927 -15065 -1911 -15048
rect -2045 -15082 -2007 -15065
rect -2127 -15120 -2007 -15082
rect -1949 -15082 -1911 -15065
rect -1867 -15065 -1851 -15048
rect -1749 -15048 -1673 -15032
rect -1749 -15065 -1733 -15048
rect -1867 -15082 -1829 -15065
rect -1949 -15120 -1829 -15082
rect -1771 -15082 -1733 -15065
rect -1689 -15065 -1673 -15048
rect -1571 -15048 -1495 -15032
rect -1571 -15065 -1555 -15048
rect -1689 -15082 -1651 -15065
rect -1771 -15120 -1651 -15082
rect -1593 -15082 -1555 -15065
rect -1511 -15065 -1495 -15048
rect -1393 -15048 -1317 -15032
rect -1393 -15065 -1377 -15048
rect -1511 -15082 -1473 -15065
rect -1593 -15120 -1473 -15082
rect -1415 -15082 -1377 -15065
rect -1333 -15065 -1317 -15048
rect -1215 -15048 -1139 -15032
rect -1215 -15065 -1199 -15048
rect -1333 -15082 -1295 -15065
rect -1415 -15120 -1295 -15082
rect -1237 -15082 -1199 -15065
rect -1155 -15065 -1139 -15048
rect -1037 -15048 -961 -15032
rect -1037 -15065 -1021 -15048
rect -1155 -15082 -1117 -15065
rect -1237 -15120 -1117 -15082
rect -1059 -15082 -1021 -15065
rect -977 -15065 -961 -15048
rect -859 -15048 -783 -15032
rect -859 -15065 -843 -15048
rect -977 -15082 -939 -15065
rect -1059 -15120 -939 -15082
rect -881 -15082 -843 -15065
rect -799 -15065 -783 -15048
rect -681 -15048 -605 -15032
rect -681 -15065 -665 -15048
rect -799 -15082 -761 -15065
rect -881 -15120 -761 -15082
rect -703 -15082 -665 -15065
rect -621 -15065 -605 -15048
rect -503 -15048 -427 -15032
rect -503 -15065 -487 -15048
rect -621 -15082 -583 -15065
rect -703 -15120 -583 -15082
rect -525 -15082 -487 -15065
rect -443 -15065 -427 -15048
rect -325 -15048 -249 -15032
rect -325 -15065 -309 -15048
rect -443 -15082 -405 -15065
rect -525 -15120 -405 -15082
rect -347 -15082 -309 -15065
rect -265 -15065 -249 -15048
rect -147 -15048 -71 -15032
rect -147 -15065 -131 -15048
rect -265 -15082 -227 -15065
rect -347 -15120 -227 -15082
rect -169 -15082 -131 -15065
rect -87 -15065 -71 -15048
rect 31 -15048 107 -15032
rect 31 -15065 47 -15048
rect -87 -15082 -49 -15065
rect -169 -15120 -49 -15082
rect 9 -15082 47 -15065
rect 91 -15065 107 -15048
rect 209 -15048 285 -15032
rect 209 -15065 225 -15048
rect 91 -15082 129 -15065
rect 9 -15120 129 -15082
rect 187 -15082 225 -15065
rect 269 -15065 285 -15048
rect 387 -15048 463 -15032
rect 387 -15065 403 -15048
rect 269 -15082 307 -15065
rect 187 -15120 307 -15082
rect 365 -15082 403 -15065
rect 447 -15065 463 -15048
rect 565 -15048 641 -15032
rect 565 -15065 581 -15048
rect 447 -15082 485 -15065
rect 365 -15120 485 -15082
rect 543 -15082 581 -15065
rect 625 -15065 641 -15048
rect 743 -15048 819 -15032
rect 743 -15065 759 -15048
rect 625 -15082 663 -15065
rect 543 -15120 663 -15082
rect 721 -15082 759 -15065
rect 803 -15065 819 -15048
rect 921 -15048 997 -15032
rect 921 -15065 937 -15048
rect 803 -15082 841 -15065
rect 721 -15120 841 -15082
rect 899 -15082 937 -15065
rect 981 -15065 997 -15048
rect 1099 -15048 1175 -15032
rect 1099 -15065 1115 -15048
rect 981 -15082 1019 -15065
rect 899 -15120 1019 -15082
rect 1077 -15082 1115 -15065
rect 1159 -15065 1175 -15048
rect 1277 -15048 1353 -15032
rect 1277 -15065 1293 -15048
rect 1159 -15082 1197 -15065
rect 1077 -15120 1197 -15082
rect 1255 -15082 1293 -15065
rect 1337 -15065 1353 -15048
rect 1455 -15048 1531 -15032
rect 1455 -15065 1471 -15048
rect 1337 -15082 1375 -15065
rect 1255 -15120 1375 -15082
rect 1433 -15082 1471 -15065
rect 1515 -15065 1531 -15048
rect 1633 -15048 1709 -15032
rect 1633 -15065 1649 -15048
rect 1515 -15082 1553 -15065
rect 1433 -15120 1553 -15082
rect 1611 -15082 1649 -15065
rect 1693 -15065 1709 -15048
rect 1811 -15048 1887 -15032
rect 1811 -15065 1827 -15048
rect 1693 -15082 1731 -15065
rect 1611 -15120 1731 -15082
rect 1789 -15082 1827 -15065
rect 1871 -15065 1887 -15048
rect 1989 -15048 2065 -15032
rect 1989 -15065 2005 -15048
rect 1871 -15082 1909 -15065
rect 1789 -15120 1909 -15082
rect 1967 -15082 2005 -15065
rect 2049 -15065 2065 -15048
rect 2167 -15048 2243 -15032
rect 2167 -15065 2183 -15048
rect 2049 -15082 2087 -15065
rect 1967 -15120 2087 -15082
rect 2145 -15082 2183 -15065
rect 2227 -15065 2243 -15048
rect 2345 -15048 2421 -15032
rect 2345 -15065 2361 -15048
rect 2227 -15082 2265 -15065
rect 2145 -15120 2265 -15082
rect 2323 -15082 2361 -15065
rect 2405 -15065 2421 -15048
rect 2523 -15048 2599 -15032
rect 2523 -15065 2539 -15048
rect 2405 -15082 2443 -15065
rect 2323 -15120 2443 -15082
rect 2501 -15082 2539 -15065
rect 2583 -15065 2599 -15048
rect 2701 -15048 2777 -15032
rect 2701 -15065 2717 -15048
rect 2583 -15082 2621 -15065
rect 2501 -15120 2621 -15082
rect 2679 -15082 2717 -15065
rect 2761 -15065 2777 -15048
rect 2879 -15048 2955 -15032
rect 2879 -15065 2895 -15048
rect 2761 -15082 2799 -15065
rect 2679 -15120 2799 -15082
rect 2857 -15082 2895 -15065
rect 2939 -15065 2955 -15048
rect 3057 -15048 3133 -15032
rect 3057 -15065 3073 -15048
rect 2939 -15082 2977 -15065
rect 2857 -15120 2977 -15082
rect 3035 -15082 3073 -15065
rect 3117 -15065 3133 -15048
rect 3235 -15048 3311 -15032
rect 3235 -15065 3251 -15048
rect 3117 -15082 3155 -15065
rect 3035 -15120 3155 -15082
rect 3213 -15082 3251 -15065
rect 3295 -15065 3311 -15048
rect 3413 -15048 3489 -15032
rect 3413 -15065 3429 -15048
rect 3295 -15082 3333 -15065
rect 3213 -15120 3333 -15082
rect 3391 -15082 3429 -15065
rect 3473 -15065 3489 -15048
rect 3591 -15048 3667 -15032
rect 3591 -15065 3607 -15048
rect 3473 -15082 3511 -15065
rect 3391 -15120 3511 -15082
rect 3569 -15082 3607 -15065
rect 3651 -15065 3667 -15048
rect 3769 -15048 3845 -15032
rect 3769 -15065 3785 -15048
rect 3651 -15082 3689 -15065
rect 3569 -15120 3689 -15082
rect 3747 -15082 3785 -15065
rect 3829 -15065 3845 -15048
rect 3947 -15048 4023 -15032
rect 3947 -15065 3963 -15048
rect 3829 -15082 3867 -15065
rect 3747 -15120 3867 -15082
rect 3925 -15082 3963 -15065
rect 4007 -15065 4023 -15048
rect 5645 -15048 5721 -15032
rect 5645 -15065 5661 -15048
rect 4007 -15082 4045 -15065
rect 3925 -15120 4045 -15082
rect 5623 -15082 5661 -15065
rect 5705 -15065 5721 -15048
rect 5823 -15048 5899 -15032
rect 5823 -15065 5839 -15048
rect 5705 -15082 5743 -15065
rect 5623 -15120 5743 -15082
rect 5801 -15082 5839 -15065
rect 5883 -15065 5899 -15048
rect 6001 -15048 6077 -15032
rect 6001 -15065 6017 -15048
rect 5883 -15082 5921 -15065
rect 5801 -15120 5921 -15082
rect 5979 -15082 6017 -15065
rect 6061 -15065 6077 -15048
rect 6179 -15048 6255 -15032
rect 6179 -15065 6195 -15048
rect 6061 -15082 6099 -15065
rect 5979 -15120 6099 -15082
rect 6157 -15082 6195 -15065
rect 6239 -15065 6255 -15048
rect 6357 -15048 6433 -15032
rect 6357 -15065 6373 -15048
rect 6239 -15082 6277 -15065
rect 6157 -15120 6277 -15082
rect 6335 -15082 6373 -15065
rect 6417 -15065 6433 -15048
rect 6535 -15048 6611 -15032
rect 6535 -15065 6551 -15048
rect 6417 -15082 6455 -15065
rect 6335 -15120 6455 -15082
rect 6513 -15082 6551 -15065
rect 6595 -15065 6611 -15048
rect 6713 -15048 6789 -15032
rect 6713 -15065 6729 -15048
rect 6595 -15082 6633 -15065
rect 6513 -15120 6633 -15082
rect 6691 -15082 6729 -15065
rect 6773 -15065 6789 -15048
rect 6891 -15048 6967 -15032
rect 6891 -15065 6907 -15048
rect 6773 -15082 6811 -15065
rect 6691 -15120 6811 -15082
rect 6869 -15082 6907 -15065
rect 6951 -15065 6967 -15048
rect 7069 -15048 7145 -15032
rect 7069 -15065 7085 -15048
rect 6951 -15082 6989 -15065
rect 6869 -15120 6989 -15082
rect 7047 -15082 7085 -15065
rect 7129 -15065 7145 -15048
rect 7247 -15048 7323 -15032
rect 7247 -15065 7263 -15048
rect 7129 -15082 7167 -15065
rect 7047 -15120 7167 -15082
rect 7225 -15082 7263 -15065
rect 7307 -15065 7323 -15048
rect 7425 -15048 7501 -15032
rect 7425 -15065 7441 -15048
rect 7307 -15082 7345 -15065
rect 7225 -15120 7345 -15082
rect 7403 -15082 7441 -15065
rect 7485 -15065 7501 -15048
rect 7603 -15048 7679 -15032
rect 7603 -15065 7619 -15048
rect 7485 -15082 7523 -15065
rect 7403 -15120 7523 -15082
rect 7581 -15082 7619 -15065
rect 7663 -15065 7679 -15048
rect 7781 -15048 7857 -15032
rect 7781 -15065 7797 -15048
rect 7663 -15082 7701 -15065
rect 7581 -15120 7701 -15082
rect 7759 -15082 7797 -15065
rect 7841 -15065 7857 -15048
rect 7959 -15048 8035 -15032
rect 7959 -15065 7975 -15048
rect 7841 -15082 7879 -15065
rect 7759 -15120 7879 -15082
rect 7937 -15082 7975 -15065
rect 8019 -15065 8035 -15048
rect 8137 -15048 8213 -15032
rect 8137 -15065 8153 -15048
rect 8019 -15082 8057 -15065
rect 7937 -15120 8057 -15082
rect 8115 -15082 8153 -15065
rect 8197 -15065 8213 -15048
rect 8315 -15048 8391 -15032
rect 8315 -15065 8331 -15048
rect 8197 -15082 8235 -15065
rect 8115 -15120 8235 -15082
rect 8293 -15082 8331 -15065
rect 8375 -15065 8391 -15048
rect 8493 -15048 8569 -15032
rect 8493 -15065 8509 -15048
rect 8375 -15082 8413 -15065
rect 8293 -15120 8413 -15082
rect 8471 -15082 8509 -15065
rect 8553 -15065 8569 -15048
rect 8671 -15048 8747 -15032
rect 8671 -15065 8687 -15048
rect 8553 -15082 8591 -15065
rect 8471 -15120 8591 -15082
rect 8649 -15082 8687 -15065
rect 8731 -15065 8747 -15048
rect 8849 -15048 8925 -15032
rect 8849 -15065 8865 -15048
rect 8731 -15082 8769 -15065
rect 8649 -15120 8769 -15082
rect 8827 -15082 8865 -15065
rect 8909 -15065 8925 -15048
rect 9027 -15048 9103 -15032
rect 9027 -15065 9043 -15048
rect 8909 -15082 8947 -15065
rect 8827 -15120 8947 -15082
rect 9005 -15082 9043 -15065
rect 9087 -15065 9103 -15048
rect 9205 -15048 9281 -15032
rect 9205 -15065 9221 -15048
rect 9087 -15082 9125 -15065
rect 9005 -15120 9125 -15082
rect 9183 -15082 9221 -15065
rect 9265 -15065 9281 -15048
rect 9383 -15048 9459 -15032
rect 9383 -15065 9399 -15048
rect 9265 -15082 9303 -15065
rect 9183 -15120 9303 -15082
rect 9361 -15082 9399 -15065
rect 9443 -15065 9459 -15048
rect 9561 -15048 9637 -15032
rect 9561 -15065 9577 -15048
rect 9443 -15082 9481 -15065
rect 9361 -15120 9481 -15082
rect 9539 -15082 9577 -15065
rect 9621 -15065 9637 -15048
rect 9739 -15048 9815 -15032
rect 9739 -15065 9755 -15048
rect 9621 -15082 9659 -15065
rect 9539 -15120 9659 -15082
rect 9717 -15082 9755 -15065
rect 9799 -15065 9815 -15048
rect 9917 -15048 9993 -15032
rect 9917 -15065 9933 -15048
rect 9799 -15082 9837 -15065
rect 9717 -15120 9837 -15082
rect 9895 -15082 9933 -15065
rect 9977 -15065 9993 -15048
rect 10095 -15048 10171 -15032
rect 10095 -15065 10111 -15048
rect 9977 -15082 10015 -15065
rect 9895 -15120 10015 -15082
rect 10073 -15082 10111 -15065
rect 10155 -15065 10171 -15048
rect 10273 -15048 10349 -15032
rect 10273 -15065 10289 -15048
rect 10155 -15082 10193 -15065
rect 10073 -15120 10193 -15082
rect 10251 -15082 10289 -15065
rect 10333 -15065 10349 -15048
rect 10451 -15048 10527 -15032
rect 10451 -15065 10467 -15048
rect 10333 -15082 10371 -15065
rect 10251 -15120 10371 -15082
rect 10429 -15082 10467 -15065
rect 10511 -15065 10527 -15048
rect 10629 -15048 10705 -15032
rect 10629 -15065 10645 -15048
rect 10511 -15082 10549 -15065
rect 10429 -15120 10549 -15082
rect 10607 -15082 10645 -15065
rect 10689 -15065 10705 -15048
rect 10807 -15048 10883 -15032
rect 10807 -15065 10823 -15048
rect 10689 -15082 10727 -15065
rect 10607 -15120 10727 -15082
rect 10785 -15082 10823 -15065
rect 10867 -15065 10883 -15048
rect 10985 -15048 11061 -15032
rect 10985 -15065 11001 -15048
rect 10867 -15082 10905 -15065
rect 10785 -15120 10905 -15082
rect 10963 -15082 11001 -15065
rect 11045 -15065 11061 -15048
rect 11163 -15048 11239 -15032
rect 11163 -15065 11179 -15048
rect 11045 -15082 11083 -15065
rect 10963 -15120 11083 -15082
rect 11141 -15082 11179 -15065
rect 11223 -15065 11239 -15048
rect 11341 -15048 11417 -15032
rect 11341 -15065 11357 -15048
rect 11223 -15082 11261 -15065
rect 11141 -15120 11261 -15082
rect 11319 -15082 11357 -15065
rect 11401 -15065 11417 -15048
rect 11519 -15048 11595 -15032
rect 11519 -15065 11535 -15048
rect 11401 -15082 11439 -15065
rect 11319 -15120 11439 -15082
rect 11497 -15082 11535 -15065
rect 11579 -15065 11595 -15048
rect 11697 -15048 11773 -15032
rect 11697 -15065 11713 -15048
rect 11579 -15082 11617 -15065
rect 11497 -15120 11617 -15082
rect 11675 -15082 11713 -15065
rect 11757 -15065 11773 -15048
rect 11875 -15048 11951 -15032
rect 11875 -15065 11891 -15048
rect 11757 -15082 11795 -15065
rect 11675 -15120 11795 -15082
rect 11853 -15082 11891 -15065
rect 11935 -15065 11951 -15048
rect 12053 -15048 12129 -15032
rect 12053 -15065 12069 -15048
rect 11935 -15082 11973 -15065
rect 11853 -15120 11973 -15082
rect 12031 -15082 12069 -15065
rect 12113 -15065 12129 -15048
rect 12231 -15048 12307 -15032
rect 12231 -15065 12247 -15048
rect 12113 -15082 12151 -15065
rect 12031 -15120 12151 -15082
rect 12209 -15082 12247 -15065
rect 12291 -15065 12307 -15048
rect 12409 -15048 12485 -15032
rect 12409 -15065 12425 -15048
rect 12291 -15082 12329 -15065
rect 12209 -15120 12329 -15082
rect 12387 -15082 12425 -15065
rect 12469 -15065 12485 -15048
rect 12587 -15048 12663 -15032
rect 12587 -15065 12603 -15048
rect 12469 -15082 12507 -15065
rect 12387 -15120 12507 -15082
rect 12565 -15082 12603 -15065
rect 12647 -15065 12663 -15048
rect 12647 -15082 12685 -15065
rect 12565 -15120 12685 -15082
rect -5982 -15400 -5862 -15362
rect -5982 -15417 -5944 -15400
rect -5960 -15434 -5944 -15417
rect -5900 -15417 -5862 -15400
rect -5804 -15400 -5684 -15362
rect -5804 -15417 -5766 -15400
rect -5900 -15434 -5884 -15417
rect -5960 -15450 -5884 -15434
rect -5782 -15434 -5766 -15417
rect -5722 -15417 -5684 -15400
rect -5626 -15400 -5506 -15362
rect -5626 -15417 -5588 -15400
rect -5722 -15434 -5706 -15417
rect -5782 -15450 -5706 -15434
rect -5604 -15434 -5588 -15417
rect -5544 -15417 -5506 -15400
rect -5448 -15400 -5328 -15362
rect -5448 -15417 -5410 -15400
rect -5544 -15434 -5528 -15417
rect -5604 -15450 -5528 -15434
rect -5426 -15434 -5410 -15417
rect -5366 -15417 -5328 -15400
rect -5270 -15400 -5150 -15362
rect -5270 -15417 -5232 -15400
rect -5366 -15434 -5350 -15417
rect -5426 -15450 -5350 -15434
rect -5248 -15434 -5232 -15417
rect -5188 -15417 -5150 -15400
rect -5092 -15400 -4972 -15362
rect -5092 -15417 -5054 -15400
rect -5188 -15434 -5172 -15417
rect -5248 -15450 -5172 -15434
rect -5070 -15434 -5054 -15417
rect -5010 -15417 -4972 -15400
rect -4914 -15400 -4794 -15362
rect -4914 -15417 -4876 -15400
rect -5010 -15434 -4994 -15417
rect -5070 -15450 -4994 -15434
rect -4892 -15434 -4876 -15417
rect -4832 -15417 -4794 -15400
rect -4736 -15400 -4616 -15362
rect -4736 -15417 -4698 -15400
rect -4832 -15434 -4816 -15417
rect -4892 -15450 -4816 -15434
rect -4714 -15434 -4698 -15417
rect -4654 -15417 -4616 -15400
rect -4558 -15400 -4438 -15362
rect -4558 -15417 -4520 -15400
rect -4654 -15434 -4638 -15417
rect -4714 -15450 -4638 -15434
rect -4536 -15434 -4520 -15417
rect -4476 -15417 -4438 -15400
rect -4380 -15400 -4260 -15362
rect -4380 -15417 -4342 -15400
rect -4476 -15434 -4460 -15417
rect -4536 -15450 -4460 -15434
rect -4358 -15434 -4342 -15417
rect -4298 -15417 -4260 -15400
rect -4202 -15400 -4082 -15362
rect -4202 -15417 -4164 -15400
rect -4298 -15434 -4282 -15417
rect -4358 -15450 -4282 -15434
rect -4180 -15434 -4164 -15417
rect -4120 -15417 -4082 -15400
rect -4120 -15434 -4104 -15417
rect -4180 -15450 -4104 -15434
rect -2127 -15438 -2007 -15400
rect -2127 -15455 -2089 -15438
rect -2105 -15472 -2089 -15455
rect -2045 -15455 -2007 -15438
rect -1949 -15438 -1829 -15400
rect -1949 -15455 -1911 -15438
rect -2045 -15472 -2029 -15455
rect -2105 -15488 -2029 -15472
rect -1927 -15472 -1911 -15455
rect -1867 -15455 -1829 -15438
rect -1771 -15438 -1651 -15400
rect -1771 -15455 -1733 -15438
rect -1867 -15472 -1851 -15455
rect -1927 -15488 -1851 -15472
rect -1749 -15472 -1733 -15455
rect -1689 -15455 -1651 -15438
rect -1593 -15438 -1473 -15400
rect -1593 -15455 -1555 -15438
rect -1689 -15472 -1673 -15455
rect -1749 -15488 -1673 -15472
rect -1571 -15472 -1555 -15455
rect -1511 -15455 -1473 -15438
rect -1415 -15438 -1295 -15400
rect -1415 -15455 -1377 -15438
rect -1511 -15472 -1495 -15455
rect -1571 -15488 -1495 -15472
rect -1393 -15472 -1377 -15455
rect -1333 -15455 -1295 -15438
rect -1237 -15438 -1117 -15400
rect -1237 -15455 -1199 -15438
rect -1333 -15472 -1317 -15455
rect -1393 -15488 -1317 -15472
rect -1215 -15472 -1199 -15455
rect -1155 -15455 -1117 -15438
rect -1059 -15438 -939 -15400
rect -1059 -15455 -1021 -15438
rect -1155 -15472 -1139 -15455
rect -1215 -15488 -1139 -15472
rect -1037 -15472 -1021 -15455
rect -977 -15455 -939 -15438
rect -881 -15438 -761 -15400
rect -881 -15455 -843 -15438
rect -977 -15472 -961 -15455
rect -1037 -15488 -961 -15472
rect -859 -15472 -843 -15455
rect -799 -15455 -761 -15438
rect -703 -15438 -583 -15400
rect -703 -15455 -665 -15438
rect -799 -15472 -783 -15455
rect -859 -15488 -783 -15472
rect -681 -15472 -665 -15455
rect -621 -15455 -583 -15438
rect -525 -15438 -405 -15400
rect -525 -15455 -487 -15438
rect -621 -15472 -605 -15455
rect -681 -15488 -605 -15472
rect -503 -15472 -487 -15455
rect -443 -15455 -405 -15438
rect -347 -15438 -227 -15400
rect -347 -15455 -309 -15438
rect -443 -15472 -427 -15455
rect -503 -15488 -427 -15472
rect -325 -15472 -309 -15455
rect -265 -15455 -227 -15438
rect -169 -15438 -49 -15400
rect -169 -15455 -131 -15438
rect -265 -15472 -249 -15455
rect -325 -15488 -249 -15472
rect -147 -15472 -131 -15455
rect -87 -15455 -49 -15438
rect 9 -15438 129 -15400
rect 9 -15455 47 -15438
rect -87 -15472 -71 -15455
rect -147 -15488 -71 -15472
rect 31 -15472 47 -15455
rect 91 -15455 129 -15438
rect 187 -15438 307 -15400
rect 187 -15455 225 -15438
rect 91 -15472 107 -15455
rect 31 -15488 107 -15472
rect 209 -15472 225 -15455
rect 269 -15455 307 -15438
rect 365 -15438 485 -15400
rect 365 -15455 403 -15438
rect 269 -15472 285 -15455
rect 209 -15488 285 -15472
rect 387 -15472 403 -15455
rect 447 -15455 485 -15438
rect 543 -15438 663 -15400
rect 543 -15455 581 -15438
rect 447 -15472 463 -15455
rect 387 -15488 463 -15472
rect 565 -15472 581 -15455
rect 625 -15455 663 -15438
rect 721 -15438 841 -15400
rect 721 -15455 759 -15438
rect 625 -15472 641 -15455
rect 565 -15488 641 -15472
rect 743 -15472 759 -15455
rect 803 -15455 841 -15438
rect 899 -15438 1019 -15400
rect 899 -15455 937 -15438
rect 803 -15472 819 -15455
rect 743 -15488 819 -15472
rect 921 -15472 937 -15455
rect 981 -15455 1019 -15438
rect 1077 -15438 1197 -15400
rect 1077 -15455 1115 -15438
rect 981 -15472 997 -15455
rect 921 -15488 997 -15472
rect 1099 -15472 1115 -15455
rect 1159 -15455 1197 -15438
rect 1255 -15438 1375 -15400
rect 1255 -15455 1293 -15438
rect 1159 -15472 1175 -15455
rect 1099 -15488 1175 -15472
rect 1277 -15472 1293 -15455
rect 1337 -15455 1375 -15438
rect 1433 -15438 1553 -15400
rect 1433 -15455 1471 -15438
rect 1337 -15472 1353 -15455
rect 1277 -15488 1353 -15472
rect 1455 -15472 1471 -15455
rect 1515 -15455 1553 -15438
rect 1611 -15438 1731 -15400
rect 1611 -15455 1649 -15438
rect 1515 -15472 1531 -15455
rect 1455 -15488 1531 -15472
rect 1633 -15472 1649 -15455
rect 1693 -15455 1731 -15438
rect 1789 -15438 1909 -15400
rect 1789 -15455 1827 -15438
rect 1693 -15472 1709 -15455
rect 1633 -15488 1709 -15472
rect 1811 -15472 1827 -15455
rect 1871 -15455 1909 -15438
rect 1967 -15438 2087 -15400
rect 1967 -15455 2005 -15438
rect 1871 -15472 1887 -15455
rect 1811 -15488 1887 -15472
rect 1989 -15472 2005 -15455
rect 2049 -15455 2087 -15438
rect 2145 -15438 2265 -15400
rect 2145 -15455 2183 -15438
rect 2049 -15472 2065 -15455
rect 1989 -15488 2065 -15472
rect 2167 -15472 2183 -15455
rect 2227 -15455 2265 -15438
rect 2323 -15438 2443 -15400
rect 2323 -15455 2361 -15438
rect 2227 -15472 2243 -15455
rect 2167 -15488 2243 -15472
rect 2345 -15472 2361 -15455
rect 2405 -15455 2443 -15438
rect 2501 -15438 2621 -15400
rect 2501 -15455 2539 -15438
rect 2405 -15472 2421 -15455
rect 2345 -15488 2421 -15472
rect 2523 -15472 2539 -15455
rect 2583 -15455 2621 -15438
rect 2679 -15438 2799 -15400
rect 2679 -15455 2717 -15438
rect 2583 -15472 2599 -15455
rect 2523 -15488 2599 -15472
rect 2701 -15472 2717 -15455
rect 2761 -15455 2799 -15438
rect 2857 -15438 2977 -15400
rect 2857 -15455 2895 -15438
rect 2761 -15472 2777 -15455
rect 2701 -15488 2777 -15472
rect 2879 -15472 2895 -15455
rect 2939 -15455 2977 -15438
rect 3035 -15438 3155 -15400
rect 3035 -15455 3073 -15438
rect 2939 -15472 2955 -15455
rect 2879 -15488 2955 -15472
rect 3057 -15472 3073 -15455
rect 3117 -15455 3155 -15438
rect 3213 -15438 3333 -15400
rect 3213 -15455 3251 -15438
rect 3117 -15472 3133 -15455
rect 3057 -15488 3133 -15472
rect 3235 -15472 3251 -15455
rect 3295 -15455 3333 -15438
rect 3391 -15438 3511 -15400
rect 3391 -15455 3429 -15438
rect 3295 -15472 3311 -15455
rect 3235 -15488 3311 -15472
rect 3413 -15472 3429 -15455
rect 3473 -15455 3511 -15438
rect 3569 -15438 3689 -15400
rect 3569 -15455 3607 -15438
rect 3473 -15472 3489 -15455
rect 3413 -15488 3489 -15472
rect 3591 -15472 3607 -15455
rect 3651 -15455 3689 -15438
rect 3747 -15438 3867 -15400
rect 3747 -15455 3785 -15438
rect 3651 -15472 3667 -15455
rect 3591 -15488 3667 -15472
rect 3769 -15472 3785 -15455
rect 3829 -15455 3867 -15438
rect 3925 -15438 4045 -15400
rect 3925 -15455 3963 -15438
rect 3829 -15472 3845 -15455
rect 3769 -15488 3845 -15472
rect 3947 -15472 3963 -15455
rect 4007 -15455 4045 -15438
rect 5623 -15438 5743 -15400
rect 5623 -15455 5661 -15438
rect 4007 -15472 4023 -15455
rect 3947 -15488 4023 -15472
rect 5645 -15472 5661 -15455
rect 5705 -15455 5743 -15438
rect 5801 -15438 5921 -15400
rect 5801 -15455 5839 -15438
rect 5705 -15472 5721 -15455
rect 5645 -15488 5721 -15472
rect 5823 -15472 5839 -15455
rect 5883 -15455 5921 -15438
rect 5979 -15438 6099 -15400
rect 5979 -15455 6017 -15438
rect 5883 -15472 5899 -15455
rect 5823 -15488 5899 -15472
rect 6001 -15472 6017 -15455
rect 6061 -15455 6099 -15438
rect 6157 -15438 6277 -15400
rect 6157 -15455 6195 -15438
rect 6061 -15472 6077 -15455
rect 6001 -15488 6077 -15472
rect 6179 -15472 6195 -15455
rect 6239 -15455 6277 -15438
rect 6335 -15438 6455 -15400
rect 6335 -15455 6373 -15438
rect 6239 -15472 6255 -15455
rect 6179 -15488 6255 -15472
rect 6357 -15472 6373 -15455
rect 6417 -15455 6455 -15438
rect 6513 -15438 6633 -15400
rect 6513 -15455 6551 -15438
rect 6417 -15472 6433 -15455
rect 6357 -15488 6433 -15472
rect 6535 -15472 6551 -15455
rect 6595 -15455 6633 -15438
rect 6691 -15438 6811 -15400
rect 6691 -15455 6729 -15438
rect 6595 -15472 6611 -15455
rect 6535 -15488 6611 -15472
rect 6713 -15472 6729 -15455
rect 6773 -15455 6811 -15438
rect 6869 -15438 6989 -15400
rect 6869 -15455 6907 -15438
rect 6773 -15472 6789 -15455
rect 6713 -15488 6789 -15472
rect 6891 -15472 6907 -15455
rect 6951 -15455 6989 -15438
rect 7047 -15438 7167 -15400
rect 7047 -15455 7085 -15438
rect 6951 -15472 6967 -15455
rect 6891 -15488 6967 -15472
rect 7069 -15472 7085 -15455
rect 7129 -15455 7167 -15438
rect 7225 -15438 7345 -15400
rect 7225 -15455 7263 -15438
rect 7129 -15472 7145 -15455
rect 7069 -15488 7145 -15472
rect 7247 -15472 7263 -15455
rect 7307 -15455 7345 -15438
rect 7403 -15438 7523 -15400
rect 7403 -15455 7441 -15438
rect 7307 -15472 7323 -15455
rect 7247 -15488 7323 -15472
rect 7425 -15472 7441 -15455
rect 7485 -15455 7523 -15438
rect 7581 -15438 7701 -15400
rect 7581 -15455 7619 -15438
rect 7485 -15472 7501 -15455
rect 7425 -15488 7501 -15472
rect 7603 -15472 7619 -15455
rect 7663 -15455 7701 -15438
rect 7759 -15438 7879 -15400
rect 7759 -15455 7797 -15438
rect 7663 -15472 7679 -15455
rect 7603 -15488 7679 -15472
rect 7781 -15472 7797 -15455
rect 7841 -15455 7879 -15438
rect 7937 -15438 8057 -15400
rect 7937 -15455 7975 -15438
rect 7841 -15472 7857 -15455
rect 7781 -15488 7857 -15472
rect 7959 -15472 7975 -15455
rect 8019 -15455 8057 -15438
rect 8115 -15438 8235 -15400
rect 8115 -15455 8153 -15438
rect 8019 -15472 8035 -15455
rect 7959 -15488 8035 -15472
rect 8137 -15472 8153 -15455
rect 8197 -15455 8235 -15438
rect 8293 -15438 8413 -15400
rect 8293 -15455 8331 -15438
rect 8197 -15472 8213 -15455
rect 8137 -15488 8213 -15472
rect 8315 -15472 8331 -15455
rect 8375 -15455 8413 -15438
rect 8471 -15438 8591 -15400
rect 8471 -15455 8509 -15438
rect 8375 -15472 8391 -15455
rect 8315 -15488 8391 -15472
rect 8493 -15472 8509 -15455
rect 8553 -15455 8591 -15438
rect 8649 -15438 8769 -15400
rect 8649 -15455 8687 -15438
rect 8553 -15472 8569 -15455
rect 8493 -15488 8569 -15472
rect 8671 -15472 8687 -15455
rect 8731 -15455 8769 -15438
rect 8827 -15438 8947 -15400
rect 8827 -15455 8865 -15438
rect 8731 -15472 8747 -15455
rect 8671 -15488 8747 -15472
rect 8849 -15472 8865 -15455
rect 8909 -15455 8947 -15438
rect 9005 -15438 9125 -15400
rect 9005 -15455 9043 -15438
rect 8909 -15472 8925 -15455
rect 8849 -15488 8925 -15472
rect 9027 -15472 9043 -15455
rect 9087 -15455 9125 -15438
rect 9183 -15438 9303 -15400
rect 9183 -15455 9221 -15438
rect 9087 -15472 9103 -15455
rect 9027 -15488 9103 -15472
rect 9205 -15472 9221 -15455
rect 9265 -15455 9303 -15438
rect 9361 -15438 9481 -15400
rect 9361 -15455 9399 -15438
rect 9265 -15472 9281 -15455
rect 9205 -15488 9281 -15472
rect 9383 -15472 9399 -15455
rect 9443 -15455 9481 -15438
rect 9539 -15438 9659 -15400
rect 9539 -15455 9577 -15438
rect 9443 -15472 9459 -15455
rect 9383 -15488 9459 -15472
rect 9561 -15472 9577 -15455
rect 9621 -15455 9659 -15438
rect 9717 -15438 9837 -15400
rect 9717 -15455 9755 -15438
rect 9621 -15472 9637 -15455
rect 9561 -15488 9637 -15472
rect 9739 -15472 9755 -15455
rect 9799 -15455 9837 -15438
rect 9895 -15438 10015 -15400
rect 9895 -15455 9933 -15438
rect 9799 -15472 9815 -15455
rect 9739 -15488 9815 -15472
rect 9917 -15472 9933 -15455
rect 9977 -15455 10015 -15438
rect 10073 -15438 10193 -15400
rect 10073 -15455 10111 -15438
rect 9977 -15472 9993 -15455
rect 9917 -15488 9993 -15472
rect 10095 -15472 10111 -15455
rect 10155 -15455 10193 -15438
rect 10251 -15438 10371 -15400
rect 10251 -15455 10289 -15438
rect 10155 -15472 10171 -15455
rect 10095 -15488 10171 -15472
rect 10273 -15472 10289 -15455
rect 10333 -15455 10371 -15438
rect 10429 -15438 10549 -15400
rect 10429 -15455 10467 -15438
rect 10333 -15472 10349 -15455
rect 10273 -15488 10349 -15472
rect 10451 -15472 10467 -15455
rect 10511 -15455 10549 -15438
rect 10607 -15438 10727 -15400
rect 10607 -15455 10645 -15438
rect 10511 -15472 10527 -15455
rect 10451 -15488 10527 -15472
rect 10629 -15472 10645 -15455
rect 10689 -15455 10727 -15438
rect 10785 -15438 10905 -15400
rect 10785 -15455 10823 -15438
rect 10689 -15472 10705 -15455
rect 10629 -15488 10705 -15472
rect 10807 -15472 10823 -15455
rect 10867 -15455 10905 -15438
rect 10963 -15438 11083 -15400
rect 10963 -15455 11001 -15438
rect 10867 -15472 10883 -15455
rect 10807 -15488 10883 -15472
rect 10985 -15472 11001 -15455
rect 11045 -15455 11083 -15438
rect 11141 -15438 11261 -15400
rect 11141 -15455 11179 -15438
rect 11045 -15472 11061 -15455
rect 10985 -15488 11061 -15472
rect 11163 -15472 11179 -15455
rect 11223 -15455 11261 -15438
rect 11319 -15438 11439 -15400
rect 11319 -15455 11357 -15438
rect 11223 -15472 11239 -15455
rect 11163 -15488 11239 -15472
rect 11341 -15472 11357 -15455
rect 11401 -15455 11439 -15438
rect 11497 -15438 11617 -15400
rect 11497 -15455 11535 -15438
rect 11401 -15472 11417 -15455
rect 11341 -15488 11417 -15472
rect 11519 -15472 11535 -15455
rect 11579 -15455 11617 -15438
rect 11675 -15438 11795 -15400
rect 11675 -15455 11713 -15438
rect 11579 -15472 11595 -15455
rect 11519 -15488 11595 -15472
rect 11697 -15472 11713 -15455
rect 11757 -15455 11795 -15438
rect 11853 -15438 11973 -15400
rect 11853 -15455 11891 -15438
rect 11757 -15472 11773 -15455
rect 11697 -15488 11773 -15472
rect 11875 -15472 11891 -15455
rect 11935 -15455 11973 -15438
rect 12031 -15438 12151 -15400
rect 12031 -15455 12069 -15438
rect 11935 -15472 11951 -15455
rect 11875 -15488 11951 -15472
rect 12053 -15472 12069 -15455
rect 12113 -15455 12151 -15438
rect 12209 -15438 12329 -15400
rect 12209 -15455 12247 -15438
rect 12113 -15472 12129 -15455
rect 12053 -15488 12129 -15472
rect 12231 -15472 12247 -15455
rect 12291 -15455 12329 -15438
rect 12387 -15438 12507 -15400
rect 12387 -15455 12425 -15438
rect 12291 -15472 12307 -15455
rect 12231 -15488 12307 -15472
rect 12409 -15472 12425 -15455
rect 12469 -15455 12507 -15438
rect 12565 -15438 12685 -15400
rect 12565 -15455 12603 -15438
rect 12469 -15472 12485 -15455
rect 12409 -15488 12485 -15472
rect 12587 -15472 12603 -15455
rect 12647 -15455 12685 -15438
rect 12647 -15472 12663 -15455
rect 12587 -15488 12663 -15472
rect -5960 -15710 -5884 -15694
rect -5960 -15727 -5944 -15710
rect -5982 -15744 -5944 -15727
rect -5900 -15727 -5884 -15710
rect -5782 -15710 -5706 -15694
rect -5782 -15727 -5766 -15710
rect -5900 -15744 -5862 -15727
rect -5982 -15782 -5862 -15744
rect -5804 -15744 -5766 -15727
rect -5722 -15727 -5706 -15710
rect -5604 -15710 -5528 -15694
rect -5604 -15727 -5588 -15710
rect -5722 -15744 -5684 -15727
rect -5804 -15782 -5684 -15744
rect -5626 -15744 -5588 -15727
rect -5544 -15727 -5528 -15710
rect -5426 -15710 -5350 -15694
rect -5426 -15727 -5410 -15710
rect -5544 -15744 -5506 -15727
rect -5626 -15782 -5506 -15744
rect -5448 -15744 -5410 -15727
rect -5366 -15727 -5350 -15710
rect -5248 -15710 -5172 -15694
rect -5248 -15727 -5232 -15710
rect -5366 -15744 -5328 -15727
rect -5448 -15782 -5328 -15744
rect -5270 -15744 -5232 -15727
rect -5188 -15727 -5172 -15710
rect -5070 -15710 -4994 -15694
rect -5070 -15727 -5054 -15710
rect -5188 -15744 -5150 -15727
rect -5270 -15782 -5150 -15744
rect -5092 -15744 -5054 -15727
rect -5010 -15727 -4994 -15710
rect -4892 -15710 -4816 -15694
rect -4892 -15727 -4876 -15710
rect -5010 -15744 -4972 -15727
rect -5092 -15782 -4972 -15744
rect -4914 -15744 -4876 -15727
rect -4832 -15727 -4816 -15710
rect -4714 -15710 -4638 -15694
rect -4714 -15727 -4698 -15710
rect -4832 -15744 -4794 -15727
rect -4914 -15782 -4794 -15744
rect -4736 -15744 -4698 -15727
rect -4654 -15727 -4638 -15710
rect -4536 -15710 -4460 -15694
rect -4536 -15727 -4520 -15710
rect -4654 -15744 -4616 -15727
rect -4736 -15782 -4616 -15744
rect -4558 -15744 -4520 -15727
rect -4476 -15727 -4460 -15710
rect -4358 -15710 -4282 -15694
rect -4358 -15727 -4342 -15710
rect -4476 -15744 -4438 -15727
rect -4558 -15782 -4438 -15744
rect -4380 -15744 -4342 -15727
rect -4298 -15727 -4282 -15710
rect -4180 -15710 -4104 -15694
rect -4180 -15727 -4164 -15710
rect -4298 -15744 -4260 -15727
rect -4380 -15782 -4260 -15744
rect -4202 -15744 -4164 -15727
rect -4120 -15727 -4104 -15710
rect -4120 -15744 -4082 -15727
rect -4202 -15782 -4082 -15744
rect -2105 -16048 -2029 -16032
rect -5982 -16100 -5862 -16062
rect -5982 -16117 -5944 -16100
rect -5960 -16134 -5944 -16117
rect -5900 -16117 -5862 -16100
rect -5804 -16100 -5684 -16062
rect -5804 -16117 -5766 -16100
rect -5900 -16134 -5884 -16117
rect -5960 -16150 -5884 -16134
rect -5782 -16134 -5766 -16117
rect -5722 -16117 -5684 -16100
rect -5626 -16100 -5506 -16062
rect -5626 -16117 -5588 -16100
rect -5722 -16134 -5706 -16117
rect -5782 -16150 -5706 -16134
rect -5604 -16134 -5588 -16117
rect -5544 -16117 -5506 -16100
rect -5448 -16100 -5328 -16062
rect -5448 -16117 -5410 -16100
rect -5544 -16134 -5528 -16117
rect -5604 -16150 -5528 -16134
rect -5426 -16134 -5410 -16117
rect -5366 -16117 -5328 -16100
rect -5270 -16100 -5150 -16062
rect -5270 -16117 -5232 -16100
rect -5366 -16134 -5350 -16117
rect -5426 -16150 -5350 -16134
rect -5248 -16134 -5232 -16117
rect -5188 -16117 -5150 -16100
rect -5092 -16100 -4972 -16062
rect -5092 -16117 -5054 -16100
rect -5188 -16134 -5172 -16117
rect -5248 -16150 -5172 -16134
rect -5070 -16134 -5054 -16117
rect -5010 -16117 -4972 -16100
rect -4914 -16100 -4794 -16062
rect -4914 -16117 -4876 -16100
rect -5010 -16134 -4994 -16117
rect -5070 -16150 -4994 -16134
rect -4892 -16134 -4876 -16117
rect -4832 -16117 -4794 -16100
rect -4736 -16100 -4616 -16062
rect -4736 -16117 -4698 -16100
rect -4832 -16134 -4816 -16117
rect -4892 -16150 -4816 -16134
rect -4714 -16134 -4698 -16117
rect -4654 -16117 -4616 -16100
rect -4558 -16100 -4438 -16062
rect -4558 -16117 -4520 -16100
rect -4654 -16134 -4638 -16117
rect -4714 -16150 -4638 -16134
rect -4536 -16134 -4520 -16117
rect -4476 -16117 -4438 -16100
rect -4380 -16100 -4260 -16062
rect -4380 -16117 -4342 -16100
rect -4476 -16134 -4460 -16117
rect -4536 -16150 -4460 -16134
rect -4358 -16134 -4342 -16117
rect -4298 -16117 -4260 -16100
rect -4202 -16100 -4082 -16062
rect -2105 -16065 -2089 -16048
rect -4202 -16117 -4164 -16100
rect -4298 -16134 -4282 -16117
rect -4358 -16150 -4282 -16134
rect -4180 -16134 -4164 -16117
rect -4120 -16117 -4082 -16100
rect -2127 -16082 -2089 -16065
rect -2045 -16065 -2029 -16048
rect -1927 -16048 -1851 -16032
rect -1927 -16065 -1911 -16048
rect -2045 -16082 -2007 -16065
rect -4120 -16134 -4104 -16117
rect -2127 -16120 -2007 -16082
rect -1949 -16082 -1911 -16065
rect -1867 -16065 -1851 -16048
rect -1749 -16048 -1673 -16032
rect -1749 -16065 -1733 -16048
rect -1867 -16082 -1829 -16065
rect -1949 -16120 -1829 -16082
rect -1771 -16082 -1733 -16065
rect -1689 -16065 -1673 -16048
rect -1571 -16048 -1495 -16032
rect -1571 -16065 -1555 -16048
rect -1689 -16082 -1651 -16065
rect -1771 -16120 -1651 -16082
rect -1593 -16082 -1555 -16065
rect -1511 -16065 -1495 -16048
rect -1393 -16048 -1317 -16032
rect -1393 -16065 -1377 -16048
rect -1511 -16082 -1473 -16065
rect -1593 -16120 -1473 -16082
rect -1415 -16082 -1377 -16065
rect -1333 -16065 -1317 -16048
rect -1215 -16048 -1139 -16032
rect -1215 -16065 -1199 -16048
rect -1333 -16082 -1295 -16065
rect -1415 -16120 -1295 -16082
rect -1237 -16082 -1199 -16065
rect -1155 -16065 -1139 -16048
rect -1037 -16048 -961 -16032
rect -1037 -16065 -1021 -16048
rect -1155 -16082 -1117 -16065
rect -1237 -16120 -1117 -16082
rect -1059 -16082 -1021 -16065
rect -977 -16065 -961 -16048
rect -859 -16048 -783 -16032
rect -859 -16065 -843 -16048
rect -977 -16082 -939 -16065
rect -1059 -16120 -939 -16082
rect -881 -16082 -843 -16065
rect -799 -16065 -783 -16048
rect -681 -16048 -605 -16032
rect -681 -16065 -665 -16048
rect -799 -16082 -761 -16065
rect -881 -16120 -761 -16082
rect -703 -16082 -665 -16065
rect -621 -16065 -605 -16048
rect -503 -16048 -427 -16032
rect -503 -16065 -487 -16048
rect -621 -16082 -583 -16065
rect -703 -16120 -583 -16082
rect -525 -16082 -487 -16065
rect -443 -16065 -427 -16048
rect -325 -16048 -249 -16032
rect -325 -16065 -309 -16048
rect -443 -16082 -405 -16065
rect -525 -16120 -405 -16082
rect -347 -16082 -309 -16065
rect -265 -16065 -249 -16048
rect -147 -16048 -71 -16032
rect -147 -16065 -131 -16048
rect -265 -16082 -227 -16065
rect -347 -16120 -227 -16082
rect -169 -16082 -131 -16065
rect -87 -16065 -71 -16048
rect 31 -16048 107 -16032
rect 31 -16065 47 -16048
rect -87 -16082 -49 -16065
rect -169 -16120 -49 -16082
rect 9 -16082 47 -16065
rect 91 -16065 107 -16048
rect 209 -16048 285 -16032
rect 209 -16065 225 -16048
rect 91 -16082 129 -16065
rect 9 -16120 129 -16082
rect 187 -16082 225 -16065
rect 269 -16065 285 -16048
rect 387 -16048 463 -16032
rect 387 -16065 403 -16048
rect 269 -16082 307 -16065
rect 187 -16120 307 -16082
rect 365 -16082 403 -16065
rect 447 -16065 463 -16048
rect 565 -16048 641 -16032
rect 565 -16065 581 -16048
rect 447 -16082 485 -16065
rect 365 -16120 485 -16082
rect 543 -16082 581 -16065
rect 625 -16065 641 -16048
rect 743 -16048 819 -16032
rect 743 -16065 759 -16048
rect 625 -16082 663 -16065
rect 543 -16120 663 -16082
rect 721 -16082 759 -16065
rect 803 -16065 819 -16048
rect 921 -16048 997 -16032
rect 921 -16065 937 -16048
rect 803 -16082 841 -16065
rect 721 -16120 841 -16082
rect 899 -16082 937 -16065
rect 981 -16065 997 -16048
rect 1099 -16048 1175 -16032
rect 1099 -16065 1115 -16048
rect 981 -16082 1019 -16065
rect 899 -16120 1019 -16082
rect 1077 -16082 1115 -16065
rect 1159 -16065 1175 -16048
rect 1277 -16048 1353 -16032
rect 1277 -16065 1293 -16048
rect 1159 -16082 1197 -16065
rect 1077 -16120 1197 -16082
rect 1255 -16082 1293 -16065
rect 1337 -16065 1353 -16048
rect 1455 -16048 1531 -16032
rect 1455 -16065 1471 -16048
rect 1337 -16082 1375 -16065
rect 1255 -16120 1375 -16082
rect 1433 -16082 1471 -16065
rect 1515 -16065 1531 -16048
rect 1633 -16048 1709 -16032
rect 1633 -16065 1649 -16048
rect 1515 -16082 1553 -16065
rect 1433 -16120 1553 -16082
rect 1611 -16082 1649 -16065
rect 1693 -16065 1709 -16048
rect 1811 -16048 1887 -16032
rect 1811 -16065 1827 -16048
rect 1693 -16082 1731 -16065
rect 1611 -16120 1731 -16082
rect 1789 -16082 1827 -16065
rect 1871 -16065 1887 -16048
rect 1989 -16048 2065 -16032
rect 1989 -16065 2005 -16048
rect 1871 -16082 1909 -16065
rect 1789 -16120 1909 -16082
rect 1967 -16082 2005 -16065
rect 2049 -16065 2065 -16048
rect 2167 -16048 2243 -16032
rect 2167 -16065 2183 -16048
rect 2049 -16082 2087 -16065
rect 1967 -16120 2087 -16082
rect 2145 -16082 2183 -16065
rect 2227 -16065 2243 -16048
rect 2345 -16048 2421 -16032
rect 2345 -16065 2361 -16048
rect 2227 -16082 2265 -16065
rect 2145 -16120 2265 -16082
rect 2323 -16082 2361 -16065
rect 2405 -16065 2421 -16048
rect 2523 -16048 2599 -16032
rect 2523 -16065 2539 -16048
rect 2405 -16082 2443 -16065
rect 2323 -16120 2443 -16082
rect 2501 -16082 2539 -16065
rect 2583 -16065 2599 -16048
rect 2701 -16048 2777 -16032
rect 2701 -16065 2717 -16048
rect 2583 -16082 2621 -16065
rect 2501 -16120 2621 -16082
rect 2679 -16082 2717 -16065
rect 2761 -16065 2777 -16048
rect 2879 -16048 2955 -16032
rect 2879 -16065 2895 -16048
rect 2761 -16082 2799 -16065
rect 2679 -16120 2799 -16082
rect 2857 -16082 2895 -16065
rect 2939 -16065 2955 -16048
rect 3057 -16048 3133 -16032
rect 3057 -16065 3073 -16048
rect 2939 -16082 2977 -16065
rect 2857 -16120 2977 -16082
rect 3035 -16082 3073 -16065
rect 3117 -16065 3133 -16048
rect 3235 -16048 3311 -16032
rect 3235 -16065 3251 -16048
rect 3117 -16082 3155 -16065
rect 3035 -16120 3155 -16082
rect 3213 -16082 3251 -16065
rect 3295 -16065 3311 -16048
rect 3413 -16048 3489 -16032
rect 3413 -16065 3429 -16048
rect 3295 -16082 3333 -16065
rect 3213 -16120 3333 -16082
rect 3391 -16082 3429 -16065
rect 3473 -16065 3489 -16048
rect 3591 -16048 3667 -16032
rect 3591 -16065 3607 -16048
rect 3473 -16082 3511 -16065
rect 3391 -16120 3511 -16082
rect 3569 -16082 3607 -16065
rect 3651 -16065 3667 -16048
rect 3769 -16048 3845 -16032
rect 3769 -16065 3785 -16048
rect 3651 -16082 3689 -16065
rect 3569 -16120 3689 -16082
rect 3747 -16082 3785 -16065
rect 3829 -16065 3845 -16048
rect 3947 -16048 4023 -16032
rect 3947 -16065 3963 -16048
rect 3829 -16082 3867 -16065
rect 3747 -16120 3867 -16082
rect 3925 -16082 3963 -16065
rect 4007 -16065 4023 -16048
rect 5645 -16048 5721 -16032
rect 5645 -16065 5661 -16048
rect 4007 -16082 4045 -16065
rect 3925 -16120 4045 -16082
rect 5623 -16082 5661 -16065
rect 5705 -16065 5721 -16048
rect 5823 -16048 5899 -16032
rect 5823 -16065 5839 -16048
rect 5705 -16082 5743 -16065
rect 5623 -16120 5743 -16082
rect 5801 -16082 5839 -16065
rect 5883 -16065 5899 -16048
rect 6001 -16048 6077 -16032
rect 6001 -16065 6017 -16048
rect 5883 -16082 5921 -16065
rect 5801 -16120 5921 -16082
rect 5979 -16082 6017 -16065
rect 6061 -16065 6077 -16048
rect 6179 -16048 6255 -16032
rect 6179 -16065 6195 -16048
rect 6061 -16082 6099 -16065
rect 5979 -16120 6099 -16082
rect 6157 -16082 6195 -16065
rect 6239 -16065 6255 -16048
rect 6357 -16048 6433 -16032
rect 6357 -16065 6373 -16048
rect 6239 -16082 6277 -16065
rect 6157 -16120 6277 -16082
rect 6335 -16082 6373 -16065
rect 6417 -16065 6433 -16048
rect 6535 -16048 6611 -16032
rect 6535 -16065 6551 -16048
rect 6417 -16082 6455 -16065
rect 6335 -16120 6455 -16082
rect 6513 -16082 6551 -16065
rect 6595 -16065 6611 -16048
rect 6713 -16048 6789 -16032
rect 6713 -16065 6729 -16048
rect 6595 -16082 6633 -16065
rect 6513 -16120 6633 -16082
rect 6691 -16082 6729 -16065
rect 6773 -16065 6789 -16048
rect 6891 -16048 6967 -16032
rect 6891 -16065 6907 -16048
rect 6773 -16082 6811 -16065
rect 6691 -16120 6811 -16082
rect 6869 -16082 6907 -16065
rect 6951 -16065 6967 -16048
rect 7069 -16048 7145 -16032
rect 7069 -16065 7085 -16048
rect 6951 -16082 6989 -16065
rect 6869 -16120 6989 -16082
rect 7047 -16082 7085 -16065
rect 7129 -16065 7145 -16048
rect 7247 -16048 7323 -16032
rect 7247 -16065 7263 -16048
rect 7129 -16082 7167 -16065
rect 7047 -16120 7167 -16082
rect 7225 -16082 7263 -16065
rect 7307 -16065 7323 -16048
rect 7425 -16048 7501 -16032
rect 7425 -16065 7441 -16048
rect 7307 -16082 7345 -16065
rect 7225 -16120 7345 -16082
rect 7403 -16082 7441 -16065
rect 7485 -16065 7501 -16048
rect 7603 -16048 7679 -16032
rect 7603 -16065 7619 -16048
rect 7485 -16082 7523 -16065
rect 7403 -16120 7523 -16082
rect 7581 -16082 7619 -16065
rect 7663 -16065 7679 -16048
rect 7781 -16048 7857 -16032
rect 7781 -16065 7797 -16048
rect 7663 -16082 7701 -16065
rect 7581 -16120 7701 -16082
rect 7759 -16082 7797 -16065
rect 7841 -16065 7857 -16048
rect 7959 -16048 8035 -16032
rect 7959 -16065 7975 -16048
rect 7841 -16082 7879 -16065
rect 7759 -16120 7879 -16082
rect 7937 -16082 7975 -16065
rect 8019 -16065 8035 -16048
rect 8137 -16048 8213 -16032
rect 8137 -16065 8153 -16048
rect 8019 -16082 8057 -16065
rect 7937 -16120 8057 -16082
rect 8115 -16082 8153 -16065
rect 8197 -16065 8213 -16048
rect 8315 -16048 8391 -16032
rect 8315 -16065 8331 -16048
rect 8197 -16082 8235 -16065
rect 8115 -16120 8235 -16082
rect 8293 -16082 8331 -16065
rect 8375 -16065 8391 -16048
rect 8493 -16048 8569 -16032
rect 8493 -16065 8509 -16048
rect 8375 -16082 8413 -16065
rect 8293 -16120 8413 -16082
rect 8471 -16082 8509 -16065
rect 8553 -16065 8569 -16048
rect 8671 -16048 8747 -16032
rect 8671 -16065 8687 -16048
rect 8553 -16082 8591 -16065
rect 8471 -16120 8591 -16082
rect 8649 -16082 8687 -16065
rect 8731 -16065 8747 -16048
rect 8849 -16048 8925 -16032
rect 8849 -16065 8865 -16048
rect 8731 -16082 8769 -16065
rect 8649 -16120 8769 -16082
rect 8827 -16082 8865 -16065
rect 8909 -16065 8925 -16048
rect 9027 -16048 9103 -16032
rect 9027 -16065 9043 -16048
rect 8909 -16082 8947 -16065
rect 8827 -16120 8947 -16082
rect 9005 -16082 9043 -16065
rect 9087 -16065 9103 -16048
rect 9205 -16048 9281 -16032
rect 9205 -16065 9221 -16048
rect 9087 -16082 9125 -16065
rect 9005 -16120 9125 -16082
rect 9183 -16082 9221 -16065
rect 9265 -16065 9281 -16048
rect 9383 -16048 9459 -16032
rect 9383 -16065 9399 -16048
rect 9265 -16082 9303 -16065
rect 9183 -16120 9303 -16082
rect 9361 -16082 9399 -16065
rect 9443 -16065 9459 -16048
rect 9561 -16048 9637 -16032
rect 9561 -16065 9577 -16048
rect 9443 -16082 9481 -16065
rect 9361 -16120 9481 -16082
rect 9539 -16082 9577 -16065
rect 9621 -16065 9637 -16048
rect 9739 -16048 9815 -16032
rect 9739 -16065 9755 -16048
rect 9621 -16082 9659 -16065
rect 9539 -16120 9659 -16082
rect 9717 -16082 9755 -16065
rect 9799 -16065 9815 -16048
rect 9917 -16048 9993 -16032
rect 9917 -16065 9933 -16048
rect 9799 -16082 9837 -16065
rect 9717 -16120 9837 -16082
rect 9895 -16082 9933 -16065
rect 9977 -16065 9993 -16048
rect 10095 -16048 10171 -16032
rect 10095 -16065 10111 -16048
rect 9977 -16082 10015 -16065
rect 9895 -16120 10015 -16082
rect 10073 -16082 10111 -16065
rect 10155 -16065 10171 -16048
rect 10273 -16048 10349 -16032
rect 10273 -16065 10289 -16048
rect 10155 -16082 10193 -16065
rect 10073 -16120 10193 -16082
rect 10251 -16082 10289 -16065
rect 10333 -16065 10349 -16048
rect 10451 -16048 10527 -16032
rect 10451 -16065 10467 -16048
rect 10333 -16082 10371 -16065
rect 10251 -16120 10371 -16082
rect 10429 -16082 10467 -16065
rect 10511 -16065 10527 -16048
rect 10629 -16048 10705 -16032
rect 10629 -16065 10645 -16048
rect 10511 -16082 10549 -16065
rect 10429 -16120 10549 -16082
rect 10607 -16082 10645 -16065
rect 10689 -16065 10705 -16048
rect 10807 -16048 10883 -16032
rect 10807 -16065 10823 -16048
rect 10689 -16082 10727 -16065
rect 10607 -16120 10727 -16082
rect 10785 -16082 10823 -16065
rect 10867 -16065 10883 -16048
rect 10985 -16048 11061 -16032
rect 10985 -16065 11001 -16048
rect 10867 -16082 10905 -16065
rect 10785 -16120 10905 -16082
rect 10963 -16082 11001 -16065
rect 11045 -16065 11061 -16048
rect 11163 -16048 11239 -16032
rect 11163 -16065 11179 -16048
rect 11045 -16082 11083 -16065
rect 10963 -16120 11083 -16082
rect 11141 -16082 11179 -16065
rect 11223 -16065 11239 -16048
rect 11341 -16048 11417 -16032
rect 11341 -16065 11357 -16048
rect 11223 -16082 11261 -16065
rect 11141 -16120 11261 -16082
rect 11319 -16082 11357 -16065
rect 11401 -16065 11417 -16048
rect 11519 -16048 11595 -16032
rect 11519 -16065 11535 -16048
rect 11401 -16082 11439 -16065
rect 11319 -16120 11439 -16082
rect 11497 -16082 11535 -16065
rect 11579 -16065 11595 -16048
rect 11697 -16048 11773 -16032
rect 11697 -16065 11713 -16048
rect 11579 -16082 11617 -16065
rect 11497 -16120 11617 -16082
rect 11675 -16082 11713 -16065
rect 11757 -16065 11773 -16048
rect 11875 -16048 11951 -16032
rect 11875 -16065 11891 -16048
rect 11757 -16082 11795 -16065
rect 11675 -16120 11795 -16082
rect 11853 -16082 11891 -16065
rect 11935 -16065 11951 -16048
rect 12053 -16048 12129 -16032
rect 12053 -16065 12069 -16048
rect 11935 -16082 11973 -16065
rect 11853 -16120 11973 -16082
rect 12031 -16082 12069 -16065
rect 12113 -16065 12129 -16048
rect 12231 -16048 12307 -16032
rect 12231 -16065 12247 -16048
rect 12113 -16082 12151 -16065
rect 12031 -16120 12151 -16082
rect 12209 -16082 12247 -16065
rect 12291 -16065 12307 -16048
rect 12409 -16048 12485 -16032
rect 12409 -16065 12425 -16048
rect 12291 -16082 12329 -16065
rect 12209 -16120 12329 -16082
rect 12387 -16082 12425 -16065
rect 12469 -16065 12485 -16048
rect 12587 -16048 12663 -16032
rect 12587 -16065 12603 -16048
rect 12469 -16082 12507 -16065
rect 12387 -16120 12507 -16082
rect 12565 -16082 12603 -16065
rect 12647 -16065 12663 -16048
rect 12647 -16082 12685 -16065
rect 12565 -16120 12685 -16082
rect -4180 -16150 -4104 -16134
rect -5960 -16410 -5884 -16394
rect -5960 -16427 -5944 -16410
rect -5982 -16444 -5944 -16427
rect -5900 -16427 -5884 -16410
rect -5782 -16410 -5706 -16394
rect -5782 -16427 -5766 -16410
rect -5900 -16444 -5862 -16427
rect -5982 -16482 -5862 -16444
rect -5804 -16444 -5766 -16427
rect -5722 -16427 -5706 -16410
rect -5604 -16410 -5528 -16394
rect -5604 -16427 -5588 -16410
rect -5722 -16444 -5684 -16427
rect -5804 -16482 -5684 -16444
rect -5626 -16444 -5588 -16427
rect -5544 -16427 -5528 -16410
rect -5426 -16410 -5350 -16394
rect -5426 -16427 -5410 -16410
rect -5544 -16444 -5506 -16427
rect -5626 -16482 -5506 -16444
rect -5448 -16444 -5410 -16427
rect -5366 -16427 -5350 -16410
rect -5248 -16410 -5172 -16394
rect -5248 -16427 -5232 -16410
rect -5366 -16444 -5328 -16427
rect -5448 -16482 -5328 -16444
rect -5270 -16444 -5232 -16427
rect -5188 -16427 -5172 -16410
rect -5070 -16410 -4994 -16394
rect -5070 -16427 -5054 -16410
rect -5188 -16444 -5150 -16427
rect -5270 -16482 -5150 -16444
rect -5092 -16444 -5054 -16427
rect -5010 -16427 -4994 -16410
rect -4892 -16410 -4816 -16394
rect -4892 -16427 -4876 -16410
rect -5010 -16444 -4972 -16427
rect -5092 -16482 -4972 -16444
rect -4914 -16444 -4876 -16427
rect -4832 -16427 -4816 -16410
rect -4714 -16410 -4638 -16394
rect -4714 -16427 -4698 -16410
rect -4832 -16444 -4794 -16427
rect -4914 -16482 -4794 -16444
rect -4736 -16444 -4698 -16427
rect -4654 -16427 -4638 -16410
rect -4536 -16410 -4460 -16394
rect -4536 -16427 -4520 -16410
rect -4654 -16444 -4616 -16427
rect -4736 -16482 -4616 -16444
rect -4558 -16444 -4520 -16427
rect -4476 -16427 -4460 -16410
rect -4358 -16410 -4282 -16394
rect -4358 -16427 -4342 -16410
rect -4476 -16444 -4438 -16427
rect -4558 -16482 -4438 -16444
rect -4380 -16444 -4342 -16427
rect -4298 -16427 -4282 -16410
rect -4180 -16410 -4104 -16394
rect -4180 -16427 -4164 -16410
rect -4298 -16444 -4260 -16427
rect -4380 -16482 -4260 -16444
rect -4202 -16444 -4164 -16427
rect -4120 -16427 -4104 -16410
rect -4120 -16444 -4082 -16427
rect -4202 -16482 -4082 -16444
rect -2127 -16438 -2007 -16400
rect -2127 -16455 -2089 -16438
rect -2105 -16472 -2089 -16455
rect -2045 -16455 -2007 -16438
rect -1949 -16438 -1829 -16400
rect -1949 -16455 -1911 -16438
rect -2045 -16472 -2029 -16455
rect -2105 -16488 -2029 -16472
rect -1927 -16472 -1911 -16455
rect -1867 -16455 -1829 -16438
rect -1771 -16438 -1651 -16400
rect -1771 -16455 -1733 -16438
rect -1867 -16472 -1851 -16455
rect -1927 -16488 -1851 -16472
rect -1749 -16472 -1733 -16455
rect -1689 -16455 -1651 -16438
rect -1593 -16438 -1473 -16400
rect -1593 -16455 -1555 -16438
rect -1689 -16472 -1673 -16455
rect -1749 -16488 -1673 -16472
rect -1571 -16472 -1555 -16455
rect -1511 -16455 -1473 -16438
rect -1415 -16438 -1295 -16400
rect -1415 -16455 -1377 -16438
rect -1511 -16472 -1495 -16455
rect -1571 -16488 -1495 -16472
rect -1393 -16472 -1377 -16455
rect -1333 -16455 -1295 -16438
rect -1237 -16438 -1117 -16400
rect -1237 -16455 -1199 -16438
rect -1333 -16472 -1317 -16455
rect -1393 -16488 -1317 -16472
rect -1215 -16472 -1199 -16455
rect -1155 -16455 -1117 -16438
rect -1059 -16438 -939 -16400
rect -1059 -16455 -1021 -16438
rect -1155 -16472 -1139 -16455
rect -1215 -16488 -1139 -16472
rect -1037 -16472 -1021 -16455
rect -977 -16455 -939 -16438
rect -881 -16438 -761 -16400
rect -881 -16455 -843 -16438
rect -977 -16472 -961 -16455
rect -1037 -16488 -961 -16472
rect -859 -16472 -843 -16455
rect -799 -16455 -761 -16438
rect -703 -16438 -583 -16400
rect -703 -16455 -665 -16438
rect -799 -16472 -783 -16455
rect -859 -16488 -783 -16472
rect -681 -16472 -665 -16455
rect -621 -16455 -583 -16438
rect -525 -16438 -405 -16400
rect -525 -16455 -487 -16438
rect -621 -16472 -605 -16455
rect -681 -16488 -605 -16472
rect -503 -16472 -487 -16455
rect -443 -16455 -405 -16438
rect -347 -16438 -227 -16400
rect -347 -16455 -309 -16438
rect -443 -16472 -427 -16455
rect -503 -16488 -427 -16472
rect -325 -16472 -309 -16455
rect -265 -16455 -227 -16438
rect -169 -16438 -49 -16400
rect -169 -16455 -131 -16438
rect -265 -16472 -249 -16455
rect -325 -16488 -249 -16472
rect -147 -16472 -131 -16455
rect -87 -16455 -49 -16438
rect 9 -16438 129 -16400
rect 9 -16455 47 -16438
rect -87 -16472 -71 -16455
rect -147 -16488 -71 -16472
rect 31 -16472 47 -16455
rect 91 -16455 129 -16438
rect 187 -16438 307 -16400
rect 187 -16455 225 -16438
rect 91 -16472 107 -16455
rect 31 -16488 107 -16472
rect 209 -16472 225 -16455
rect 269 -16455 307 -16438
rect 365 -16438 485 -16400
rect 365 -16455 403 -16438
rect 269 -16472 285 -16455
rect 209 -16488 285 -16472
rect 387 -16472 403 -16455
rect 447 -16455 485 -16438
rect 543 -16438 663 -16400
rect 543 -16455 581 -16438
rect 447 -16472 463 -16455
rect 387 -16488 463 -16472
rect 565 -16472 581 -16455
rect 625 -16455 663 -16438
rect 721 -16438 841 -16400
rect 721 -16455 759 -16438
rect 625 -16472 641 -16455
rect 565 -16488 641 -16472
rect 743 -16472 759 -16455
rect 803 -16455 841 -16438
rect 899 -16438 1019 -16400
rect 899 -16455 937 -16438
rect 803 -16472 819 -16455
rect 743 -16488 819 -16472
rect 921 -16472 937 -16455
rect 981 -16455 1019 -16438
rect 1077 -16438 1197 -16400
rect 1077 -16455 1115 -16438
rect 981 -16472 997 -16455
rect 921 -16488 997 -16472
rect 1099 -16472 1115 -16455
rect 1159 -16455 1197 -16438
rect 1255 -16438 1375 -16400
rect 1255 -16455 1293 -16438
rect 1159 -16472 1175 -16455
rect 1099 -16488 1175 -16472
rect 1277 -16472 1293 -16455
rect 1337 -16455 1375 -16438
rect 1433 -16438 1553 -16400
rect 1433 -16455 1471 -16438
rect 1337 -16472 1353 -16455
rect 1277 -16488 1353 -16472
rect 1455 -16472 1471 -16455
rect 1515 -16455 1553 -16438
rect 1611 -16438 1731 -16400
rect 1611 -16455 1649 -16438
rect 1515 -16472 1531 -16455
rect 1455 -16488 1531 -16472
rect 1633 -16472 1649 -16455
rect 1693 -16455 1731 -16438
rect 1789 -16438 1909 -16400
rect 1789 -16455 1827 -16438
rect 1693 -16472 1709 -16455
rect 1633 -16488 1709 -16472
rect 1811 -16472 1827 -16455
rect 1871 -16455 1909 -16438
rect 1967 -16438 2087 -16400
rect 1967 -16455 2005 -16438
rect 1871 -16472 1887 -16455
rect 1811 -16488 1887 -16472
rect 1989 -16472 2005 -16455
rect 2049 -16455 2087 -16438
rect 2145 -16438 2265 -16400
rect 2145 -16455 2183 -16438
rect 2049 -16472 2065 -16455
rect 1989 -16488 2065 -16472
rect 2167 -16472 2183 -16455
rect 2227 -16455 2265 -16438
rect 2323 -16438 2443 -16400
rect 2323 -16455 2361 -16438
rect 2227 -16472 2243 -16455
rect 2167 -16488 2243 -16472
rect 2345 -16472 2361 -16455
rect 2405 -16455 2443 -16438
rect 2501 -16438 2621 -16400
rect 2501 -16455 2539 -16438
rect 2405 -16472 2421 -16455
rect 2345 -16488 2421 -16472
rect 2523 -16472 2539 -16455
rect 2583 -16455 2621 -16438
rect 2679 -16438 2799 -16400
rect 2679 -16455 2717 -16438
rect 2583 -16472 2599 -16455
rect 2523 -16488 2599 -16472
rect 2701 -16472 2717 -16455
rect 2761 -16455 2799 -16438
rect 2857 -16438 2977 -16400
rect 2857 -16455 2895 -16438
rect 2761 -16472 2777 -16455
rect 2701 -16488 2777 -16472
rect 2879 -16472 2895 -16455
rect 2939 -16455 2977 -16438
rect 3035 -16438 3155 -16400
rect 3035 -16455 3073 -16438
rect 2939 -16472 2955 -16455
rect 2879 -16488 2955 -16472
rect 3057 -16472 3073 -16455
rect 3117 -16455 3155 -16438
rect 3213 -16438 3333 -16400
rect 3213 -16455 3251 -16438
rect 3117 -16472 3133 -16455
rect 3057 -16488 3133 -16472
rect 3235 -16472 3251 -16455
rect 3295 -16455 3333 -16438
rect 3391 -16438 3511 -16400
rect 3391 -16455 3429 -16438
rect 3295 -16472 3311 -16455
rect 3235 -16488 3311 -16472
rect 3413 -16472 3429 -16455
rect 3473 -16455 3511 -16438
rect 3569 -16438 3689 -16400
rect 3569 -16455 3607 -16438
rect 3473 -16472 3489 -16455
rect 3413 -16488 3489 -16472
rect 3591 -16472 3607 -16455
rect 3651 -16455 3689 -16438
rect 3747 -16438 3867 -16400
rect 3747 -16455 3785 -16438
rect 3651 -16472 3667 -16455
rect 3591 -16488 3667 -16472
rect 3769 -16472 3785 -16455
rect 3829 -16455 3867 -16438
rect 3925 -16438 4045 -16400
rect 3925 -16455 3963 -16438
rect 3829 -16472 3845 -16455
rect 3769 -16488 3845 -16472
rect 3947 -16472 3963 -16455
rect 4007 -16455 4045 -16438
rect 5623 -16438 5743 -16400
rect 5623 -16455 5661 -16438
rect 4007 -16472 4023 -16455
rect 3947 -16488 4023 -16472
rect 5645 -16472 5661 -16455
rect 5705 -16455 5743 -16438
rect 5801 -16438 5921 -16400
rect 5801 -16455 5839 -16438
rect 5705 -16472 5721 -16455
rect 5645 -16488 5721 -16472
rect 5823 -16472 5839 -16455
rect 5883 -16455 5921 -16438
rect 5979 -16438 6099 -16400
rect 5979 -16455 6017 -16438
rect 5883 -16472 5899 -16455
rect 5823 -16488 5899 -16472
rect 6001 -16472 6017 -16455
rect 6061 -16455 6099 -16438
rect 6157 -16438 6277 -16400
rect 6157 -16455 6195 -16438
rect 6061 -16472 6077 -16455
rect 6001 -16488 6077 -16472
rect 6179 -16472 6195 -16455
rect 6239 -16455 6277 -16438
rect 6335 -16438 6455 -16400
rect 6335 -16455 6373 -16438
rect 6239 -16472 6255 -16455
rect 6179 -16488 6255 -16472
rect 6357 -16472 6373 -16455
rect 6417 -16455 6455 -16438
rect 6513 -16438 6633 -16400
rect 6513 -16455 6551 -16438
rect 6417 -16472 6433 -16455
rect 6357 -16488 6433 -16472
rect 6535 -16472 6551 -16455
rect 6595 -16455 6633 -16438
rect 6691 -16438 6811 -16400
rect 6691 -16455 6729 -16438
rect 6595 -16472 6611 -16455
rect 6535 -16488 6611 -16472
rect 6713 -16472 6729 -16455
rect 6773 -16455 6811 -16438
rect 6869 -16438 6989 -16400
rect 6869 -16455 6907 -16438
rect 6773 -16472 6789 -16455
rect 6713 -16488 6789 -16472
rect 6891 -16472 6907 -16455
rect 6951 -16455 6989 -16438
rect 7047 -16438 7167 -16400
rect 7047 -16455 7085 -16438
rect 6951 -16472 6967 -16455
rect 6891 -16488 6967 -16472
rect 7069 -16472 7085 -16455
rect 7129 -16455 7167 -16438
rect 7225 -16438 7345 -16400
rect 7225 -16455 7263 -16438
rect 7129 -16472 7145 -16455
rect 7069 -16488 7145 -16472
rect 7247 -16472 7263 -16455
rect 7307 -16455 7345 -16438
rect 7403 -16438 7523 -16400
rect 7403 -16455 7441 -16438
rect 7307 -16472 7323 -16455
rect 7247 -16488 7323 -16472
rect 7425 -16472 7441 -16455
rect 7485 -16455 7523 -16438
rect 7581 -16438 7701 -16400
rect 7581 -16455 7619 -16438
rect 7485 -16472 7501 -16455
rect 7425 -16488 7501 -16472
rect 7603 -16472 7619 -16455
rect 7663 -16455 7701 -16438
rect 7759 -16438 7879 -16400
rect 7759 -16455 7797 -16438
rect 7663 -16472 7679 -16455
rect 7603 -16488 7679 -16472
rect 7781 -16472 7797 -16455
rect 7841 -16455 7879 -16438
rect 7937 -16438 8057 -16400
rect 7937 -16455 7975 -16438
rect 7841 -16472 7857 -16455
rect 7781 -16488 7857 -16472
rect 7959 -16472 7975 -16455
rect 8019 -16455 8057 -16438
rect 8115 -16438 8235 -16400
rect 8115 -16455 8153 -16438
rect 8019 -16472 8035 -16455
rect 7959 -16488 8035 -16472
rect 8137 -16472 8153 -16455
rect 8197 -16455 8235 -16438
rect 8293 -16438 8413 -16400
rect 8293 -16455 8331 -16438
rect 8197 -16472 8213 -16455
rect 8137 -16488 8213 -16472
rect 8315 -16472 8331 -16455
rect 8375 -16455 8413 -16438
rect 8471 -16438 8591 -16400
rect 8471 -16455 8509 -16438
rect 8375 -16472 8391 -16455
rect 8315 -16488 8391 -16472
rect 8493 -16472 8509 -16455
rect 8553 -16455 8591 -16438
rect 8649 -16438 8769 -16400
rect 8649 -16455 8687 -16438
rect 8553 -16472 8569 -16455
rect 8493 -16488 8569 -16472
rect 8671 -16472 8687 -16455
rect 8731 -16455 8769 -16438
rect 8827 -16438 8947 -16400
rect 8827 -16455 8865 -16438
rect 8731 -16472 8747 -16455
rect 8671 -16488 8747 -16472
rect 8849 -16472 8865 -16455
rect 8909 -16455 8947 -16438
rect 9005 -16438 9125 -16400
rect 9005 -16455 9043 -16438
rect 8909 -16472 8925 -16455
rect 8849 -16488 8925 -16472
rect 9027 -16472 9043 -16455
rect 9087 -16455 9125 -16438
rect 9183 -16438 9303 -16400
rect 9183 -16455 9221 -16438
rect 9087 -16472 9103 -16455
rect 9027 -16488 9103 -16472
rect 9205 -16472 9221 -16455
rect 9265 -16455 9303 -16438
rect 9361 -16438 9481 -16400
rect 9361 -16455 9399 -16438
rect 9265 -16472 9281 -16455
rect 9205 -16488 9281 -16472
rect 9383 -16472 9399 -16455
rect 9443 -16455 9481 -16438
rect 9539 -16438 9659 -16400
rect 9539 -16455 9577 -16438
rect 9443 -16472 9459 -16455
rect 9383 -16488 9459 -16472
rect 9561 -16472 9577 -16455
rect 9621 -16455 9659 -16438
rect 9717 -16438 9837 -16400
rect 9717 -16455 9755 -16438
rect 9621 -16472 9637 -16455
rect 9561 -16488 9637 -16472
rect 9739 -16472 9755 -16455
rect 9799 -16455 9837 -16438
rect 9895 -16438 10015 -16400
rect 9895 -16455 9933 -16438
rect 9799 -16472 9815 -16455
rect 9739 -16488 9815 -16472
rect 9917 -16472 9933 -16455
rect 9977 -16455 10015 -16438
rect 10073 -16438 10193 -16400
rect 10073 -16455 10111 -16438
rect 9977 -16472 9993 -16455
rect 9917 -16488 9993 -16472
rect 10095 -16472 10111 -16455
rect 10155 -16455 10193 -16438
rect 10251 -16438 10371 -16400
rect 10251 -16455 10289 -16438
rect 10155 -16472 10171 -16455
rect 10095 -16488 10171 -16472
rect 10273 -16472 10289 -16455
rect 10333 -16455 10371 -16438
rect 10429 -16438 10549 -16400
rect 10429 -16455 10467 -16438
rect 10333 -16472 10349 -16455
rect 10273 -16488 10349 -16472
rect 10451 -16472 10467 -16455
rect 10511 -16455 10549 -16438
rect 10607 -16438 10727 -16400
rect 10607 -16455 10645 -16438
rect 10511 -16472 10527 -16455
rect 10451 -16488 10527 -16472
rect 10629 -16472 10645 -16455
rect 10689 -16455 10727 -16438
rect 10785 -16438 10905 -16400
rect 10785 -16455 10823 -16438
rect 10689 -16472 10705 -16455
rect 10629 -16488 10705 -16472
rect 10807 -16472 10823 -16455
rect 10867 -16455 10905 -16438
rect 10963 -16438 11083 -16400
rect 10963 -16455 11001 -16438
rect 10867 -16472 10883 -16455
rect 10807 -16488 10883 -16472
rect 10985 -16472 11001 -16455
rect 11045 -16455 11083 -16438
rect 11141 -16438 11261 -16400
rect 11141 -16455 11179 -16438
rect 11045 -16472 11061 -16455
rect 10985 -16488 11061 -16472
rect 11163 -16472 11179 -16455
rect 11223 -16455 11261 -16438
rect 11319 -16438 11439 -16400
rect 11319 -16455 11357 -16438
rect 11223 -16472 11239 -16455
rect 11163 -16488 11239 -16472
rect 11341 -16472 11357 -16455
rect 11401 -16455 11439 -16438
rect 11497 -16438 11617 -16400
rect 11497 -16455 11535 -16438
rect 11401 -16472 11417 -16455
rect 11341 -16488 11417 -16472
rect 11519 -16472 11535 -16455
rect 11579 -16455 11617 -16438
rect 11675 -16438 11795 -16400
rect 11675 -16455 11713 -16438
rect 11579 -16472 11595 -16455
rect 11519 -16488 11595 -16472
rect 11697 -16472 11713 -16455
rect 11757 -16455 11795 -16438
rect 11853 -16438 11973 -16400
rect 11853 -16455 11891 -16438
rect 11757 -16472 11773 -16455
rect 11697 -16488 11773 -16472
rect 11875 -16472 11891 -16455
rect 11935 -16455 11973 -16438
rect 12031 -16438 12151 -16400
rect 12031 -16455 12069 -16438
rect 11935 -16472 11951 -16455
rect 11875 -16488 11951 -16472
rect 12053 -16472 12069 -16455
rect 12113 -16455 12151 -16438
rect 12209 -16438 12329 -16400
rect 12209 -16455 12247 -16438
rect 12113 -16472 12129 -16455
rect 12053 -16488 12129 -16472
rect 12231 -16472 12247 -16455
rect 12291 -16455 12329 -16438
rect 12387 -16438 12507 -16400
rect 12387 -16455 12425 -16438
rect 12291 -16472 12307 -16455
rect 12231 -16488 12307 -16472
rect 12409 -16472 12425 -16455
rect 12469 -16455 12507 -16438
rect 12565 -16438 12685 -16400
rect 12565 -16455 12603 -16438
rect 12469 -16472 12485 -16455
rect 12409 -16488 12485 -16472
rect 12587 -16472 12603 -16455
rect 12647 -16455 12685 -16438
rect 12647 -16472 12663 -16455
rect 12587 -16488 12663 -16472
rect -5982 -16800 -5862 -16762
rect -5982 -16817 -5944 -16800
rect -5960 -16834 -5944 -16817
rect -5900 -16817 -5862 -16800
rect -5804 -16800 -5684 -16762
rect -5804 -16817 -5766 -16800
rect -5900 -16834 -5884 -16817
rect -5960 -16850 -5884 -16834
rect -5782 -16834 -5766 -16817
rect -5722 -16817 -5684 -16800
rect -5626 -16800 -5506 -16762
rect -5626 -16817 -5588 -16800
rect -5722 -16834 -5706 -16817
rect -5782 -16850 -5706 -16834
rect -5604 -16834 -5588 -16817
rect -5544 -16817 -5506 -16800
rect -5448 -16800 -5328 -16762
rect -5448 -16817 -5410 -16800
rect -5544 -16834 -5528 -16817
rect -5604 -16850 -5528 -16834
rect -5426 -16834 -5410 -16817
rect -5366 -16817 -5328 -16800
rect -5270 -16800 -5150 -16762
rect -5270 -16817 -5232 -16800
rect -5366 -16834 -5350 -16817
rect -5426 -16850 -5350 -16834
rect -5248 -16834 -5232 -16817
rect -5188 -16817 -5150 -16800
rect -5092 -16800 -4972 -16762
rect -5092 -16817 -5054 -16800
rect -5188 -16834 -5172 -16817
rect -5248 -16850 -5172 -16834
rect -5070 -16834 -5054 -16817
rect -5010 -16817 -4972 -16800
rect -4914 -16800 -4794 -16762
rect -4914 -16817 -4876 -16800
rect -5010 -16834 -4994 -16817
rect -5070 -16850 -4994 -16834
rect -4892 -16834 -4876 -16817
rect -4832 -16817 -4794 -16800
rect -4736 -16800 -4616 -16762
rect -4736 -16817 -4698 -16800
rect -4832 -16834 -4816 -16817
rect -4892 -16850 -4816 -16834
rect -4714 -16834 -4698 -16817
rect -4654 -16817 -4616 -16800
rect -4558 -16800 -4438 -16762
rect -4558 -16817 -4520 -16800
rect -4654 -16834 -4638 -16817
rect -4714 -16850 -4638 -16834
rect -4536 -16834 -4520 -16817
rect -4476 -16817 -4438 -16800
rect -4380 -16800 -4260 -16762
rect -4380 -16817 -4342 -16800
rect -4476 -16834 -4460 -16817
rect -4536 -16850 -4460 -16834
rect -4358 -16834 -4342 -16817
rect -4298 -16817 -4260 -16800
rect -4202 -16800 -4082 -16762
rect -4202 -16817 -4164 -16800
rect -4298 -16834 -4282 -16817
rect -4358 -16850 -4282 -16834
rect -4180 -16834 -4164 -16817
rect -4120 -16817 -4082 -16800
rect -4120 -16834 -4104 -16817
rect -4180 -16850 -4104 -16834
<< polycont >>
rect -6218 -2073 -6174 -2039
rect -6040 -2073 -5996 -2039
rect -5862 -2073 -5818 -2039
rect -5684 -2073 -5640 -2039
rect -5506 -2073 -5462 -2039
rect -5328 -2073 -5284 -2039
rect -5150 -2073 -5106 -2039
rect -4972 -2073 -4928 -2039
rect -4794 -2073 -4750 -2039
rect -4616 -2073 -4572 -2039
rect -4438 -2073 -4394 -2039
rect -4260 -2073 -4216 -2039
rect -4082 -2073 -4038 -2039
rect -3904 -2073 -3860 -2039
rect -3726 -2073 -3682 -2039
rect -3548 -2073 -3504 -2039
rect -6218 -2481 -6174 -2447
rect -6040 -2481 -5996 -2447
rect -5862 -2481 -5818 -2447
rect -5684 -2481 -5640 -2447
rect -5506 -2481 -5462 -2447
rect -5328 -2481 -5284 -2447
rect -5150 -2481 -5106 -2447
rect -4972 -2481 -4928 -2447
rect -4794 -2481 -4750 -2447
rect -4616 -2481 -4572 -2447
rect -4438 -2481 -4394 -2447
rect -4260 -2481 -4216 -2447
rect -4082 -2481 -4038 -2447
rect -3904 -2481 -3860 -2447
rect -3726 -2481 -3682 -2447
rect -3548 -2481 -3504 -2447
rect -1370 -2825 -1326 -2791
rect -1192 -2825 -1148 -2791
rect -1014 -2825 -970 -2791
rect -836 -2825 -792 -2791
rect -658 -2825 -614 -2791
rect -480 -2825 -436 -2791
rect -302 -2825 -258 -2791
rect -124 -2825 -80 -2791
rect 54 -2825 98 -2791
rect 232 -2825 276 -2791
rect 410 -2825 454 -2791
rect 588 -2825 632 -2791
rect 766 -2825 810 -2791
rect 944 -2825 988 -2791
rect 1122 -2825 1166 -2791
rect 1300 -2825 1344 -2791
rect 1478 -2825 1522 -2791
rect 1656 -2825 1700 -2791
rect 1834 -2825 1878 -2791
rect 2012 -2825 2056 -2791
rect 2190 -2825 2234 -2791
rect 2368 -2825 2412 -2791
rect 2546 -2825 2590 -2791
rect -6218 -2943 -6174 -2909
rect -6040 -2943 -5996 -2909
rect -5862 -2943 -5818 -2909
rect -5684 -2943 -5640 -2909
rect -5506 -2943 -5462 -2909
rect -5328 -2943 -5284 -2909
rect -5150 -2943 -5106 -2909
rect -4972 -2943 -4928 -2909
rect -4794 -2943 -4750 -2909
rect -4616 -2943 -4572 -2909
rect -4438 -2943 -4394 -2909
rect -4260 -2943 -4216 -2909
rect -4082 -2943 -4038 -2909
rect -3904 -2943 -3860 -2909
rect -3726 -2943 -3682 -2909
rect -3548 -2943 -3504 -2909
rect -1370 -3233 -1326 -3199
rect -1192 -3233 -1148 -3199
rect -1014 -3233 -970 -3199
rect -836 -3233 -792 -3199
rect -658 -3233 -614 -3199
rect -480 -3233 -436 -3199
rect -302 -3233 -258 -3199
rect -124 -3233 -80 -3199
rect 54 -3233 98 -3199
rect 232 -3233 276 -3199
rect 410 -3233 454 -3199
rect 588 -3233 632 -3199
rect 766 -3233 810 -3199
rect 944 -3233 988 -3199
rect 1122 -3233 1166 -3199
rect 1300 -3233 1344 -3199
rect 1478 -3233 1522 -3199
rect 1656 -3233 1700 -3199
rect 1834 -3233 1878 -3199
rect 2012 -3233 2056 -3199
rect 2190 -3233 2234 -3199
rect 2368 -3233 2412 -3199
rect 2546 -3233 2590 -3199
rect -6218 -3351 -6174 -3317
rect -6040 -3351 -5996 -3317
rect -5862 -3351 -5818 -3317
rect -5684 -3351 -5640 -3317
rect -5506 -3351 -5462 -3317
rect -5328 -3351 -5284 -3317
rect -5150 -3351 -5106 -3317
rect -4972 -3351 -4928 -3317
rect -4794 -3351 -4750 -3317
rect -4616 -3351 -4572 -3317
rect -4438 -3351 -4394 -3317
rect -4260 -3351 -4216 -3317
rect -4082 -3351 -4038 -3317
rect -3904 -3351 -3860 -3317
rect -3726 -3351 -3682 -3317
rect -3548 -3351 -3504 -3317
rect -1370 -3725 -1326 -3691
rect -6218 -3813 -6174 -3779
rect -6040 -3813 -5996 -3779
rect -5862 -3813 -5818 -3779
rect -5684 -3813 -5640 -3779
rect -5506 -3813 -5462 -3779
rect -5328 -3813 -5284 -3779
rect -5150 -3813 -5106 -3779
rect -4972 -3813 -4928 -3779
rect -4794 -3813 -4750 -3779
rect -4616 -3813 -4572 -3779
rect -4438 -3813 -4394 -3779
rect -4260 -3813 -4216 -3779
rect -4082 -3813 -4038 -3779
rect -3904 -3813 -3860 -3779
rect -3726 -3813 -3682 -3779
rect -1192 -3725 -1148 -3691
rect -1014 -3725 -970 -3691
rect -836 -3725 -792 -3691
rect -658 -3725 -614 -3691
rect -480 -3725 -436 -3691
rect -302 -3725 -258 -3691
rect -124 -3725 -80 -3691
rect 54 -3725 98 -3691
rect 232 -3725 276 -3691
rect 410 -3725 454 -3691
rect 588 -3725 632 -3691
rect 766 -3725 810 -3691
rect 944 -3725 988 -3691
rect 1122 -3725 1166 -3691
rect 1300 -3725 1344 -3691
rect 1478 -3725 1522 -3691
rect 1656 -3725 1700 -3691
rect 1834 -3725 1878 -3691
rect 2012 -3725 2056 -3691
rect 2190 -3725 2234 -3691
rect 2368 -3725 2412 -3691
rect 2546 -3725 2590 -3691
rect -3548 -3813 -3504 -3779
rect -1370 -4133 -1326 -4099
rect -6218 -4221 -6174 -4187
rect -6040 -4221 -5996 -4187
rect -5862 -4221 -5818 -4187
rect -5684 -4221 -5640 -4187
rect -5506 -4221 -5462 -4187
rect -5328 -4221 -5284 -4187
rect -5150 -4221 -5106 -4187
rect -4972 -4221 -4928 -4187
rect -4794 -4221 -4750 -4187
rect -4616 -4221 -4572 -4187
rect -4438 -4221 -4394 -4187
rect -4260 -4221 -4216 -4187
rect -4082 -4221 -4038 -4187
rect -3904 -4221 -3860 -4187
rect -3726 -4221 -3682 -4187
rect -1192 -4133 -1148 -4099
rect -1014 -4133 -970 -4099
rect -836 -4133 -792 -4099
rect -658 -4133 -614 -4099
rect -480 -4133 -436 -4099
rect -302 -4133 -258 -4099
rect -124 -4133 -80 -4099
rect 54 -4133 98 -4099
rect 232 -4133 276 -4099
rect 410 -4133 454 -4099
rect 588 -4133 632 -4099
rect 766 -4133 810 -4099
rect 944 -4133 988 -4099
rect 1122 -4133 1166 -4099
rect 1300 -4133 1344 -4099
rect 1478 -4133 1522 -4099
rect 1656 -4133 1700 -4099
rect 1834 -4133 1878 -4099
rect 2012 -4133 2056 -4099
rect 2190 -4133 2234 -4099
rect 2368 -4133 2412 -4099
rect 2546 -4133 2590 -4099
rect -3548 -4221 -3504 -4187
rect -1370 -4625 -1326 -4591
rect -6218 -4683 -6174 -4649
rect -6040 -4683 -5996 -4649
rect -5862 -4683 -5818 -4649
rect -5684 -4683 -5640 -4649
rect -5506 -4683 -5462 -4649
rect -5328 -4683 -5284 -4649
rect -5150 -4683 -5106 -4649
rect -4972 -4683 -4928 -4649
rect -4794 -4683 -4750 -4649
rect -4616 -4683 -4572 -4649
rect -4438 -4683 -4394 -4649
rect -4260 -4683 -4216 -4649
rect -4082 -4683 -4038 -4649
rect -3904 -4683 -3860 -4649
rect -3726 -4683 -3682 -4649
rect -3548 -4683 -3504 -4649
rect -1192 -4625 -1148 -4591
rect -1014 -4625 -970 -4591
rect -836 -4625 -792 -4591
rect -658 -4625 -614 -4591
rect -480 -4625 -436 -4591
rect -302 -4625 -258 -4591
rect -124 -4625 -80 -4591
rect 54 -4625 98 -4591
rect 232 -4625 276 -4591
rect 410 -4625 454 -4591
rect 588 -4625 632 -4591
rect 766 -4625 810 -4591
rect 944 -4625 988 -4591
rect 1122 -4625 1166 -4591
rect 1300 -4625 1344 -4591
rect 1478 -4625 1522 -4591
rect 1656 -4625 1700 -4591
rect 1834 -4625 1878 -4591
rect 2012 -4625 2056 -4591
rect 2190 -4625 2234 -4591
rect 2368 -4625 2412 -4591
rect 2546 -4625 2590 -4591
rect -6218 -5091 -6174 -5057
rect -6040 -5091 -5996 -5057
rect -5862 -5091 -5818 -5057
rect -5684 -5091 -5640 -5057
rect -5506 -5091 -5462 -5057
rect -5328 -5091 -5284 -5057
rect -5150 -5091 -5106 -5057
rect -4972 -5091 -4928 -5057
rect -4794 -5091 -4750 -5057
rect -4616 -5091 -4572 -5057
rect -4438 -5091 -4394 -5057
rect -4260 -5091 -4216 -5057
rect -4082 -5091 -4038 -5057
rect -3904 -5091 -3860 -5057
rect -3726 -5091 -3682 -5057
rect -1370 -5033 -1326 -4999
rect -1192 -5033 -1148 -4999
rect -1014 -5033 -970 -4999
rect -836 -5033 -792 -4999
rect -658 -5033 -614 -4999
rect -480 -5033 -436 -4999
rect -302 -5033 -258 -4999
rect -124 -5033 -80 -4999
rect 54 -5033 98 -4999
rect 232 -5033 276 -4999
rect 410 -5033 454 -4999
rect 588 -5033 632 -4999
rect 766 -5033 810 -4999
rect 944 -5033 988 -4999
rect 1122 -5033 1166 -4999
rect 1300 -5033 1344 -4999
rect 1478 -5033 1522 -4999
rect 1656 -5033 1700 -4999
rect 1834 -5033 1878 -4999
rect 2012 -5033 2056 -4999
rect 2190 -5033 2234 -4999
rect 2368 -5033 2412 -4999
rect 2546 -5033 2590 -4999
rect -3548 -5091 -3504 -5057
rect -6218 -5553 -6174 -5519
rect -6040 -5553 -5996 -5519
rect -5862 -5553 -5818 -5519
rect -5684 -5553 -5640 -5519
rect -5506 -5553 -5462 -5519
rect -5328 -5553 -5284 -5519
rect -5150 -5553 -5106 -5519
rect -4972 -5553 -4928 -5519
rect -4794 -5553 -4750 -5519
rect -4616 -5553 -4572 -5519
rect -4438 -5553 -4394 -5519
rect -4260 -5553 -4216 -5519
rect -4082 -5553 -4038 -5519
rect -3904 -5553 -3860 -5519
rect -3726 -5553 -3682 -5519
rect -3548 -5553 -3504 -5519
rect -1370 -5525 -1326 -5491
rect -1192 -5525 -1148 -5491
rect -1014 -5525 -970 -5491
rect -836 -5525 -792 -5491
rect -658 -5525 -614 -5491
rect -480 -5525 -436 -5491
rect -302 -5525 -258 -5491
rect -124 -5525 -80 -5491
rect 54 -5525 98 -5491
rect 232 -5525 276 -5491
rect 410 -5525 454 -5491
rect 588 -5525 632 -5491
rect 766 -5525 810 -5491
rect 944 -5525 988 -5491
rect 1122 -5525 1166 -5491
rect 1300 -5525 1344 -5491
rect 1478 -5525 1522 -5491
rect 1656 -5525 1700 -5491
rect 1834 -5525 1878 -5491
rect 2012 -5525 2056 -5491
rect 2190 -5525 2234 -5491
rect 2368 -5525 2412 -5491
rect 2546 -5525 2590 -5491
rect -6218 -5961 -6174 -5927
rect -6040 -5961 -5996 -5927
rect -5862 -5961 -5818 -5927
rect -5684 -5961 -5640 -5927
rect -5506 -5961 -5462 -5927
rect -5328 -5961 -5284 -5927
rect -5150 -5961 -5106 -5927
rect -4972 -5961 -4928 -5927
rect -4794 -5961 -4750 -5927
rect -4616 -5961 -4572 -5927
rect -4438 -5961 -4394 -5927
rect -4260 -5961 -4216 -5927
rect -4082 -5961 -4038 -5927
rect -3904 -5961 -3860 -5927
rect -3726 -5961 -3682 -5927
rect -3548 -5961 -3504 -5927
rect -1370 -5933 -1326 -5899
rect -1192 -5933 -1148 -5899
rect -1014 -5933 -970 -5899
rect -836 -5933 -792 -5899
rect -658 -5933 -614 -5899
rect -480 -5933 -436 -5899
rect -302 -5933 -258 -5899
rect -124 -5933 -80 -5899
rect 54 -5933 98 -5899
rect 232 -5933 276 -5899
rect 410 -5933 454 -5899
rect 588 -5933 632 -5899
rect 766 -5933 810 -5899
rect 944 -5933 988 -5899
rect 1122 -5933 1166 -5899
rect 1300 -5933 1344 -5899
rect 1478 -5933 1522 -5899
rect 1656 -5933 1700 -5899
rect 1834 -5933 1878 -5899
rect 2012 -5933 2056 -5899
rect 2190 -5933 2234 -5899
rect 2368 -5933 2412 -5899
rect 2546 -5933 2590 -5899
rect -5544 -7824 -5500 -7790
rect -5366 -7824 -5322 -7790
rect -5188 -7824 -5144 -7790
rect -5010 -7824 -4966 -7790
rect -4832 -7824 -4788 -7790
rect -4654 -7824 -4610 -7790
rect -4476 -7824 -4432 -7790
rect -4298 -7824 -4254 -7790
rect -4120 -7824 -4076 -7790
rect -2089 -8082 -2045 -8048
rect -1911 -8082 -1867 -8048
rect -1733 -8082 -1689 -8048
rect -1555 -8082 -1511 -8048
rect -1377 -8082 -1333 -8048
rect -1199 -8082 -1155 -8048
rect -1021 -8082 -977 -8048
rect -843 -8082 -799 -8048
rect -665 -8082 -621 -8048
rect -487 -8082 -443 -8048
rect -309 -8082 -265 -8048
rect -131 -8082 -87 -8048
rect 47 -8082 91 -8048
rect 225 -8082 269 -8048
rect 403 -8082 447 -8048
rect 581 -8082 625 -8048
rect 759 -8082 803 -8048
rect 937 -8082 981 -8048
rect 1115 -8082 1159 -8048
rect 1293 -8082 1337 -8048
rect 1471 -8082 1515 -8048
rect 1649 -8082 1693 -8048
rect 1827 -8082 1871 -8048
rect 2005 -8082 2049 -8048
rect 2183 -8082 2227 -8048
rect 2361 -8082 2405 -8048
rect 2539 -8082 2583 -8048
rect 2717 -8082 2761 -8048
rect 2895 -8082 2939 -8048
rect 3073 -8082 3117 -8048
rect 3251 -8082 3295 -8048
rect 3429 -8082 3473 -8048
rect 3607 -8082 3651 -8048
rect 3785 -8082 3829 -8048
rect 3963 -8082 4007 -8048
rect -5544 -8214 -5500 -8180
rect -5366 -8214 -5322 -8180
rect -5188 -8214 -5144 -8180
rect -5010 -8214 -4966 -8180
rect -4832 -8214 -4788 -8180
rect -4654 -8214 -4610 -8180
rect -4476 -8214 -4432 -8180
rect -4298 -8214 -4254 -8180
rect -4120 -8214 -4076 -8180
rect -5544 -8374 -5500 -8340
rect -5366 -8374 -5322 -8340
rect -5188 -8374 -5144 -8340
rect -5010 -8374 -4966 -8340
rect -4832 -8374 -4788 -8340
rect -4654 -8374 -4610 -8340
rect -4476 -8374 -4432 -8340
rect -4298 -8374 -4254 -8340
rect -4120 -8374 -4076 -8340
rect -2089 -8472 -2045 -8438
rect -1911 -8472 -1867 -8438
rect -1733 -8472 -1689 -8438
rect -1555 -8472 -1511 -8438
rect -1377 -8472 -1333 -8438
rect -1199 -8472 -1155 -8438
rect -1021 -8472 -977 -8438
rect -843 -8472 -799 -8438
rect -665 -8472 -621 -8438
rect -487 -8472 -443 -8438
rect -309 -8472 -265 -8438
rect -131 -8472 -87 -8438
rect 47 -8472 91 -8438
rect 225 -8472 269 -8438
rect 403 -8472 447 -8438
rect 581 -8472 625 -8438
rect 759 -8472 803 -8438
rect 937 -8472 981 -8438
rect 1115 -8472 1159 -8438
rect 1293 -8472 1337 -8438
rect 1471 -8472 1515 -8438
rect 1649 -8472 1693 -8438
rect 1827 -8472 1871 -8438
rect 2005 -8472 2049 -8438
rect 2183 -8472 2227 -8438
rect 2361 -8472 2405 -8438
rect 2539 -8472 2583 -8438
rect 2717 -8472 2761 -8438
rect 2895 -8472 2939 -8438
rect 3073 -8472 3117 -8438
rect 3251 -8472 3295 -8438
rect 3429 -8472 3473 -8438
rect 3607 -8472 3651 -8438
rect 3785 -8472 3829 -8438
rect 3963 -8472 4007 -8438
rect -5544 -8764 -5500 -8730
rect -5366 -8764 -5322 -8730
rect -5188 -8764 -5144 -8730
rect -5010 -8764 -4966 -8730
rect -4832 -8764 -4788 -8730
rect -4654 -8764 -4610 -8730
rect -4476 -8764 -4432 -8730
rect -4298 -8764 -4254 -8730
rect -4120 -8764 -4076 -8730
rect 6596 -8844 6640 -8810
rect -5544 -8924 -5500 -8890
rect -5366 -8924 -5322 -8890
rect -5188 -8924 -5144 -8890
rect -5010 -8924 -4966 -8890
rect -4832 -8924 -4788 -8890
rect -4654 -8924 -4610 -8890
rect -4476 -8924 -4432 -8890
rect -4298 -8924 -4254 -8890
rect 6774 -8844 6818 -8810
rect 6952 -8844 6996 -8810
rect 7130 -8844 7174 -8810
rect 7308 -8844 7352 -8810
rect 7486 -8844 7530 -8810
rect 7664 -8844 7708 -8810
rect 7842 -8844 7886 -8810
rect 8020 -8844 8064 -8810
rect 8198 -8844 8242 -8810
rect 8376 -8844 8420 -8810
rect 8554 -8844 8598 -8810
rect 8732 -8844 8776 -8810
rect 8910 -8844 8954 -8810
rect 9088 -8844 9132 -8810
rect 9266 -8844 9310 -8810
rect 10856 -8874 10900 -8840
rect -4120 -8924 -4076 -8890
rect -2089 -9082 -2045 -9048
rect -1911 -9082 -1867 -9048
rect -1733 -9082 -1689 -9048
rect -1555 -9082 -1511 -9048
rect -1377 -9082 -1333 -9048
rect -1199 -9082 -1155 -9048
rect -1021 -9082 -977 -9048
rect -843 -9082 -799 -9048
rect -665 -9082 -621 -9048
rect -487 -9082 -443 -9048
rect -309 -9082 -265 -9048
rect -131 -9082 -87 -9048
rect 47 -9082 91 -9048
rect 225 -9082 269 -9048
rect 403 -9082 447 -9048
rect 581 -9082 625 -9048
rect 759 -9082 803 -9048
rect 937 -9082 981 -9048
rect 1115 -9082 1159 -9048
rect 1293 -9082 1337 -9048
rect 1471 -9082 1515 -9048
rect 1649 -9082 1693 -9048
rect 1827 -9082 1871 -9048
rect 2005 -9082 2049 -9048
rect 2183 -9082 2227 -9048
rect 2361 -9082 2405 -9048
rect 2539 -9082 2583 -9048
rect 2717 -9082 2761 -9048
rect 2895 -9082 2939 -9048
rect 3073 -9082 3117 -9048
rect 3251 -9082 3295 -9048
rect 3429 -9082 3473 -9048
rect 3607 -9082 3651 -9048
rect 3785 -9082 3829 -9048
rect 3963 -9082 4007 -9048
rect -5544 -9314 -5500 -9280
rect -5366 -9314 -5322 -9280
rect -5188 -9314 -5144 -9280
rect -5010 -9314 -4966 -9280
rect -4832 -9314 -4788 -9280
rect -4654 -9314 -4610 -9280
rect -4476 -9314 -4432 -9280
rect -4298 -9314 -4254 -9280
rect -4120 -9314 -4076 -9280
rect 11148 -8874 11192 -8840
rect 11440 -8874 11484 -8840
rect 11732 -8874 11776 -8840
rect 12024 -8874 12068 -8840
rect 12316 -8874 12360 -8840
rect 12608 -8874 12652 -8840
rect 6596 -9234 6640 -9200
rect 6774 -9234 6818 -9200
rect 6952 -9234 6996 -9200
rect 7130 -9234 7174 -9200
rect 7308 -9234 7352 -9200
rect 7486 -9234 7530 -9200
rect 7664 -9234 7708 -9200
rect 7842 -9234 7886 -9200
rect 8020 -9234 8064 -9200
rect 8198 -9234 8242 -9200
rect 8376 -9234 8420 -9200
rect 8554 -9234 8598 -9200
rect 8732 -9234 8776 -9200
rect 8910 -9234 8954 -9200
rect 9088 -9234 9132 -9200
rect 9266 -9234 9310 -9200
rect 10856 -9264 10900 -9230
rect 11148 -9264 11192 -9230
rect 11440 -9264 11484 -9230
rect 11732 -9264 11776 -9230
rect 12024 -9264 12068 -9230
rect 12316 -9264 12360 -9230
rect 12608 -9264 12652 -9230
rect -5544 -9474 -5500 -9440
rect -5366 -9474 -5322 -9440
rect -5188 -9474 -5144 -9440
rect -5010 -9474 -4966 -9440
rect -4832 -9474 -4788 -9440
rect -4654 -9474 -4610 -9440
rect -4476 -9474 -4432 -9440
rect -4298 -9474 -4254 -9440
rect -4120 -9474 -4076 -9440
rect -2089 -9472 -2045 -9438
rect -1911 -9472 -1867 -9438
rect -1733 -9472 -1689 -9438
rect -1555 -9472 -1511 -9438
rect -1377 -9472 -1333 -9438
rect -1199 -9472 -1155 -9438
rect -1021 -9472 -977 -9438
rect -843 -9472 -799 -9438
rect -665 -9472 -621 -9438
rect -487 -9472 -443 -9438
rect -309 -9472 -265 -9438
rect -131 -9472 -87 -9438
rect 47 -9472 91 -9438
rect 225 -9472 269 -9438
rect 403 -9472 447 -9438
rect 581 -9472 625 -9438
rect 759 -9472 803 -9438
rect 937 -9472 981 -9438
rect 1115 -9472 1159 -9438
rect 1293 -9472 1337 -9438
rect 1471 -9472 1515 -9438
rect 1649 -9472 1693 -9438
rect 1827 -9472 1871 -9438
rect 2005 -9472 2049 -9438
rect 2183 -9472 2227 -9438
rect 2361 -9472 2405 -9438
rect 2539 -9472 2583 -9438
rect 2717 -9472 2761 -9438
rect 2895 -9472 2939 -9438
rect 3073 -9472 3117 -9438
rect 3251 -9472 3295 -9438
rect 3429 -9472 3473 -9438
rect 3607 -9472 3651 -9438
rect 3785 -9472 3829 -9438
rect 3963 -9472 4007 -9438
rect 10856 -9644 10900 -9610
rect 11148 -9644 11192 -9610
rect 11440 -9644 11484 -9610
rect 11732 -9644 11776 -9610
rect 12024 -9644 12068 -9610
rect 12316 -9644 12360 -9610
rect 12608 -9644 12652 -9610
rect 6596 -9744 6640 -9710
rect 6774 -9744 6818 -9710
rect 6952 -9744 6996 -9710
rect 7130 -9744 7174 -9710
rect 7308 -9744 7352 -9710
rect 7486 -9744 7530 -9710
rect 7664 -9744 7708 -9710
rect 7842 -9744 7886 -9710
rect 8020 -9744 8064 -9710
rect 8198 -9744 8242 -9710
rect 8376 -9744 8420 -9710
rect 8554 -9744 8598 -9710
rect 8732 -9744 8776 -9710
rect 8910 -9744 8954 -9710
rect 9088 -9744 9132 -9710
rect 9266 -9744 9310 -9710
rect -5544 -9864 -5500 -9830
rect -5366 -9864 -5322 -9830
rect -5188 -9864 -5144 -9830
rect -5010 -9864 -4966 -9830
rect -4832 -9864 -4788 -9830
rect -4654 -9864 -4610 -9830
rect -4476 -9864 -4432 -9830
rect -4298 -9864 -4254 -9830
rect -4120 -9864 -4076 -9830
rect -5544 -10024 -5500 -9990
rect -5366 -10024 -5322 -9990
rect -5188 -10024 -5144 -9990
rect -5010 -10024 -4966 -9990
rect -4832 -10024 -4788 -9990
rect -4654 -10024 -4610 -9990
rect -4476 -10024 -4432 -9990
rect -4298 -10024 -4254 -9990
rect -4120 -10024 -4076 -9990
rect -2089 -10082 -2045 -10048
rect -1911 -10082 -1867 -10048
rect -1733 -10082 -1689 -10048
rect -1555 -10082 -1511 -10048
rect -1377 -10082 -1333 -10048
rect -1199 -10082 -1155 -10048
rect -1021 -10082 -977 -10048
rect -843 -10082 -799 -10048
rect -665 -10082 -621 -10048
rect -487 -10082 -443 -10048
rect -309 -10082 -265 -10048
rect -131 -10082 -87 -10048
rect 47 -10082 91 -10048
rect 225 -10082 269 -10048
rect 403 -10082 447 -10048
rect 581 -10082 625 -10048
rect 759 -10082 803 -10048
rect 937 -10082 981 -10048
rect 1115 -10082 1159 -10048
rect 1293 -10082 1337 -10048
rect 1471 -10082 1515 -10048
rect 1649 -10082 1693 -10048
rect 1827 -10082 1871 -10048
rect 2005 -10082 2049 -10048
rect 2183 -10082 2227 -10048
rect 2361 -10082 2405 -10048
rect 2539 -10082 2583 -10048
rect 2717 -10082 2761 -10048
rect 2895 -10082 2939 -10048
rect 3073 -10082 3117 -10048
rect 3251 -10082 3295 -10048
rect 3429 -10082 3473 -10048
rect 3607 -10082 3651 -10048
rect 3785 -10082 3829 -10048
rect 3963 -10082 4007 -10048
rect 10856 -10034 10900 -10000
rect 11148 -10034 11192 -10000
rect 11440 -10034 11484 -10000
rect 11732 -10034 11776 -10000
rect 12024 -10034 12068 -10000
rect 12316 -10034 12360 -10000
rect 12608 -10034 12652 -10000
rect -5544 -10414 -5500 -10380
rect -5366 -10414 -5322 -10380
rect -5188 -10414 -5144 -10380
rect -5010 -10414 -4966 -10380
rect -4832 -10414 -4788 -10380
rect -4654 -10414 -4610 -10380
rect -4476 -10414 -4432 -10380
rect -4298 -10414 -4254 -10380
rect -4120 -10414 -4076 -10380
rect 6596 -10134 6640 -10100
rect 6774 -10134 6818 -10100
rect 6952 -10134 6996 -10100
rect 7130 -10134 7174 -10100
rect 7308 -10134 7352 -10100
rect 7486 -10134 7530 -10100
rect 7664 -10134 7708 -10100
rect 7842 -10134 7886 -10100
rect 8020 -10134 8064 -10100
rect 8198 -10134 8242 -10100
rect 8376 -10134 8420 -10100
rect 8554 -10134 8598 -10100
rect 8732 -10134 8776 -10100
rect 8910 -10134 8954 -10100
rect 9088 -10134 9132 -10100
rect 9266 -10134 9310 -10100
rect -2089 -10472 -2045 -10438
rect -1911 -10472 -1867 -10438
rect -1733 -10472 -1689 -10438
rect -1555 -10472 -1511 -10438
rect -1377 -10472 -1333 -10438
rect -1199 -10472 -1155 -10438
rect -1021 -10472 -977 -10438
rect -843 -10472 -799 -10438
rect -665 -10472 -621 -10438
rect -487 -10472 -443 -10438
rect -309 -10472 -265 -10438
rect -131 -10472 -87 -10438
rect 47 -10472 91 -10438
rect 225 -10472 269 -10438
rect 403 -10472 447 -10438
rect 581 -10472 625 -10438
rect 759 -10472 803 -10438
rect 937 -10472 981 -10438
rect 1115 -10472 1159 -10438
rect 1293 -10472 1337 -10438
rect 1471 -10472 1515 -10438
rect 1649 -10472 1693 -10438
rect 1827 -10472 1871 -10438
rect 2005 -10472 2049 -10438
rect 2183 -10472 2227 -10438
rect 2361 -10472 2405 -10438
rect 2539 -10472 2583 -10438
rect 2717 -10472 2761 -10438
rect 2895 -10472 2939 -10438
rect 3073 -10472 3117 -10438
rect 3251 -10472 3295 -10438
rect 3429 -10472 3473 -10438
rect 3607 -10472 3651 -10438
rect 3785 -10472 3829 -10438
rect 3963 -10472 4007 -10438
rect 10856 -10414 10900 -10380
rect 11148 -10414 11192 -10380
rect 11440 -10414 11484 -10380
rect 11732 -10414 11776 -10380
rect 12024 -10414 12068 -10380
rect 12316 -10414 12360 -10380
rect 12608 -10414 12652 -10380
rect -5544 -10574 -5500 -10540
rect -5366 -10574 -5322 -10540
rect -5188 -10574 -5144 -10540
rect -5010 -10574 -4966 -10540
rect -4832 -10574 -4788 -10540
rect -4654 -10574 -4610 -10540
rect -4476 -10574 -4432 -10540
rect -4298 -10574 -4254 -10540
rect -4120 -10574 -4076 -10540
rect 6596 -10644 6640 -10610
rect 6774 -10644 6818 -10610
rect 6952 -10644 6996 -10610
rect 7130 -10644 7174 -10610
rect 7308 -10644 7352 -10610
rect 7486 -10644 7530 -10610
rect 7664 -10644 7708 -10610
rect 7842 -10644 7886 -10610
rect 8020 -10644 8064 -10610
rect 8198 -10644 8242 -10610
rect 8376 -10644 8420 -10610
rect 8554 -10644 8598 -10610
rect 8732 -10644 8776 -10610
rect 8910 -10644 8954 -10610
rect 9088 -10644 9132 -10610
rect 9266 -10644 9310 -10610
rect -5544 -10964 -5500 -10930
rect -5366 -10964 -5322 -10930
rect -5188 -10964 -5144 -10930
rect -5010 -10964 -4966 -10930
rect -4832 -10964 -4788 -10930
rect -4654 -10964 -4610 -10930
rect -4476 -10964 -4432 -10930
rect -4298 -10964 -4254 -10930
rect -4120 -10964 -4076 -10930
rect 10856 -10804 10900 -10770
rect 11148 -10804 11192 -10770
rect 11440 -10804 11484 -10770
rect 11732 -10804 11776 -10770
rect 12024 -10804 12068 -10770
rect 12316 -10804 12360 -10770
rect 12608 -10804 12652 -10770
rect -5544 -11124 -5500 -11090
rect -5366 -11124 -5322 -11090
rect -5188 -11124 -5144 -11090
rect -5010 -11124 -4966 -11090
rect -4832 -11124 -4788 -11090
rect -4654 -11124 -4610 -11090
rect -4476 -11124 -4432 -11090
rect -4298 -11124 -4254 -11090
rect -4120 -11124 -4076 -11090
rect -2089 -11082 -2045 -11048
rect -1911 -11082 -1867 -11048
rect -1733 -11082 -1689 -11048
rect -1555 -11082 -1511 -11048
rect -1377 -11082 -1333 -11048
rect -1199 -11082 -1155 -11048
rect -1021 -11082 -977 -11048
rect -843 -11082 -799 -11048
rect -665 -11082 -621 -11048
rect -487 -11082 -443 -11048
rect -309 -11082 -265 -11048
rect -131 -11082 -87 -11048
rect 47 -11082 91 -11048
rect 225 -11082 269 -11048
rect 403 -11082 447 -11048
rect 581 -11082 625 -11048
rect 759 -11082 803 -11048
rect 937 -11082 981 -11048
rect 1115 -11082 1159 -11048
rect 1293 -11082 1337 -11048
rect 1471 -11082 1515 -11048
rect 1649 -11082 1693 -11048
rect 1827 -11082 1871 -11048
rect 2005 -11082 2049 -11048
rect 2183 -11082 2227 -11048
rect 2361 -11082 2405 -11048
rect 2539 -11082 2583 -11048
rect 2717 -11082 2761 -11048
rect 2895 -11082 2939 -11048
rect 3073 -11082 3117 -11048
rect 3251 -11082 3295 -11048
rect 3429 -11082 3473 -11048
rect 3607 -11082 3651 -11048
rect 3785 -11082 3829 -11048
rect 3963 -11082 4007 -11048
rect 6596 -11034 6640 -11000
rect 6774 -11034 6818 -11000
rect 6952 -11034 6996 -11000
rect 7130 -11034 7174 -11000
rect 7308 -11034 7352 -11000
rect 7486 -11034 7530 -11000
rect 7664 -11034 7708 -11000
rect 7842 -11034 7886 -11000
rect 8020 -11034 8064 -11000
rect 8198 -11034 8242 -11000
rect 8376 -11034 8420 -11000
rect 8554 -11034 8598 -11000
rect 8732 -11034 8776 -11000
rect 8910 -11034 8954 -11000
rect 9088 -11034 9132 -11000
rect 9266 -11034 9310 -11000
rect 10856 -11184 10900 -11150
rect 11148 -11184 11192 -11150
rect 11440 -11184 11484 -11150
rect 11732 -11184 11776 -11150
rect 12024 -11184 12068 -11150
rect 12316 -11184 12360 -11150
rect 12608 -11184 12652 -11150
rect -5544 -11514 -5500 -11480
rect -5366 -11514 -5322 -11480
rect -5188 -11514 -5144 -11480
rect -5010 -11514 -4966 -11480
rect -4832 -11514 -4788 -11480
rect -4654 -11514 -4610 -11480
rect -4476 -11514 -4432 -11480
rect -4298 -11514 -4254 -11480
rect -4120 -11514 -4076 -11480
rect -2089 -11472 -2045 -11438
rect -1911 -11472 -1867 -11438
rect -1733 -11472 -1689 -11438
rect -1555 -11472 -1511 -11438
rect -1377 -11472 -1333 -11438
rect -1199 -11472 -1155 -11438
rect -1021 -11472 -977 -11438
rect -843 -11472 -799 -11438
rect -665 -11472 -621 -11438
rect -487 -11472 -443 -11438
rect -309 -11472 -265 -11438
rect -131 -11472 -87 -11438
rect 47 -11472 91 -11438
rect 225 -11472 269 -11438
rect 403 -11472 447 -11438
rect 581 -11472 625 -11438
rect 759 -11472 803 -11438
rect 937 -11472 981 -11438
rect 1115 -11472 1159 -11438
rect 1293 -11472 1337 -11438
rect 1471 -11472 1515 -11438
rect 1649 -11472 1693 -11438
rect 1827 -11472 1871 -11438
rect 2005 -11472 2049 -11438
rect 2183 -11472 2227 -11438
rect 2361 -11472 2405 -11438
rect 2539 -11472 2583 -11438
rect 2717 -11472 2761 -11438
rect 2895 -11472 2939 -11438
rect 3073 -11472 3117 -11438
rect 3251 -11472 3295 -11438
rect 3429 -11472 3473 -11438
rect 3607 -11472 3651 -11438
rect 3785 -11472 3829 -11438
rect 3963 -11472 4007 -11438
rect 6596 -11544 6640 -11510
rect 6774 -11544 6818 -11510
rect 6952 -11544 6996 -11510
rect 7130 -11544 7174 -11510
rect 7308 -11544 7352 -11510
rect 7486 -11544 7530 -11510
rect 7664 -11544 7708 -11510
rect 7842 -11544 7886 -11510
rect 8020 -11544 8064 -11510
rect 8198 -11544 8242 -11510
rect 8376 -11544 8420 -11510
rect 8554 -11544 8598 -11510
rect 8732 -11544 8776 -11510
rect 8910 -11544 8954 -11510
rect 9088 -11544 9132 -11510
rect 9266 -11544 9310 -11510
rect 10856 -11574 10900 -11540
rect -5544 -11674 -5500 -11640
rect -5366 -11674 -5322 -11640
rect -5188 -11674 -5144 -11640
rect -5010 -11674 -4966 -11640
rect -4832 -11674 -4788 -11640
rect -4654 -11674 -4610 -11640
rect -4476 -11674 -4432 -11640
rect -4298 -11674 -4254 -11640
rect -4120 -11674 -4076 -11640
rect 11148 -11574 11192 -11540
rect 11440 -11574 11484 -11540
rect 11732 -11574 11776 -11540
rect 12024 -11574 12068 -11540
rect 12316 -11574 12360 -11540
rect 12608 -11574 12652 -11540
rect 6596 -11934 6640 -11900
rect 6774 -11934 6818 -11900
rect 6952 -11934 6996 -11900
rect 7130 -11934 7174 -11900
rect 7308 -11934 7352 -11900
rect 7486 -11934 7530 -11900
rect 7664 -11934 7708 -11900
rect 7842 -11934 7886 -11900
rect 8020 -11934 8064 -11900
rect 8198 -11934 8242 -11900
rect 8376 -11934 8420 -11900
rect 8554 -11934 8598 -11900
rect 8732 -11934 8776 -11900
rect 8910 -11934 8954 -11900
rect 9088 -11934 9132 -11900
rect 9266 -11934 9310 -11900
rect -5544 -12064 -5500 -12030
rect -5366 -12064 -5322 -12030
rect -5188 -12064 -5144 -12030
rect -5010 -12064 -4966 -12030
rect -4832 -12064 -4788 -12030
rect -4654 -12064 -4610 -12030
rect -4476 -12064 -4432 -12030
rect -4298 -12064 -4254 -12030
rect -4120 -12064 -4076 -12030
rect -2089 -12082 -2045 -12048
rect -1911 -12082 -1867 -12048
rect -1733 -12082 -1689 -12048
rect -1555 -12082 -1511 -12048
rect -1377 -12082 -1333 -12048
rect -1199 -12082 -1155 -12048
rect -1021 -12082 -977 -12048
rect -843 -12082 -799 -12048
rect -665 -12082 -621 -12048
rect -487 -12082 -443 -12048
rect -309 -12082 -265 -12048
rect -131 -12082 -87 -12048
rect 47 -12082 91 -12048
rect 225 -12082 269 -12048
rect 403 -12082 447 -12048
rect 581 -12082 625 -12048
rect 759 -12082 803 -12048
rect 937 -12082 981 -12048
rect 1115 -12082 1159 -12048
rect 1293 -12082 1337 -12048
rect 1471 -12082 1515 -12048
rect 1649 -12082 1693 -12048
rect 1827 -12082 1871 -12048
rect 2005 -12082 2049 -12048
rect 2183 -12082 2227 -12048
rect 2361 -12082 2405 -12048
rect 2539 -12082 2583 -12048
rect 2717 -12082 2761 -12048
rect 2895 -12082 2939 -12048
rect 3073 -12082 3117 -12048
rect 3251 -12082 3295 -12048
rect 3429 -12082 3473 -12048
rect 3607 -12082 3651 -12048
rect 3785 -12082 3829 -12048
rect 3963 -12082 4007 -12048
rect -2089 -12472 -2045 -12438
rect -1911 -12472 -1867 -12438
rect -1733 -12472 -1689 -12438
rect -1555 -12472 -1511 -12438
rect -1377 -12472 -1333 -12438
rect -1199 -12472 -1155 -12438
rect -1021 -12472 -977 -12438
rect -843 -12472 -799 -12438
rect -665 -12472 -621 -12438
rect -487 -12472 -443 -12438
rect -309 -12472 -265 -12438
rect -131 -12472 -87 -12438
rect 47 -12472 91 -12438
rect 225 -12472 269 -12438
rect 403 -12472 447 -12438
rect 581 -12472 625 -12438
rect 759 -12472 803 -12438
rect 937 -12472 981 -12438
rect 1115 -12472 1159 -12438
rect 1293 -12472 1337 -12438
rect 1471 -12472 1515 -12438
rect 1649 -12472 1693 -12438
rect 1827 -12472 1871 -12438
rect 2005 -12472 2049 -12438
rect 2183 -12472 2227 -12438
rect 2361 -12472 2405 -12438
rect 2539 -12472 2583 -12438
rect 2717 -12472 2761 -12438
rect 2895 -12472 2939 -12438
rect 3073 -12472 3117 -12438
rect 3251 -12472 3295 -12438
rect 3429 -12472 3473 -12438
rect 3607 -12472 3651 -12438
rect 3785 -12472 3829 -12438
rect 3963 -12472 4007 -12438
rect -5867 -12662 -5833 -12628
rect -5617 -12662 -5583 -12628
rect -5367 -12662 -5333 -12628
rect -5117 -12662 -5083 -12628
rect -4867 -12662 -4833 -12628
rect -4617 -12662 -4583 -12628
rect -4367 -12662 -4333 -12628
rect -4117 -12662 -4083 -12628
rect -5867 -13012 -5833 -12978
rect -5617 -13012 -5583 -12978
rect -5367 -13012 -5333 -12978
rect -5117 -13012 -5083 -12978
rect -4867 -13012 -4833 -12978
rect -4617 -13012 -4583 -12978
rect -4367 -13012 -4333 -12978
rect -4117 -13012 -4083 -12978
rect -2089 -13082 -2045 -13048
rect -1911 -13082 -1867 -13048
rect -1733 -13082 -1689 -13048
rect -1555 -13082 -1511 -13048
rect -1377 -13082 -1333 -13048
rect -1199 -13082 -1155 -13048
rect -1021 -13082 -977 -13048
rect -843 -13082 -799 -13048
rect -665 -13082 -621 -13048
rect -487 -13082 -443 -13048
rect -309 -13082 -265 -13048
rect -131 -13082 -87 -13048
rect 47 -13082 91 -13048
rect 225 -13082 269 -13048
rect 403 -13082 447 -13048
rect 581 -13082 625 -13048
rect 759 -13082 803 -13048
rect 937 -13082 981 -13048
rect 1115 -13082 1159 -13048
rect 1293 -13082 1337 -13048
rect 1471 -13082 1515 -13048
rect 1649 -13082 1693 -13048
rect 1827 -13082 1871 -13048
rect 2005 -13082 2049 -13048
rect 2183 -13082 2227 -13048
rect 2361 -13082 2405 -13048
rect 2539 -13082 2583 -13048
rect 2717 -13082 2761 -13048
rect 2895 -13082 2939 -13048
rect 3073 -13082 3117 -13048
rect 3251 -13082 3295 -13048
rect 3429 -13082 3473 -13048
rect 3607 -13082 3651 -13048
rect 3785 -13082 3829 -13048
rect 3963 -13082 4007 -13048
rect -5867 -13342 -5833 -13308
rect -5617 -13342 -5583 -13308
rect -5367 -13342 -5333 -13308
rect -5117 -13342 -5083 -13308
rect -4867 -13342 -4833 -13308
rect -4617 -13342 -4583 -13308
rect -4367 -13342 -4333 -13308
rect -4117 -13342 -4083 -13308
rect -2089 -13472 -2045 -13438
rect -1911 -13472 -1867 -13438
rect -1733 -13472 -1689 -13438
rect -1555 -13472 -1511 -13438
rect -1377 -13472 -1333 -13438
rect -1199 -13472 -1155 -13438
rect -1021 -13472 -977 -13438
rect -843 -13472 -799 -13438
rect -665 -13472 -621 -13438
rect -487 -13472 -443 -13438
rect -309 -13472 -265 -13438
rect -131 -13472 -87 -13438
rect 47 -13472 91 -13438
rect 225 -13472 269 -13438
rect 403 -13472 447 -13438
rect 581 -13472 625 -13438
rect 759 -13472 803 -13438
rect 937 -13472 981 -13438
rect 1115 -13472 1159 -13438
rect 1293 -13472 1337 -13438
rect 1471 -13472 1515 -13438
rect 1649 -13472 1693 -13438
rect 1827 -13472 1871 -13438
rect 2005 -13472 2049 -13438
rect 2183 -13472 2227 -13438
rect 2361 -13472 2405 -13438
rect 2539 -13472 2583 -13438
rect 2717 -13472 2761 -13438
rect 2895 -13472 2939 -13438
rect 3073 -13472 3117 -13438
rect 3251 -13472 3295 -13438
rect 3429 -13472 3473 -13438
rect 3607 -13472 3651 -13438
rect 3785 -13472 3829 -13438
rect 3963 -13472 4007 -13438
rect -5867 -13692 -5833 -13658
rect -5617 -13692 -5583 -13658
rect -5367 -13692 -5333 -13658
rect -5117 -13692 -5083 -13658
rect -4867 -13692 -4833 -13658
rect -4617 -13692 -4583 -13658
rect -4367 -13692 -4333 -13658
rect -4117 -13692 -4083 -13658
rect -2089 -14082 -2045 -14048
rect -1911 -14082 -1867 -14048
rect -1733 -14082 -1689 -14048
rect -1555 -14082 -1511 -14048
rect -1377 -14082 -1333 -14048
rect -1199 -14082 -1155 -14048
rect -1021 -14082 -977 -14048
rect -843 -14082 -799 -14048
rect -665 -14082 -621 -14048
rect -487 -14082 -443 -14048
rect -309 -14082 -265 -14048
rect -131 -14082 -87 -14048
rect 47 -14082 91 -14048
rect 225 -14082 269 -14048
rect 403 -14082 447 -14048
rect 581 -14082 625 -14048
rect 759 -14082 803 -14048
rect 937 -14082 981 -14048
rect 1115 -14082 1159 -14048
rect 1293 -14082 1337 -14048
rect 1471 -14082 1515 -14048
rect 1649 -14082 1693 -14048
rect 1827 -14082 1871 -14048
rect 2005 -14082 2049 -14048
rect 2183 -14082 2227 -14048
rect 2361 -14082 2405 -14048
rect 2539 -14082 2583 -14048
rect 2717 -14082 2761 -14048
rect 2895 -14082 2939 -14048
rect 3073 -14082 3117 -14048
rect 3251 -14082 3295 -14048
rect 3429 -14082 3473 -14048
rect 3607 -14082 3651 -14048
rect 3785 -14082 3829 -14048
rect 3963 -14082 4007 -14048
rect 5661 -14082 5705 -14048
rect 5839 -14082 5883 -14048
rect 6017 -14082 6061 -14048
rect 6195 -14082 6239 -14048
rect 6373 -14082 6417 -14048
rect 6551 -14082 6595 -14048
rect 6729 -14082 6773 -14048
rect 6907 -14082 6951 -14048
rect 7085 -14082 7129 -14048
rect 7263 -14082 7307 -14048
rect 7441 -14082 7485 -14048
rect 7619 -14082 7663 -14048
rect 7797 -14082 7841 -14048
rect 7975 -14082 8019 -14048
rect 8153 -14082 8197 -14048
rect 8331 -14082 8375 -14048
rect 8509 -14082 8553 -14048
rect 8687 -14082 8731 -14048
rect 8865 -14082 8909 -14048
rect 9043 -14082 9087 -14048
rect 9221 -14082 9265 -14048
rect 9399 -14082 9443 -14048
rect 9577 -14082 9621 -14048
rect 9755 -14082 9799 -14048
rect 9933 -14082 9977 -14048
rect 10111 -14082 10155 -14048
rect 10289 -14082 10333 -14048
rect 10467 -14082 10511 -14048
rect 10645 -14082 10689 -14048
rect 10823 -14082 10867 -14048
rect 11001 -14082 11045 -14048
rect 11179 -14082 11223 -14048
rect 11357 -14082 11401 -14048
rect 11535 -14082 11579 -14048
rect 11713 -14082 11757 -14048
rect 11891 -14082 11935 -14048
rect 12069 -14082 12113 -14048
rect 12247 -14082 12291 -14048
rect 12425 -14082 12469 -14048
rect 12603 -14082 12647 -14048
rect -5944 -14344 -5900 -14310
rect -5766 -14344 -5722 -14310
rect -5588 -14344 -5544 -14310
rect -5410 -14344 -5366 -14310
rect -5232 -14344 -5188 -14310
rect -5054 -14344 -5010 -14310
rect -4876 -14344 -4832 -14310
rect -4698 -14344 -4654 -14310
rect -4520 -14344 -4476 -14310
rect -4342 -14344 -4298 -14310
rect -4164 -14344 -4120 -14310
rect -2089 -14472 -2045 -14438
rect -1911 -14472 -1867 -14438
rect -1733 -14472 -1689 -14438
rect -1555 -14472 -1511 -14438
rect -1377 -14472 -1333 -14438
rect -1199 -14472 -1155 -14438
rect -1021 -14472 -977 -14438
rect -843 -14472 -799 -14438
rect -665 -14472 -621 -14438
rect -487 -14472 -443 -14438
rect -309 -14472 -265 -14438
rect -131 -14472 -87 -14438
rect 47 -14472 91 -14438
rect 225 -14472 269 -14438
rect 403 -14472 447 -14438
rect 581 -14472 625 -14438
rect 759 -14472 803 -14438
rect 937 -14472 981 -14438
rect 1115 -14472 1159 -14438
rect 1293 -14472 1337 -14438
rect 1471 -14472 1515 -14438
rect 1649 -14472 1693 -14438
rect 1827 -14472 1871 -14438
rect 2005 -14472 2049 -14438
rect 2183 -14472 2227 -14438
rect 2361 -14472 2405 -14438
rect 2539 -14472 2583 -14438
rect 2717 -14472 2761 -14438
rect 2895 -14472 2939 -14438
rect 3073 -14472 3117 -14438
rect 3251 -14472 3295 -14438
rect 3429 -14472 3473 -14438
rect 3607 -14472 3651 -14438
rect 3785 -14472 3829 -14438
rect 3963 -14472 4007 -14438
rect 5661 -14472 5705 -14438
rect 5839 -14472 5883 -14438
rect 6017 -14472 6061 -14438
rect 6195 -14472 6239 -14438
rect 6373 -14472 6417 -14438
rect 6551 -14472 6595 -14438
rect 6729 -14472 6773 -14438
rect 6907 -14472 6951 -14438
rect 7085 -14472 7129 -14438
rect 7263 -14472 7307 -14438
rect 7441 -14472 7485 -14438
rect 7619 -14472 7663 -14438
rect 7797 -14472 7841 -14438
rect 7975 -14472 8019 -14438
rect 8153 -14472 8197 -14438
rect 8331 -14472 8375 -14438
rect 8509 -14472 8553 -14438
rect 8687 -14472 8731 -14438
rect 8865 -14472 8909 -14438
rect 9043 -14472 9087 -14438
rect 9221 -14472 9265 -14438
rect 9399 -14472 9443 -14438
rect 9577 -14472 9621 -14438
rect 9755 -14472 9799 -14438
rect 9933 -14472 9977 -14438
rect 10111 -14472 10155 -14438
rect 10289 -14472 10333 -14438
rect 10467 -14472 10511 -14438
rect 10645 -14472 10689 -14438
rect 10823 -14472 10867 -14438
rect 11001 -14472 11045 -14438
rect 11179 -14472 11223 -14438
rect 11357 -14472 11401 -14438
rect 11535 -14472 11579 -14438
rect 11713 -14472 11757 -14438
rect 11891 -14472 11935 -14438
rect 12069 -14472 12113 -14438
rect 12247 -14472 12291 -14438
rect 12425 -14472 12469 -14438
rect 12603 -14472 12647 -14438
rect -5944 -14734 -5900 -14700
rect -5766 -14734 -5722 -14700
rect -5588 -14734 -5544 -14700
rect -5410 -14734 -5366 -14700
rect -5232 -14734 -5188 -14700
rect -5054 -14734 -5010 -14700
rect -4876 -14734 -4832 -14700
rect -4698 -14734 -4654 -14700
rect -4520 -14734 -4476 -14700
rect -4342 -14734 -4298 -14700
rect -4164 -14734 -4120 -14700
rect -5944 -15044 -5900 -15010
rect -5766 -15044 -5722 -15010
rect -5588 -15044 -5544 -15010
rect -5410 -15044 -5366 -15010
rect -5232 -15044 -5188 -15010
rect -5054 -15044 -5010 -15010
rect -4876 -15044 -4832 -15010
rect -4698 -15044 -4654 -15010
rect -4520 -15044 -4476 -15010
rect -4342 -15044 -4298 -15010
rect -4164 -15044 -4120 -15010
rect -2089 -15082 -2045 -15048
rect -1911 -15082 -1867 -15048
rect -1733 -15082 -1689 -15048
rect -1555 -15082 -1511 -15048
rect -1377 -15082 -1333 -15048
rect -1199 -15082 -1155 -15048
rect -1021 -15082 -977 -15048
rect -843 -15082 -799 -15048
rect -665 -15082 -621 -15048
rect -487 -15082 -443 -15048
rect -309 -15082 -265 -15048
rect -131 -15082 -87 -15048
rect 47 -15082 91 -15048
rect 225 -15082 269 -15048
rect 403 -15082 447 -15048
rect 581 -15082 625 -15048
rect 759 -15082 803 -15048
rect 937 -15082 981 -15048
rect 1115 -15082 1159 -15048
rect 1293 -15082 1337 -15048
rect 1471 -15082 1515 -15048
rect 1649 -15082 1693 -15048
rect 1827 -15082 1871 -15048
rect 2005 -15082 2049 -15048
rect 2183 -15082 2227 -15048
rect 2361 -15082 2405 -15048
rect 2539 -15082 2583 -15048
rect 2717 -15082 2761 -15048
rect 2895 -15082 2939 -15048
rect 3073 -15082 3117 -15048
rect 3251 -15082 3295 -15048
rect 3429 -15082 3473 -15048
rect 3607 -15082 3651 -15048
rect 3785 -15082 3829 -15048
rect 3963 -15082 4007 -15048
rect 5661 -15082 5705 -15048
rect 5839 -15082 5883 -15048
rect 6017 -15082 6061 -15048
rect 6195 -15082 6239 -15048
rect 6373 -15082 6417 -15048
rect 6551 -15082 6595 -15048
rect 6729 -15082 6773 -15048
rect 6907 -15082 6951 -15048
rect 7085 -15082 7129 -15048
rect 7263 -15082 7307 -15048
rect 7441 -15082 7485 -15048
rect 7619 -15082 7663 -15048
rect 7797 -15082 7841 -15048
rect 7975 -15082 8019 -15048
rect 8153 -15082 8197 -15048
rect 8331 -15082 8375 -15048
rect 8509 -15082 8553 -15048
rect 8687 -15082 8731 -15048
rect 8865 -15082 8909 -15048
rect 9043 -15082 9087 -15048
rect 9221 -15082 9265 -15048
rect 9399 -15082 9443 -15048
rect 9577 -15082 9621 -15048
rect 9755 -15082 9799 -15048
rect 9933 -15082 9977 -15048
rect 10111 -15082 10155 -15048
rect 10289 -15082 10333 -15048
rect 10467 -15082 10511 -15048
rect 10645 -15082 10689 -15048
rect 10823 -15082 10867 -15048
rect 11001 -15082 11045 -15048
rect 11179 -15082 11223 -15048
rect 11357 -15082 11401 -15048
rect 11535 -15082 11579 -15048
rect 11713 -15082 11757 -15048
rect 11891 -15082 11935 -15048
rect 12069 -15082 12113 -15048
rect 12247 -15082 12291 -15048
rect 12425 -15082 12469 -15048
rect 12603 -15082 12647 -15048
rect -5944 -15434 -5900 -15400
rect -5766 -15434 -5722 -15400
rect -5588 -15434 -5544 -15400
rect -5410 -15434 -5366 -15400
rect -5232 -15434 -5188 -15400
rect -5054 -15434 -5010 -15400
rect -4876 -15434 -4832 -15400
rect -4698 -15434 -4654 -15400
rect -4520 -15434 -4476 -15400
rect -4342 -15434 -4298 -15400
rect -4164 -15434 -4120 -15400
rect -2089 -15472 -2045 -15438
rect -1911 -15472 -1867 -15438
rect -1733 -15472 -1689 -15438
rect -1555 -15472 -1511 -15438
rect -1377 -15472 -1333 -15438
rect -1199 -15472 -1155 -15438
rect -1021 -15472 -977 -15438
rect -843 -15472 -799 -15438
rect -665 -15472 -621 -15438
rect -487 -15472 -443 -15438
rect -309 -15472 -265 -15438
rect -131 -15472 -87 -15438
rect 47 -15472 91 -15438
rect 225 -15472 269 -15438
rect 403 -15472 447 -15438
rect 581 -15472 625 -15438
rect 759 -15472 803 -15438
rect 937 -15472 981 -15438
rect 1115 -15472 1159 -15438
rect 1293 -15472 1337 -15438
rect 1471 -15472 1515 -15438
rect 1649 -15472 1693 -15438
rect 1827 -15472 1871 -15438
rect 2005 -15472 2049 -15438
rect 2183 -15472 2227 -15438
rect 2361 -15472 2405 -15438
rect 2539 -15472 2583 -15438
rect 2717 -15472 2761 -15438
rect 2895 -15472 2939 -15438
rect 3073 -15472 3117 -15438
rect 3251 -15472 3295 -15438
rect 3429 -15472 3473 -15438
rect 3607 -15472 3651 -15438
rect 3785 -15472 3829 -15438
rect 3963 -15472 4007 -15438
rect 5661 -15472 5705 -15438
rect 5839 -15472 5883 -15438
rect 6017 -15472 6061 -15438
rect 6195 -15472 6239 -15438
rect 6373 -15472 6417 -15438
rect 6551 -15472 6595 -15438
rect 6729 -15472 6773 -15438
rect 6907 -15472 6951 -15438
rect 7085 -15472 7129 -15438
rect 7263 -15472 7307 -15438
rect 7441 -15472 7485 -15438
rect 7619 -15472 7663 -15438
rect 7797 -15472 7841 -15438
rect 7975 -15472 8019 -15438
rect 8153 -15472 8197 -15438
rect 8331 -15472 8375 -15438
rect 8509 -15472 8553 -15438
rect 8687 -15472 8731 -15438
rect 8865 -15472 8909 -15438
rect 9043 -15472 9087 -15438
rect 9221 -15472 9265 -15438
rect 9399 -15472 9443 -15438
rect 9577 -15472 9621 -15438
rect 9755 -15472 9799 -15438
rect 9933 -15472 9977 -15438
rect 10111 -15472 10155 -15438
rect 10289 -15472 10333 -15438
rect 10467 -15472 10511 -15438
rect 10645 -15472 10689 -15438
rect 10823 -15472 10867 -15438
rect 11001 -15472 11045 -15438
rect 11179 -15472 11223 -15438
rect 11357 -15472 11401 -15438
rect 11535 -15472 11579 -15438
rect 11713 -15472 11757 -15438
rect 11891 -15472 11935 -15438
rect 12069 -15472 12113 -15438
rect 12247 -15472 12291 -15438
rect 12425 -15472 12469 -15438
rect 12603 -15472 12647 -15438
rect -5944 -15744 -5900 -15710
rect -5766 -15744 -5722 -15710
rect -5588 -15744 -5544 -15710
rect -5410 -15744 -5366 -15710
rect -5232 -15744 -5188 -15710
rect -5054 -15744 -5010 -15710
rect -4876 -15744 -4832 -15710
rect -4698 -15744 -4654 -15710
rect -4520 -15744 -4476 -15710
rect -4342 -15744 -4298 -15710
rect -4164 -15744 -4120 -15710
rect -5944 -16134 -5900 -16100
rect -5766 -16134 -5722 -16100
rect -5588 -16134 -5544 -16100
rect -5410 -16134 -5366 -16100
rect -5232 -16134 -5188 -16100
rect -5054 -16134 -5010 -16100
rect -4876 -16134 -4832 -16100
rect -4698 -16134 -4654 -16100
rect -4520 -16134 -4476 -16100
rect -4342 -16134 -4298 -16100
rect -4164 -16134 -4120 -16100
rect -2089 -16082 -2045 -16048
rect -1911 -16082 -1867 -16048
rect -1733 -16082 -1689 -16048
rect -1555 -16082 -1511 -16048
rect -1377 -16082 -1333 -16048
rect -1199 -16082 -1155 -16048
rect -1021 -16082 -977 -16048
rect -843 -16082 -799 -16048
rect -665 -16082 -621 -16048
rect -487 -16082 -443 -16048
rect -309 -16082 -265 -16048
rect -131 -16082 -87 -16048
rect 47 -16082 91 -16048
rect 225 -16082 269 -16048
rect 403 -16082 447 -16048
rect 581 -16082 625 -16048
rect 759 -16082 803 -16048
rect 937 -16082 981 -16048
rect 1115 -16082 1159 -16048
rect 1293 -16082 1337 -16048
rect 1471 -16082 1515 -16048
rect 1649 -16082 1693 -16048
rect 1827 -16082 1871 -16048
rect 2005 -16082 2049 -16048
rect 2183 -16082 2227 -16048
rect 2361 -16082 2405 -16048
rect 2539 -16082 2583 -16048
rect 2717 -16082 2761 -16048
rect 2895 -16082 2939 -16048
rect 3073 -16082 3117 -16048
rect 3251 -16082 3295 -16048
rect 3429 -16082 3473 -16048
rect 3607 -16082 3651 -16048
rect 3785 -16082 3829 -16048
rect 3963 -16082 4007 -16048
rect 5661 -16082 5705 -16048
rect 5839 -16082 5883 -16048
rect 6017 -16082 6061 -16048
rect 6195 -16082 6239 -16048
rect 6373 -16082 6417 -16048
rect 6551 -16082 6595 -16048
rect 6729 -16082 6773 -16048
rect 6907 -16082 6951 -16048
rect 7085 -16082 7129 -16048
rect 7263 -16082 7307 -16048
rect 7441 -16082 7485 -16048
rect 7619 -16082 7663 -16048
rect 7797 -16082 7841 -16048
rect 7975 -16082 8019 -16048
rect 8153 -16082 8197 -16048
rect 8331 -16082 8375 -16048
rect 8509 -16082 8553 -16048
rect 8687 -16082 8731 -16048
rect 8865 -16082 8909 -16048
rect 9043 -16082 9087 -16048
rect 9221 -16082 9265 -16048
rect 9399 -16082 9443 -16048
rect 9577 -16082 9621 -16048
rect 9755 -16082 9799 -16048
rect 9933 -16082 9977 -16048
rect 10111 -16082 10155 -16048
rect 10289 -16082 10333 -16048
rect 10467 -16082 10511 -16048
rect 10645 -16082 10689 -16048
rect 10823 -16082 10867 -16048
rect 11001 -16082 11045 -16048
rect 11179 -16082 11223 -16048
rect 11357 -16082 11401 -16048
rect 11535 -16082 11579 -16048
rect 11713 -16082 11757 -16048
rect 11891 -16082 11935 -16048
rect 12069 -16082 12113 -16048
rect 12247 -16082 12291 -16048
rect 12425 -16082 12469 -16048
rect 12603 -16082 12647 -16048
rect -5944 -16444 -5900 -16410
rect -5766 -16444 -5722 -16410
rect -5588 -16444 -5544 -16410
rect -5410 -16444 -5366 -16410
rect -5232 -16444 -5188 -16410
rect -5054 -16444 -5010 -16410
rect -4876 -16444 -4832 -16410
rect -4698 -16444 -4654 -16410
rect -4520 -16444 -4476 -16410
rect -4342 -16444 -4298 -16410
rect -4164 -16444 -4120 -16410
rect -2089 -16472 -2045 -16438
rect -1911 -16472 -1867 -16438
rect -1733 -16472 -1689 -16438
rect -1555 -16472 -1511 -16438
rect -1377 -16472 -1333 -16438
rect -1199 -16472 -1155 -16438
rect -1021 -16472 -977 -16438
rect -843 -16472 -799 -16438
rect -665 -16472 -621 -16438
rect -487 -16472 -443 -16438
rect -309 -16472 -265 -16438
rect -131 -16472 -87 -16438
rect 47 -16472 91 -16438
rect 225 -16472 269 -16438
rect 403 -16472 447 -16438
rect 581 -16472 625 -16438
rect 759 -16472 803 -16438
rect 937 -16472 981 -16438
rect 1115 -16472 1159 -16438
rect 1293 -16472 1337 -16438
rect 1471 -16472 1515 -16438
rect 1649 -16472 1693 -16438
rect 1827 -16472 1871 -16438
rect 2005 -16472 2049 -16438
rect 2183 -16472 2227 -16438
rect 2361 -16472 2405 -16438
rect 2539 -16472 2583 -16438
rect 2717 -16472 2761 -16438
rect 2895 -16472 2939 -16438
rect 3073 -16472 3117 -16438
rect 3251 -16472 3295 -16438
rect 3429 -16472 3473 -16438
rect 3607 -16472 3651 -16438
rect 3785 -16472 3829 -16438
rect 3963 -16472 4007 -16438
rect 5661 -16472 5705 -16438
rect 5839 -16472 5883 -16438
rect 6017 -16472 6061 -16438
rect 6195 -16472 6239 -16438
rect 6373 -16472 6417 -16438
rect 6551 -16472 6595 -16438
rect 6729 -16472 6773 -16438
rect 6907 -16472 6951 -16438
rect 7085 -16472 7129 -16438
rect 7263 -16472 7307 -16438
rect 7441 -16472 7485 -16438
rect 7619 -16472 7663 -16438
rect 7797 -16472 7841 -16438
rect 7975 -16472 8019 -16438
rect 8153 -16472 8197 -16438
rect 8331 -16472 8375 -16438
rect 8509 -16472 8553 -16438
rect 8687 -16472 8731 -16438
rect 8865 -16472 8909 -16438
rect 9043 -16472 9087 -16438
rect 9221 -16472 9265 -16438
rect 9399 -16472 9443 -16438
rect 9577 -16472 9621 -16438
rect 9755 -16472 9799 -16438
rect 9933 -16472 9977 -16438
rect 10111 -16472 10155 -16438
rect 10289 -16472 10333 -16438
rect 10467 -16472 10511 -16438
rect 10645 -16472 10689 -16438
rect 10823 -16472 10867 -16438
rect 11001 -16472 11045 -16438
rect 11179 -16472 11223 -16438
rect 11357 -16472 11401 -16438
rect 11535 -16472 11579 -16438
rect 11713 -16472 11757 -16438
rect 11891 -16472 11935 -16438
rect 12069 -16472 12113 -16438
rect 12247 -16472 12291 -16438
rect 12425 -16472 12469 -16438
rect 12603 -16472 12647 -16438
rect -5944 -16834 -5900 -16800
rect -5766 -16834 -5722 -16800
rect -5588 -16834 -5544 -16800
rect -5410 -16834 -5366 -16800
rect -5232 -16834 -5188 -16800
rect -5054 -16834 -5010 -16800
rect -4876 -16834 -4832 -16800
rect -4698 -16834 -4654 -16800
rect -4520 -16834 -4476 -16800
rect -4342 -16834 -4298 -16800
rect -4164 -16834 -4120 -16800
<< locali >>
rect -7606 -1353 -7379 -1260
rect 3329 -1353 3703 -1260
rect -7605 -1507 -7512 -1353
rect 3610 -1520 3703 -1353
rect -6234 -2073 -6218 -2039
rect -6174 -2073 -6158 -2039
rect -6056 -2073 -6040 -2039
rect -5996 -2073 -5980 -2039
rect -5878 -2073 -5862 -2039
rect -5818 -2073 -5802 -2039
rect -5700 -2073 -5684 -2039
rect -5640 -2073 -5624 -2039
rect -5522 -2073 -5506 -2039
rect -5462 -2073 -5446 -2039
rect -5344 -2073 -5328 -2039
rect -5284 -2073 -5268 -2039
rect -5166 -2073 -5150 -2039
rect -5106 -2073 -5090 -2039
rect -4988 -2073 -4972 -2039
rect -4928 -2073 -4912 -2039
rect -4810 -2073 -4794 -2039
rect -4750 -2073 -4734 -2039
rect -4632 -2073 -4616 -2039
rect -4572 -2073 -4556 -2039
rect -4454 -2073 -4438 -2039
rect -4394 -2073 -4378 -2039
rect -4276 -2073 -4260 -2039
rect -4216 -2073 -4200 -2039
rect -4098 -2073 -4082 -2039
rect -4038 -2073 -4022 -2039
rect -3920 -2073 -3904 -2039
rect -3860 -2073 -3844 -2039
rect -3742 -2073 -3726 -2039
rect -3682 -2073 -3666 -2039
rect -3564 -2073 -3548 -2039
rect -3504 -2073 -3488 -2039
rect -6302 -2132 -6268 -2116
rect -6302 -2404 -6268 -2388
rect -6124 -2132 -6090 -2116
rect -6124 -2404 -6090 -2388
rect -5946 -2132 -5912 -2116
rect -5946 -2404 -5912 -2388
rect -5768 -2132 -5734 -2116
rect -5768 -2404 -5734 -2388
rect -5590 -2132 -5556 -2116
rect -5590 -2404 -5556 -2388
rect -5412 -2132 -5378 -2116
rect -5412 -2404 -5378 -2388
rect -5234 -2132 -5200 -2116
rect -5234 -2404 -5200 -2388
rect -5056 -2132 -5022 -2116
rect -5056 -2404 -5022 -2388
rect -4878 -2132 -4844 -2116
rect -4878 -2404 -4844 -2388
rect -4700 -2132 -4666 -2116
rect -4700 -2404 -4666 -2388
rect -4522 -2132 -4488 -2116
rect -4522 -2404 -4488 -2388
rect -4344 -2132 -4310 -2116
rect -4344 -2404 -4310 -2388
rect -4166 -2132 -4132 -2116
rect -4166 -2404 -4132 -2388
rect -3988 -2132 -3954 -2116
rect -3988 -2404 -3954 -2388
rect -3810 -2132 -3776 -2116
rect -3810 -2404 -3776 -2388
rect -3632 -2132 -3598 -2116
rect -3632 -2404 -3598 -2388
rect -3454 -2132 -3420 -2116
rect -3454 -2404 -3420 -2388
rect -6234 -2481 -6218 -2447
rect -6174 -2481 -6158 -2447
rect -6056 -2481 -6040 -2447
rect -5996 -2481 -5980 -2447
rect -5878 -2481 -5862 -2447
rect -5818 -2481 -5802 -2447
rect -5700 -2481 -5684 -2447
rect -5640 -2481 -5624 -2447
rect -5522 -2481 -5506 -2447
rect -5462 -2481 -5446 -2447
rect -5344 -2481 -5328 -2447
rect -5284 -2481 -5268 -2447
rect -5166 -2481 -5150 -2447
rect -5106 -2481 -5090 -2447
rect -4988 -2481 -4972 -2447
rect -4928 -2481 -4912 -2447
rect -4810 -2481 -4794 -2447
rect -4750 -2481 -4734 -2447
rect -4632 -2481 -4616 -2447
rect -4572 -2481 -4556 -2447
rect -4454 -2481 -4438 -2447
rect -4394 -2481 -4378 -2447
rect -4276 -2481 -4260 -2447
rect -4216 -2481 -4200 -2447
rect -4098 -2481 -4082 -2447
rect -4038 -2481 -4022 -2447
rect -3920 -2481 -3904 -2447
rect -3860 -2481 -3844 -2447
rect -3742 -2481 -3726 -2447
rect -3682 -2481 -3666 -2447
rect -3564 -2481 -3548 -2447
rect -3504 -2481 -3488 -2447
rect -1386 -2825 -1370 -2791
rect -1326 -2825 -1310 -2791
rect -1208 -2825 -1192 -2791
rect -1148 -2825 -1132 -2791
rect -1030 -2825 -1014 -2791
rect -970 -2825 -954 -2791
rect -852 -2825 -836 -2791
rect -792 -2825 -776 -2791
rect -674 -2825 -658 -2791
rect -614 -2825 -598 -2791
rect -496 -2825 -480 -2791
rect -436 -2825 -420 -2791
rect -318 -2825 -302 -2791
rect -258 -2825 -242 -2791
rect -140 -2825 -124 -2791
rect -80 -2825 -64 -2791
rect 38 -2825 54 -2791
rect 98 -2825 114 -2791
rect 216 -2825 232 -2791
rect 276 -2825 292 -2791
rect 394 -2825 410 -2791
rect 454 -2825 470 -2791
rect 572 -2825 588 -2791
rect 632 -2825 648 -2791
rect 750 -2825 766 -2791
rect 810 -2825 826 -2791
rect 928 -2825 944 -2791
rect 988 -2825 1004 -2791
rect 1106 -2825 1122 -2791
rect 1166 -2825 1182 -2791
rect 1284 -2825 1300 -2791
rect 1344 -2825 1360 -2791
rect 1462 -2825 1478 -2791
rect 1522 -2825 1538 -2791
rect 1640 -2825 1656 -2791
rect 1700 -2825 1716 -2791
rect 1818 -2825 1834 -2791
rect 1878 -2825 1894 -2791
rect 1996 -2825 2012 -2791
rect 2056 -2825 2072 -2791
rect 2174 -2825 2190 -2791
rect 2234 -2825 2250 -2791
rect 2352 -2825 2368 -2791
rect 2412 -2825 2428 -2791
rect 2530 -2825 2546 -2791
rect 2590 -2825 2606 -2791
rect -1454 -2884 -1420 -2868
rect -6234 -2943 -6218 -2909
rect -6174 -2943 -6158 -2909
rect -6056 -2943 -6040 -2909
rect -5996 -2943 -5980 -2909
rect -5878 -2943 -5862 -2909
rect -5818 -2943 -5802 -2909
rect -5700 -2943 -5684 -2909
rect -5640 -2943 -5624 -2909
rect -5522 -2943 -5506 -2909
rect -5462 -2943 -5446 -2909
rect -5344 -2943 -5328 -2909
rect -5284 -2943 -5268 -2909
rect -5166 -2943 -5150 -2909
rect -5106 -2943 -5090 -2909
rect -4988 -2943 -4972 -2909
rect -4928 -2943 -4912 -2909
rect -4810 -2943 -4794 -2909
rect -4750 -2943 -4734 -2909
rect -4632 -2943 -4616 -2909
rect -4572 -2943 -4556 -2909
rect -4454 -2943 -4438 -2909
rect -4394 -2943 -4378 -2909
rect -4276 -2943 -4260 -2909
rect -4216 -2943 -4200 -2909
rect -4098 -2943 -4082 -2909
rect -4038 -2943 -4022 -2909
rect -3920 -2943 -3904 -2909
rect -3860 -2943 -3844 -2909
rect -3742 -2943 -3726 -2909
rect -3682 -2943 -3666 -2909
rect -3564 -2943 -3548 -2909
rect -3504 -2943 -3488 -2909
rect -6302 -3002 -6268 -2986
rect -6302 -3274 -6268 -3258
rect -6124 -3002 -6090 -2986
rect -6124 -3274 -6090 -3258
rect -5946 -3002 -5912 -2986
rect -5946 -3274 -5912 -3258
rect -5768 -3002 -5734 -2986
rect -5768 -3274 -5734 -3258
rect -5590 -3002 -5556 -2986
rect -5590 -3274 -5556 -3258
rect -5412 -3002 -5378 -2986
rect -5412 -3274 -5378 -3258
rect -5234 -3002 -5200 -2986
rect -5234 -3274 -5200 -3258
rect -5056 -3002 -5022 -2986
rect -5056 -3274 -5022 -3258
rect -4878 -3002 -4844 -2986
rect -4878 -3274 -4844 -3258
rect -4700 -3002 -4666 -2986
rect -4700 -3274 -4666 -3258
rect -4522 -3002 -4488 -2986
rect -4522 -3274 -4488 -3258
rect -4344 -3002 -4310 -2986
rect -4344 -3274 -4310 -3258
rect -4166 -3002 -4132 -2986
rect -4166 -3274 -4132 -3258
rect -3988 -3002 -3954 -2986
rect -3988 -3274 -3954 -3258
rect -3810 -3002 -3776 -2986
rect -3810 -3274 -3776 -3258
rect -3632 -3002 -3598 -2986
rect -3632 -3274 -3598 -3258
rect -3454 -3002 -3420 -2986
rect -1454 -3156 -1420 -3140
rect -1276 -2884 -1242 -2868
rect -1276 -3156 -1242 -3140
rect -1098 -2884 -1064 -2868
rect -1098 -3156 -1064 -3140
rect -920 -2884 -886 -2868
rect -920 -3156 -886 -3140
rect -742 -2884 -708 -2868
rect -742 -3156 -708 -3140
rect -564 -2884 -530 -2868
rect -564 -3156 -530 -3140
rect -386 -2884 -352 -2868
rect -386 -3156 -352 -3140
rect -208 -2884 -174 -2868
rect -208 -3156 -174 -3140
rect -30 -2884 4 -2868
rect -30 -3156 4 -3140
rect 148 -2884 182 -2868
rect 148 -3156 182 -3140
rect 326 -2884 360 -2868
rect 326 -3156 360 -3140
rect 504 -2884 538 -2868
rect 504 -3156 538 -3140
rect 682 -2884 716 -2868
rect 682 -3156 716 -3140
rect 860 -2884 894 -2868
rect 860 -3156 894 -3140
rect 1038 -2884 1072 -2868
rect 1038 -3156 1072 -3140
rect 1216 -2884 1250 -2868
rect 1216 -3156 1250 -3140
rect 1394 -2884 1428 -2868
rect 1394 -3156 1428 -3140
rect 1572 -2884 1606 -2868
rect 1572 -3156 1606 -3140
rect 1750 -2884 1784 -2868
rect 1750 -3156 1784 -3140
rect 1928 -2884 1962 -2868
rect 1928 -3156 1962 -3140
rect 2106 -2884 2140 -2868
rect 2106 -3156 2140 -3140
rect 2284 -2884 2318 -2868
rect 2284 -3156 2318 -3140
rect 2462 -2884 2496 -2868
rect 2462 -3156 2496 -3140
rect 2640 -2884 2674 -2868
rect 2640 -3156 2674 -3140
rect -1386 -3233 -1370 -3199
rect -1326 -3233 -1310 -3199
rect -1208 -3233 -1192 -3199
rect -1148 -3233 -1132 -3199
rect -1030 -3233 -1014 -3199
rect -970 -3233 -954 -3199
rect -852 -3233 -836 -3199
rect -792 -3233 -776 -3199
rect -674 -3233 -658 -3199
rect -614 -3233 -598 -3199
rect -496 -3233 -480 -3199
rect -436 -3233 -420 -3199
rect -318 -3233 -302 -3199
rect -258 -3233 -242 -3199
rect -140 -3233 -124 -3199
rect -80 -3233 -64 -3199
rect 38 -3233 54 -3199
rect 98 -3233 114 -3199
rect 216 -3233 232 -3199
rect 276 -3233 292 -3199
rect 394 -3233 410 -3199
rect 454 -3233 470 -3199
rect 572 -3233 588 -3199
rect 632 -3233 648 -3199
rect 750 -3233 766 -3199
rect 810 -3233 826 -3199
rect 928 -3233 944 -3199
rect 988 -3233 1004 -3199
rect 1106 -3233 1122 -3199
rect 1166 -3233 1182 -3199
rect 1284 -3233 1300 -3199
rect 1344 -3233 1360 -3199
rect 1462 -3233 1478 -3199
rect 1522 -3233 1538 -3199
rect 1640 -3233 1656 -3199
rect 1700 -3233 1716 -3199
rect 1818 -3233 1834 -3199
rect 1878 -3233 1894 -3199
rect 1996 -3233 2012 -3199
rect 2056 -3233 2072 -3199
rect 2174 -3233 2190 -3199
rect 2234 -3233 2250 -3199
rect 2352 -3233 2368 -3199
rect 2412 -3233 2428 -3199
rect 2530 -3233 2546 -3199
rect 2590 -3233 2606 -3199
rect -3454 -3274 -3420 -3258
rect -6234 -3351 -6218 -3317
rect -6174 -3351 -6158 -3317
rect -6056 -3351 -6040 -3317
rect -5996 -3351 -5980 -3317
rect -5878 -3351 -5862 -3317
rect -5818 -3351 -5802 -3317
rect -5700 -3351 -5684 -3317
rect -5640 -3351 -5624 -3317
rect -5522 -3351 -5506 -3317
rect -5462 -3351 -5446 -3317
rect -5344 -3351 -5328 -3317
rect -5284 -3351 -5268 -3317
rect -5166 -3351 -5150 -3317
rect -5106 -3351 -5090 -3317
rect -4988 -3351 -4972 -3317
rect -4928 -3351 -4912 -3317
rect -4810 -3351 -4794 -3317
rect -4750 -3351 -4734 -3317
rect -4632 -3351 -4616 -3317
rect -4572 -3351 -4556 -3317
rect -4454 -3351 -4438 -3317
rect -4394 -3351 -4378 -3317
rect -4276 -3351 -4260 -3317
rect -4216 -3351 -4200 -3317
rect -4098 -3351 -4082 -3317
rect -4038 -3351 -4022 -3317
rect -3920 -3351 -3904 -3317
rect -3860 -3351 -3844 -3317
rect -3742 -3351 -3726 -3317
rect -3682 -3351 -3666 -3317
rect -3564 -3351 -3548 -3317
rect -3504 -3351 -3488 -3317
rect -1386 -3725 -1370 -3691
rect -1326 -3725 -1310 -3691
rect -1208 -3725 -1192 -3691
rect -1148 -3725 -1132 -3691
rect -1030 -3725 -1014 -3691
rect -970 -3725 -954 -3691
rect -852 -3725 -836 -3691
rect -792 -3725 -776 -3691
rect -674 -3725 -658 -3691
rect -614 -3725 -598 -3691
rect -496 -3725 -480 -3691
rect -436 -3725 -420 -3691
rect -318 -3725 -302 -3691
rect -258 -3725 -242 -3691
rect -140 -3725 -124 -3691
rect -80 -3725 -64 -3691
rect 38 -3725 54 -3691
rect 98 -3725 114 -3691
rect 216 -3725 232 -3691
rect 276 -3725 292 -3691
rect 394 -3725 410 -3691
rect 454 -3725 470 -3691
rect 572 -3725 588 -3691
rect 632 -3725 648 -3691
rect 750 -3725 766 -3691
rect 810 -3725 826 -3691
rect 928 -3725 944 -3691
rect 988 -3725 1004 -3691
rect 1106 -3725 1122 -3691
rect 1166 -3725 1182 -3691
rect 1284 -3725 1300 -3691
rect 1344 -3725 1360 -3691
rect 1462 -3725 1478 -3691
rect 1522 -3725 1538 -3691
rect 1640 -3725 1656 -3691
rect 1700 -3725 1716 -3691
rect 1818 -3725 1834 -3691
rect 1878 -3725 1894 -3691
rect 1996 -3725 2012 -3691
rect 2056 -3725 2072 -3691
rect 2174 -3725 2190 -3691
rect 2234 -3725 2250 -3691
rect 2352 -3725 2368 -3691
rect 2412 -3725 2428 -3691
rect 2530 -3725 2546 -3691
rect 2590 -3725 2606 -3691
rect -6234 -3813 -6218 -3779
rect -6174 -3813 -6158 -3779
rect -6056 -3813 -6040 -3779
rect -5996 -3813 -5980 -3779
rect -5878 -3813 -5862 -3779
rect -5818 -3813 -5802 -3779
rect -5700 -3813 -5684 -3779
rect -5640 -3813 -5624 -3779
rect -5522 -3813 -5506 -3779
rect -5462 -3813 -5446 -3779
rect -5344 -3813 -5328 -3779
rect -5284 -3813 -5268 -3779
rect -5166 -3813 -5150 -3779
rect -5106 -3813 -5090 -3779
rect -4988 -3813 -4972 -3779
rect -4928 -3813 -4912 -3779
rect -4810 -3813 -4794 -3779
rect -4750 -3813 -4734 -3779
rect -4632 -3813 -4616 -3779
rect -4572 -3813 -4556 -3779
rect -4454 -3813 -4438 -3779
rect -4394 -3813 -4378 -3779
rect -4276 -3813 -4260 -3779
rect -4216 -3813 -4200 -3779
rect -4098 -3813 -4082 -3779
rect -4038 -3813 -4022 -3779
rect -3920 -3813 -3904 -3779
rect -3860 -3813 -3844 -3779
rect -3742 -3813 -3726 -3779
rect -3682 -3813 -3666 -3779
rect -3564 -3813 -3548 -3779
rect -3504 -3813 -3488 -3779
rect -1454 -3784 -1420 -3768
rect -6302 -3872 -6268 -3856
rect -6302 -4144 -6268 -4128
rect -6124 -3872 -6090 -3856
rect -6124 -4144 -6090 -4128
rect -5946 -3872 -5912 -3856
rect -5946 -4144 -5912 -4128
rect -5768 -3872 -5734 -3856
rect -5768 -4144 -5734 -4128
rect -5590 -3872 -5556 -3856
rect -5590 -4144 -5556 -4128
rect -5412 -3872 -5378 -3856
rect -5412 -4144 -5378 -4128
rect -5234 -3872 -5200 -3856
rect -5234 -4144 -5200 -4128
rect -5056 -3872 -5022 -3856
rect -5056 -4144 -5022 -4128
rect -4878 -3872 -4844 -3856
rect -4878 -4144 -4844 -4128
rect -4700 -3872 -4666 -3856
rect -4700 -4144 -4666 -4128
rect -4522 -3872 -4488 -3856
rect -4522 -4144 -4488 -4128
rect -4344 -3872 -4310 -3856
rect -4344 -4144 -4310 -4128
rect -4166 -3872 -4132 -3856
rect -4166 -4144 -4132 -4128
rect -3988 -3872 -3954 -3856
rect -3988 -4144 -3954 -4128
rect -3810 -3872 -3776 -3856
rect -3810 -4144 -3776 -4128
rect -3632 -3872 -3598 -3856
rect -3632 -4144 -3598 -4128
rect -3454 -3872 -3420 -3856
rect -1454 -4056 -1420 -4040
rect -1276 -3784 -1242 -3768
rect -1276 -4056 -1242 -4040
rect -1098 -3784 -1064 -3768
rect -1098 -4056 -1064 -4040
rect -920 -3784 -886 -3768
rect -920 -4056 -886 -4040
rect -742 -3784 -708 -3768
rect -742 -4056 -708 -4040
rect -564 -3784 -530 -3768
rect -564 -4056 -530 -4040
rect -386 -3784 -352 -3768
rect -386 -4056 -352 -4040
rect -208 -3784 -174 -3768
rect -208 -4056 -174 -4040
rect -30 -3784 4 -3768
rect -30 -4056 4 -4040
rect 148 -3784 182 -3768
rect 148 -4056 182 -4040
rect 326 -3784 360 -3768
rect 326 -4056 360 -4040
rect 504 -3784 538 -3768
rect 504 -4056 538 -4040
rect 682 -3784 716 -3768
rect 682 -4056 716 -4040
rect 860 -3784 894 -3768
rect 860 -4056 894 -4040
rect 1038 -3784 1072 -3768
rect 1038 -4056 1072 -4040
rect 1216 -3784 1250 -3768
rect 1216 -4056 1250 -4040
rect 1394 -3784 1428 -3768
rect 1394 -4056 1428 -4040
rect 1572 -3784 1606 -3768
rect 1572 -4056 1606 -4040
rect 1750 -3784 1784 -3768
rect 1750 -4056 1784 -4040
rect 1928 -3784 1962 -3768
rect 1928 -4056 1962 -4040
rect 2106 -3784 2140 -3768
rect 2106 -4056 2140 -4040
rect 2284 -3784 2318 -3768
rect 2284 -4056 2318 -4040
rect 2462 -3784 2496 -3768
rect 2462 -4056 2496 -4040
rect 2640 -3784 2674 -3768
rect 2640 -4056 2674 -4040
rect -3454 -4144 -3420 -4128
rect -1386 -4133 -1370 -4099
rect -1326 -4133 -1310 -4099
rect -1208 -4133 -1192 -4099
rect -1148 -4133 -1132 -4099
rect -1030 -4133 -1014 -4099
rect -970 -4133 -954 -4099
rect -852 -4133 -836 -4099
rect -792 -4133 -776 -4099
rect -674 -4133 -658 -4099
rect -614 -4133 -598 -4099
rect -496 -4133 -480 -4099
rect -436 -4133 -420 -4099
rect -318 -4133 -302 -4099
rect -258 -4133 -242 -4099
rect -140 -4133 -124 -4099
rect -80 -4133 -64 -4099
rect 38 -4133 54 -4099
rect 98 -4133 114 -4099
rect 216 -4133 232 -4099
rect 276 -4133 292 -4099
rect 394 -4133 410 -4099
rect 454 -4133 470 -4099
rect 572 -4133 588 -4099
rect 632 -4133 648 -4099
rect 750 -4133 766 -4099
rect 810 -4133 826 -4099
rect 928 -4133 944 -4099
rect 988 -4133 1004 -4099
rect 1106 -4133 1122 -4099
rect 1166 -4133 1182 -4099
rect 1284 -4133 1300 -4099
rect 1344 -4133 1360 -4099
rect 1462 -4133 1478 -4099
rect 1522 -4133 1538 -4099
rect 1640 -4133 1656 -4099
rect 1700 -4133 1716 -4099
rect 1818 -4133 1834 -4099
rect 1878 -4133 1894 -4099
rect 1996 -4133 2012 -4099
rect 2056 -4133 2072 -4099
rect 2174 -4133 2190 -4099
rect 2234 -4133 2250 -4099
rect 2352 -4133 2368 -4099
rect 2412 -4133 2428 -4099
rect 2530 -4133 2546 -4099
rect 2590 -4133 2606 -4099
rect -6234 -4221 -6218 -4187
rect -6174 -4221 -6158 -4187
rect -6056 -4221 -6040 -4187
rect -5996 -4221 -5980 -4187
rect -5878 -4221 -5862 -4187
rect -5818 -4221 -5802 -4187
rect -5700 -4221 -5684 -4187
rect -5640 -4221 -5624 -4187
rect -5522 -4221 -5506 -4187
rect -5462 -4221 -5446 -4187
rect -5344 -4221 -5328 -4187
rect -5284 -4221 -5268 -4187
rect -5166 -4221 -5150 -4187
rect -5106 -4221 -5090 -4187
rect -4988 -4221 -4972 -4187
rect -4928 -4221 -4912 -4187
rect -4810 -4221 -4794 -4187
rect -4750 -4221 -4734 -4187
rect -4632 -4221 -4616 -4187
rect -4572 -4221 -4556 -4187
rect -4454 -4221 -4438 -4187
rect -4394 -4221 -4378 -4187
rect -4276 -4221 -4260 -4187
rect -4216 -4221 -4200 -4187
rect -4098 -4221 -4082 -4187
rect -4038 -4221 -4022 -4187
rect -3920 -4221 -3904 -4187
rect -3860 -4221 -3844 -4187
rect -3742 -4221 -3726 -4187
rect -3682 -4221 -3666 -4187
rect -3564 -4221 -3548 -4187
rect -3504 -4221 -3488 -4187
rect -1386 -4625 -1370 -4591
rect -1326 -4625 -1310 -4591
rect -1208 -4625 -1192 -4591
rect -1148 -4625 -1132 -4591
rect -1030 -4625 -1014 -4591
rect -970 -4625 -954 -4591
rect -852 -4625 -836 -4591
rect -792 -4625 -776 -4591
rect -674 -4625 -658 -4591
rect -614 -4625 -598 -4591
rect -496 -4625 -480 -4591
rect -436 -4625 -420 -4591
rect -318 -4625 -302 -4591
rect -258 -4625 -242 -4591
rect -140 -4625 -124 -4591
rect -80 -4625 -64 -4591
rect 38 -4625 54 -4591
rect 98 -4625 114 -4591
rect 216 -4625 232 -4591
rect 276 -4625 292 -4591
rect 394 -4625 410 -4591
rect 454 -4625 470 -4591
rect 572 -4625 588 -4591
rect 632 -4625 648 -4591
rect 750 -4625 766 -4591
rect 810 -4625 826 -4591
rect 928 -4625 944 -4591
rect 988 -4625 1004 -4591
rect 1106 -4625 1122 -4591
rect 1166 -4625 1182 -4591
rect 1284 -4625 1300 -4591
rect 1344 -4625 1360 -4591
rect 1462 -4625 1478 -4591
rect 1522 -4625 1538 -4591
rect 1640 -4625 1656 -4591
rect 1700 -4625 1716 -4591
rect 1818 -4625 1834 -4591
rect 1878 -4625 1894 -4591
rect 1996 -4625 2012 -4591
rect 2056 -4625 2072 -4591
rect 2174 -4625 2190 -4591
rect 2234 -4625 2250 -4591
rect 2352 -4625 2368 -4591
rect 2412 -4625 2428 -4591
rect 2530 -4625 2546 -4591
rect 2590 -4625 2606 -4591
rect -6234 -4683 -6218 -4649
rect -6174 -4683 -6158 -4649
rect -6056 -4683 -6040 -4649
rect -5996 -4683 -5980 -4649
rect -5878 -4683 -5862 -4649
rect -5818 -4683 -5802 -4649
rect -5700 -4683 -5684 -4649
rect -5640 -4683 -5624 -4649
rect -5522 -4683 -5506 -4649
rect -5462 -4683 -5446 -4649
rect -5344 -4683 -5328 -4649
rect -5284 -4683 -5268 -4649
rect -5166 -4683 -5150 -4649
rect -5106 -4683 -5090 -4649
rect -4988 -4683 -4972 -4649
rect -4928 -4683 -4912 -4649
rect -4810 -4683 -4794 -4649
rect -4750 -4683 -4734 -4649
rect -4632 -4683 -4616 -4649
rect -4572 -4683 -4556 -4649
rect -4454 -4683 -4438 -4649
rect -4394 -4683 -4378 -4649
rect -4276 -4683 -4260 -4649
rect -4216 -4683 -4200 -4649
rect -4098 -4683 -4082 -4649
rect -4038 -4683 -4022 -4649
rect -3920 -4683 -3904 -4649
rect -3860 -4683 -3844 -4649
rect -3742 -4683 -3726 -4649
rect -3682 -4683 -3666 -4649
rect -3564 -4683 -3548 -4649
rect -3504 -4683 -3488 -4649
rect -1454 -4684 -1420 -4668
rect -6302 -4742 -6268 -4726
rect -6302 -5014 -6268 -4998
rect -6124 -4742 -6090 -4726
rect -6124 -5014 -6090 -4998
rect -5946 -4742 -5912 -4726
rect -5946 -5014 -5912 -4998
rect -5768 -4742 -5734 -4726
rect -5768 -5014 -5734 -4998
rect -5590 -4742 -5556 -4726
rect -5590 -5014 -5556 -4998
rect -5412 -4742 -5378 -4726
rect -5412 -5014 -5378 -4998
rect -5234 -4742 -5200 -4726
rect -5234 -5014 -5200 -4998
rect -5056 -4742 -5022 -4726
rect -5056 -5014 -5022 -4998
rect -4878 -4742 -4844 -4726
rect -4878 -5014 -4844 -4998
rect -4700 -4742 -4666 -4726
rect -4700 -5014 -4666 -4998
rect -4522 -4742 -4488 -4726
rect -4522 -5014 -4488 -4998
rect -4344 -4742 -4310 -4726
rect -4344 -5014 -4310 -4998
rect -4166 -4742 -4132 -4726
rect -4166 -5014 -4132 -4998
rect -3988 -4742 -3954 -4726
rect -3988 -5014 -3954 -4998
rect -3810 -4742 -3776 -4726
rect -3810 -5014 -3776 -4998
rect -3632 -4742 -3598 -4726
rect -3632 -5014 -3598 -4998
rect -3454 -4742 -3420 -4726
rect -1454 -4956 -1420 -4940
rect -1276 -4684 -1242 -4668
rect -1276 -4956 -1242 -4940
rect -1098 -4684 -1064 -4668
rect -1098 -4956 -1064 -4940
rect -920 -4684 -886 -4668
rect -920 -4956 -886 -4940
rect -742 -4684 -708 -4668
rect -742 -4956 -708 -4940
rect -564 -4684 -530 -4668
rect -564 -4956 -530 -4940
rect -386 -4684 -352 -4668
rect -386 -4956 -352 -4940
rect -208 -4684 -174 -4668
rect -208 -4956 -174 -4940
rect -30 -4684 4 -4668
rect -30 -4956 4 -4940
rect 148 -4684 182 -4668
rect 148 -4956 182 -4940
rect 326 -4684 360 -4668
rect 326 -4956 360 -4940
rect 504 -4684 538 -4668
rect 504 -4956 538 -4940
rect 682 -4684 716 -4668
rect 682 -4956 716 -4940
rect 860 -4684 894 -4668
rect 860 -4956 894 -4940
rect 1038 -4684 1072 -4668
rect 1038 -4956 1072 -4940
rect 1216 -4684 1250 -4668
rect 1216 -4956 1250 -4940
rect 1394 -4684 1428 -4668
rect 1394 -4956 1428 -4940
rect 1572 -4684 1606 -4668
rect 1572 -4956 1606 -4940
rect 1750 -4684 1784 -4668
rect 1750 -4956 1784 -4940
rect 1928 -4684 1962 -4668
rect 1928 -4956 1962 -4940
rect 2106 -4684 2140 -4668
rect 2106 -4956 2140 -4940
rect 2284 -4684 2318 -4668
rect 2284 -4956 2318 -4940
rect 2462 -4684 2496 -4668
rect 2462 -4956 2496 -4940
rect 2640 -4684 2674 -4668
rect 2640 -4956 2674 -4940
rect -3454 -5014 -3420 -4998
rect -1386 -5033 -1370 -4999
rect -1326 -5033 -1310 -4999
rect -1208 -5033 -1192 -4999
rect -1148 -5033 -1132 -4999
rect -1030 -5033 -1014 -4999
rect -970 -5033 -954 -4999
rect -852 -5033 -836 -4999
rect -792 -5033 -776 -4999
rect -674 -5033 -658 -4999
rect -614 -5033 -598 -4999
rect -496 -5033 -480 -4999
rect -436 -5033 -420 -4999
rect -318 -5033 -302 -4999
rect -258 -5033 -242 -4999
rect -140 -5033 -124 -4999
rect -80 -5033 -64 -4999
rect 38 -5033 54 -4999
rect 98 -5033 114 -4999
rect 216 -5033 232 -4999
rect 276 -5033 292 -4999
rect 394 -5033 410 -4999
rect 454 -5033 470 -4999
rect 572 -5033 588 -4999
rect 632 -5033 648 -4999
rect 750 -5033 766 -4999
rect 810 -5033 826 -4999
rect 928 -5033 944 -4999
rect 988 -5033 1004 -4999
rect 1106 -5033 1122 -4999
rect 1166 -5033 1182 -4999
rect 1284 -5033 1300 -4999
rect 1344 -5033 1360 -4999
rect 1462 -5033 1478 -4999
rect 1522 -5033 1538 -4999
rect 1640 -5033 1656 -4999
rect 1700 -5033 1716 -4999
rect 1818 -5033 1834 -4999
rect 1878 -5033 1894 -4999
rect 1996 -5033 2012 -4999
rect 2056 -5033 2072 -4999
rect 2174 -5033 2190 -4999
rect 2234 -5033 2250 -4999
rect 2352 -5033 2368 -4999
rect 2412 -5033 2428 -4999
rect 2530 -5033 2546 -4999
rect 2590 -5033 2606 -4999
rect -6234 -5091 -6218 -5057
rect -6174 -5091 -6158 -5057
rect -6056 -5091 -6040 -5057
rect -5996 -5091 -5980 -5057
rect -5878 -5091 -5862 -5057
rect -5818 -5091 -5802 -5057
rect -5700 -5091 -5684 -5057
rect -5640 -5091 -5624 -5057
rect -5522 -5091 -5506 -5057
rect -5462 -5091 -5446 -5057
rect -5344 -5091 -5328 -5057
rect -5284 -5091 -5268 -5057
rect -5166 -5091 -5150 -5057
rect -5106 -5091 -5090 -5057
rect -4988 -5091 -4972 -5057
rect -4928 -5091 -4912 -5057
rect -4810 -5091 -4794 -5057
rect -4750 -5091 -4734 -5057
rect -4632 -5091 -4616 -5057
rect -4572 -5091 -4556 -5057
rect -4454 -5091 -4438 -5057
rect -4394 -5091 -4378 -5057
rect -4276 -5091 -4260 -5057
rect -4216 -5091 -4200 -5057
rect -4098 -5091 -4082 -5057
rect -4038 -5091 -4022 -5057
rect -3920 -5091 -3904 -5057
rect -3860 -5091 -3844 -5057
rect -3742 -5091 -3726 -5057
rect -3682 -5091 -3666 -5057
rect -3564 -5091 -3548 -5057
rect -3504 -5091 -3488 -5057
rect -6234 -5553 -6218 -5519
rect -6174 -5553 -6158 -5519
rect -6056 -5553 -6040 -5519
rect -5996 -5553 -5980 -5519
rect -5878 -5553 -5862 -5519
rect -5818 -5553 -5802 -5519
rect -5700 -5553 -5684 -5519
rect -5640 -5553 -5624 -5519
rect -5522 -5553 -5506 -5519
rect -5462 -5553 -5446 -5519
rect -5344 -5553 -5328 -5519
rect -5284 -5553 -5268 -5519
rect -5166 -5553 -5150 -5519
rect -5106 -5553 -5090 -5519
rect -4988 -5553 -4972 -5519
rect -4928 -5553 -4912 -5519
rect -4810 -5553 -4794 -5519
rect -4750 -5553 -4734 -5519
rect -4632 -5553 -4616 -5519
rect -4572 -5553 -4556 -5519
rect -4454 -5553 -4438 -5519
rect -4394 -5553 -4378 -5519
rect -4276 -5553 -4260 -5519
rect -4216 -5553 -4200 -5519
rect -4098 -5553 -4082 -5519
rect -4038 -5553 -4022 -5519
rect -3920 -5553 -3904 -5519
rect -3860 -5553 -3844 -5519
rect -3742 -5553 -3726 -5519
rect -3682 -5553 -3666 -5519
rect -3564 -5553 -3548 -5519
rect -3504 -5553 -3488 -5519
rect -1386 -5525 -1370 -5491
rect -1326 -5525 -1310 -5491
rect -1208 -5525 -1192 -5491
rect -1148 -5525 -1132 -5491
rect -1030 -5525 -1014 -5491
rect -970 -5525 -954 -5491
rect -852 -5525 -836 -5491
rect -792 -5525 -776 -5491
rect -674 -5525 -658 -5491
rect -614 -5525 -598 -5491
rect -496 -5525 -480 -5491
rect -436 -5525 -420 -5491
rect -318 -5525 -302 -5491
rect -258 -5525 -242 -5491
rect -140 -5525 -124 -5491
rect -80 -5525 -64 -5491
rect 38 -5525 54 -5491
rect 98 -5525 114 -5491
rect 216 -5525 232 -5491
rect 276 -5525 292 -5491
rect 394 -5525 410 -5491
rect 454 -5525 470 -5491
rect 572 -5525 588 -5491
rect 632 -5525 648 -5491
rect 750 -5525 766 -5491
rect 810 -5525 826 -5491
rect 928 -5525 944 -5491
rect 988 -5525 1004 -5491
rect 1106 -5525 1122 -5491
rect 1166 -5525 1182 -5491
rect 1284 -5525 1300 -5491
rect 1344 -5525 1360 -5491
rect 1462 -5525 1478 -5491
rect 1522 -5525 1538 -5491
rect 1640 -5525 1656 -5491
rect 1700 -5525 1716 -5491
rect 1818 -5525 1834 -5491
rect 1878 -5525 1894 -5491
rect 1996 -5525 2012 -5491
rect 2056 -5525 2072 -5491
rect 2174 -5525 2190 -5491
rect 2234 -5525 2250 -5491
rect 2352 -5525 2368 -5491
rect 2412 -5525 2428 -5491
rect 2530 -5525 2546 -5491
rect 2590 -5525 2606 -5491
rect -1454 -5584 -1420 -5568
rect -6302 -5612 -6268 -5596
rect -6302 -5884 -6268 -5868
rect -6124 -5612 -6090 -5596
rect -6124 -5884 -6090 -5868
rect -5946 -5612 -5912 -5596
rect -5946 -5884 -5912 -5868
rect -5768 -5612 -5734 -5596
rect -5768 -5884 -5734 -5868
rect -5590 -5612 -5556 -5596
rect -5590 -5884 -5556 -5868
rect -5412 -5612 -5378 -5596
rect -5412 -5884 -5378 -5868
rect -5234 -5612 -5200 -5596
rect -5234 -5884 -5200 -5868
rect -5056 -5612 -5022 -5596
rect -5056 -5884 -5022 -5868
rect -4878 -5612 -4844 -5596
rect -4878 -5884 -4844 -5868
rect -4700 -5612 -4666 -5596
rect -4700 -5884 -4666 -5868
rect -4522 -5612 -4488 -5596
rect -4522 -5884 -4488 -5868
rect -4344 -5612 -4310 -5596
rect -4344 -5884 -4310 -5868
rect -4166 -5612 -4132 -5596
rect -4166 -5884 -4132 -5868
rect -3988 -5612 -3954 -5596
rect -3988 -5884 -3954 -5868
rect -3810 -5612 -3776 -5596
rect -3810 -5884 -3776 -5868
rect -3632 -5612 -3598 -5596
rect -3632 -5884 -3598 -5868
rect -3454 -5612 -3420 -5596
rect -1454 -5856 -1420 -5840
rect -1276 -5584 -1242 -5568
rect -1276 -5856 -1242 -5840
rect -1098 -5584 -1064 -5568
rect -1098 -5856 -1064 -5840
rect -920 -5584 -886 -5568
rect -920 -5856 -886 -5840
rect -742 -5584 -708 -5568
rect -742 -5856 -708 -5840
rect -564 -5584 -530 -5568
rect -564 -5856 -530 -5840
rect -386 -5584 -352 -5568
rect -386 -5856 -352 -5840
rect -208 -5584 -174 -5568
rect -208 -5856 -174 -5840
rect -30 -5584 4 -5568
rect -30 -5856 4 -5840
rect 148 -5584 182 -5568
rect 148 -5856 182 -5840
rect 326 -5584 360 -5568
rect 326 -5856 360 -5840
rect 504 -5584 538 -5568
rect 504 -5856 538 -5840
rect 682 -5584 716 -5568
rect 682 -5856 716 -5840
rect 860 -5584 894 -5568
rect 860 -5856 894 -5840
rect 1038 -5584 1072 -5568
rect 1038 -5856 1072 -5840
rect 1216 -5584 1250 -5568
rect 1216 -5856 1250 -5840
rect 1394 -5584 1428 -5568
rect 1394 -5856 1428 -5840
rect 1572 -5584 1606 -5568
rect 1572 -5856 1606 -5840
rect 1750 -5584 1784 -5568
rect 1750 -5856 1784 -5840
rect 1928 -5584 1962 -5568
rect 1928 -5856 1962 -5840
rect 2106 -5584 2140 -5568
rect 2106 -5856 2140 -5840
rect 2284 -5584 2318 -5568
rect 2284 -5856 2318 -5840
rect 2462 -5584 2496 -5568
rect 2462 -5856 2496 -5840
rect 2640 -5584 2674 -5568
rect 2640 -5856 2674 -5840
rect -3454 -5884 -3420 -5868
rect -6234 -5961 -6218 -5927
rect -6174 -5961 -6158 -5927
rect -6056 -5961 -6040 -5927
rect -5996 -5961 -5980 -5927
rect -5878 -5961 -5862 -5927
rect -5818 -5961 -5802 -5927
rect -5700 -5961 -5684 -5927
rect -5640 -5961 -5624 -5927
rect -5522 -5961 -5506 -5927
rect -5462 -5961 -5446 -5927
rect -5344 -5961 -5328 -5927
rect -5284 -5961 -5268 -5927
rect -5166 -5961 -5150 -5927
rect -5106 -5961 -5090 -5927
rect -4988 -5961 -4972 -5927
rect -4928 -5961 -4912 -5927
rect -4810 -5961 -4794 -5927
rect -4750 -5961 -4734 -5927
rect -4632 -5961 -4616 -5927
rect -4572 -5961 -4556 -5927
rect -4454 -5961 -4438 -5927
rect -4394 -5961 -4378 -5927
rect -4276 -5961 -4260 -5927
rect -4216 -5961 -4200 -5927
rect -4098 -5961 -4082 -5927
rect -4038 -5961 -4022 -5927
rect -3920 -5961 -3904 -5927
rect -3860 -5961 -3844 -5927
rect -3742 -5961 -3726 -5927
rect -3682 -5961 -3666 -5927
rect -3564 -5961 -3548 -5927
rect -3504 -5961 -3488 -5927
rect -1386 -5933 -1370 -5899
rect -1326 -5933 -1310 -5899
rect -1208 -5933 -1192 -5899
rect -1148 -5933 -1132 -5899
rect -1030 -5933 -1014 -5899
rect -970 -5933 -954 -5899
rect -852 -5933 -836 -5899
rect -792 -5933 -776 -5899
rect -674 -5933 -658 -5899
rect -614 -5933 -598 -5899
rect -496 -5933 -480 -5899
rect -436 -5933 -420 -5899
rect -318 -5933 -302 -5899
rect -258 -5933 -242 -5899
rect -140 -5933 -124 -5899
rect -80 -5933 -64 -5899
rect 38 -5933 54 -5899
rect 98 -5933 114 -5899
rect 216 -5933 232 -5899
rect 276 -5933 292 -5899
rect 394 -5933 410 -5899
rect 454 -5933 470 -5899
rect 572 -5933 588 -5899
rect 632 -5933 648 -5899
rect 750 -5933 766 -5899
rect 810 -5933 826 -5899
rect 928 -5933 944 -5899
rect 988 -5933 1004 -5899
rect 1106 -5933 1122 -5899
rect 1166 -5933 1182 -5899
rect 1284 -5933 1300 -5899
rect 1344 -5933 1360 -5899
rect 1462 -5933 1478 -5899
rect 1522 -5933 1538 -5899
rect 1640 -5933 1656 -5899
rect 1700 -5933 1716 -5899
rect 1818 -5933 1834 -5899
rect 1878 -5933 1894 -5899
rect 1996 -5933 2012 -5899
rect 2056 -5933 2072 -5899
rect 2174 -5933 2190 -5899
rect 2234 -5933 2250 -5899
rect 2352 -5933 2368 -5899
rect 2412 -5933 2428 -5899
rect 2530 -5933 2546 -5899
rect 2590 -5933 2606 -5899
rect -7605 -7140 -7512 -6976
rect 3610 -7140 3703 -6989
rect -7605 -7233 -7282 -7140
rect 3426 -7233 3703 -7140
rect -7605 -7621 -7264 -7521
rect 13443 -7621 13719 -7521
rect -7605 -7850 -7505 -7621
rect 13619 -7731 13719 -7621
rect -5560 -7824 -5544 -7790
rect -5500 -7824 -5484 -7790
rect -5382 -7824 -5366 -7790
rect -5322 -7824 -5306 -7790
rect -5204 -7824 -5188 -7790
rect -5144 -7824 -5128 -7790
rect -5026 -7824 -5010 -7790
rect -4966 -7824 -4950 -7790
rect -4848 -7824 -4832 -7790
rect -4788 -7824 -4772 -7790
rect -4670 -7824 -4654 -7790
rect -4610 -7824 -4594 -7790
rect -4492 -7824 -4476 -7790
rect -4432 -7824 -4416 -7790
rect -4314 -7824 -4298 -7790
rect -4254 -7824 -4238 -7790
rect -4136 -7824 -4120 -7790
rect -4076 -7824 -4060 -7790
rect -5628 -7874 -5594 -7858
rect -5628 -8146 -5594 -8130
rect -5450 -7874 -5416 -7858
rect -5450 -8146 -5416 -8130
rect -5272 -7874 -5238 -7858
rect -5272 -8146 -5238 -8130
rect -5094 -7874 -5060 -7858
rect -5094 -8146 -5060 -8130
rect -4916 -7874 -4882 -7858
rect -4916 -8146 -4882 -8130
rect -4738 -7874 -4704 -7858
rect -4738 -8146 -4704 -8130
rect -4560 -7874 -4526 -7858
rect -4560 -8146 -4526 -8130
rect -4382 -7874 -4348 -7858
rect -4382 -8146 -4348 -8130
rect -4204 -7874 -4170 -7858
rect -4204 -8146 -4170 -8130
rect -4026 -7874 -3992 -7858
rect -2105 -8082 -2089 -8048
rect -2045 -8082 -2029 -8048
rect -1927 -8082 -1911 -8048
rect -1867 -8082 -1851 -8048
rect -1749 -8082 -1733 -8048
rect -1689 -8082 -1673 -8048
rect -1571 -8082 -1555 -8048
rect -1511 -8082 -1495 -8048
rect -1393 -8082 -1377 -8048
rect -1333 -8082 -1317 -8048
rect -1215 -8082 -1199 -8048
rect -1155 -8082 -1139 -8048
rect -1037 -8082 -1021 -8048
rect -977 -8082 -961 -8048
rect -859 -8082 -843 -8048
rect -799 -8082 -783 -8048
rect -681 -8082 -665 -8048
rect -621 -8082 -605 -8048
rect -503 -8082 -487 -8048
rect -443 -8082 -427 -8048
rect -325 -8082 -309 -8048
rect -265 -8082 -249 -8048
rect -147 -8082 -131 -8048
rect -87 -8082 -71 -8048
rect 31 -8082 47 -8048
rect 91 -8082 107 -8048
rect 209 -8082 225 -8048
rect 269 -8082 285 -8048
rect 387 -8082 403 -8048
rect 447 -8082 463 -8048
rect 565 -8082 581 -8048
rect 625 -8082 641 -8048
rect 743 -8082 759 -8048
rect 803 -8082 819 -8048
rect 921 -8082 937 -8048
rect 981 -8082 997 -8048
rect 1099 -8082 1115 -8048
rect 1159 -8082 1175 -8048
rect 1277 -8082 1293 -8048
rect 1337 -8082 1353 -8048
rect 1455 -8082 1471 -8048
rect 1515 -8082 1531 -8048
rect 1633 -8082 1649 -8048
rect 1693 -8082 1709 -8048
rect 1811 -8082 1827 -8048
rect 1871 -8082 1887 -8048
rect 1989 -8082 2005 -8048
rect 2049 -8082 2065 -8048
rect 2167 -8082 2183 -8048
rect 2227 -8082 2243 -8048
rect 2345 -8082 2361 -8048
rect 2405 -8082 2421 -8048
rect 2523 -8082 2539 -8048
rect 2583 -8082 2599 -8048
rect 2701 -8082 2717 -8048
rect 2761 -8082 2777 -8048
rect 2879 -8082 2895 -8048
rect 2939 -8082 2955 -8048
rect 3057 -8082 3073 -8048
rect 3117 -8082 3133 -8048
rect 3235 -8082 3251 -8048
rect 3295 -8082 3311 -8048
rect 3413 -8082 3429 -8048
rect 3473 -8082 3489 -8048
rect 3591 -8082 3607 -8048
rect 3651 -8082 3667 -8048
rect 3769 -8082 3785 -8048
rect 3829 -8082 3845 -8048
rect 3947 -8082 3963 -8048
rect 4007 -8082 4023 -8048
rect -4026 -8146 -3992 -8130
rect -2173 -8132 -2139 -8116
rect -5560 -8214 -5544 -8180
rect -5500 -8214 -5484 -8180
rect -5382 -8214 -5366 -8180
rect -5322 -8214 -5306 -8180
rect -5204 -8214 -5188 -8180
rect -5144 -8214 -5128 -8180
rect -5026 -8214 -5010 -8180
rect -4966 -8214 -4950 -8180
rect -4848 -8214 -4832 -8180
rect -4788 -8214 -4772 -8180
rect -4670 -8214 -4654 -8180
rect -4610 -8214 -4594 -8180
rect -4492 -8214 -4476 -8180
rect -4432 -8214 -4416 -8180
rect -4314 -8214 -4298 -8180
rect -4254 -8214 -4238 -8180
rect -4136 -8214 -4120 -8180
rect -4076 -8214 -4060 -8180
rect -5560 -8374 -5544 -8340
rect -5500 -8374 -5484 -8340
rect -5382 -8374 -5366 -8340
rect -5322 -8374 -5306 -8340
rect -5204 -8374 -5188 -8340
rect -5144 -8374 -5128 -8340
rect -5026 -8374 -5010 -8340
rect -4966 -8374 -4950 -8340
rect -4848 -8374 -4832 -8340
rect -4788 -8374 -4772 -8340
rect -4670 -8374 -4654 -8340
rect -4610 -8374 -4594 -8340
rect -4492 -8374 -4476 -8340
rect -4432 -8374 -4416 -8340
rect -4314 -8374 -4298 -8340
rect -4254 -8374 -4238 -8340
rect -4136 -8374 -4120 -8340
rect -4076 -8374 -4060 -8340
rect -2173 -8404 -2139 -8388
rect -1995 -8132 -1961 -8116
rect -1995 -8404 -1961 -8388
rect -1817 -8132 -1783 -8116
rect -1817 -8404 -1783 -8388
rect -1639 -8132 -1605 -8116
rect -1639 -8404 -1605 -8388
rect -1461 -8132 -1427 -8116
rect -1461 -8404 -1427 -8388
rect -1283 -8132 -1249 -8116
rect -1283 -8404 -1249 -8388
rect -1105 -8132 -1071 -8116
rect -1105 -8404 -1071 -8388
rect -927 -8132 -893 -8116
rect -927 -8404 -893 -8388
rect -749 -8132 -715 -8116
rect -749 -8404 -715 -8388
rect -571 -8132 -537 -8116
rect -571 -8404 -537 -8388
rect -393 -8132 -359 -8116
rect -393 -8404 -359 -8388
rect -215 -8132 -181 -8116
rect -215 -8404 -181 -8388
rect -37 -8132 -3 -8116
rect -37 -8404 -3 -8388
rect 141 -8132 175 -8116
rect 141 -8404 175 -8388
rect 319 -8132 353 -8116
rect 319 -8404 353 -8388
rect 497 -8132 531 -8116
rect 497 -8404 531 -8388
rect 675 -8132 709 -8116
rect 675 -8404 709 -8388
rect 853 -8132 887 -8116
rect 853 -8404 887 -8388
rect 1031 -8132 1065 -8116
rect 1031 -8404 1065 -8388
rect 1209 -8132 1243 -8116
rect 1209 -8404 1243 -8388
rect 1387 -8132 1421 -8116
rect 1387 -8404 1421 -8388
rect 1565 -8132 1599 -8116
rect 1565 -8404 1599 -8388
rect 1743 -8132 1777 -8116
rect 1743 -8404 1777 -8388
rect 1921 -8132 1955 -8116
rect 1921 -8404 1955 -8388
rect 2099 -8132 2133 -8116
rect 2099 -8404 2133 -8388
rect 2277 -8132 2311 -8116
rect 2277 -8404 2311 -8388
rect 2455 -8132 2489 -8116
rect 2455 -8404 2489 -8388
rect 2633 -8132 2667 -8116
rect 2633 -8404 2667 -8388
rect 2811 -8132 2845 -8116
rect 2811 -8404 2845 -8388
rect 2989 -8132 3023 -8116
rect 2989 -8404 3023 -8388
rect 3167 -8132 3201 -8116
rect 3167 -8404 3201 -8388
rect 3345 -8132 3379 -8116
rect 3345 -8404 3379 -8388
rect 3523 -8132 3557 -8116
rect 3523 -8404 3557 -8388
rect 3701 -8132 3735 -8116
rect 3701 -8404 3735 -8388
rect 3879 -8132 3913 -8116
rect 3879 -8404 3913 -8388
rect 4057 -8132 4091 -8116
rect 4057 -8404 4091 -8388
rect -5628 -8424 -5594 -8408
rect -5628 -8696 -5594 -8680
rect -5450 -8424 -5416 -8408
rect -5450 -8696 -5416 -8680
rect -5272 -8424 -5238 -8408
rect -5272 -8696 -5238 -8680
rect -5094 -8424 -5060 -8408
rect -5094 -8696 -5060 -8680
rect -4916 -8424 -4882 -8408
rect -4916 -8696 -4882 -8680
rect -4738 -8424 -4704 -8408
rect -4738 -8696 -4704 -8680
rect -4560 -8424 -4526 -8408
rect -4560 -8696 -4526 -8680
rect -4382 -8424 -4348 -8408
rect -4382 -8696 -4348 -8680
rect -4204 -8424 -4170 -8408
rect -4204 -8696 -4170 -8680
rect -4026 -8424 -3992 -8408
rect -2105 -8472 -2089 -8438
rect -2045 -8472 -2029 -8438
rect -1927 -8472 -1911 -8438
rect -1867 -8472 -1851 -8438
rect -1749 -8472 -1733 -8438
rect -1689 -8472 -1673 -8438
rect -1571 -8472 -1555 -8438
rect -1511 -8472 -1495 -8438
rect -1393 -8472 -1377 -8438
rect -1333 -8472 -1317 -8438
rect -1215 -8472 -1199 -8438
rect -1155 -8472 -1139 -8438
rect -1037 -8472 -1021 -8438
rect -977 -8472 -961 -8438
rect -859 -8472 -843 -8438
rect -799 -8472 -783 -8438
rect -681 -8472 -665 -8438
rect -621 -8472 -605 -8438
rect -503 -8472 -487 -8438
rect -443 -8472 -427 -8438
rect -325 -8472 -309 -8438
rect -265 -8472 -249 -8438
rect -147 -8472 -131 -8438
rect -87 -8472 -71 -8438
rect 31 -8472 47 -8438
rect 91 -8472 107 -8438
rect 209 -8472 225 -8438
rect 269 -8472 285 -8438
rect 387 -8472 403 -8438
rect 447 -8472 463 -8438
rect 565 -8472 581 -8438
rect 625 -8472 641 -8438
rect 743 -8472 759 -8438
rect 803 -8472 819 -8438
rect 921 -8472 937 -8438
rect 981 -8472 997 -8438
rect 1099 -8472 1115 -8438
rect 1159 -8472 1175 -8438
rect 1277 -8472 1293 -8438
rect 1337 -8472 1353 -8438
rect 1455 -8472 1471 -8438
rect 1515 -8472 1531 -8438
rect 1633 -8472 1649 -8438
rect 1693 -8472 1709 -8438
rect 1811 -8472 1827 -8438
rect 1871 -8472 1887 -8438
rect 1989 -8472 2005 -8438
rect 2049 -8472 2065 -8438
rect 2167 -8472 2183 -8438
rect 2227 -8472 2243 -8438
rect 2345 -8472 2361 -8438
rect 2405 -8472 2421 -8438
rect 2523 -8472 2539 -8438
rect 2583 -8472 2599 -8438
rect 2701 -8472 2717 -8438
rect 2761 -8472 2777 -8438
rect 2879 -8472 2895 -8438
rect 2939 -8472 2955 -8438
rect 3057 -8472 3073 -8438
rect 3117 -8472 3133 -8438
rect 3235 -8472 3251 -8438
rect 3295 -8472 3311 -8438
rect 3413 -8472 3429 -8438
rect 3473 -8472 3489 -8438
rect 3591 -8472 3607 -8438
rect 3651 -8472 3667 -8438
rect 3769 -8472 3785 -8438
rect 3829 -8472 3845 -8438
rect 3947 -8472 3963 -8438
rect 4007 -8472 4023 -8438
rect -4026 -8696 -3992 -8680
rect -5560 -8764 -5544 -8730
rect -5500 -8764 -5484 -8730
rect -5382 -8764 -5366 -8730
rect -5322 -8764 -5306 -8730
rect -5204 -8764 -5188 -8730
rect -5144 -8764 -5128 -8730
rect -5026 -8764 -5010 -8730
rect -4966 -8764 -4950 -8730
rect -4848 -8764 -4832 -8730
rect -4788 -8764 -4772 -8730
rect -4670 -8764 -4654 -8730
rect -4610 -8764 -4594 -8730
rect -4492 -8764 -4476 -8730
rect -4432 -8764 -4416 -8730
rect -4314 -8764 -4298 -8730
rect -4254 -8764 -4238 -8730
rect -4136 -8764 -4120 -8730
rect -4076 -8764 -4060 -8730
rect 6580 -8844 6596 -8810
rect 6640 -8844 6656 -8810
rect 6758 -8844 6774 -8810
rect 6818 -8844 6834 -8810
rect 6936 -8844 6952 -8810
rect 6996 -8844 7012 -8810
rect 7114 -8844 7130 -8810
rect 7174 -8844 7190 -8810
rect 7292 -8844 7308 -8810
rect 7352 -8844 7368 -8810
rect 7470 -8844 7486 -8810
rect 7530 -8844 7546 -8810
rect 7648 -8844 7664 -8810
rect 7708 -8844 7724 -8810
rect 7826 -8844 7842 -8810
rect 7886 -8844 7902 -8810
rect 8004 -8844 8020 -8810
rect 8064 -8844 8080 -8810
rect 8182 -8844 8198 -8810
rect 8242 -8844 8258 -8810
rect 8360 -8844 8376 -8810
rect 8420 -8844 8436 -8810
rect 8538 -8844 8554 -8810
rect 8598 -8844 8614 -8810
rect 8716 -8844 8732 -8810
rect 8776 -8844 8792 -8810
rect 8894 -8844 8910 -8810
rect 8954 -8844 8970 -8810
rect 9072 -8844 9088 -8810
rect 9132 -8844 9148 -8810
rect 9250 -8844 9266 -8810
rect 9310 -8844 9326 -8810
rect 10840 -8874 10856 -8840
rect 10900 -8874 10916 -8840
rect 11132 -8874 11148 -8840
rect 11192 -8874 11208 -8840
rect 11424 -8874 11440 -8840
rect 11484 -8874 11500 -8840
rect 11716 -8874 11732 -8840
rect 11776 -8874 11792 -8840
rect 12008 -8874 12024 -8840
rect 12068 -8874 12084 -8840
rect 12300 -8874 12316 -8840
rect 12360 -8874 12376 -8840
rect 12592 -8874 12608 -8840
rect 12652 -8874 12668 -8840
rect -5560 -8924 -5544 -8890
rect -5500 -8924 -5484 -8890
rect -5382 -8924 -5366 -8890
rect -5322 -8924 -5306 -8890
rect -5204 -8924 -5188 -8890
rect -5144 -8924 -5128 -8890
rect -5026 -8924 -5010 -8890
rect -4966 -8924 -4950 -8890
rect -4848 -8924 -4832 -8890
rect -4788 -8924 -4772 -8890
rect -4670 -8924 -4654 -8890
rect -4610 -8924 -4594 -8890
rect -4492 -8924 -4476 -8890
rect -4432 -8924 -4416 -8890
rect -4314 -8924 -4298 -8890
rect -4254 -8924 -4238 -8890
rect -4136 -8924 -4120 -8890
rect -4076 -8924 -4060 -8890
rect 6512 -8894 6546 -8878
rect -5628 -8974 -5594 -8958
rect -5628 -9246 -5594 -9230
rect -5450 -8974 -5416 -8958
rect -5450 -9246 -5416 -9230
rect -5272 -8974 -5238 -8958
rect -5272 -9246 -5238 -9230
rect -5094 -8974 -5060 -8958
rect -5094 -9246 -5060 -9230
rect -4916 -8974 -4882 -8958
rect -4916 -9246 -4882 -9230
rect -4738 -8974 -4704 -8958
rect -4738 -9246 -4704 -9230
rect -4560 -8974 -4526 -8958
rect -4560 -9246 -4526 -9230
rect -4382 -8974 -4348 -8958
rect -4382 -9246 -4348 -9230
rect -4204 -8974 -4170 -8958
rect -4204 -9246 -4170 -9230
rect -4026 -8974 -3992 -8958
rect -2105 -9082 -2089 -9048
rect -2045 -9082 -2029 -9048
rect -1927 -9082 -1911 -9048
rect -1867 -9082 -1851 -9048
rect -1749 -9082 -1733 -9048
rect -1689 -9082 -1673 -9048
rect -1571 -9082 -1555 -9048
rect -1511 -9082 -1495 -9048
rect -1393 -9082 -1377 -9048
rect -1333 -9082 -1317 -9048
rect -1215 -9082 -1199 -9048
rect -1155 -9082 -1139 -9048
rect -1037 -9082 -1021 -9048
rect -977 -9082 -961 -9048
rect -859 -9082 -843 -9048
rect -799 -9082 -783 -9048
rect -681 -9082 -665 -9048
rect -621 -9082 -605 -9048
rect -503 -9082 -487 -9048
rect -443 -9082 -427 -9048
rect -325 -9082 -309 -9048
rect -265 -9082 -249 -9048
rect -147 -9082 -131 -9048
rect -87 -9082 -71 -9048
rect 31 -9082 47 -9048
rect 91 -9082 107 -9048
rect 209 -9082 225 -9048
rect 269 -9082 285 -9048
rect 387 -9082 403 -9048
rect 447 -9082 463 -9048
rect 565 -9082 581 -9048
rect 625 -9082 641 -9048
rect 743 -9082 759 -9048
rect 803 -9082 819 -9048
rect 921 -9082 937 -9048
rect 981 -9082 997 -9048
rect 1099 -9082 1115 -9048
rect 1159 -9082 1175 -9048
rect 1277 -9082 1293 -9048
rect 1337 -9082 1353 -9048
rect 1455 -9082 1471 -9048
rect 1515 -9082 1531 -9048
rect 1633 -9082 1649 -9048
rect 1693 -9082 1709 -9048
rect 1811 -9082 1827 -9048
rect 1871 -9082 1887 -9048
rect 1989 -9082 2005 -9048
rect 2049 -9082 2065 -9048
rect 2167 -9082 2183 -9048
rect 2227 -9082 2243 -9048
rect 2345 -9082 2361 -9048
rect 2405 -9082 2421 -9048
rect 2523 -9082 2539 -9048
rect 2583 -9082 2599 -9048
rect 2701 -9082 2717 -9048
rect 2761 -9082 2777 -9048
rect 2879 -9082 2895 -9048
rect 2939 -9082 2955 -9048
rect 3057 -9082 3073 -9048
rect 3117 -9082 3133 -9048
rect 3235 -9082 3251 -9048
rect 3295 -9082 3311 -9048
rect 3413 -9082 3429 -9048
rect 3473 -9082 3489 -9048
rect 3591 -9082 3607 -9048
rect 3651 -9082 3667 -9048
rect 3769 -9082 3785 -9048
rect 3829 -9082 3845 -9048
rect 3947 -9082 3963 -9048
rect 4007 -9082 4023 -9048
rect -4026 -9246 -3992 -9230
rect -2173 -9132 -2139 -9116
rect -5560 -9314 -5544 -9280
rect -5500 -9314 -5484 -9280
rect -5382 -9314 -5366 -9280
rect -5322 -9314 -5306 -9280
rect -5204 -9314 -5188 -9280
rect -5144 -9314 -5128 -9280
rect -5026 -9314 -5010 -9280
rect -4966 -9314 -4950 -9280
rect -4848 -9314 -4832 -9280
rect -4788 -9314 -4772 -9280
rect -4670 -9314 -4654 -9280
rect -4610 -9314 -4594 -9280
rect -4492 -9314 -4476 -9280
rect -4432 -9314 -4416 -9280
rect -4314 -9314 -4298 -9280
rect -4254 -9314 -4238 -9280
rect -4136 -9314 -4120 -9280
rect -4076 -9314 -4060 -9280
rect -2173 -9404 -2139 -9388
rect -1995 -9132 -1961 -9116
rect -1995 -9404 -1961 -9388
rect -1817 -9132 -1783 -9116
rect -1817 -9404 -1783 -9388
rect -1639 -9132 -1605 -9116
rect -1639 -9404 -1605 -9388
rect -1461 -9132 -1427 -9116
rect -1461 -9404 -1427 -9388
rect -1283 -9132 -1249 -9116
rect -1283 -9404 -1249 -9388
rect -1105 -9132 -1071 -9116
rect -1105 -9404 -1071 -9388
rect -927 -9132 -893 -9116
rect -927 -9404 -893 -9388
rect -749 -9132 -715 -9116
rect -749 -9404 -715 -9388
rect -571 -9132 -537 -9116
rect -571 -9404 -537 -9388
rect -393 -9132 -359 -9116
rect -393 -9404 -359 -9388
rect -215 -9132 -181 -9116
rect -215 -9404 -181 -9388
rect -37 -9132 -3 -9116
rect -37 -9404 -3 -9388
rect 141 -9132 175 -9116
rect 141 -9404 175 -9388
rect 319 -9132 353 -9116
rect 319 -9404 353 -9388
rect 497 -9132 531 -9116
rect 497 -9404 531 -9388
rect 675 -9132 709 -9116
rect 675 -9404 709 -9388
rect 853 -9132 887 -9116
rect 853 -9404 887 -9388
rect 1031 -9132 1065 -9116
rect 1031 -9404 1065 -9388
rect 1209 -9132 1243 -9116
rect 1209 -9404 1243 -9388
rect 1387 -9132 1421 -9116
rect 1387 -9404 1421 -9388
rect 1565 -9132 1599 -9116
rect 1565 -9404 1599 -9388
rect 1743 -9132 1777 -9116
rect 1743 -9404 1777 -9388
rect 1921 -9132 1955 -9116
rect 1921 -9404 1955 -9388
rect 2099 -9132 2133 -9116
rect 2099 -9404 2133 -9388
rect 2277 -9132 2311 -9116
rect 2277 -9404 2311 -9388
rect 2455 -9132 2489 -9116
rect 2455 -9404 2489 -9388
rect 2633 -9132 2667 -9116
rect 2633 -9404 2667 -9388
rect 2811 -9132 2845 -9116
rect 2811 -9404 2845 -9388
rect 2989 -9132 3023 -9116
rect 2989 -9404 3023 -9388
rect 3167 -9132 3201 -9116
rect 3167 -9404 3201 -9388
rect 3345 -9132 3379 -9116
rect 3345 -9404 3379 -9388
rect 3523 -9132 3557 -9116
rect 3523 -9404 3557 -9388
rect 3701 -9132 3735 -9116
rect 3701 -9404 3735 -9388
rect 3879 -9132 3913 -9116
rect 3879 -9404 3913 -9388
rect 4057 -9132 4091 -9116
rect 6512 -9166 6546 -9150
rect 6690 -8894 6724 -8878
rect 6690 -9166 6724 -9150
rect 6868 -8894 6902 -8878
rect 6868 -9166 6902 -9150
rect 7046 -8894 7080 -8878
rect 7046 -9166 7080 -9150
rect 7224 -8894 7258 -8878
rect 7224 -9166 7258 -9150
rect 7402 -8894 7436 -8878
rect 7402 -9166 7436 -9150
rect 7580 -8894 7614 -8878
rect 7580 -9166 7614 -9150
rect 7758 -8894 7792 -8878
rect 7758 -9166 7792 -9150
rect 7936 -8894 7970 -8878
rect 7936 -9166 7970 -9150
rect 8114 -8894 8148 -8878
rect 8114 -9166 8148 -9150
rect 8292 -8894 8326 -8878
rect 8292 -9166 8326 -9150
rect 8470 -8894 8504 -8878
rect 8470 -9166 8504 -9150
rect 8648 -8894 8682 -8878
rect 8648 -9166 8682 -9150
rect 8826 -8894 8860 -8878
rect 8826 -9166 8860 -9150
rect 9004 -8894 9038 -8878
rect 9004 -9166 9038 -9150
rect 9182 -8894 9216 -8878
rect 9182 -9166 9216 -9150
rect 9360 -8894 9394 -8878
rect 9360 -9166 9394 -9150
rect 10772 -8924 10806 -8908
rect 10772 -9196 10806 -9180
rect 10950 -8924 10984 -8908
rect 10950 -9196 10984 -9180
rect 11064 -8924 11098 -8908
rect 11064 -9196 11098 -9180
rect 11242 -8924 11276 -8908
rect 11242 -9196 11276 -9180
rect 11356 -8924 11390 -8908
rect 11356 -9196 11390 -9180
rect 11534 -8924 11568 -8908
rect 11534 -9196 11568 -9180
rect 11648 -8924 11682 -8908
rect 11648 -9196 11682 -9180
rect 11826 -8924 11860 -8908
rect 11826 -9196 11860 -9180
rect 11940 -8924 11974 -8908
rect 11940 -9196 11974 -9180
rect 12118 -8924 12152 -8908
rect 12118 -9196 12152 -9180
rect 12232 -8924 12266 -8908
rect 12232 -9196 12266 -9180
rect 12410 -8924 12444 -8908
rect 12410 -9196 12444 -9180
rect 12524 -8924 12558 -8908
rect 12524 -9196 12558 -9180
rect 12702 -8924 12736 -8908
rect 12702 -9196 12736 -9180
rect 6580 -9234 6596 -9200
rect 6640 -9234 6656 -9200
rect 6758 -9234 6774 -9200
rect 6818 -9234 6834 -9200
rect 6936 -9234 6952 -9200
rect 6996 -9234 7012 -9200
rect 7114 -9234 7130 -9200
rect 7174 -9234 7190 -9200
rect 7292 -9234 7308 -9200
rect 7352 -9234 7368 -9200
rect 7470 -9234 7486 -9200
rect 7530 -9234 7546 -9200
rect 7648 -9234 7664 -9200
rect 7708 -9234 7724 -9200
rect 7826 -9234 7842 -9200
rect 7886 -9234 7902 -9200
rect 8004 -9234 8020 -9200
rect 8064 -9234 8080 -9200
rect 8182 -9234 8198 -9200
rect 8242 -9234 8258 -9200
rect 8360 -9234 8376 -9200
rect 8420 -9234 8436 -9200
rect 8538 -9234 8554 -9200
rect 8598 -9234 8614 -9200
rect 8716 -9234 8732 -9200
rect 8776 -9234 8792 -9200
rect 8894 -9234 8910 -9200
rect 8954 -9234 8970 -9200
rect 9072 -9234 9088 -9200
rect 9132 -9234 9148 -9200
rect 9250 -9234 9266 -9200
rect 9310 -9234 9326 -9200
rect 10840 -9264 10856 -9230
rect 10900 -9264 10916 -9230
rect 11132 -9264 11148 -9230
rect 11192 -9264 11208 -9230
rect 11424 -9264 11440 -9230
rect 11484 -9264 11500 -9230
rect 11716 -9264 11732 -9230
rect 11776 -9264 11792 -9230
rect 12008 -9264 12024 -9230
rect 12068 -9264 12084 -9230
rect 12300 -9264 12316 -9230
rect 12360 -9264 12376 -9230
rect 12592 -9264 12608 -9230
rect 12652 -9264 12668 -9230
rect 4057 -9404 4091 -9388
rect -5560 -9474 -5544 -9440
rect -5500 -9474 -5484 -9440
rect -5382 -9474 -5366 -9440
rect -5322 -9474 -5306 -9440
rect -5204 -9474 -5188 -9440
rect -5144 -9474 -5128 -9440
rect -5026 -9474 -5010 -9440
rect -4966 -9474 -4950 -9440
rect -4848 -9474 -4832 -9440
rect -4788 -9474 -4772 -9440
rect -4670 -9474 -4654 -9440
rect -4610 -9474 -4594 -9440
rect -4492 -9474 -4476 -9440
rect -4432 -9474 -4416 -9440
rect -4314 -9474 -4298 -9440
rect -4254 -9474 -4238 -9440
rect -4136 -9474 -4120 -9440
rect -4076 -9474 -4060 -9440
rect -2105 -9472 -2089 -9438
rect -2045 -9472 -2029 -9438
rect -1927 -9472 -1911 -9438
rect -1867 -9472 -1851 -9438
rect -1749 -9472 -1733 -9438
rect -1689 -9472 -1673 -9438
rect -1571 -9472 -1555 -9438
rect -1511 -9472 -1495 -9438
rect -1393 -9472 -1377 -9438
rect -1333 -9472 -1317 -9438
rect -1215 -9472 -1199 -9438
rect -1155 -9472 -1139 -9438
rect -1037 -9472 -1021 -9438
rect -977 -9472 -961 -9438
rect -859 -9472 -843 -9438
rect -799 -9472 -783 -9438
rect -681 -9472 -665 -9438
rect -621 -9472 -605 -9438
rect -503 -9472 -487 -9438
rect -443 -9472 -427 -9438
rect -325 -9472 -309 -9438
rect -265 -9472 -249 -9438
rect -147 -9472 -131 -9438
rect -87 -9472 -71 -9438
rect 31 -9472 47 -9438
rect 91 -9472 107 -9438
rect 209 -9472 225 -9438
rect 269 -9472 285 -9438
rect 387 -9472 403 -9438
rect 447 -9472 463 -9438
rect 565 -9472 581 -9438
rect 625 -9472 641 -9438
rect 743 -9472 759 -9438
rect 803 -9472 819 -9438
rect 921 -9472 937 -9438
rect 981 -9472 997 -9438
rect 1099 -9472 1115 -9438
rect 1159 -9472 1175 -9438
rect 1277 -9472 1293 -9438
rect 1337 -9472 1353 -9438
rect 1455 -9472 1471 -9438
rect 1515 -9472 1531 -9438
rect 1633 -9472 1649 -9438
rect 1693 -9472 1709 -9438
rect 1811 -9472 1827 -9438
rect 1871 -9472 1887 -9438
rect 1989 -9472 2005 -9438
rect 2049 -9472 2065 -9438
rect 2167 -9472 2183 -9438
rect 2227 -9472 2243 -9438
rect 2345 -9472 2361 -9438
rect 2405 -9472 2421 -9438
rect 2523 -9472 2539 -9438
rect 2583 -9472 2599 -9438
rect 2701 -9472 2717 -9438
rect 2761 -9472 2777 -9438
rect 2879 -9472 2895 -9438
rect 2939 -9472 2955 -9438
rect 3057 -9472 3073 -9438
rect 3117 -9472 3133 -9438
rect 3235 -9472 3251 -9438
rect 3295 -9472 3311 -9438
rect 3413 -9472 3429 -9438
rect 3473 -9472 3489 -9438
rect 3591 -9472 3607 -9438
rect 3651 -9472 3667 -9438
rect 3769 -9472 3785 -9438
rect 3829 -9472 3845 -9438
rect 3947 -9472 3963 -9438
rect 4007 -9472 4023 -9438
rect -5628 -9524 -5594 -9508
rect -5628 -9796 -5594 -9780
rect -5450 -9524 -5416 -9508
rect -5450 -9796 -5416 -9780
rect -5272 -9524 -5238 -9508
rect -5272 -9796 -5238 -9780
rect -5094 -9524 -5060 -9508
rect -5094 -9796 -5060 -9780
rect -4916 -9524 -4882 -9508
rect -4916 -9796 -4882 -9780
rect -4738 -9524 -4704 -9508
rect -4738 -9796 -4704 -9780
rect -4560 -9524 -4526 -9508
rect -4560 -9796 -4526 -9780
rect -4382 -9524 -4348 -9508
rect -4382 -9796 -4348 -9780
rect -4204 -9524 -4170 -9508
rect -4204 -9796 -4170 -9780
rect -4026 -9524 -3992 -9508
rect 10840 -9644 10856 -9610
rect 10900 -9644 10916 -9610
rect 11132 -9644 11148 -9610
rect 11192 -9644 11208 -9610
rect 11424 -9644 11440 -9610
rect 11484 -9644 11500 -9610
rect 11716 -9644 11732 -9610
rect 11776 -9644 11792 -9610
rect 12008 -9644 12024 -9610
rect 12068 -9644 12084 -9610
rect 12300 -9644 12316 -9610
rect 12360 -9644 12376 -9610
rect 12592 -9644 12608 -9610
rect 12652 -9644 12668 -9610
rect 10772 -9694 10806 -9678
rect 6580 -9744 6596 -9710
rect 6640 -9744 6656 -9710
rect 6758 -9744 6774 -9710
rect 6818 -9744 6834 -9710
rect 6936 -9744 6952 -9710
rect 6996 -9744 7012 -9710
rect 7114 -9744 7130 -9710
rect 7174 -9744 7190 -9710
rect 7292 -9744 7308 -9710
rect 7352 -9744 7368 -9710
rect 7470 -9744 7486 -9710
rect 7530 -9744 7546 -9710
rect 7648 -9744 7664 -9710
rect 7708 -9744 7724 -9710
rect 7826 -9744 7842 -9710
rect 7886 -9744 7902 -9710
rect 8004 -9744 8020 -9710
rect 8064 -9744 8080 -9710
rect 8182 -9744 8198 -9710
rect 8242 -9744 8258 -9710
rect 8360 -9744 8376 -9710
rect 8420 -9744 8436 -9710
rect 8538 -9744 8554 -9710
rect 8598 -9744 8614 -9710
rect 8716 -9744 8732 -9710
rect 8776 -9744 8792 -9710
rect 8894 -9744 8910 -9710
rect 8954 -9744 8970 -9710
rect 9072 -9744 9088 -9710
rect 9132 -9744 9148 -9710
rect 9250 -9744 9266 -9710
rect 9310 -9744 9326 -9710
rect -4026 -9796 -3992 -9780
rect 6512 -9794 6546 -9778
rect -5560 -9864 -5544 -9830
rect -5500 -9864 -5484 -9830
rect -5382 -9864 -5366 -9830
rect -5322 -9864 -5306 -9830
rect -5204 -9864 -5188 -9830
rect -5144 -9864 -5128 -9830
rect -5026 -9864 -5010 -9830
rect -4966 -9864 -4950 -9830
rect -4848 -9864 -4832 -9830
rect -4788 -9864 -4772 -9830
rect -4670 -9864 -4654 -9830
rect -4610 -9864 -4594 -9830
rect -4492 -9864 -4476 -9830
rect -4432 -9864 -4416 -9830
rect -4314 -9864 -4298 -9830
rect -4254 -9864 -4238 -9830
rect -4136 -9864 -4120 -9830
rect -4076 -9864 -4060 -9830
rect -5560 -10024 -5544 -9990
rect -5500 -10024 -5484 -9990
rect -5382 -10024 -5366 -9990
rect -5322 -10024 -5306 -9990
rect -5204 -10024 -5188 -9990
rect -5144 -10024 -5128 -9990
rect -5026 -10024 -5010 -9990
rect -4966 -10024 -4950 -9990
rect -4848 -10024 -4832 -9990
rect -4788 -10024 -4772 -9990
rect -4670 -10024 -4654 -9990
rect -4610 -10024 -4594 -9990
rect -4492 -10024 -4476 -9990
rect -4432 -10024 -4416 -9990
rect -4314 -10024 -4298 -9990
rect -4254 -10024 -4238 -9990
rect -4136 -10024 -4120 -9990
rect -4076 -10024 -4060 -9990
rect -5628 -10074 -5594 -10058
rect -5628 -10346 -5594 -10330
rect -5450 -10074 -5416 -10058
rect -5450 -10346 -5416 -10330
rect -5272 -10074 -5238 -10058
rect -5272 -10346 -5238 -10330
rect -5094 -10074 -5060 -10058
rect -5094 -10346 -5060 -10330
rect -4916 -10074 -4882 -10058
rect -4916 -10346 -4882 -10330
rect -4738 -10074 -4704 -10058
rect -4738 -10346 -4704 -10330
rect -4560 -10074 -4526 -10058
rect -4560 -10346 -4526 -10330
rect -4382 -10074 -4348 -10058
rect -4382 -10346 -4348 -10330
rect -4204 -10074 -4170 -10058
rect -4204 -10346 -4170 -10330
rect -4026 -10074 -3992 -10058
rect -2105 -10082 -2089 -10048
rect -2045 -10082 -2029 -10048
rect -1927 -10082 -1911 -10048
rect -1867 -10082 -1851 -10048
rect -1749 -10082 -1733 -10048
rect -1689 -10082 -1673 -10048
rect -1571 -10082 -1555 -10048
rect -1511 -10082 -1495 -10048
rect -1393 -10082 -1377 -10048
rect -1333 -10082 -1317 -10048
rect -1215 -10082 -1199 -10048
rect -1155 -10082 -1139 -10048
rect -1037 -10082 -1021 -10048
rect -977 -10082 -961 -10048
rect -859 -10082 -843 -10048
rect -799 -10082 -783 -10048
rect -681 -10082 -665 -10048
rect -621 -10082 -605 -10048
rect -503 -10082 -487 -10048
rect -443 -10082 -427 -10048
rect -325 -10082 -309 -10048
rect -265 -10082 -249 -10048
rect -147 -10082 -131 -10048
rect -87 -10082 -71 -10048
rect 31 -10082 47 -10048
rect 91 -10082 107 -10048
rect 209 -10082 225 -10048
rect 269 -10082 285 -10048
rect 387 -10082 403 -10048
rect 447 -10082 463 -10048
rect 565 -10082 581 -10048
rect 625 -10082 641 -10048
rect 743 -10082 759 -10048
rect 803 -10082 819 -10048
rect 921 -10082 937 -10048
rect 981 -10082 997 -10048
rect 1099 -10082 1115 -10048
rect 1159 -10082 1175 -10048
rect 1277 -10082 1293 -10048
rect 1337 -10082 1353 -10048
rect 1455 -10082 1471 -10048
rect 1515 -10082 1531 -10048
rect 1633 -10082 1649 -10048
rect 1693 -10082 1709 -10048
rect 1811 -10082 1827 -10048
rect 1871 -10082 1887 -10048
rect 1989 -10082 2005 -10048
rect 2049 -10082 2065 -10048
rect 2167 -10082 2183 -10048
rect 2227 -10082 2243 -10048
rect 2345 -10082 2361 -10048
rect 2405 -10082 2421 -10048
rect 2523 -10082 2539 -10048
rect 2583 -10082 2599 -10048
rect 2701 -10082 2717 -10048
rect 2761 -10082 2777 -10048
rect 2879 -10082 2895 -10048
rect 2939 -10082 2955 -10048
rect 3057 -10082 3073 -10048
rect 3117 -10082 3133 -10048
rect 3235 -10082 3251 -10048
rect 3295 -10082 3311 -10048
rect 3413 -10082 3429 -10048
rect 3473 -10082 3489 -10048
rect 3591 -10082 3607 -10048
rect 3651 -10082 3667 -10048
rect 3769 -10082 3785 -10048
rect 3829 -10082 3845 -10048
rect 3947 -10082 3963 -10048
rect 4007 -10082 4023 -10048
rect 6512 -10066 6546 -10050
rect 6690 -9794 6724 -9778
rect 6690 -10066 6724 -10050
rect 6868 -9794 6902 -9778
rect 6868 -10066 6902 -10050
rect 7046 -9794 7080 -9778
rect 7046 -10066 7080 -10050
rect 7224 -9794 7258 -9778
rect 7224 -10066 7258 -10050
rect 7402 -9794 7436 -9778
rect 7402 -10066 7436 -10050
rect 7580 -9794 7614 -9778
rect 7580 -10066 7614 -10050
rect 7758 -9794 7792 -9778
rect 7758 -10066 7792 -10050
rect 7936 -9794 7970 -9778
rect 7936 -10066 7970 -10050
rect 8114 -9794 8148 -9778
rect 8114 -10066 8148 -10050
rect 8292 -9794 8326 -9778
rect 8292 -10066 8326 -10050
rect 8470 -9794 8504 -9778
rect 8470 -10066 8504 -10050
rect 8648 -9794 8682 -9778
rect 8648 -10066 8682 -10050
rect 8826 -9794 8860 -9778
rect 8826 -10066 8860 -10050
rect 9004 -9794 9038 -9778
rect 9004 -10066 9038 -10050
rect 9182 -9794 9216 -9778
rect 9182 -10066 9216 -10050
rect 9360 -9794 9394 -9778
rect 10772 -9966 10806 -9950
rect 10950 -9694 10984 -9678
rect 10950 -9966 10984 -9950
rect 11064 -9694 11098 -9678
rect 11064 -9966 11098 -9950
rect 11242 -9694 11276 -9678
rect 11242 -9966 11276 -9950
rect 11356 -9694 11390 -9678
rect 11356 -9966 11390 -9950
rect 11534 -9694 11568 -9678
rect 11534 -9966 11568 -9950
rect 11648 -9694 11682 -9678
rect 11648 -9966 11682 -9950
rect 11826 -9694 11860 -9678
rect 11826 -9966 11860 -9950
rect 11940 -9694 11974 -9678
rect 11940 -9966 11974 -9950
rect 12118 -9694 12152 -9678
rect 12118 -9966 12152 -9950
rect 12232 -9694 12266 -9678
rect 12232 -9966 12266 -9950
rect 12410 -9694 12444 -9678
rect 12410 -9966 12444 -9950
rect 12524 -9694 12558 -9678
rect 12524 -9966 12558 -9950
rect 12702 -9694 12736 -9678
rect 12702 -9966 12736 -9950
rect 10840 -10034 10856 -10000
rect 10900 -10034 10916 -10000
rect 11132 -10034 11148 -10000
rect 11192 -10034 11208 -10000
rect 11424 -10034 11440 -10000
rect 11484 -10034 11500 -10000
rect 11716 -10034 11732 -10000
rect 11776 -10034 11792 -10000
rect 12008 -10034 12024 -10000
rect 12068 -10034 12084 -10000
rect 12300 -10034 12316 -10000
rect 12360 -10034 12376 -10000
rect 12592 -10034 12608 -10000
rect 12652 -10034 12668 -10000
rect 9360 -10066 9394 -10050
rect -4026 -10346 -3992 -10330
rect -2173 -10132 -2139 -10116
rect -5560 -10414 -5544 -10380
rect -5500 -10414 -5484 -10380
rect -5382 -10414 -5366 -10380
rect -5322 -10414 -5306 -10380
rect -5204 -10414 -5188 -10380
rect -5144 -10414 -5128 -10380
rect -5026 -10414 -5010 -10380
rect -4966 -10414 -4950 -10380
rect -4848 -10414 -4832 -10380
rect -4788 -10414 -4772 -10380
rect -4670 -10414 -4654 -10380
rect -4610 -10414 -4594 -10380
rect -4492 -10414 -4476 -10380
rect -4432 -10414 -4416 -10380
rect -4314 -10414 -4298 -10380
rect -4254 -10414 -4238 -10380
rect -4136 -10414 -4120 -10380
rect -4076 -10414 -4060 -10380
rect -2173 -10404 -2139 -10388
rect -1995 -10132 -1961 -10116
rect -1995 -10404 -1961 -10388
rect -1817 -10132 -1783 -10116
rect -1817 -10404 -1783 -10388
rect -1639 -10132 -1605 -10116
rect -1639 -10404 -1605 -10388
rect -1461 -10132 -1427 -10116
rect -1461 -10404 -1427 -10388
rect -1283 -10132 -1249 -10116
rect -1283 -10404 -1249 -10388
rect -1105 -10132 -1071 -10116
rect -1105 -10404 -1071 -10388
rect -927 -10132 -893 -10116
rect -927 -10404 -893 -10388
rect -749 -10132 -715 -10116
rect -749 -10404 -715 -10388
rect -571 -10132 -537 -10116
rect -571 -10404 -537 -10388
rect -393 -10132 -359 -10116
rect -393 -10404 -359 -10388
rect -215 -10132 -181 -10116
rect -215 -10404 -181 -10388
rect -37 -10132 -3 -10116
rect -37 -10404 -3 -10388
rect 141 -10132 175 -10116
rect 141 -10404 175 -10388
rect 319 -10132 353 -10116
rect 319 -10404 353 -10388
rect 497 -10132 531 -10116
rect 497 -10404 531 -10388
rect 675 -10132 709 -10116
rect 675 -10404 709 -10388
rect 853 -10132 887 -10116
rect 853 -10404 887 -10388
rect 1031 -10132 1065 -10116
rect 1031 -10404 1065 -10388
rect 1209 -10132 1243 -10116
rect 1209 -10404 1243 -10388
rect 1387 -10132 1421 -10116
rect 1387 -10404 1421 -10388
rect 1565 -10132 1599 -10116
rect 1565 -10404 1599 -10388
rect 1743 -10132 1777 -10116
rect 1743 -10404 1777 -10388
rect 1921 -10132 1955 -10116
rect 1921 -10404 1955 -10388
rect 2099 -10132 2133 -10116
rect 2099 -10404 2133 -10388
rect 2277 -10132 2311 -10116
rect 2277 -10404 2311 -10388
rect 2455 -10132 2489 -10116
rect 2455 -10404 2489 -10388
rect 2633 -10132 2667 -10116
rect 2633 -10404 2667 -10388
rect 2811 -10132 2845 -10116
rect 2811 -10404 2845 -10388
rect 2989 -10132 3023 -10116
rect 2989 -10404 3023 -10388
rect 3167 -10132 3201 -10116
rect 3167 -10404 3201 -10388
rect 3345 -10132 3379 -10116
rect 3345 -10404 3379 -10388
rect 3523 -10132 3557 -10116
rect 3523 -10404 3557 -10388
rect 3701 -10132 3735 -10116
rect 3701 -10404 3735 -10388
rect 3879 -10132 3913 -10116
rect 3879 -10404 3913 -10388
rect 4057 -10132 4091 -10116
rect 6580 -10134 6596 -10100
rect 6640 -10134 6656 -10100
rect 6758 -10134 6774 -10100
rect 6818 -10134 6834 -10100
rect 6936 -10134 6952 -10100
rect 6996 -10134 7012 -10100
rect 7114 -10134 7130 -10100
rect 7174 -10134 7190 -10100
rect 7292 -10134 7308 -10100
rect 7352 -10134 7368 -10100
rect 7470 -10134 7486 -10100
rect 7530 -10134 7546 -10100
rect 7648 -10134 7664 -10100
rect 7708 -10134 7724 -10100
rect 7826 -10134 7842 -10100
rect 7886 -10134 7902 -10100
rect 8004 -10134 8020 -10100
rect 8064 -10134 8080 -10100
rect 8182 -10134 8198 -10100
rect 8242 -10134 8258 -10100
rect 8360 -10134 8376 -10100
rect 8420 -10134 8436 -10100
rect 8538 -10134 8554 -10100
rect 8598 -10134 8614 -10100
rect 8716 -10134 8732 -10100
rect 8776 -10134 8792 -10100
rect 8894 -10134 8910 -10100
rect 8954 -10134 8970 -10100
rect 9072 -10134 9088 -10100
rect 9132 -10134 9148 -10100
rect 9250 -10134 9266 -10100
rect 9310 -10134 9326 -10100
rect 4057 -10404 4091 -10388
rect 10840 -10414 10856 -10380
rect 10900 -10414 10916 -10380
rect 11132 -10414 11148 -10380
rect 11192 -10414 11208 -10380
rect 11424 -10414 11440 -10380
rect 11484 -10414 11500 -10380
rect 11716 -10414 11732 -10380
rect 11776 -10414 11792 -10380
rect 12008 -10414 12024 -10380
rect 12068 -10414 12084 -10380
rect 12300 -10414 12316 -10380
rect 12360 -10414 12376 -10380
rect 12592 -10414 12608 -10380
rect 12652 -10414 12668 -10380
rect -2105 -10472 -2089 -10438
rect -2045 -10472 -2029 -10438
rect -1927 -10472 -1911 -10438
rect -1867 -10472 -1851 -10438
rect -1749 -10472 -1733 -10438
rect -1689 -10472 -1673 -10438
rect -1571 -10472 -1555 -10438
rect -1511 -10472 -1495 -10438
rect -1393 -10472 -1377 -10438
rect -1333 -10472 -1317 -10438
rect -1215 -10472 -1199 -10438
rect -1155 -10472 -1139 -10438
rect -1037 -10472 -1021 -10438
rect -977 -10472 -961 -10438
rect -859 -10472 -843 -10438
rect -799 -10472 -783 -10438
rect -681 -10472 -665 -10438
rect -621 -10472 -605 -10438
rect -503 -10472 -487 -10438
rect -443 -10472 -427 -10438
rect -325 -10472 -309 -10438
rect -265 -10472 -249 -10438
rect -147 -10472 -131 -10438
rect -87 -10472 -71 -10438
rect 31 -10472 47 -10438
rect 91 -10472 107 -10438
rect 209 -10472 225 -10438
rect 269 -10472 285 -10438
rect 387 -10472 403 -10438
rect 447 -10472 463 -10438
rect 565 -10472 581 -10438
rect 625 -10472 641 -10438
rect 743 -10472 759 -10438
rect 803 -10472 819 -10438
rect 921 -10472 937 -10438
rect 981 -10472 997 -10438
rect 1099 -10472 1115 -10438
rect 1159 -10472 1175 -10438
rect 1277 -10472 1293 -10438
rect 1337 -10472 1353 -10438
rect 1455 -10472 1471 -10438
rect 1515 -10472 1531 -10438
rect 1633 -10472 1649 -10438
rect 1693 -10472 1709 -10438
rect 1811 -10472 1827 -10438
rect 1871 -10472 1887 -10438
rect 1989 -10472 2005 -10438
rect 2049 -10472 2065 -10438
rect 2167 -10472 2183 -10438
rect 2227 -10472 2243 -10438
rect 2345 -10472 2361 -10438
rect 2405 -10472 2421 -10438
rect 2523 -10472 2539 -10438
rect 2583 -10472 2599 -10438
rect 2701 -10472 2717 -10438
rect 2761 -10472 2777 -10438
rect 2879 -10472 2895 -10438
rect 2939 -10472 2955 -10438
rect 3057 -10472 3073 -10438
rect 3117 -10472 3133 -10438
rect 3235 -10472 3251 -10438
rect 3295 -10472 3311 -10438
rect 3413 -10472 3429 -10438
rect 3473 -10472 3489 -10438
rect 3591 -10472 3607 -10438
rect 3651 -10472 3667 -10438
rect 3769 -10472 3785 -10438
rect 3829 -10472 3845 -10438
rect 3947 -10472 3963 -10438
rect 4007 -10472 4023 -10438
rect 10772 -10464 10806 -10448
rect -5560 -10574 -5544 -10540
rect -5500 -10574 -5484 -10540
rect -5382 -10574 -5366 -10540
rect -5322 -10574 -5306 -10540
rect -5204 -10574 -5188 -10540
rect -5144 -10574 -5128 -10540
rect -5026 -10574 -5010 -10540
rect -4966 -10574 -4950 -10540
rect -4848 -10574 -4832 -10540
rect -4788 -10574 -4772 -10540
rect -4670 -10574 -4654 -10540
rect -4610 -10574 -4594 -10540
rect -4492 -10574 -4476 -10540
rect -4432 -10574 -4416 -10540
rect -4314 -10574 -4298 -10540
rect -4254 -10574 -4238 -10540
rect -4136 -10574 -4120 -10540
rect -4076 -10574 -4060 -10540
rect -5628 -10624 -5594 -10608
rect -5628 -10896 -5594 -10880
rect -5450 -10624 -5416 -10608
rect -5450 -10896 -5416 -10880
rect -5272 -10624 -5238 -10608
rect -5272 -10896 -5238 -10880
rect -5094 -10624 -5060 -10608
rect -5094 -10896 -5060 -10880
rect -4916 -10624 -4882 -10608
rect -4916 -10896 -4882 -10880
rect -4738 -10624 -4704 -10608
rect -4738 -10896 -4704 -10880
rect -4560 -10624 -4526 -10608
rect -4560 -10896 -4526 -10880
rect -4382 -10624 -4348 -10608
rect -4382 -10896 -4348 -10880
rect -4204 -10624 -4170 -10608
rect -4204 -10896 -4170 -10880
rect -4026 -10624 -3992 -10608
rect 6580 -10644 6596 -10610
rect 6640 -10644 6656 -10610
rect 6758 -10644 6774 -10610
rect 6818 -10644 6834 -10610
rect 6936 -10644 6952 -10610
rect 6996 -10644 7012 -10610
rect 7114 -10644 7130 -10610
rect 7174 -10644 7190 -10610
rect 7292 -10644 7308 -10610
rect 7352 -10644 7368 -10610
rect 7470 -10644 7486 -10610
rect 7530 -10644 7546 -10610
rect 7648 -10644 7664 -10610
rect 7708 -10644 7724 -10610
rect 7826 -10644 7842 -10610
rect 7886 -10644 7902 -10610
rect 8004 -10644 8020 -10610
rect 8064 -10644 8080 -10610
rect 8182 -10644 8198 -10610
rect 8242 -10644 8258 -10610
rect 8360 -10644 8376 -10610
rect 8420 -10644 8436 -10610
rect 8538 -10644 8554 -10610
rect 8598 -10644 8614 -10610
rect 8716 -10644 8732 -10610
rect 8776 -10644 8792 -10610
rect 8894 -10644 8910 -10610
rect 8954 -10644 8970 -10610
rect 9072 -10644 9088 -10610
rect 9132 -10644 9148 -10610
rect 9250 -10644 9266 -10610
rect 9310 -10644 9326 -10610
rect -4026 -10896 -3992 -10880
rect 6512 -10694 6546 -10678
rect -5560 -10964 -5544 -10930
rect -5500 -10964 -5484 -10930
rect -5382 -10964 -5366 -10930
rect -5322 -10964 -5306 -10930
rect -5204 -10964 -5188 -10930
rect -5144 -10964 -5128 -10930
rect -5026 -10964 -5010 -10930
rect -4966 -10964 -4950 -10930
rect -4848 -10964 -4832 -10930
rect -4788 -10964 -4772 -10930
rect -4670 -10964 -4654 -10930
rect -4610 -10964 -4594 -10930
rect -4492 -10964 -4476 -10930
rect -4432 -10964 -4416 -10930
rect -4314 -10964 -4298 -10930
rect -4254 -10964 -4238 -10930
rect -4136 -10964 -4120 -10930
rect -4076 -10964 -4060 -10930
rect 6512 -10966 6546 -10950
rect 6690 -10694 6724 -10678
rect 6690 -10966 6724 -10950
rect 6868 -10694 6902 -10678
rect 6868 -10966 6902 -10950
rect 7046 -10694 7080 -10678
rect 7046 -10966 7080 -10950
rect 7224 -10694 7258 -10678
rect 7224 -10966 7258 -10950
rect 7402 -10694 7436 -10678
rect 7402 -10966 7436 -10950
rect 7580 -10694 7614 -10678
rect 7580 -10966 7614 -10950
rect 7758 -10694 7792 -10678
rect 7758 -10966 7792 -10950
rect 7936 -10694 7970 -10678
rect 7936 -10966 7970 -10950
rect 8114 -10694 8148 -10678
rect 8114 -10966 8148 -10950
rect 8292 -10694 8326 -10678
rect 8292 -10966 8326 -10950
rect 8470 -10694 8504 -10678
rect 8470 -10966 8504 -10950
rect 8648 -10694 8682 -10678
rect 8648 -10966 8682 -10950
rect 8826 -10694 8860 -10678
rect 8826 -10966 8860 -10950
rect 9004 -10694 9038 -10678
rect 9004 -10966 9038 -10950
rect 9182 -10694 9216 -10678
rect 9182 -10966 9216 -10950
rect 9360 -10694 9394 -10678
rect 10772 -10736 10806 -10720
rect 10950 -10464 10984 -10448
rect 10950 -10736 10984 -10720
rect 11064 -10464 11098 -10448
rect 11064 -10736 11098 -10720
rect 11242 -10464 11276 -10448
rect 11242 -10736 11276 -10720
rect 11356 -10464 11390 -10448
rect 11356 -10736 11390 -10720
rect 11534 -10464 11568 -10448
rect 11534 -10736 11568 -10720
rect 11648 -10464 11682 -10448
rect 11648 -10736 11682 -10720
rect 11826 -10464 11860 -10448
rect 11826 -10736 11860 -10720
rect 11940 -10464 11974 -10448
rect 11940 -10736 11974 -10720
rect 12118 -10464 12152 -10448
rect 12118 -10736 12152 -10720
rect 12232 -10464 12266 -10448
rect 12232 -10736 12266 -10720
rect 12410 -10464 12444 -10448
rect 12410 -10736 12444 -10720
rect 12524 -10464 12558 -10448
rect 12524 -10736 12558 -10720
rect 12702 -10464 12736 -10448
rect 12702 -10736 12736 -10720
rect 10840 -10804 10856 -10770
rect 10900 -10804 10916 -10770
rect 11132 -10804 11148 -10770
rect 11192 -10804 11208 -10770
rect 11424 -10804 11440 -10770
rect 11484 -10804 11500 -10770
rect 11716 -10804 11732 -10770
rect 11776 -10804 11792 -10770
rect 12008 -10804 12024 -10770
rect 12068 -10804 12084 -10770
rect 12300 -10804 12316 -10770
rect 12360 -10804 12376 -10770
rect 12592 -10804 12608 -10770
rect 12652 -10804 12668 -10770
rect 9360 -10966 9394 -10950
rect 6580 -11034 6596 -11000
rect 6640 -11034 6656 -11000
rect 6758 -11034 6774 -11000
rect 6818 -11034 6834 -11000
rect 6936 -11034 6952 -11000
rect 6996 -11034 7012 -11000
rect 7114 -11034 7130 -11000
rect 7174 -11034 7190 -11000
rect 7292 -11034 7308 -11000
rect 7352 -11034 7368 -11000
rect 7470 -11034 7486 -11000
rect 7530 -11034 7546 -11000
rect 7648 -11034 7664 -11000
rect 7708 -11034 7724 -11000
rect 7826 -11034 7842 -11000
rect 7886 -11034 7902 -11000
rect 8004 -11034 8020 -11000
rect 8064 -11034 8080 -11000
rect 8182 -11034 8198 -11000
rect 8242 -11034 8258 -11000
rect 8360 -11034 8376 -11000
rect 8420 -11034 8436 -11000
rect 8538 -11034 8554 -11000
rect 8598 -11034 8614 -11000
rect 8716 -11034 8732 -11000
rect 8776 -11034 8792 -11000
rect 8894 -11034 8910 -11000
rect 8954 -11034 8970 -11000
rect 9072 -11034 9088 -11000
rect 9132 -11034 9148 -11000
rect 9250 -11034 9266 -11000
rect 9310 -11034 9326 -11000
rect -2105 -11082 -2089 -11048
rect -2045 -11082 -2029 -11048
rect -1927 -11082 -1911 -11048
rect -1867 -11082 -1851 -11048
rect -1749 -11082 -1733 -11048
rect -1689 -11082 -1673 -11048
rect -1571 -11082 -1555 -11048
rect -1511 -11082 -1495 -11048
rect -1393 -11082 -1377 -11048
rect -1333 -11082 -1317 -11048
rect -1215 -11082 -1199 -11048
rect -1155 -11082 -1139 -11048
rect -1037 -11082 -1021 -11048
rect -977 -11082 -961 -11048
rect -859 -11082 -843 -11048
rect -799 -11082 -783 -11048
rect -681 -11082 -665 -11048
rect -621 -11082 -605 -11048
rect -503 -11082 -487 -11048
rect -443 -11082 -427 -11048
rect -325 -11082 -309 -11048
rect -265 -11082 -249 -11048
rect -147 -11082 -131 -11048
rect -87 -11082 -71 -11048
rect 31 -11082 47 -11048
rect 91 -11082 107 -11048
rect 209 -11082 225 -11048
rect 269 -11082 285 -11048
rect 387 -11082 403 -11048
rect 447 -11082 463 -11048
rect 565 -11082 581 -11048
rect 625 -11082 641 -11048
rect 743 -11082 759 -11048
rect 803 -11082 819 -11048
rect 921 -11082 937 -11048
rect 981 -11082 997 -11048
rect 1099 -11082 1115 -11048
rect 1159 -11082 1175 -11048
rect 1277 -11082 1293 -11048
rect 1337 -11082 1353 -11048
rect 1455 -11082 1471 -11048
rect 1515 -11082 1531 -11048
rect 1633 -11082 1649 -11048
rect 1693 -11082 1709 -11048
rect 1811 -11082 1827 -11048
rect 1871 -11082 1887 -11048
rect 1989 -11082 2005 -11048
rect 2049 -11082 2065 -11048
rect 2167 -11082 2183 -11048
rect 2227 -11082 2243 -11048
rect 2345 -11082 2361 -11048
rect 2405 -11082 2421 -11048
rect 2523 -11082 2539 -11048
rect 2583 -11082 2599 -11048
rect 2701 -11082 2717 -11048
rect 2761 -11082 2777 -11048
rect 2879 -11082 2895 -11048
rect 2939 -11082 2955 -11048
rect 3057 -11082 3073 -11048
rect 3117 -11082 3133 -11048
rect 3235 -11082 3251 -11048
rect 3295 -11082 3311 -11048
rect 3413 -11082 3429 -11048
rect 3473 -11082 3489 -11048
rect 3591 -11082 3607 -11048
rect 3651 -11082 3667 -11048
rect 3769 -11082 3785 -11048
rect 3829 -11082 3845 -11048
rect 3947 -11082 3963 -11048
rect 4007 -11082 4023 -11048
rect -5560 -11124 -5544 -11090
rect -5500 -11124 -5484 -11090
rect -5382 -11124 -5366 -11090
rect -5322 -11124 -5306 -11090
rect -5204 -11124 -5188 -11090
rect -5144 -11124 -5128 -11090
rect -5026 -11124 -5010 -11090
rect -4966 -11124 -4950 -11090
rect -4848 -11124 -4832 -11090
rect -4788 -11124 -4772 -11090
rect -4670 -11124 -4654 -11090
rect -4610 -11124 -4594 -11090
rect -4492 -11124 -4476 -11090
rect -4432 -11124 -4416 -11090
rect -4314 -11124 -4298 -11090
rect -4254 -11124 -4238 -11090
rect -4136 -11124 -4120 -11090
rect -4076 -11124 -4060 -11090
rect -2173 -11132 -2139 -11116
rect -5628 -11174 -5594 -11158
rect -5628 -11446 -5594 -11430
rect -5450 -11174 -5416 -11158
rect -5450 -11446 -5416 -11430
rect -5272 -11174 -5238 -11158
rect -5272 -11446 -5238 -11430
rect -5094 -11174 -5060 -11158
rect -5094 -11446 -5060 -11430
rect -4916 -11174 -4882 -11158
rect -4916 -11446 -4882 -11430
rect -4738 -11174 -4704 -11158
rect -4738 -11446 -4704 -11430
rect -4560 -11174 -4526 -11158
rect -4560 -11446 -4526 -11430
rect -4382 -11174 -4348 -11158
rect -4382 -11446 -4348 -11430
rect -4204 -11174 -4170 -11158
rect -4204 -11446 -4170 -11430
rect -4026 -11174 -3992 -11158
rect -2173 -11404 -2139 -11388
rect -1995 -11132 -1961 -11116
rect -1995 -11404 -1961 -11388
rect -1817 -11132 -1783 -11116
rect -1817 -11404 -1783 -11388
rect -1639 -11132 -1605 -11116
rect -1639 -11404 -1605 -11388
rect -1461 -11132 -1427 -11116
rect -1461 -11404 -1427 -11388
rect -1283 -11132 -1249 -11116
rect -1283 -11404 -1249 -11388
rect -1105 -11132 -1071 -11116
rect -1105 -11404 -1071 -11388
rect -927 -11132 -893 -11116
rect -927 -11404 -893 -11388
rect -749 -11132 -715 -11116
rect -749 -11404 -715 -11388
rect -571 -11132 -537 -11116
rect -571 -11404 -537 -11388
rect -393 -11132 -359 -11116
rect -393 -11404 -359 -11388
rect -215 -11132 -181 -11116
rect -215 -11404 -181 -11388
rect -37 -11132 -3 -11116
rect -37 -11404 -3 -11388
rect 141 -11132 175 -11116
rect 141 -11404 175 -11388
rect 319 -11132 353 -11116
rect 319 -11404 353 -11388
rect 497 -11132 531 -11116
rect 497 -11404 531 -11388
rect 675 -11132 709 -11116
rect 675 -11404 709 -11388
rect 853 -11132 887 -11116
rect 853 -11404 887 -11388
rect 1031 -11132 1065 -11116
rect 1031 -11404 1065 -11388
rect 1209 -11132 1243 -11116
rect 1209 -11404 1243 -11388
rect 1387 -11132 1421 -11116
rect 1387 -11404 1421 -11388
rect 1565 -11132 1599 -11116
rect 1565 -11404 1599 -11388
rect 1743 -11132 1777 -11116
rect 1743 -11404 1777 -11388
rect 1921 -11132 1955 -11116
rect 1921 -11404 1955 -11388
rect 2099 -11132 2133 -11116
rect 2099 -11404 2133 -11388
rect 2277 -11132 2311 -11116
rect 2277 -11404 2311 -11388
rect 2455 -11132 2489 -11116
rect 2455 -11404 2489 -11388
rect 2633 -11132 2667 -11116
rect 2633 -11404 2667 -11388
rect 2811 -11132 2845 -11116
rect 2811 -11404 2845 -11388
rect 2989 -11132 3023 -11116
rect 2989 -11404 3023 -11388
rect 3167 -11132 3201 -11116
rect 3167 -11404 3201 -11388
rect 3345 -11132 3379 -11116
rect 3345 -11404 3379 -11388
rect 3523 -11132 3557 -11116
rect 3523 -11404 3557 -11388
rect 3701 -11132 3735 -11116
rect 3701 -11404 3735 -11388
rect 3879 -11132 3913 -11116
rect 3879 -11404 3913 -11388
rect 4057 -11132 4091 -11116
rect 10840 -11184 10856 -11150
rect 10900 -11184 10916 -11150
rect 11132 -11184 11148 -11150
rect 11192 -11184 11208 -11150
rect 11424 -11184 11440 -11150
rect 11484 -11184 11500 -11150
rect 11716 -11184 11732 -11150
rect 11776 -11184 11792 -11150
rect 12008 -11184 12024 -11150
rect 12068 -11184 12084 -11150
rect 12300 -11184 12316 -11150
rect 12360 -11184 12376 -11150
rect 12592 -11184 12608 -11150
rect 12652 -11184 12668 -11150
rect 4057 -11404 4091 -11388
rect 10772 -11234 10806 -11218
rect -4026 -11446 -3992 -11430
rect -2105 -11472 -2089 -11438
rect -2045 -11472 -2029 -11438
rect -1927 -11472 -1911 -11438
rect -1867 -11472 -1851 -11438
rect -1749 -11472 -1733 -11438
rect -1689 -11472 -1673 -11438
rect -1571 -11472 -1555 -11438
rect -1511 -11472 -1495 -11438
rect -1393 -11472 -1377 -11438
rect -1333 -11472 -1317 -11438
rect -1215 -11472 -1199 -11438
rect -1155 -11472 -1139 -11438
rect -1037 -11472 -1021 -11438
rect -977 -11472 -961 -11438
rect -859 -11472 -843 -11438
rect -799 -11472 -783 -11438
rect -681 -11472 -665 -11438
rect -621 -11472 -605 -11438
rect -503 -11472 -487 -11438
rect -443 -11472 -427 -11438
rect -325 -11472 -309 -11438
rect -265 -11472 -249 -11438
rect -147 -11472 -131 -11438
rect -87 -11472 -71 -11438
rect 31 -11472 47 -11438
rect 91 -11472 107 -11438
rect 209 -11472 225 -11438
rect 269 -11472 285 -11438
rect 387 -11472 403 -11438
rect 447 -11472 463 -11438
rect 565 -11472 581 -11438
rect 625 -11472 641 -11438
rect 743 -11472 759 -11438
rect 803 -11472 819 -11438
rect 921 -11472 937 -11438
rect 981 -11472 997 -11438
rect 1099 -11472 1115 -11438
rect 1159 -11472 1175 -11438
rect 1277 -11472 1293 -11438
rect 1337 -11472 1353 -11438
rect 1455 -11472 1471 -11438
rect 1515 -11472 1531 -11438
rect 1633 -11472 1649 -11438
rect 1693 -11472 1709 -11438
rect 1811 -11472 1827 -11438
rect 1871 -11472 1887 -11438
rect 1989 -11472 2005 -11438
rect 2049 -11472 2065 -11438
rect 2167 -11472 2183 -11438
rect 2227 -11472 2243 -11438
rect 2345 -11472 2361 -11438
rect 2405 -11472 2421 -11438
rect 2523 -11472 2539 -11438
rect 2583 -11472 2599 -11438
rect 2701 -11472 2717 -11438
rect 2761 -11472 2777 -11438
rect 2879 -11472 2895 -11438
rect 2939 -11472 2955 -11438
rect 3057 -11472 3073 -11438
rect 3117 -11472 3133 -11438
rect 3235 -11472 3251 -11438
rect 3295 -11472 3311 -11438
rect 3413 -11472 3429 -11438
rect 3473 -11472 3489 -11438
rect 3591 -11472 3607 -11438
rect 3651 -11472 3667 -11438
rect 3769 -11472 3785 -11438
rect 3829 -11472 3845 -11438
rect 3947 -11472 3963 -11438
rect 4007 -11472 4023 -11438
rect -5560 -11514 -5544 -11480
rect -5500 -11514 -5484 -11480
rect -5382 -11514 -5366 -11480
rect -5322 -11514 -5306 -11480
rect -5204 -11514 -5188 -11480
rect -5144 -11514 -5128 -11480
rect -5026 -11514 -5010 -11480
rect -4966 -11514 -4950 -11480
rect -4848 -11514 -4832 -11480
rect -4788 -11514 -4772 -11480
rect -4670 -11514 -4654 -11480
rect -4610 -11514 -4594 -11480
rect -4492 -11514 -4476 -11480
rect -4432 -11514 -4416 -11480
rect -4314 -11514 -4298 -11480
rect -4254 -11514 -4238 -11480
rect -4136 -11514 -4120 -11480
rect -4076 -11514 -4060 -11480
rect 10772 -11506 10806 -11490
rect 10950 -11234 10984 -11218
rect 10950 -11506 10984 -11490
rect 11064 -11234 11098 -11218
rect 11064 -11506 11098 -11490
rect 11242 -11234 11276 -11218
rect 11242 -11506 11276 -11490
rect 11356 -11234 11390 -11218
rect 11356 -11506 11390 -11490
rect 11534 -11234 11568 -11218
rect 11534 -11506 11568 -11490
rect 11648 -11234 11682 -11218
rect 11648 -11506 11682 -11490
rect 11826 -11234 11860 -11218
rect 11826 -11506 11860 -11490
rect 11940 -11234 11974 -11218
rect 11940 -11506 11974 -11490
rect 12118 -11234 12152 -11218
rect 12118 -11506 12152 -11490
rect 12232 -11234 12266 -11218
rect 12232 -11506 12266 -11490
rect 12410 -11234 12444 -11218
rect 12410 -11506 12444 -11490
rect 12524 -11234 12558 -11218
rect 12524 -11506 12558 -11490
rect 12702 -11234 12736 -11218
rect 12702 -11506 12736 -11490
rect 6580 -11544 6596 -11510
rect 6640 -11544 6656 -11510
rect 6758 -11544 6774 -11510
rect 6818 -11544 6834 -11510
rect 6936 -11544 6952 -11510
rect 6996 -11544 7012 -11510
rect 7114 -11544 7130 -11510
rect 7174 -11544 7190 -11510
rect 7292 -11544 7308 -11510
rect 7352 -11544 7368 -11510
rect 7470 -11544 7486 -11510
rect 7530 -11544 7546 -11510
rect 7648 -11544 7664 -11510
rect 7708 -11544 7724 -11510
rect 7826 -11544 7842 -11510
rect 7886 -11544 7902 -11510
rect 8004 -11544 8020 -11510
rect 8064 -11544 8080 -11510
rect 8182 -11544 8198 -11510
rect 8242 -11544 8258 -11510
rect 8360 -11544 8376 -11510
rect 8420 -11544 8436 -11510
rect 8538 -11544 8554 -11510
rect 8598 -11544 8614 -11510
rect 8716 -11544 8732 -11510
rect 8776 -11544 8792 -11510
rect 8894 -11544 8910 -11510
rect 8954 -11544 8970 -11510
rect 9072 -11544 9088 -11510
rect 9132 -11544 9148 -11510
rect 9250 -11544 9266 -11510
rect 9310 -11544 9326 -11510
rect 10840 -11574 10856 -11540
rect 10900 -11574 10916 -11540
rect 11132 -11574 11148 -11540
rect 11192 -11574 11208 -11540
rect 11424 -11574 11440 -11540
rect 11484 -11574 11500 -11540
rect 11716 -11574 11732 -11540
rect 11776 -11574 11792 -11540
rect 12008 -11574 12024 -11540
rect 12068 -11574 12084 -11540
rect 12300 -11574 12316 -11540
rect 12360 -11574 12376 -11540
rect 12592 -11574 12608 -11540
rect 12652 -11574 12668 -11540
rect 6512 -11594 6546 -11578
rect -5560 -11674 -5544 -11640
rect -5500 -11674 -5484 -11640
rect -5382 -11674 -5366 -11640
rect -5322 -11674 -5306 -11640
rect -5204 -11674 -5188 -11640
rect -5144 -11674 -5128 -11640
rect -5026 -11674 -5010 -11640
rect -4966 -11674 -4950 -11640
rect -4848 -11674 -4832 -11640
rect -4788 -11674 -4772 -11640
rect -4670 -11674 -4654 -11640
rect -4610 -11674 -4594 -11640
rect -4492 -11674 -4476 -11640
rect -4432 -11674 -4416 -11640
rect -4314 -11674 -4298 -11640
rect -4254 -11674 -4238 -11640
rect -4136 -11674 -4120 -11640
rect -4076 -11674 -4060 -11640
rect -5628 -11724 -5594 -11708
rect -5628 -11996 -5594 -11980
rect -5450 -11724 -5416 -11708
rect -5450 -11996 -5416 -11980
rect -5272 -11724 -5238 -11708
rect -5272 -11996 -5238 -11980
rect -5094 -11724 -5060 -11708
rect -5094 -11996 -5060 -11980
rect -4916 -11724 -4882 -11708
rect -4916 -11996 -4882 -11980
rect -4738 -11724 -4704 -11708
rect -4738 -11996 -4704 -11980
rect -4560 -11724 -4526 -11708
rect -4560 -11996 -4526 -11980
rect -4382 -11724 -4348 -11708
rect -4382 -11996 -4348 -11980
rect -4204 -11724 -4170 -11708
rect -4204 -11996 -4170 -11980
rect -4026 -11724 -3992 -11708
rect 6512 -11866 6546 -11850
rect 6690 -11594 6724 -11578
rect 6690 -11866 6724 -11850
rect 6868 -11594 6902 -11578
rect 6868 -11866 6902 -11850
rect 7046 -11594 7080 -11578
rect 7046 -11866 7080 -11850
rect 7224 -11594 7258 -11578
rect 7224 -11866 7258 -11850
rect 7402 -11594 7436 -11578
rect 7402 -11866 7436 -11850
rect 7580 -11594 7614 -11578
rect 7580 -11866 7614 -11850
rect 7758 -11594 7792 -11578
rect 7758 -11866 7792 -11850
rect 7936 -11594 7970 -11578
rect 7936 -11866 7970 -11850
rect 8114 -11594 8148 -11578
rect 8114 -11866 8148 -11850
rect 8292 -11594 8326 -11578
rect 8292 -11866 8326 -11850
rect 8470 -11594 8504 -11578
rect 8470 -11866 8504 -11850
rect 8648 -11594 8682 -11578
rect 8648 -11866 8682 -11850
rect 8826 -11594 8860 -11578
rect 8826 -11866 8860 -11850
rect 9004 -11594 9038 -11578
rect 9004 -11866 9038 -11850
rect 9182 -11594 9216 -11578
rect 9182 -11866 9216 -11850
rect 9360 -11594 9394 -11578
rect 9360 -11866 9394 -11850
rect 6580 -11934 6596 -11900
rect 6640 -11934 6656 -11900
rect 6758 -11934 6774 -11900
rect 6818 -11934 6834 -11900
rect 6936 -11934 6952 -11900
rect 6996 -11934 7012 -11900
rect 7114 -11934 7130 -11900
rect 7174 -11934 7190 -11900
rect 7292 -11934 7308 -11900
rect 7352 -11934 7368 -11900
rect 7470 -11934 7486 -11900
rect 7530 -11934 7546 -11900
rect 7648 -11934 7664 -11900
rect 7708 -11934 7724 -11900
rect 7826 -11934 7842 -11900
rect 7886 -11934 7902 -11900
rect 8004 -11934 8020 -11900
rect 8064 -11934 8080 -11900
rect 8182 -11934 8198 -11900
rect 8242 -11934 8258 -11900
rect 8360 -11934 8376 -11900
rect 8420 -11934 8436 -11900
rect 8538 -11934 8554 -11900
rect 8598 -11934 8614 -11900
rect 8716 -11934 8732 -11900
rect 8776 -11934 8792 -11900
rect 8894 -11934 8910 -11900
rect 8954 -11934 8970 -11900
rect 9072 -11934 9088 -11900
rect 9132 -11934 9148 -11900
rect 9250 -11934 9266 -11900
rect 9310 -11934 9326 -11900
rect -4026 -11996 -3992 -11980
rect -5560 -12064 -5544 -12030
rect -5500 -12064 -5484 -12030
rect -5382 -12064 -5366 -12030
rect -5322 -12064 -5306 -12030
rect -5204 -12064 -5188 -12030
rect -5144 -12064 -5128 -12030
rect -5026 -12064 -5010 -12030
rect -4966 -12064 -4950 -12030
rect -4848 -12064 -4832 -12030
rect -4788 -12064 -4772 -12030
rect -4670 -12064 -4654 -12030
rect -4610 -12064 -4594 -12030
rect -4492 -12064 -4476 -12030
rect -4432 -12064 -4416 -12030
rect -4314 -12064 -4298 -12030
rect -4254 -12064 -4238 -12030
rect -4136 -12064 -4120 -12030
rect -4076 -12064 -4060 -12030
rect -2105 -12082 -2089 -12048
rect -2045 -12082 -2029 -12048
rect -1927 -12082 -1911 -12048
rect -1867 -12082 -1851 -12048
rect -1749 -12082 -1733 -12048
rect -1689 -12082 -1673 -12048
rect -1571 -12082 -1555 -12048
rect -1511 -12082 -1495 -12048
rect -1393 -12082 -1377 -12048
rect -1333 -12082 -1317 -12048
rect -1215 -12082 -1199 -12048
rect -1155 -12082 -1139 -12048
rect -1037 -12082 -1021 -12048
rect -977 -12082 -961 -12048
rect -859 -12082 -843 -12048
rect -799 -12082 -783 -12048
rect -681 -12082 -665 -12048
rect -621 -12082 -605 -12048
rect -503 -12082 -487 -12048
rect -443 -12082 -427 -12048
rect -325 -12082 -309 -12048
rect -265 -12082 -249 -12048
rect -147 -12082 -131 -12048
rect -87 -12082 -71 -12048
rect 31 -12082 47 -12048
rect 91 -12082 107 -12048
rect 209 -12082 225 -12048
rect 269 -12082 285 -12048
rect 387 -12082 403 -12048
rect 447 -12082 463 -12048
rect 565 -12082 581 -12048
rect 625 -12082 641 -12048
rect 743 -12082 759 -12048
rect 803 -12082 819 -12048
rect 921 -12082 937 -12048
rect 981 -12082 997 -12048
rect 1099 -12082 1115 -12048
rect 1159 -12082 1175 -12048
rect 1277 -12082 1293 -12048
rect 1337 -12082 1353 -12048
rect 1455 -12082 1471 -12048
rect 1515 -12082 1531 -12048
rect 1633 -12082 1649 -12048
rect 1693 -12082 1709 -12048
rect 1811 -12082 1827 -12048
rect 1871 -12082 1887 -12048
rect 1989 -12082 2005 -12048
rect 2049 -12082 2065 -12048
rect 2167 -12082 2183 -12048
rect 2227 -12082 2243 -12048
rect 2345 -12082 2361 -12048
rect 2405 -12082 2421 -12048
rect 2523 -12082 2539 -12048
rect 2583 -12082 2599 -12048
rect 2701 -12082 2717 -12048
rect 2761 -12082 2777 -12048
rect 2879 -12082 2895 -12048
rect 2939 -12082 2955 -12048
rect 3057 -12082 3073 -12048
rect 3117 -12082 3133 -12048
rect 3235 -12082 3251 -12048
rect 3295 -12082 3311 -12048
rect 3413 -12082 3429 -12048
rect 3473 -12082 3489 -12048
rect 3591 -12082 3607 -12048
rect 3651 -12082 3667 -12048
rect 3769 -12082 3785 -12048
rect 3829 -12082 3845 -12048
rect 3947 -12082 3963 -12048
rect 4007 -12082 4023 -12048
rect -2173 -12132 -2139 -12116
rect -2173 -12404 -2139 -12388
rect -1995 -12132 -1961 -12116
rect -1995 -12404 -1961 -12388
rect -1817 -12132 -1783 -12116
rect -1817 -12404 -1783 -12388
rect -1639 -12132 -1605 -12116
rect -1639 -12404 -1605 -12388
rect -1461 -12132 -1427 -12116
rect -1461 -12404 -1427 -12388
rect -1283 -12132 -1249 -12116
rect -1283 -12404 -1249 -12388
rect -1105 -12132 -1071 -12116
rect -1105 -12404 -1071 -12388
rect -927 -12132 -893 -12116
rect -927 -12404 -893 -12388
rect -749 -12132 -715 -12116
rect -749 -12404 -715 -12388
rect -571 -12132 -537 -12116
rect -571 -12404 -537 -12388
rect -393 -12132 -359 -12116
rect -393 -12404 -359 -12388
rect -215 -12132 -181 -12116
rect -215 -12404 -181 -12388
rect -37 -12132 -3 -12116
rect -37 -12404 -3 -12388
rect 141 -12132 175 -12116
rect 141 -12404 175 -12388
rect 319 -12132 353 -12116
rect 319 -12404 353 -12388
rect 497 -12132 531 -12116
rect 497 -12404 531 -12388
rect 675 -12132 709 -12116
rect 675 -12404 709 -12388
rect 853 -12132 887 -12116
rect 853 -12404 887 -12388
rect 1031 -12132 1065 -12116
rect 1031 -12404 1065 -12388
rect 1209 -12132 1243 -12116
rect 1209 -12404 1243 -12388
rect 1387 -12132 1421 -12116
rect 1387 -12404 1421 -12388
rect 1565 -12132 1599 -12116
rect 1565 -12404 1599 -12388
rect 1743 -12132 1777 -12116
rect 1743 -12404 1777 -12388
rect 1921 -12132 1955 -12116
rect 1921 -12404 1955 -12388
rect 2099 -12132 2133 -12116
rect 2099 -12404 2133 -12388
rect 2277 -12132 2311 -12116
rect 2277 -12404 2311 -12388
rect 2455 -12132 2489 -12116
rect 2455 -12404 2489 -12388
rect 2633 -12132 2667 -12116
rect 2633 -12404 2667 -12388
rect 2811 -12132 2845 -12116
rect 2811 -12404 2845 -12388
rect 2989 -12132 3023 -12116
rect 2989 -12404 3023 -12388
rect 3167 -12132 3201 -12116
rect 3167 -12404 3201 -12388
rect 3345 -12132 3379 -12116
rect 3345 -12404 3379 -12388
rect 3523 -12132 3557 -12116
rect 3523 -12404 3557 -12388
rect 3701 -12132 3735 -12116
rect 3701 -12404 3735 -12388
rect 3879 -12132 3913 -12116
rect 3879 -12404 3913 -12388
rect 4057 -12132 4091 -12116
rect 4057 -12404 4091 -12388
rect -2105 -12472 -2089 -12438
rect -2045 -12472 -2029 -12438
rect -1927 -12472 -1911 -12438
rect -1867 -12472 -1851 -12438
rect -1749 -12472 -1733 -12438
rect -1689 -12472 -1673 -12438
rect -1571 -12472 -1555 -12438
rect -1511 -12472 -1495 -12438
rect -1393 -12472 -1377 -12438
rect -1333 -12472 -1317 -12438
rect -1215 -12472 -1199 -12438
rect -1155 -12472 -1139 -12438
rect -1037 -12472 -1021 -12438
rect -977 -12472 -961 -12438
rect -859 -12472 -843 -12438
rect -799 -12472 -783 -12438
rect -681 -12472 -665 -12438
rect -621 -12472 -605 -12438
rect -503 -12472 -487 -12438
rect -443 -12472 -427 -12438
rect -325 -12472 -309 -12438
rect -265 -12472 -249 -12438
rect -147 -12472 -131 -12438
rect -87 -12472 -71 -12438
rect 31 -12472 47 -12438
rect 91 -12472 107 -12438
rect 209 -12472 225 -12438
rect 269 -12472 285 -12438
rect 387 -12472 403 -12438
rect 447 -12472 463 -12438
rect 565 -12472 581 -12438
rect 625 -12472 641 -12438
rect 743 -12472 759 -12438
rect 803 -12472 819 -12438
rect 921 -12472 937 -12438
rect 981 -12472 997 -12438
rect 1099 -12472 1115 -12438
rect 1159 -12472 1175 -12438
rect 1277 -12472 1293 -12438
rect 1337 -12472 1353 -12438
rect 1455 -12472 1471 -12438
rect 1515 -12472 1531 -12438
rect 1633 -12472 1649 -12438
rect 1693 -12472 1709 -12438
rect 1811 -12472 1827 -12438
rect 1871 -12472 1887 -12438
rect 1989 -12472 2005 -12438
rect 2049 -12472 2065 -12438
rect 2167 -12472 2183 -12438
rect 2227 -12472 2243 -12438
rect 2345 -12472 2361 -12438
rect 2405 -12472 2421 -12438
rect 2523 -12472 2539 -12438
rect 2583 -12472 2599 -12438
rect 2701 -12472 2717 -12438
rect 2761 -12472 2777 -12438
rect 2879 -12472 2895 -12438
rect 2939 -12472 2955 -12438
rect 3057 -12472 3073 -12438
rect 3117 -12472 3133 -12438
rect 3235 -12472 3251 -12438
rect 3295 -12472 3311 -12438
rect 3413 -12472 3429 -12438
rect 3473 -12472 3489 -12438
rect 3591 -12472 3607 -12438
rect 3651 -12472 3667 -12438
rect 3769 -12472 3785 -12438
rect 3829 -12472 3845 -12438
rect 3947 -12472 3963 -12438
rect 4007 -12472 4023 -12438
rect -5883 -12662 -5867 -12628
rect -5833 -12662 -5817 -12628
rect -5633 -12662 -5617 -12628
rect -5583 -12662 -5567 -12628
rect -5383 -12662 -5367 -12628
rect -5333 -12662 -5317 -12628
rect -5133 -12662 -5117 -12628
rect -5083 -12662 -5067 -12628
rect -4883 -12662 -4867 -12628
rect -4833 -12662 -4817 -12628
rect -4633 -12662 -4617 -12628
rect -4583 -12662 -4567 -12628
rect -4383 -12662 -4367 -12628
rect -4333 -12662 -4317 -12628
rect -4133 -12662 -4117 -12628
rect -4083 -12662 -4067 -12628
rect -5916 -12712 -5882 -12696
rect -5916 -12944 -5882 -12928
rect -5818 -12712 -5784 -12696
rect -5818 -12944 -5784 -12928
rect -5666 -12712 -5632 -12696
rect -5666 -12944 -5632 -12928
rect -5568 -12712 -5534 -12696
rect -5568 -12944 -5534 -12928
rect -5416 -12712 -5382 -12696
rect -5416 -12944 -5382 -12928
rect -5318 -12712 -5284 -12696
rect -5318 -12944 -5284 -12928
rect -5166 -12712 -5132 -12696
rect -5166 -12944 -5132 -12928
rect -5068 -12712 -5034 -12696
rect -5068 -12944 -5034 -12928
rect -4916 -12712 -4882 -12696
rect -4916 -12944 -4882 -12928
rect -4818 -12712 -4784 -12696
rect -4818 -12944 -4784 -12928
rect -4666 -12712 -4632 -12696
rect -4666 -12944 -4632 -12928
rect -4568 -12712 -4534 -12696
rect -4568 -12944 -4534 -12928
rect -4416 -12712 -4382 -12696
rect -4416 -12944 -4382 -12928
rect -4318 -12712 -4284 -12696
rect -4318 -12944 -4284 -12928
rect -4166 -12712 -4132 -12696
rect -4166 -12944 -4132 -12928
rect -4068 -12712 -4034 -12696
rect -4068 -12944 -4034 -12928
rect -5883 -13012 -5867 -12978
rect -5833 -13012 -5817 -12978
rect -5633 -13012 -5617 -12978
rect -5583 -13012 -5567 -12978
rect -5383 -13012 -5367 -12978
rect -5333 -13012 -5317 -12978
rect -5133 -13012 -5117 -12978
rect -5083 -13012 -5067 -12978
rect -4883 -13012 -4867 -12978
rect -4833 -13012 -4817 -12978
rect -4633 -13012 -4617 -12978
rect -4583 -13012 -4567 -12978
rect -4383 -13012 -4367 -12978
rect -4333 -13012 -4317 -12978
rect -4133 -13012 -4117 -12978
rect -4083 -13012 -4067 -12978
rect -2105 -13082 -2089 -13048
rect -2045 -13082 -2029 -13048
rect -1927 -13082 -1911 -13048
rect -1867 -13082 -1851 -13048
rect -1749 -13082 -1733 -13048
rect -1689 -13082 -1673 -13048
rect -1571 -13082 -1555 -13048
rect -1511 -13082 -1495 -13048
rect -1393 -13082 -1377 -13048
rect -1333 -13082 -1317 -13048
rect -1215 -13082 -1199 -13048
rect -1155 -13082 -1139 -13048
rect -1037 -13082 -1021 -13048
rect -977 -13082 -961 -13048
rect -859 -13082 -843 -13048
rect -799 -13082 -783 -13048
rect -681 -13082 -665 -13048
rect -621 -13082 -605 -13048
rect -503 -13082 -487 -13048
rect -443 -13082 -427 -13048
rect -325 -13082 -309 -13048
rect -265 -13082 -249 -13048
rect -147 -13082 -131 -13048
rect -87 -13082 -71 -13048
rect 31 -13082 47 -13048
rect 91 -13082 107 -13048
rect 209 -13082 225 -13048
rect 269 -13082 285 -13048
rect 387 -13082 403 -13048
rect 447 -13082 463 -13048
rect 565 -13082 581 -13048
rect 625 -13082 641 -13048
rect 743 -13082 759 -13048
rect 803 -13082 819 -13048
rect 921 -13082 937 -13048
rect 981 -13082 997 -13048
rect 1099 -13082 1115 -13048
rect 1159 -13082 1175 -13048
rect 1277 -13082 1293 -13048
rect 1337 -13082 1353 -13048
rect 1455 -13082 1471 -13048
rect 1515 -13082 1531 -13048
rect 1633 -13082 1649 -13048
rect 1693 -13082 1709 -13048
rect 1811 -13082 1827 -13048
rect 1871 -13082 1887 -13048
rect 1989 -13082 2005 -13048
rect 2049 -13082 2065 -13048
rect 2167 -13082 2183 -13048
rect 2227 -13082 2243 -13048
rect 2345 -13082 2361 -13048
rect 2405 -13082 2421 -13048
rect 2523 -13082 2539 -13048
rect 2583 -13082 2599 -13048
rect 2701 -13082 2717 -13048
rect 2761 -13082 2777 -13048
rect 2879 -13082 2895 -13048
rect 2939 -13082 2955 -13048
rect 3057 -13082 3073 -13048
rect 3117 -13082 3133 -13048
rect 3235 -13082 3251 -13048
rect 3295 -13082 3311 -13048
rect 3413 -13082 3429 -13048
rect 3473 -13082 3489 -13048
rect 3591 -13082 3607 -13048
rect 3651 -13082 3667 -13048
rect 3769 -13082 3785 -13048
rect 3829 -13082 3845 -13048
rect 3947 -13082 3963 -13048
rect 4007 -13082 4023 -13048
rect -2173 -13132 -2139 -13116
rect -5883 -13342 -5867 -13308
rect -5833 -13342 -5817 -13308
rect -5633 -13342 -5617 -13308
rect -5583 -13342 -5567 -13308
rect -5383 -13342 -5367 -13308
rect -5333 -13342 -5317 -13308
rect -5133 -13342 -5117 -13308
rect -5083 -13342 -5067 -13308
rect -4883 -13342 -4867 -13308
rect -4833 -13342 -4817 -13308
rect -4633 -13342 -4617 -13308
rect -4583 -13342 -4567 -13308
rect -4383 -13342 -4367 -13308
rect -4333 -13342 -4317 -13308
rect -4133 -13342 -4117 -13308
rect -4083 -13342 -4067 -13308
rect -5916 -13392 -5882 -13376
rect -5916 -13624 -5882 -13608
rect -5818 -13392 -5784 -13376
rect -5818 -13624 -5784 -13608
rect -5666 -13392 -5632 -13376
rect -5666 -13624 -5632 -13608
rect -5568 -13392 -5534 -13376
rect -5568 -13624 -5534 -13608
rect -5416 -13392 -5382 -13376
rect -5416 -13624 -5382 -13608
rect -5318 -13392 -5284 -13376
rect -5318 -13624 -5284 -13608
rect -5166 -13392 -5132 -13376
rect -5166 -13624 -5132 -13608
rect -5068 -13392 -5034 -13376
rect -5068 -13624 -5034 -13608
rect -4916 -13392 -4882 -13376
rect -4916 -13624 -4882 -13608
rect -4818 -13392 -4784 -13376
rect -4818 -13624 -4784 -13608
rect -4666 -13392 -4632 -13376
rect -4666 -13624 -4632 -13608
rect -4568 -13392 -4534 -13376
rect -4568 -13624 -4534 -13608
rect -4416 -13392 -4382 -13376
rect -4416 -13624 -4382 -13608
rect -4318 -13392 -4284 -13376
rect -4318 -13624 -4284 -13608
rect -4166 -13392 -4132 -13376
rect -4166 -13624 -4132 -13608
rect -4068 -13392 -4034 -13376
rect -2173 -13404 -2139 -13388
rect -1995 -13132 -1961 -13116
rect -1995 -13404 -1961 -13388
rect -1817 -13132 -1783 -13116
rect -1817 -13404 -1783 -13388
rect -1639 -13132 -1605 -13116
rect -1639 -13404 -1605 -13388
rect -1461 -13132 -1427 -13116
rect -1461 -13404 -1427 -13388
rect -1283 -13132 -1249 -13116
rect -1283 -13404 -1249 -13388
rect -1105 -13132 -1071 -13116
rect -1105 -13404 -1071 -13388
rect -927 -13132 -893 -13116
rect -927 -13404 -893 -13388
rect -749 -13132 -715 -13116
rect -749 -13404 -715 -13388
rect -571 -13132 -537 -13116
rect -571 -13404 -537 -13388
rect -393 -13132 -359 -13116
rect -393 -13404 -359 -13388
rect -215 -13132 -181 -13116
rect -215 -13404 -181 -13388
rect -37 -13132 -3 -13116
rect -37 -13404 -3 -13388
rect 141 -13132 175 -13116
rect 141 -13404 175 -13388
rect 319 -13132 353 -13116
rect 319 -13404 353 -13388
rect 497 -13132 531 -13116
rect 497 -13404 531 -13388
rect 675 -13132 709 -13116
rect 675 -13404 709 -13388
rect 853 -13132 887 -13116
rect 853 -13404 887 -13388
rect 1031 -13132 1065 -13116
rect 1031 -13404 1065 -13388
rect 1209 -13132 1243 -13116
rect 1209 -13404 1243 -13388
rect 1387 -13132 1421 -13116
rect 1387 -13404 1421 -13388
rect 1565 -13132 1599 -13116
rect 1565 -13404 1599 -13388
rect 1743 -13132 1777 -13116
rect 1743 -13404 1777 -13388
rect 1921 -13132 1955 -13116
rect 1921 -13404 1955 -13388
rect 2099 -13132 2133 -13116
rect 2099 -13404 2133 -13388
rect 2277 -13132 2311 -13116
rect 2277 -13404 2311 -13388
rect 2455 -13132 2489 -13116
rect 2455 -13404 2489 -13388
rect 2633 -13132 2667 -13116
rect 2633 -13404 2667 -13388
rect 2811 -13132 2845 -13116
rect 2811 -13404 2845 -13388
rect 2989 -13132 3023 -13116
rect 2989 -13404 3023 -13388
rect 3167 -13132 3201 -13116
rect 3167 -13404 3201 -13388
rect 3345 -13132 3379 -13116
rect 3345 -13404 3379 -13388
rect 3523 -13132 3557 -13116
rect 3523 -13404 3557 -13388
rect 3701 -13132 3735 -13116
rect 3701 -13404 3735 -13388
rect 3879 -13132 3913 -13116
rect 3879 -13404 3913 -13388
rect 4057 -13132 4091 -13116
rect 4057 -13404 4091 -13388
rect -2105 -13472 -2089 -13438
rect -2045 -13472 -2029 -13438
rect -1927 -13472 -1911 -13438
rect -1867 -13472 -1851 -13438
rect -1749 -13472 -1733 -13438
rect -1689 -13472 -1673 -13438
rect -1571 -13472 -1555 -13438
rect -1511 -13472 -1495 -13438
rect -1393 -13472 -1377 -13438
rect -1333 -13472 -1317 -13438
rect -1215 -13472 -1199 -13438
rect -1155 -13472 -1139 -13438
rect -1037 -13472 -1021 -13438
rect -977 -13472 -961 -13438
rect -859 -13472 -843 -13438
rect -799 -13472 -783 -13438
rect -681 -13472 -665 -13438
rect -621 -13472 -605 -13438
rect -503 -13472 -487 -13438
rect -443 -13472 -427 -13438
rect -325 -13472 -309 -13438
rect -265 -13472 -249 -13438
rect -147 -13472 -131 -13438
rect -87 -13472 -71 -13438
rect 31 -13472 47 -13438
rect 91 -13472 107 -13438
rect 209 -13472 225 -13438
rect 269 -13472 285 -13438
rect 387 -13472 403 -13438
rect 447 -13472 463 -13438
rect 565 -13472 581 -13438
rect 625 -13472 641 -13438
rect 743 -13472 759 -13438
rect 803 -13472 819 -13438
rect 921 -13472 937 -13438
rect 981 -13472 997 -13438
rect 1099 -13472 1115 -13438
rect 1159 -13472 1175 -13438
rect 1277 -13472 1293 -13438
rect 1337 -13472 1353 -13438
rect 1455 -13472 1471 -13438
rect 1515 -13472 1531 -13438
rect 1633 -13472 1649 -13438
rect 1693 -13472 1709 -13438
rect 1811 -13472 1827 -13438
rect 1871 -13472 1887 -13438
rect 1989 -13472 2005 -13438
rect 2049 -13472 2065 -13438
rect 2167 -13472 2183 -13438
rect 2227 -13472 2243 -13438
rect 2345 -13472 2361 -13438
rect 2405 -13472 2421 -13438
rect 2523 -13472 2539 -13438
rect 2583 -13472 2599 -13438
rect 2701 -13472 2717 -13438
rect 2761 -13472 2777 -13438
rect 2879 -13472 2895 -13438
rect 2939 -13472 2955 -13438
rect 3057 -13472 3073 -13438
rect 3117 -13472 3133 -13438
rect 3235 -13472 3251 -13438
rect 3295 -13472 3311 -13438
rect 3413 -13472 3429 -13438
rect 3473 -13472 3489 -13438
rect 3591 -13472 3607 -13438
rect 3651 -13472 3667 -13438
rect 3769 -13472 3785 -13438
rect 3829 -13472 3845 -13438
rect 3947 -13472 3963 -13438
rect 4007 -13472 4023 -13438
rect -4068 -13624 -4034 -13608
rect -5883 -13692 -5867 -13658
rect -5833 -13692 -5817 -13658
rect -5633 -13692 -5617 -13658
rect -5583 -13692 -5567 -13658
rect -5383 -13692 -5367 -13658
rect -5333 -13692 -5317 -13658
rect -5133 -13692 -5117 -13658
rect -5083 -13692 -5067 -13658
rect -4883 -13692 -4867 -13658
rect -4833 -13692 -4817 -13658
rect -4633 -13692 -4617 -13658
rect -4583 -13692 -4567 -13658
rect -4383 -13692 -4367 -13658
rect -4333 -13692 -4317 -13658
rect -4133 -13692 -4117 -13658
rect -4083 -13692 -4067 -13658
rect -2105 -14082 -2089 -14048
rect -2045 -14082 -2029 -14048
rect -1927 -14082 -1911 -14048
rect -1867 -14082 -1851 -14048
rect -1749 -14082 -1733 -14048
rect -1689 -14082 -1673 -14048
rect -1571 -14082 -1555 -14048
rect -1511 -14082 -1495 -14048
rect -1393 -14082 -1377 -14048
rect -1333 -14082 -1317 -14048
rect -1215 -14082 -1199 -14048
rect -1155 -14082 -1139 -14048
rect -1037 -14082 -1021 -14048
rect -977 -14082 -961 -14048
rect -859 -14082 -843 -14048
rect -799 -14082 -783 -14048
rect -681 -14082 -665 -14048
rect -621 -14082 -605 -14048
rect -503 -14082 -487 -14048
rect -443 -14082 -427 -14048
rect -325 -14082 -309 -14048
rect -265 -14082 -249 -14048
rect -147 -14082 -131 -14048
rect -87 -14082 -71 -14048
rect 31 -14082 47 -14048
rect 91 -14082 107 -14048
rect 209 -14082 225 -14048
rect 269 -14082 285 -14048
rect 387 -14082 403 -14048
rect 447 -14082 463 -14048
rect 565 -14082 581 -14048
rect 625 -14082 641 -14048
rect 743 -14082 759 -14048
rect 803 -14082 819 -14048
rect 921 -14082 937 -14048
rect 981 -14082 997 -14048
rect 1099 -14082 1115 -14048
rect 1159 -14082 1175 -14048
rect 1277 -14082 1293 -14048
rect 1337 -14082 1353 -14048
rect 1455 -14082 1471 -14048
rect 1515 -14082 1531 -14048
rect 1633 -14082 1649 -14048
rect 1693 -14082 1709 -14048
rect 1811 -14082 1827 -14048
rect 1871 -14082 1887 -14048
rect 1989 -14082 2005 -14048
rect 2049 -14082 2065 -14048
rect 2167 -14082 2183 -14048
rect 2227 -14082 2243 -14048
rect 2345 -14082 2361 -14048
rect 2405 -14082 2421 -14048
rect 2523 -14082 2539 -14048
rect 2583 -14082 2599 -14048
rect 2701 -14082 2717 -14048
rect 2761 -14082 2777 -14048
rect 2879 -14082 2895 -14048
rect 2939 -14082 2955 -14048
rect 3057 -14082 3073 -14048
rect 3117 -14082 3133 -14048
rect 3235 -14082 3251 -14048
rect 3295 -14082 3311 -14048
rect 3413 -14082 3429 -14048
rect 3473 -14082 3489 -14048
rect 3591 -14082 3607 -14048
rect 3651 -14082 3667 -14048
rect 3769 -14082 3785 -14048
rect 3829 -14082 3845 -14048
rect 3947 -14082 3963 -14048
rect 4007 -14082 4023 -14048
rect 5645 -14082 5661 -14048
rect 5705 -14082 5721 -14048
rect 5823 -14082 5839 -14048
rect 5883 -14082 5899 -14048
rect 6001 -14082 6017 -14048
rect 6061 -14082 6077 -14048
rect 6179 -14082 6195 -14048
rect 6239 -14082 6255 -14048
rect 6357 -14082 6373 -14048
rect 6417 -14082 6433 -14048
rect 6535 -14082 6551 -14048
rect 6595 -14082 6611 -14048
rect 6713 -14082 6729 -14048
rect 6773 -14082 6789 -14048
rect 6891 -14082 6907 -14048
rect 6951 -14082 6967 -14048
rect 7069 -14082 7085 -14048
rect 7129 -14082 7145 -14048
rect 7247 -14082 7263 -14048
rect 7307 -14082 7323 -14048
rect 7425 -14082 7441 -14048
rect 7485 -14082 7501 -14048
rect 7603 -14082 7619 -14048
rect 7663 -14082 7679 -14048
rect 7781 -14082 7797 -14048
rect 7841 -14082 7857 -14048
rect 7959 -14082 7975 -14048
rect 8019 -14082 8035 -14048
rect 8137 -14082 8153 -14048
rect 8197 -14082 8213 -14048
rect 8315 -14082 8331 -14048
rect 8375 -14082 8391 -14048
rect 8493 -14082 8509 -14048
rect 8553 -14082 8569 -14048
rect 8671 -14082 8687 -14048
rect 8731 -14082 8747 -14048
rect 8849 -14082 8865 -14048
rect 8909 -14082 8925 -14048
rect 9027 -14082 9043 -14048
rect 9087 -14082 9103 -14048
rect 9205 -14082 9221 -14048
rect 9265 -14082 9281 -14048
rect 9383 -14082 9399 -14048
rect 9443 -14082 9459 -14048
rect 9561 -14082 9577 -14048
rect 9621 -14082 9637 -14048
rect 9739 -14082 9755 -14048
rect 9799 -14082 9815 -14048
rect 9917 -14082 9933 -14048
rect 9977 -14082 9993 -14048
rect 10095 -14082 10111 -14048
rect 10155 -14082 10171 -14048
rect 10273 -14082 10289 -14048
rect 10333 -14082 10349 -14048
rect 10451 -14082 10467 -14048
rect 10511 -14082 10527 -14048
rect 10629 -14082 10645 -14048
rect 10689 -14082 10705 -14048
rect 10807 -14082 10823 -14048
rect 10867 -14082 10883 -14048
rect 10985 -14082 11001 -14048
rect 11045 -14082 11061 -14048
rect 11163 -14082 11179 -14048
rect 11223 -14082 11239 -14048
rect 11341 -14082 11357 -14048
rect 11401 -14082 11417 -14048
rect 11519 -14082 11535 -14048
rect 11579 -14082 11595 -14048
rect 11697 -14082 11713 -14048
rect 11757 -14082 11773 -14048
rect 11875 -14082 11891 -14048
rect 11935 -14082 11951 -14048
rect 12053 -14082 12069 -14048
rect 12113 -14082 12129 -14048
rect 12231 -14082 12247 -14048
rect 12291 -14082 12307 -14048
rect 12409 -14082 12425 -14048
rect 12469 -14082 12485 -14048
rect 12587 -14082 12603 -14048
rect 12647 -14082 12663 -14048
rect -2173 -14132 -2139 -14116
rect -5960 -14344 -5944 -14310
rect -5900 -14344 -5884 -14310
rect -5782 -14344 -5766 -14310
rect -5722 -14344 -5706 -14310
rect -5604 -14344 -5588 -14310
rect -5544 -14344 -5528 -14310
rect -5426 -14344 -5410 -14310
rect -5366 -14344 -5350 -14310
rect -5248 -14344 -5232 -14310
rect -5188 -14344 -5172 -14310
rect -5070 -14344 -5054 -14310
rect -5010 -14344 -4994 -14310
rect -4892 -14344 -4876 -14310
rect -4832 -14344 -4816 -14310
rect -4714 -14344 -4698 -14310
rect -4654 -14344 -4638 -14310
rect -4536 -14344 -4520 -14310
rect -4476 -14344 -4460 -14310
rect -4358 -14344 -4342 -14310
rect -4298 -14344 -4282 -14310
rect -4180 -14344 -4164 -14310
rect -4120 -14344 -4104 -14310
rect -6028 -14394 -5994 -14378
rect -6028 -14666 -5994 -14650
rect -5850 -14394 -5816 -14378
rect -5850 -14666 -5816 -14650
rect -5672 -14394 -5638 -14378
rect -5672 -14666 -5638 -14650
rect -5494 -14394 -5460 -14378
rect -5494 -14666 -5460 -14650
rect -5316 -14394 -5282 -14378
rect -5316 -14666 -5282 -14650
rect -5138 -14394 -5104 -14378
rect -5138 -14666 -5104 -14650
rect -4960 -14394 -4926 -14378
rect -4960 -14666 -4926 -14650
rect -4782 -14394 -4748 -14378
rect -4782 -14666 -4748 -14650
rect -4604 -14394 -4570 -14378
rect -4604 -14666 -4570 -14650
rect -4426 -14394 -4392 -14378
rect -4426 -14666 -4392 -14650
rect -4248 -14394 -4214 -14378
rect -4248 -14666 -4214 -14650
rect -4070 -14394 -4036 -14378
rect -2173 -14404 -2139 -14388
rect -1995 -14132 -1961 -14116
rect -1995 -14404 -1961 -14388
rect -1817 -14132 -1783 -14116
rect -1817 -14404 -1783 -14388
rect -1639 -14132 -1605 -14116
rect -1639 -14404 -1605 -14388
rect -1461 -14132 -1427 -14116
rect -1461 -14404 -1427 -14388
rect -1283 -14132 -1249 -14116
rect -1283 -14404 -1249 -14388
rect -1105 -14132 -1071 -14116
rect -1105 -14404 -1071 -14388
rect -927 -14132 -893 -14116
rect -927 -14404 -893 -14388
rect -749 -14132 -715 -14116
rect -749 -14404 -715 -14388
rect -571 -14132 -537 -14116
rect -571 -14404 -537 -14388
rect -393 -14132 -359 -14116
rect -393 -14404 -359 -14388
rect -215 -14132 -181 -14116
rect -215 -14404 -181 -14388
rect -37 -14132 -3 -14116
rect -37 -14404 -3 -14388
rect 141 -14132 175 -14116
rect 141 -14404 175 -14388
rect 319 -14132 353 -14116
rect 319 -14404 353 -14388
rect 497 -14132 531 -14116
rect 497 -14404 531 -14388
rect 675 -14132 709 -14116
rect 675 -14404 709 -14388
rect 853 -14132 887 -14116
rect 853 -14404 887 -14388
rect 1031 -14132 1065 -14116
rect 1031 -14404 1065 -14388
rect 1209 -14132 1243 -14116
rect 1209 -14404 1243 -14388
rect 1387 -14132 1421 -14116
rect 1387 -14404 1421 -14388
rect 1565 -14132 1599 -14116
rect 1565 -14404 1599 -14388
rect 1743 -14132 1777 -14116
rect 1743 -14404 1777 -14388
rect 1921 -14132 1955 -14116
rect 1921 -14404 1955 -14388
rect 2099 -14132 2133 -14116
rect 2099 -14404 2133 -14388
rect 2277 -14132 2311 -14116
rect 2277 -14404 2311 -14388
rect 2455 -14132 2489 -14116
rect 2455 -14404 2489 -14388
rect 2633 -14132 2667 -14116
rect 2633 -14404 2667 -14388
rect 2811 -14132 2845 -14116
rect 2811 -14404 2845 -14388
rect 2989 -14132 3023 -14116
rect 2989 -14404 3023 -14388
rect 3167 -14132 3201 -14116
rect 3167 -14404 3201 -14388
rect 3345 -14132 3379 -14116
rect 3345 -14404 3379 -14388
rect 3523 -14132 3557 -14116
rect 3523 -14404 3557 -14388
rect 3701 -14132 3735 -14116
rect 3701 -14404 3735 -14388
rect 3879 -14132 3913 -14116
rect 3879 -14404 3913 -14388
rect 4057 -14132 4091 -14116
rect 4057 -14404 4091 -14388
rect 5577 -14132 5611 -14116
rect 5577 -14404 5611 -14388
rect 5755 -14132 5789 -14116
rect 5755 -14404 5789 -14388
rect 5933 -14132 5967 -14116
rect 5933 -14404 5967 -14388
rect 6111 -14132 6145 -14116
rect 6111 -14404 6145 -14388
rect 6289 -14132 6323 -14116
rect 6289 -14404 6323 -14388
rect 6467 -14132 6501 -14116
rect 6467 -14404 6501 -14388
rect 6645 -14132 6679 -14116
rect 6645 -14404 6679 -14388
rect 6823 -14132 6857 -14116
rect 6823 -14404 6857 -14388
rect 7001 -14132 7035 -14116
rect 7001 -14404 7035 -14388
rect 7179 -14132 7213 -14116
rect 7179 -14404 7213 -14388
rect 7357 -14132 7391 -14116
rect 7357 -14404 7391 -14388
rect 7535 -14132 7569 -14116
rect 7535 -14404 7569 -14388
rect 7713 -14132 7747 -14116
rect 7713 -14404 7747 -14388
rect 7891 -14132 7925 -14116
rect 7891 -14404 7925 -14388
rect 8069 -14132 8103 -14116
rect 8069 -14404 8103 -14388
rect 8247 -14132 8281 -14116
rect 8247 -14404 8281 -14388
rect 8425 -14132 8459 -14116
rect 8425 -14404 8459 -14388
rect 8603 -14132 8637 -14116
rect 8603 -14404 8637 -14388
rect 8781 -14132 8815 -14116
rect 8781 -14404 8815 -14388
rect 8959 -14132 8993 -14116
rect 8959 -14404 8993 -14388
rect 9137 -14132 9171 -14116
rect 9137 -14404 9171 -14388
rect 9315 -14132 9349 -14116
rect 9315 -14404 9349 -14388
rect 9493 -14132 9527 -14116
rect 9493 -14404 9527 -14388
rect 9671 -14132 9705 -14116
rect 9671 -14404 9705 -14388
rect 9849 -14132 9883 -14116
rect 9849 -14404 9883 -14388
rect 10027 -14132 10061 -14116
rect 10027 -14404 10061 -14388
rect 10205 -14132 10239 -14116
rect 10205 -14404 10239 -14388
rect 10383 -14132 10417 -14116
rect 10383 -14404 10417 -14388
rect 10561 -14132 10595 -14116
rect 10561 -14404 10595 -14388
rect 10739 -14132 10773 -14116
rect 10739 -14404 10773 -14388
rect 10917 -14132 10951 -14116
rect 10917 -14404 10951 -14388
rect 11095 -14132 11129 -14116
rect 11095 -14404 11129 -14388
rect 11273 -14132 11307 -14116
rect 11273 -14404 11307 -14388
rect 11451 -14132 11485 -14116
rect 11451 -14404 11485 -14388
rect 11629 -14132 11663 -14116
rect 11629 -14404 11663 -14388
rect 11807 -14132 11841 -14116
rect 11807 -14404 11841 -14388
rect 11985 -14132 12019 -14116
rect 11985 -14404 12019 -14388
rect 12163 -14132 12197 -14116
rect 12163 -14404 12197 -14388
rect 12341 -14132 12375 -14116
rect 12341 -14404 12375 -14388
rect 12519 -14132 12553 -14116
rect 12519 -14404 12553 -14388
rect 12697 -14132 12731 -14116
rect 12697 -14404 12731 -14388
rect -2105 -14472 -2089 -14438
rect -2045 -14472 -2029 -14438
rect -1927 -14472 -1911 -14438
rect -1867 -14472 -1851 -14438
rect -1749 -14472 -1733 -14438
rect -1689 -14472 -1673 -14438
rect -1571 -14472 -1555 -14438
rect -1511 -14472 -1495 -14438
rect -1393 -14472 -1377 -14438
rect -1333 -14472 -1317 -14438
rect -1215 -14472 -1199 -14438
rect -1155 -14472 -1139 -14438
rect -1037 -14472 -1021 -14438
rect -977 -14472 -961 -14438
rect -859 -14472 -843 -14438
rect -799 -14472 -783 -14438
rect -681 -14472 -665 -14438
rect -621 -14472 -605 -14438
rect -503 -14472 -487 -14438
rect -443 -14472 -427 -14438
rect -325 -14472 -309 -14438
rect -265 -14472 -249 -14438
rect -147 -14472 -131 -14438
rect -87 -14472 -71 -14438
rect 31 -14472 47 -14438
rect 91 -14472 107 -14438
rect 209 -14472 225 -14438
rect 269 -14472 285 -14438
rect 387 -14472 403 -14438
rect 447 -14472 463 -14438
rect 565 -14472 581 -14438
rect 625 -14472 641 -14438
rect 743 -14472 759 -14438
rect 803 -14472 819 -14438
rect 921 -14472 937 -14438
rect 981 -14472 997 -14438
rect 1099 -14472 1115 -14438
rect 1159 -14472 1175 -14438
rect 1277 -14472 1293 -14438
rect 1337 -14472 1353 -14438
rect 1455 -14472 1471 -14438
rect 1515 -14472 1531 -14438
rect 1633 -14472 1649 -14438
rect 1693 -14472 1709 -14438
rect 1811 -14472 1827 -14438
rect 1871 -14472 1887 -14438
rect 1989 -14472 2005 -14438
rect 2049 -14472 2065 -14438
rect 2167 -14472 2183 -14438
rect 2227 -14472 2243 -14438
rect 2345 -14472 2361 -14438
rect 2405 -14472 2421 -14438
rect 2523 -14472 2539 -14438
rect 2583 -14472 2599 -14438
rect 2701 -14472 2717 -14438
rect 2761 -14472 2777 -14438
rect 2879 -14472 2895 -14438
rect 2939 -14472 2955 -14438
rect 3057 -14472 3073 -14438
rect 3117 -14472 3133 -14438
rect 3235 -14472 3251 -14438
rect 3295 -14472 3311 -14438
rect 3413 -14472 3429 -14438
rect 3473 -14472 3489 -14438
rect 3591 -14472 3607 -14438
rect 3651 -14472 3667 -14438
rect 3769 -14472 3785 -14438
rect 3829 -14472 3845 -14438
rect 3947 -14472 3963 -14438
rect 4007 -14472 4023 -14438
rect 5645 -14472 5661 -14438
rect 5705 -14472 5721 -14438
rect 5823 -14472 5839 -14438
rect 5883 -14472 5899 -14438
rect 6001 -14472 6017 -14438
rect 6061 -14472 6077 -14438
rect 6179 -14472 6195 -14438
rect 6239 -14472 6255 -14438
rect 6357 -14472 6373 -14438
rect 6417 -14472 6433 -14438
rect 6535 -14472 6551 -14438
rect 6595 -14472 6611 -14438
rect 6713 -14472 6729 -14438
rect 6773 -14472 6789 -14438
rect 6891 -14472 6907 -14438
rect 6951 -14472 6967 -14438
rect 7069 -14472 7085 -14438
rect 7129 -14472 7145 -14438
rect 7247 -14472 7263 -14438
rect 7307 -14472 7323 -14438
rect 7425 -14472 7441 -14438
rect 7485 -14472 7501 -14438
rect 7603 -14472 7619 -14438
rect 7663 -14472 7679 -14438
rect 7781 -14472 7797 -14438
rect 7841 -14472 7857 -14438
rect 7959 -14472 7975 -14438
rect 8019 -14472 8035 -14438
rect 8137 -14472 8153 -14438
rect 8197 -14472 8213 -14438
rect 8315 -14472 8331 -14438
rect 8375 -14472 8391 -14438
rect 8493 -14472 8509 -14438
rect 8553 -14472 8569 -14438
rect 8671 -14472 8687 -14438
rect 8731 -14472 8747 -14438
rect 8849 -14472 8865 -14438
rect 8909 -14472 8925 -14438
rect 9027 -14472 9043 -14438
rect 9087 -14472 9103 -14438
rect 9205 -14472 9221 -14438
rect 9265 -14472 9281 -14438
rect 9383 -14472 9399 -14438
rect 9443 -14472 9459 -14438
rect 9561 -14472 9577 -14438
rect 9621 -14472 9637 -14438
rect 9739 -14472 9755 -14438
rect 9799 -14472 9815 -14438
rect 9917 -14472 9933 -14438
rect 9977 -14472 9993 -14438
rect 10095 -14472 10111 -14438
rect 10155 -14472 10171 -14438
rect 10273 -14472 10289 -14438
rect 10333 -14472 10349 -14438
rect 10451 -14472 10467 -14438
rect 10511 -14472 10527 -14438
rect 10629 -14472 10645 -14438
rect 10689 -14472 10705 -14438
rect 10807 -14472 10823 -14438
rect 10867 -14472 10883 -14438
rect 10985 -14472 11001 -14438
rect 11045 -14472 11061 -14438
rect 11163 -14472 11179 -14438
rect 11223 -14472 11239 -14438
rect 11341 -14472 11357 -14438
rect 11401 -14472 11417 -14438
rect 11519 -14472 11535 -14438
rect 11579 -14472 11595 -14438
rect 11697 -14472 11713 -14438
rect 11757 -14472 11773 -14438
rect 11875 -14472 11891 -14438
rect 11935 -14472 11951 -14438
rect 12053 -14472 12069 -14438
rect 12113 -14472 12129 -14438
rect 12231 -14472 12247 -14438
rect 12291 -14472 12307 -14438
rect 12409 -14472 12425 -14438
rect 12469 -14472 12485 -14438
rect 12587 -14472 12603 -14438
rect 12647 -14472 12663 -14438
rect -4070 -14666 -4036 -14650
rect -5960 -14734 -5944 -14700
rect -5900 -14734 -5884 -14700
rect -5782 -14734 -5766 -14700
rect -5722 -14734 -5706 -14700
rect -5604 -14734 -5588 -14700
rect -5544 -14734 -5528 -14700
rect -5426 -14734 -5410 -14700
rect -5366 -14734 -5350 -14700
rect -5248 -14734 -5232 -14700
rect -5188 -14734 -5172 -14700
rect -5070 -14734 -5054 -14700
rect -5010 -14734 -4994 -14700
rect -4892 -14734 -4876 -14700
rect -4832 -14734 -4816 -14700
rect -4714 -14734 -4698 -14700
rect -4654 -14734 -4638 -14700
rect -4536 -14734 -4520 -14700
rect -4476 -14734 -4460 -14700
rect -4358 -14734 -4342 -14700
rect -4298 -14734 -4282 -14700
rect -4180 -14734 -4164 -14700
rect -4120 -14734 -4104 -14700
rect -5960 -15044 -5944 -15010
rect -5900 -15044 -5884 -15010
rect -5782 -15044 -5766 -15010
rect -5722 -15044 -5706 -15010
rect -5604 -15044 -5588 -15010
rect -5544 -15044 -5528 -15010
rect -5426 -15044 -5410 -15010
rect -5366 -15044 -5350 -15010
rect -5248 -15044 -5232 -15010
rect -5188 -15044 -5172 -15010
rect -5070 -15044 -5054 -15010
rect -5010 -15044 -4994 -15010
rect -4892 -15044 -4876 -15010
rect -4832 -15044 -4816 -15010
rect -4714 -15044 -4698 -15010
rect -4654 -15044 -4638 -15010
rect -4536 -15044 -4520 -15010
rect -4476 -15044 -4460 -15010
rect -4358 -15044 -4342 -15010
rect -4298 -15044 -4282 -15010
rect -4180 -15044 -4164 -15010
rect -4120 -15044 -4104 -15010
rect -6028 -15094 -5994 -15078
rect -6028 -15366 -5994 -15350
rect -5850 -15094 -5816 -15078
rect -5850 -15366 -5816 -15350
rect -5672 -15094 -5638 -15078
rect -5672 -15366 -5638 -15350
rect -5494 -15094 -5460 -15078
rect -5494 -15366 -5460 -15350
rect -5316 -15094 -5282 -15078
rect -5316 -15366 -5282 -15350
rect -5138 -15094 -5104 -15078
rect -5138 -15366 -5104 -15350
rect -4960 -15094 -4926 -15078
rect -4960 -15366 -4926 -15350
rect -4782 -15094 -4748 -15078
rect -4782 -15366 -4748 -15350
rect -4604 -15094 -4570 -15078
rect -4604 -15366 -4570 -15350
rect -4426 -15094 -4392 -15078
rect -4426 -15366 -4392 -15350
rect -4248 -15094 -4214 -15078
rect -4248 -15366 -4214 -15350
rect -4070 -15094 -4036 -15078
rect -2105 -15082 -2089 -15048
rect -2045 -15082 -2029 -15048
rect -1927 -15082 -1911 -15048
rect -1867 -15082 -1851 -15048
rect -1749 -15082 -1733 -15048
rect -1689 -15082 -1673 -15048
rect -1571 -15082 -1555 -15048
rect -1511 -15082 -1495 -15048
rect -1393 -15082 -1377 -15048
rect -1333 -15082 -1317 -15048
rect -1215 -15082 -1199 -15048
rect -1155 -15082 -1139 -15048
rect -1037 -15082 -1021 -15048
rect -977 -15082 -961 -15048
rect -859 -15082 -843 -15048
rect -799 -15082 -783 -15048
rect -681 -15082 -665 -15048
rect -621 -15082 -605 -15048
rect -503 -15082 -487 -15048
rect -443 -15082 -427 -15048
rect -325 -15082 -309 -15048
rect -265 -15082 -249 -15048
rect -147 -15082 -131 -15048
rect -87 -15082 -71 -15048
rect 31 -15082 47 -15048
rect 91 -15082 107 -15048
rect 209 -15082 225 -15048
rect 269 -15082 285 -15048
rect 387 -15082 403 -15048
rect 447 -15082 463 -15048
rect 565 -15082 581 -15048
rect 625 -15082 641 -15048
rect 743 -15082 759 -15048
rect 803 -15082 819 -15048
rect 921 -15082 937 -15048
rect 981 -15082 997 -15048
rect 1099 -15082 1115 -15048
rect 1159 -15082 1175 -15048
rect 1277 -15082 1293 -15048
rect 1337 -15082 1353 -15048
rect 1455 -15082 1471 -15048
rect 1515 -15082 1531 -15048
rect 1633 -15082 1649 -15048
rect 1693 -15082 1709 -15048
rect 1811 -15082 1827 -15048
rect 1871 -15082 1887 -15048
rect 1989 -15082 2005 -15048
rect 2049 -15082 2065 -15048
rect 2167 -15082 2183 -15048
rect 2227 -15082 2243 -15048
rect 2345 -15082 2361 -15048
rect 2405 -15082 2421 -15048
rect 2523 -15082 2539 -15048
rect 2583 -15082 2599 -15048
rect 2701 -15082 2717 -15048
rect 2761 -15082 2777 -15048
rect 2879 -15082 2895 -15048
rect 2939 -15082 2955 -15048
rect 3057 -15082 3073 -15048
rect 3117 -15082 3133 -15048
rect 3235 -15082 3251 -15048
rect 3295 -15082 3311 -15048
rect 3413 -15082 3429 -15048
rect 3473 -15082 3489 -15048
rect 3591 -15082 3607 -15048
rect 3651 -15082 3667 -15048
rect 3769 -15082 3785 -15048
rect 3829 -15082 3845 -15048
rect 3947 -15082 3963 -15048
rect 4007 -15082 4023 -15048
rect 5645 -15082 5661 -15048
rect 5705 -15082 5721 -15048
rect 5823 -15082 5839 -15048
rect 5883 -15082 5899 -15048
rect 6001 -15082 6017 -15048
rect 6061 -15082 6077 -15048
rect 6179 -15082 6195 -15048
rect 6239 -15082 6255 -15048
rect 6357 -15082 6373 -15048
rect 6417 -15082 6433 -15048
rect 6535 -15082 6551 -15048
rect 6595 -15082 6611 -15048
rect 6713 -15082 6729 -15048
rect 6773 -15082 6789 -15048
rect 6891 -15082 6907 -15048
rect 6951 -15082 6967 -15048
rect 7069 -15082 7085 -15048
rect 7129 -15082 7145 -15048
rect 7247 -15082 7263 -15048
rect 7307 -15082 7323 -15048
rect 7425 -15082 7441 -15048
rect 7485 -15082 7501 -15048
rect 7603 -15082 7619 -15048
rect 7663 -15082 7679 -15048
rect 7781 -15082 7797 -15048
rect 7841 -15082 7857 -15048
rect 7959 -15082 7975 -15048
rect 8019 -15082 8035 -15048
rect 8137 -15082 8153 -15048
rect 8197 -15082 8213 -15048
rect 8315 -15082 8331 -15048
rect 8375 -15082 8391 -15048
rect 8493 -15082 8509 -15048
rect 8553 -15082 8569 -15048
rect 8671 -15082 8687 -15048
rect 8731 -15082 8747 -15048
rect 8849 -15082 8865 -15048
rect 8909 -15082 8925 -15048
rect 9027 -15082 9043 -15048
rect 9087 -15082 9103 -15048
rect 9205 -15082 9221 -15048
rect 9265 -15082 9281 -15048
rect 9383 -15082 9399 -15048
rect 9443 -15082 9459 -15048
rect 9561 -15082 9577 -15048
rect 9621 -15082 9637 -15048
rect 9739 -15082 9755 -15048
rect 9799 -15082 9815 -15048
rect 9917 -15082 9933 -15048
rect 9977 -15082 9993 -15048
rect 10095 -15082 10111 -15048
rect 10155 -15082 10171 -15048
rect 10273 -15082 10289 -15048
rect 10333 -15082 10349 -15048
rect 10451 -15082 10467 -15048
rect 10511 -15082 10527 -15048
rect 10629 -15082 10645 -15048
rect 10689 -15082 10705 -15048
rect 10807 -15082 10823 -15048
rect 10867 -15082 10883 -15048
rect 10985 -15082 11001 -15048
rect 11045 -15082 11061 -15048
rect 11163 -15082 11179 -15048
rect 11223 -15082 11239 -15048
rect 11341 -15082 11357 -15048
rect 11401 -15082 11417 -15048
rect 11519 -15082 11535 -15048
rect 11579 -15082 11595 -15048
rect 11697 -15082 11713 -15048
rect 11757 -15082 11773 -15048
rect 11875 -15082 11891 -15048
rect 11935 -15082 11951 -15048
rect 12053 -15082 12069 -15048
rect 12113 -15082 12129 -15048
rect 12231 -15082 12247 -15048
rect 12291 -15082 12307 -15048
rect 12409 -15082 12425 -15048
rect 12469 -15082 12485 -15048
rect 12587 -15082 12603 -15048
rect 12647 -15082 12663 -15048
rect -4070 -15366 -4036 -15350
rect -2173 -15132 -2139 -15116
rect -5960 -15434 -5944 -15400
rect -5900 -15434 -5884 -15400
rect -5782 -15434 -5766 -15400
rect -5722 -15434 -5706 -15400
rect -5604 -15434 -5588 -15400
rect -5544 -15434 -5528 -15400
rect -5426 -15434 -5410 -15400
rect -5366 -15434 -5350 -15400
rect -5248 -15434 -5232 -15400
rect -5188 -15434 -5172 -15400
rect -5070 -15434 -5054 -15400
rect -5010 -15434 -4994 -15400
rect -4892 -15434 -4876 -15400
rect -4832 -15434 -4816 -15400
rect -4714 -15434 -4698 -15400
rect -4654 -15434 -4638 -15400
rect -4536 -15434 -4520 -15400
rect -4476 -15434 -4460 -15400
rect -4358 -15434 -4342 -15400
rect -4298 -15434 -4282 -15400
rect -4180 -15434 -4164 -15400
rect -4120 -15434 -4104 -15400
rect -2173 -15404 -2139 -15388
rect -1995 -15132 -1961 -15116
rect -1995 -15404 -1961 -15388
rect -1817 -15132 -1783 -15116
rect -1817 -15404 -1783 -15388
rect -1639 -15132 -1605 -15116
rect -1639 -15404 -1605 -15388
rect -1461 -15132 -1427 -15116
rect -1461 -15404 -1427 -15388
rect -1283 -15132 -1249 -15116
rect -1283 -15404 -1249 -15388
rect -1105 -15132 -1071 -15116
rect -1105 -15404 -1071 -15388
rect -927 -15132 -893 -15116
rect -927 -15404 -893 -15388
rect -749 -15132 -715 -15116
rect -749 -15404 -715 -15388
rect -571 -15132 -537 -15116
rect -571 -15404 -537 -15388
rect -393 -15132 -359 -15116
rect -393 -15404 -359 -15388
rect -215 -15132 -181 -15116
rect -215 -15404 -181 -15388
rect -37 -15132 -3 -15116
rect -37 -15404 -3 -15388
rect 141 -15132 175 -15116
rect 141 -15404 175 -15388
rect 319 -15132 353 -15116
rect 319 -15404 353 -15388
rect 497 -15132 531 -15116
rect 497 -15404 531 -15388
rect 675 -15132 709 -15116
rect 675 -15404 709 -15388
rect 853 -15132 887 -15116
rect 853 -15404 887 -15388
rect 1031 -15132 1065 -15116
rect 1031 -15404 1065 -15388
rect 1209 -15132 1243 -15116
rect 1209 -15404 1243 -15388
rect 1387 -15132 1421 -15116
rect 1387 -15404 1421 -15388
rect 1565 -15132 1599 -15116
rect 1565 -15404 1599 -15388
rect 1743 -15132 1777 -15116
rect 1743 -15404 1777 -15388
rect 1921 -15132 1955 -15116
rect 1921 -15404 1955 -15388
rect 2099 -15132 2133 -15116
rect 2099 -15404 2133 -15388
rect 2277 -15132 2311 -15116
rect 2277 -15404 2311 -15388
rect 2455 -15132 2489 -15116
rect 2455 -15404 2489 -15388
rect 2633 -15132 2667 -15116
rect 2633 -15404 2667 -15388
rect 2811 -15132 2845 -15116
rect 2811 -15404 2845 -15388
rect 2989 -15132 3023 -15116
rect 2989 -15404 3023 -15388
rect 3167 -15132 3201 -15116
rect 3167 -15404 3201 -15388
rect 3345 -15132 3379 -15116
rect 3345 -15404 3379 -15388
rect 3523 -15132 3557 -15116
rect 3523 -15404 3557 -15388
rect 3701 -15132 3735 -15116
rect 3701 -15404 3735 -15388
rect 3879 -15132 3913 -15116
rect 3879 -15404 3913 -15388
rect 4057 -15132 4091 -15116
rect 4057 -15404 4091 -15388
rect 5577 -15132 5611 -15116
rect 5577 -15404 5611 -15388
rect 5755 -15132 5789 -15116
rect 5755 -15404 5789 -15388
rect 5933 -15132 5967 -15116
rect 5933 -15404 5967 -15388
rect 6111 -15132 6145 -15116
rect 6111 -15404 6145 -15388
rect 6289 -15132 6323 -15116
rect 6289 -15404 6323 -15388
rect 6467 -15132 6501 -15116
rect 6467 -15404 6501 -15388
rect 6645 -15132 6679 -15116
rect 6645 -15404 6679 -15388
rect 6823 -15132 6857 -15116
rect 6823 -15404 6857 -15388
rect 7001 -15132 7035 -15116
rect 7001 -15404 7035 -15388
rect 7179 -15132 7213 -15116
rect 7179 -15404 7213 -15388
rect 7357 -15132 7391 -15116
rect 7357 -15404 7391 -15388
rect 7535 -15132 7569 -15116
rect 7535 -15404 7569 -15388
rect 7713 -15132 7747 -15116
rect 7713 -15404 7747 -15388
rect 7891 -15132 7925 -15116
rect 7891 -15404 7925 -15388
rect 8069 -15132 8103 -15116
rect 8069 -15404 8103 -15388
rect 8247 -15132 8281 -15116
rect 8247 -15404 8281 -15388
rect 8425 -15132 8459 -15116
rect 8425 -15404 8459 -15388
rect 8603 -15132 8637 -15116
rect 8603 -15404 8637 -15388
rect 8781 -15132 8815 -15116
rect 8781 -15404 8815 -15388
rect 8959 -15132 8993 -15116
rect 8959 -15404 8993 -15388
rect 9137 -15132 9171 -15116
rect 9137 -15404 9171 -15388
rect 9315 -15132 9349 -15116
rect 9315 -15404 9349 -15388
rect 9493 -15132 9527 -15116
rect 9493 -15404 9527 -15388
rect 9671 -15132 9705 -15116
rect 9671 -15404 9705 -15388
rect 9849 -15132 9883 -15116
rect 9849 -15404 9883 -15388
rect 10027 -15132 10061 -15116
rect 10027 -15404 10061 -15388
rect 10205 -15132 10239 -15116
rect 10205 -15404 10239 -15388
rect 10383 -15132 10417 -15116
rect 10383 -15404 10417 -15388
rect 10561 -15132 10595 -15116
rect 10561 -15404 10595 -15388
rect 10739 -15132 10773 -15116
rect 10739 -15404 10773 -15388
rect 10917 -15132 10951 -15116
rect 10917 -15404 10951 -15388
rect 11095 -15132 11129 -15116
rect 11095 -15404 11129 -15388
rect 11273 -15132 11307 -15116
rect 11273 -15404 11307 -15388
rect 11451 -15132 11485 -15116
rect 11451 -15404 11485 -15388
rect 11629 -15132 11663 -15116
rect 11629 -15404 11663 -15388
rect 11807 -15132 11841 -15116
rect 11807 -15404 11841 -15388
rect 11985 -15132 12019 -15116
rect 11985 -15404 12019 -15388
rect 12163 -15132 12197 -15116
rect 12163 -15404 12197 -15388
rect 12341 -15132 12375 -15116
rect 12341 -15404 12375 -15388
rect 12519 -15132 12553 -15116
rect 12519 -15404 12553 -15388
rect 12697 -15132 12731 -15116
rect 12697 -15404 12731 -15388
rect -2105 -15472 -2089 -15438
rect -2045 -15472 -2029 -15438
rect -1927 -15472 -1911 -15438
rect -1867 -15472 -1851 -15438
rect -1749 -15472 -1733 -15438
rect -1689 -15472 -1673 -15438
rect -1571 -15472 -1555 -15438
rect -1511 -15472 -1495 -15438
rect -1393 -15472 -1377 -15438
rect -1333 -15472 -1317 -15438
rect -1215 -15472 -1199 -15438
rect -1155 -15472 -1139 -15438
rect -1037 -15472 -1021 -15438
rect -977 -15472 -961 -15438
rect -859 -15472 -843 -15438
rect -799 -15472 -783 -15438
rect -681 -15472 -665 -15438
rect -621 -15472 -605 -15438
rect -503 -15472 -487 -15438
rect -443 -15472 -427 -15438
rect -325 -15472 -309 -15438
rect -265 -15472 -249 -15438
rect -147 -15472 -131 -15438
rect -87 -15472 -71 -15438
rect 31 -15472 47 -15438
rect 91 -15472 107 -15438
rect 209 -15472 225 -15438
rect 269 -15472 285 -15438
rect 387 -15472 403 -15438
rect 447 -15472 463 -15438
rect 565 -15472 581 -15438
rect 625 -15472 641 -15438
rect 743 -15472 759 -15438
rect 803 -15472 819 -15438
rect 921 -15472 937 -15438
rect 981 -15472 997 -15438
rect 1099 -15472 1115 -15438
rect 1159 -15472 1175 -15438
rect 1277 -15472 1293 -15438
rect 1337 -15472 1353 -15438
rect 1455 -15472 1471 -15438
rect 1515 -15472 1531 -15438
rect 1633 -15472 1649 -15438
rect 1693 -15472 1709 -15438
rect 1811 -15472 1827 -15438
rect 1871 -15472 1887 -15438
rect 1989 -15472 2005 -15438
rect 2049 -15472 2065 -15438
rect 2167 -15472 2183 -15438
rect 2227 -15472 2243 -15438
rect 2345 -15472 2361 -15438
rect 2405 -15472 2421 -15438
rect 2523 -15472 2539 -15438
rect 2583 -15472 2599 -15438
rect 2701 -15472 2717 -15438
rect 2761 -15472 2777 -15438
rect 2879 -15472 2895 -15438
rect 2939 -15472 2955 -15438
rect 3057 -15472 3073 -15438
rect 3117 -15472 3133 -15438
rect 3235 -15472 3251 -15438
rect 3295 -15472 3311 -15438
rect 3413 -15472 3429 -15438
rect 3473 -15472 3489 -15438
rect 3591 -15472 3607 -15438
rect 3651 -15472 3667 -15438
rect 3769 -15472 3785 -15438
rect 3829 -15472 3845 -15438
rect 3947 -15472 3963 -15438
rect 4007 -15472 4023 -15438
rect 5645 -15472 5661 -15438
rect 5705 -15472 5721 -15438
rect 5823 -15472 5839 -15438
rect 5883 -15472 5899 -15438
rect 6001 -15472 6017 -15438
rect 6061 -15472 6077 -15438
rect 6179 -15472 6195 -15438
rect 6239 -15472 6255 -15438
rect 6357 -15472 6373 -15438
rect 6417 -15472 6433 -15438
rect 6535 -15472 6551 -15438
rect 6595 -15472 6611 -15438
rect 6713 -15472 6729 -15438
rect 6773 -15472 6789 -15438
rect 6891 -15472 6907 -15438
rect 6951 -15472 6967 -15438
rect 7069 -15472 7085 -15438
rect 7129 -15472 7145 -15438
rect 7247 -15472 7263 -15438
rect 7307 -15472 7323 -15438
rect 7425 -15472 7441 -15438
rect 7485 -15472 7501 -15438
rect 7603 -15472 7619 -15438
rect 7663 -15472 7679 -15438
rect 7781 -15472 7797 -15438
rect 7841 -15472 7857 -15438
rect 7959 -15472 7975 -15438
rect 8019 -15472 8035 -15438
rect 8137 -15472 8153 -15438
rect 8197 -15472 8213 -15438
rect 8315 -15472 8331 -15438
rect 8375 -15472 8391 -15438
rect 8493 -15472 8509 -15438
rect 8553 -15472 8569 -15438
rect 8671 -15472 8687 -15438
rect 8731 -15472 8747 -15438
rect 8849 -15472 8865 -15438
rect 8909 -15472 8925 -15438
rect 9027 -15472 9043 -15438
rect 9087 -15472 9103 -15438
rect 9205 -15472 9221 -15438
rect 9265 -15472 9281 -15438
rect 9383 -15472 9399 -15438
rect 9443 -15472 9459 -15438
rect 9561 -15472 9577 -15438
rect 9621 -15472 9637 -15438
rect 9739 -15472 9755 -15438
rect 9799 -15472 9815 -15438
rect 9917 -15472 9933 -15438
rect 9977 -15472 9993 -15438
rect 10095 -15472 10111 -15438
rect 10155 -15472 10171 -15438
rect 10273 -15472 10289 -15438
rect 10333 -15472 10349 -15438
rect 10451 -15472 10467 -15438
rect 10511 -15472 10527 -15438
rect 10629 -15472 10645 -15438
rect 10689 -15472 10705 -15438
rect 10807 -15472 10823 -15438
rect 10867 -15472 10883 -15438
rect 10985 -15472 11001 -15438
rect 11045 -15472 11061 -15438
rect 11163 -15472 11179 -15438
rect 11223 -15472 11239 -15438
rect 11341 -15472 11357 -15438
rect 11401 -15472 11417 -15438
rect 11519 -15472 11535 -15438
rect 11579 -15472 11595 -15438
rect 11697 -15472 11713 -15438
rect 11757 -15472 11773 -15438
rect 11875 -15472 11891 -15438
rect 11935 -15472 11951 -15438
rect 12053 -15472 12069 -15438
rect 12113 -15472 12129 -15438
rect 12231 -15472 12247 -15438
rect 12291 -15472 12307 -15438
rect 12409 -15472 12425 -15438
rect 12469 -15472 12485 -15438
rect 12587 -15472 12603 -15438
rect 12647 -15472 12663 -15438
rect -5960 -15744 -5944 -15710
rect -5900 -15744 -5884 -15710
rect -5782 -15744 -5766 -15710
rect -5722 -15744 -5706 -15710
rect -5604 -15744 -5588 -15710
rect -5544 -15744 -5528 -15710
rect -5426 -15744 -5410 -15710
rect -5366 -15744 -5350 -15710
rect -5248 -15744 -5232 -15710
rect -5188 -15744 -5172 -15710
rect -5070 -15744 -5054 -15710
rect -5010 -15744 -4994 -15710
rect -4892 -15744 -4876 -15710
rect -4832 -15744 -4816 -15710
rect -4714 -15744 -4698 -15710
rect -4654 -15744 -4638 -15710
rect -4536 -15744 -4520 -15710
rect -4476 -15744 -4460 -15710
rect -4358 -15744 -4342 -15710
rect -4298 -15744 -4282 -15710
rect -4180 -15744 -4164 -15710
rect -4120 -15744 -4104 -15710
rect -6028 -15794 -5994 -15778
rect -6028 -16066 -5994 -16050
rect -5850 -15794 -5816 -15778
rect -5850 -16066 -5816 -16050
rect -5672 -15794 -5638 -15778
rect -5672 -16066 -5638 -16050
rect -5494 -15794 -5460 -15778
rect -5494 -16066 -5460 -16050
rect -5316 -15794 -5282 -15778
rect -5316 -16066 -5282 -16050
rect -5138 -15794 -5104 -15778
rect -5138 -16066 -5104 -16050
rect -4960 -15794 -4926 -15778
rect -4960 -16066 -4926 -16050
rect -4782 -15794 -4748 -15778
rect -4782 -16066 -4748 -16050
rect -4604 -15794 -4570 -15778
rect -4604 -16066 -4570 -16050
rect -4426 -15794 -4392 -15778
rect -4426 -16066 -4392 -16050
rect -4248 -15794 -4214 -15778
rect -4248 -16066 -4214 -16050
rect -4070 -15794 -4036 -15778
rect -4070 -16066 -4036 -16050
rect -2105 -16082 -2089 -16048
rect -2045 -16082 -2029 -16048
rect -1927 -16082 -1911 -16048
rect -1867 -16082 -1851 -16048
rect -1749 -16082 -1733 -16048
rect -1689 -16082 -1673 -16048
rect -1571 -16082 -1555 -16048
rect -1511 -16082 -1495 -16048
rect -1393 -16082 -1377 -16048
rect -1333 -16082 -1317 -16048
rect -1215 -16082 -1199 -16048
rect -1155 -16082 -1139 -16048
rect -1037 -16082 -1021 -16048
rect -977 -16082 -961 -16048
rect -859 -16082 -843 -16048
rect -799 -16082 -783 -16048
rect -681 -16082 -665 -16048
rect -621 -16082 -605 -16048
rect -503 -16082 -487 -16048
rect -443 -16082 -427 -16048
rect -325 -16082 -309 -16048
rect -265 -16082 -249 -16048
rect -147 -16082 -131 -16048
rect -87 -16082 -71 -16048
rect 31 -16082 47 -16048
rect 91 -16082 107 -16048
rect 209 -16082 225 -16048
rect 269 -16082 285 -16048
rect 387 -16082 403 -16048
rect 447 -16082 463 -16048
rect 565 -16082 581 -16048
rect 625 -16082 641 -16048
rect 743 -16082 759 -16048
rect 803 -16082 819 -16048
rect 921 -16082 937 -16048
rect 981 -16082 997 -16048
rect 1099 -16082 1115 -16048
rect 1159 -16082 1175 -16048
rect 1277 -16082 1293 -16048
rect 1337 -16082 1353 -16048
rect 1455 -16082 1471 -16048
rect 1515 -16082 1531 -16048
rect 1633 -16082 1649 -16048
rect 1693 -16082 1709 -16048
rect 1811 -16082 1827 -16048
rect 1871 -16082 1887 -16048
rect 1989 -16082 2005 -16048
rect 2049 -16082 2065 -16048
rect 2167 -16082 2183 -16048
rect 2227 -16082 2243 -16048
rect 2345 -16082 2361 -16048
rect 2405 -16082 2421 -16048
rect 2523 -16082 2539 -16048
rect 2583 -16082 2599 -16048
rect 2701 -16082 2717 -16048
rect 2761 -16082 2777 -16048
rect 2879 -16082 2895 -16048
rect 2939 -16082 2955 -16048
rect 3057 -16082 3073 -16048
rect 3117 -16082 3133 -16048
rect 3235 -16082 3251 -16048
rect 3295 -16082 3311 -16048
rect 3413 -16082 3429 -16048
rect 3473 -16082 3489 -16048
rect 3591 -16082 3607 -16048
rect 3651 -16082 3667 -16048
rect 3769 -16082 3785 -16048
rect 3829 -16082 3845 -16048
rect 3947 -16082 3963 -16048
rect 4007 -16082 4023 -16048
rect 5645 -16082 5661 -16048
rect 5705 -16082 5721 -16048
rect 5823 -16082 5839 -16048
rect 5883 -16082 5899 -16048
rect 6001 -16082 6017 -16048
rect 6061 -16082 6077 -16048
rect 6179 -16082 6195 -16048
rect 6239 -16082 6255 -16048
rect 6357 -16082 6373 -16048
rect 6417 -16082 6433 -16048
rect 6535 -16082 6551 -16048
rect 6595 -16082 6611 -16048
rect 6713 -16082 6729 -16048
rect 6773 -16082 6789 -16048
rect 6891 -16082 6907 -16048
rect 6951 -16082 6967 -16048
rect 7069 -16082 7085 -16048
rect 7129 -16082 7145 -16048
rect 7247 -16082 7263 -16048
rect 7307 -16082 7323 -16048
rect 7425 -16082 7441 -16048
rect 7485 -16082 7501 -16048
rect 7603 -16082 7619 -16048
rect 7663 -16082 7679 -16048
rect 7781 -16082 7797 -16048
rect 7841 -16082 7857 -16048
rect 7959 -16082 7975 -16048
rect 8019 -16082 8035 -16048
rect 8137 -16082 8153 -16048
rect 8197 -16082 8213 -16048
rect 8315 -16082 8331 -16048
rect 8375 -16082 8391 -16048
rect 8493 -16082 8509 -16048
rect 8553 -16082 8569 -16048
rect 8671 -16082 8687 -16048
rect 8731 -16082 8747 -16048
rect 8849 -16082 8865 -16048
rect 8909 -16082 8925 -16048
rect 9027 -16082 9043 -16048
rect 9087 -16082 9103 -16048
rect 9205 -16082 9221 -16048
rect 9265 -16082 9281 -16048
rect 9383 -16082 9399 -16048
rect 9443 -16082 9459 -16048
rect 9561 -16082 9577 -16048
rect 9621 -16082 9637 -16048
rect 9739 -16082 9755 -16048
rect 9799 -16082 9815 -16048
rect 9917 -16082 9933 -16048
rect 9977 -16082 9993 -16048
rect 10095 -16082 10111 -16048
rect 10155 -16082 10171 -16048
rect 10273 -16082 10289 -16048
rect 10333 -16082 10349 -16048
rect 10451 -16082 10467 -16048
rect 10511 -16082 10527 -16048
rect 10629 -16082 10645 -16048
rect 10689 -16082 10705 -16048
rect 10807 -16082 10823 -16048
rect 10867 -16082 10883 -16048
rect 10985 -16082 11001 -16048
rect 11045 -16082 11061 -16048
rect 11163 -16082 11179 -16048
rect 11223 -16082 11239 -16048
rect 11341 -16082 11357 -16048
rect 11401 -16082 11417 -16048
rect 11519 -16082 11535 -16048
rect 11579 -16082 11595 -16048
rect 11697 -16082 11713 -16048
rect 11757 -16082 11773 -16048
rect 11875 -16082 11891 -16048
rect 11935 -16082 11951 -16048
rect 12053 -16082 12069 -16048
rect 12113 -16082 12129 -16048
rect 12231 -16082 12247 -16048
rect 12291 -16082 12307 -16048
rect 12409 -16082 12425 -16048
rect 12469 -16082 12485 -16048
rect 12587 -16082 12603 -16048
rect 12647 -16082 12663 -16048
rect -5960 -16134 -5944 -16100
rect -5900 -16134 -5884 -16100
rect -5782 -16134 -5766 -16100
rect -5722 -16134 -5706 -16100
rect -5604 -16134 -5588 -16100
rect -5544 -16134 -5528 -16100
rect -5426 -16134 -5410 -16100
rect -5366 -16134 -5350 -16100
rect -5248 -16134 -5232 -16100
rect -5188 -16134 -5172 -16100
rect -5070 -16134 -5054 -16100
rect -5010 -16134 -4994 -16100
rect -4892 -16134 -4876 -16100
rect -4832 -16134 -4816 -16100
rect -4714 -16134 -4698 -16100
rect -4654 -16134 -4638 -16100
rect -4536 -16134 -4520 -16100
rect -4476 -16134 -4460 -16100
rect -4358 -16134 -4342 -16100
rect -4298 -16134 -4282 -16100
rect -4180 -16134 -4164 -16100
rect -4120 -16134 -4104 -16100
rect -2173 -16132 -2139 -16116
rect -2173 -16404 -2139 -16388
rect -1995 -16132 -1961 -16116
rect -1995 -16404 -1961 -16388
rect -1817 -16132 -1783 -16116
rect -1817 -16404 -1783 -16388
rect -1639 -16132 -1605 -16116
rect -1639 -16404 -1605 -16388
rect -1461 -16132 -1427 -16116
rect -1461 -16404 -1427 -16388
rect -1283 -16132 -1249 -16116
rect -1283 -16404 -1249 -16388
rect -1105 -16132 -1071 -16116
rect -1105 -16404 -1071 -16388
rect -927 -16132 -893 -16116
rect -927 -16404 -893 -16388
rect -749 -16132 -715 -16116
rect -749 -16404 -715 -16388
rect -571 -16132 -537 -16116
rect -571 -16404 -537 -16388
rect -393 -16132 -359 -16116
rect -393 -16404 -359 -16388
rect -215 -16132 -181 -16116
rect -215 -16404 -181 -16388
rect -37 -16132 -3 -16116
rect -37 -16404 -3 -16388
rect 141 -16132 175 -16116
rect 141 -16404 175 -16388
rect 319 -16132 353 -16116
rect 319 -16404 353 -16388
rect 497 -16132 531 -16116
rect 497 -16404 531 -16388
rect 675 -16132 709 -16116
rect 675 -16404 709 -16388
rect 853 -16132 887 -16116
rect 853 -16404 887 -16388
rect 1031 -16132 1065 -16116
rect 1031 -16404 1065 -16388
rect 1209 -16132 1243 -16116
rect 1209 -16404 1243 -16388
rect 1387 -16132 1421 -16116
rect 1387 -16404 1421 -16388
rect 1565 -16132 1599 -16116
rect 1565 -16404 1599 -16388
rect 1743 -16132 1777 -16116
rect 1743 -16404 1777 -16388
rect 1921 -16132 1955 -16116
rect 1921 -16404 1955 -16388
rect 2099 -16132 2133 -16116
rect 2099 -16404 2133 -16388
rect 2277 -16132 2311 -16116
rect 2277 -16404 2311 -16388
rect 2455 -16132 2489 -16116
rect 2455 -16404 2489 -16388
rect 2633 -16132 2667 -16116
rect 2633 -16404 2667 -16388
rect 2811 -16132 2845 -16116
rect 2811 -16404 2845 -16388
rect 2989 -16132 3023 -16116
rect 2989 -16404 3023 -16388
rect 3167 -16132 3201 -16116
rect 3167 -16404 3201 -16388
rect 3345 -16132 3379 -16116
rect 3345 -16404 3379 -16388
rect 3523 -16132 3557 -16116
rect 3523 -16404 3557 -16388
rect 3701 -16132 3735 -16116
rect 3701 -16404 3735 -16388
rect 3879 -16132 3913 -16116
rect 3879 -16404 3913 -16388
rect 4057 -16132 4091 -16116
rect 4057 -16404 4091 -16388
rect 5577 -16132 5611 -16116
rect 5577 -16404 5611 -16388
rect 5755 -16132 5789 -16116
rect 5755 -16404 5789 -16388
rect 5933 -16132 5967 -16116
rect 5933 -16404 5967 -16388
rect 6111 -16132 6145 -16116
rect 6111 -16404 6145 -16388
rect 6289 -16132 6323 -16116
rect 6289 -16404 6323 -16388
rect 6467 -16132 6501 -16116
rect 6467 -16404 6501 -16388
rect 6645 -16132 6679 -16116
rect 6645 -16404 6679 -16388
rect 6823 -16132 6857 -16116
rect 6823 -16404 6857 -16388
rect 7001 -16132 7035 -16116
rect 7001 -16404 7035 -16388
rect 7179 -16132 7213 -16116
rect 7179 -16404 7213 -16388
rect 7357 -16132 7391 -16116
rect 7357 -16404 7391 -16388
rect 7535 -16132 7569 -16116
rect 7535 -16404 7569 -16388
rect 7713 -16132 7747 -16116
rect 7713 -16404 7747 -16388
rect 7891 -16132 7925 -16116
rect 7891 -16404 7925 -16388
rect 8069 -16132 8103 -16116
rect 8069 -16404 8103 -16388
rect 8247 -16132 8281 -16116
rect 8247 -16404 8281 -16388
rect 8425 -16132 8459 -16116
rect 8425 -16404 8459 -16388
rect 8603 -16132 8637 -16116
rect 8603 -16404 8637 -16388
rect 8781 -16132 8815 -16116
rect 8781 -16404 8815 -16388
rect 8959 -16132 8993 -16116
rect 8959 -16404 8993 -16388
rect 9137 -16132 9171 -16116
rect 9137 -16404 9171 -16388
rect 9315 -16132 9349 -16116
rect 9315 -16404 9349 -16388
rect 9493 -16132 9527 -16116
rect 9493 -16404 9527 -16388
rect 9671 -16132 9705 -16116
rect 9671 -16404 9705 -16388
rect 9849 -16132 9883 -16116
rect 9849 -16404 9883 -16388
rect 10027 -16132 10061 -16116
rect 10027 -16404 10061 -16388
rect 10205 -16132 10239 -16116
rect 10205 -16404 10239 -16388
rect 10383 -16132 10417 -16116
rect 10383 -16404 10417 -16388
rect 10561 -16132 10595 -16116
rect 10561 -16404 10595 -16388
rect 10739 -16132 10773 -16116
rect 10739 -16404 10773 -16388
rect 10917 -16132 10951 -16116
rect 10917 -16404 10951 -16388
rect 11095 -16132 11129 -16116
rect 11095 -16404 11129 -16388
rect 11273 -16132 11307 -16116
rect 11273 -16404 11307 -16388
rect 11451 -16132 11485 -16116
rect 11451 -16404 11485 -16388
rect 11629 -16132 11663 -16116
rect 11629 -16404 11663 -16388
rect 11807 -16132 11841 -16116
rect 11807 -16404 11841 -16388
rect 11985 -16132 12019 -16116
rect 11985 -16404 12019 -16388
rect 12163 -16132 12197 -16116
rect 12163 -16404 12197 -16388
rect 12341 -16132 12375 -16116
rect 12341 -16404 12375 -16388
rect 12519 -16132 12553 -16116
rect 12519 -16404 12553 -16388
rect 12697 -16132 12731 -16116
rect 12697 -16404 12731 -16388
rect -5960 -16444 -5944 -16410
rect -5900 -16444 -5884 -16410
rect -5782 -16444 -5766 -16410
rect -5722 -16444 -5706 -16410
rect -5604 -16444 -5588 -16410
rect -5544 -16444 -5528 -16410
rect -5426 -16444 -5410 -16410
rect -5366 -16444 -5350 -16410
rect -5248 -16444 -5232 -16410
rect -5188 -16444 -5172 -16410
rect -5070 -16444 -5054 -16410
rect -5010 -16444 -4994 -16410
rect -4892 -16444 -4876 -16410
rect -4832 -16444 -4816 -16410
rect -4714 -16444 -4698 -16410
rect -4654 -16444 -4638 -16410
rect -4536 -16444 -4520 -16410
rect -4476 -16444 -4460 -16410
rect -4358 -16444 -4342 -16410
rect -4298 -16444 -4282 -16410
rect -4180 -16444 -4164 -16410
rect -4120 -16444 -4104 -16410
rect -2105 -16472 -2089 -16438
rect -2045 -16472 -2029 -16438
rect -1927 -16472 -1911 -16438
rect -1867 -16472 -1851 -16438
rect -1749 -16472 -1733 -16438
rect -1689 -16472 -1673 -16438
rect -1571 -16472 -1555 -16438
rect -1511 -16472 -1495 -16438
rect -1393 -16472 -1377 -16438
rect -1333 -16472 -1317 -16438
rect -1215 -16472 -1199 -16438
rect -1155 -16472 -1139 -16438
rect -1037 -16472 -1021 -16438
rect -977 -16472 -961 -16438
rect -859 -16472 -843 -16438
rect -799 -16472 -783 -16438
rect -681 -16472 -665 -16438
rect -621 -16472 -605 -16438
rect -503 -16472 -487 -16438
rect -443 -16472 -427 -16438
rect -325 -16472 -309 -16438
rect -265 -16472 -249 -16438
rect -147 -16472 -131 -16438
rect -87 -16472 -71 -16438
rect 31 -16472 47 -16438
rect 91 -16472 107 -16438
rect 209 -16472 225 -16438
rect 269 -16472 285 -16438
rect 387 -16472 403 -16438
rect 447 -16472 463 -16438
rect 565 -16472 581 -16438
rect 625 -16472 641 -16438
rect 743 -16472 759 -16438
rect 803 -16472 819 -16438
rect 921 -16472 937 -16438
rect 981 -16472 997 -16438
rect 1099 -16472 1115 -16438
rect 1159 -16472 1175 -16438
rect 1277 -16472 1293 -16438
rect 1337 -16472 1353 -16438
rect 1455 -16472 1471 -16438
rect 1515 -16472 1531 -16438
rect 1633 -16472 1649 -16438
rect 1693 -16472 1709 -16438
rect 1811 -16472 1827 -16438
rect 1871 -16472 1887 -16438
rect 1989 -16472 2005 -16438
rect 2049 -16472 2065 -16438
rect 2167 -16472 2183 -16438
rect 2227 -16472 2243 -16438
rect 2345 -16472 2361 -16438
rect 2405 -16472 2421 -16438
rect 2523 -16472 2539 -16438
rect 2583 -16472 2599 -16438
rect 2701 -16472 2717 -16438
rect 2761 -16472 2777 -16438
rect 2879 -16472 2895 -16438
rect 2939 -16472 2955 -16438
rect 3057 -16472 3073 -16438
rect 3117 -16472 3133 -16438
rect 3235 -16472 3251 -16438
rect 3295 -16472 3311 -16438
rect 3413 -16472 3429 -16438
rect 3473 -16472 3489 -16438
rect 3591 -16472 3607 -16438
rect 3651 -16472 3667 -16438
rect 3769 -16472 3785 -16438
rect 3829 -16472 3845 -16438
rect 3947 -16472 3963 -16438
rect 4007 -16472 4023 -16438
rect 5645 -16472 5661 -16438
rect 5705 -16472 5721 -16438
rect 5823 -16472 5839 -16438
rect 5883 -16472 5899 -16438
rect 6001 -16472 6017 -16438
rect 6061 -16472 6077 -16438
rect 6179 -16472 6195 -16438
rect 6239 -16472 6255 -16438
rect 6357 -16472 6373 -16438
rect 6417 -16472 6433 -16438
rect 6535 -16472 6551 -16438
rect 6595 -16472 6611 -16438
rect 6713 -16472 6729 -16438
rect 6773 -16472 6789 -16438
rect 6891 -16472 6907 -16438
rect 6951 -16472 6967 -16438
rect 7069 -16472 7085 -16438
rect 7129 -16472 7145 -16438
rect 7247 -16472 7263 -16438
rect 7307 -16472 7323 -16438
rect 7425 -16472 7441 -16438
rect 7485 -16472 7501 -16438
rect 7603 -16472 7619 -16438
rect 7663 -16472 7679 -16438
rect 7781 -16472 7797 -16438
rect 7841 -16472 7857 -16438
rect 7959 -16472 7975 -16438
rect 8019 -16472 8035 -16438
rect 8137 -16472 8153 -16438
rect 8197 -16472 8213 -16438
rect 8315 -16472 8331 -16438
rect 8375 -16472 8391 -16438
rect 8493 -16472 8509 -16438
rect 8553 -16472 8569 -16438
rect 8671 -16472 8687 -16438
rect 8731 -16472 8747 -16438
rect 8849 -16472 8865 -16438
rect 8909 -16472 8925 -16438
rect 9027 -16472 9043 -16438
rect 9087 -16472 9103 -16438
rect 9205 -16472 9221 -16438
rect 9265 -16472 9281 -16438
rect 9383 -16472 9399 -16438
rect 9443 -16472 9459 -16438
rect 9561 -16472 9577 -16438
rect 9621 -16472 9637 -16438
rect 9739 -16472 9755 -16438
rect 9799 -16472 9815 -16438
rect 9917 -16472 9933 -16438
rect 9977 -16472 9993 -16438
rect 10095 -16472 10111 -16438
rect 10155 -16472 10171 -16438
rect 10273 -16472 10289 -16438
rect 10333 -16472 10349 -16438
rect 10451 -16472 10467 -16438
rect 10511 -16472 10527 -16438
rect 10629 -16472 10645 -16438
rect 10689 -16472 10705 -16438
rect 10807 -16472 10823 -16438
rect 10867 -16472 10883 -16438
rect 10985 -16472 11001 -16438
rect 11045 -16472 11061 -16438
rect 11163 -16472 11179 -16438
rect 11223 -16472 11239 -16438
rect 11341 -16472 11357 -16438
rect 11401 -16472 11417 -16438
rect 11519 -16472 11535 -16438
rect 11579 -16472 11595 -16438
rect 11697 -16472 11713 -16438
rect 11757 -16472 11773 -16438
rect 11875 -16472 11891 -16438
rect 11935 -16472 11951 -16438
rect 12053 -16472 12069 -16438
rect 12113 -16472 12129 -16438
rect 12231 -16472 12247 -16438
rect 12291 -16472 12307 -16438
rect 12409 -16472 12425 -16438
rect 12469 -16472 12485 -16438
rect 12587 -16472 12603 -16438
rect 12647 -16472 12663 -16438
rect -6028 -16494 -5994 -16478
rect -6028 -16766 -5994 -16750
rect -5850 -16494 -5816 -16478
rect -5850 -16766 -5816 -16750
rect -5672 -16494 -5638 -16478
rect -5672 -16766 -5638 -16750
rect -5494 -16494 -5460 -16478
rect -5494 -16766 -5460 -16750
rect -5316 -16494 -5282 -16478
rect -5316 -16766 -5282 -16750
rect -5138 -16494 -5104 -16478
rect -5138 -16766 -5104 -16750
rect -4960 -16494 -4926 -16478
rect -4960 -16766 -4926 -16750
rect -4782 -16494 -4748 -16478
rect -4782 -16766 -4748 -16750
rect -4604 -16494 -4570 -16478
rect -4604 -16766 -4570 -16750
rect -4426 -16494 -4392 -16478
rect -4426 -16766 -4392 -16750
rect -4248 -16494 -4214 -16478
rect -4248 -16766 -4214 -16750
rect -4070 -16494 -4036 -16478
rect -4070 -16766 -4036 -16750
rect -5960 -16834 -5944 -16800
rect -5900 -16834 -5884 -16800
rect -5782 -16834 -5766 -16800
rect -5722 -16834 -5706 -16800
rect -5604 -16834 -5588 -16800
rect -5544 -16834 -5528 -16800
rect -5426 -16834 -5410 -16800
rect -5366 -16834 -5350 -16800
rect -5248 -16834 -5232 -16800
rect -5188 -16834 -5172 -16800
rect -5070 -16834 -5054 -16800
rect -5010 -16834 -4994 -16800
rect -4892 -16834 -4876 -16800
rect -4832 -16834 -4816 -16800
rect -4714 -16834 -4698 -16800
rect -4654 -16834 -4638 -16800
rect -4536 -16834 -4520 -16800
rect -4476 -16834 -4460 -16800
rect -4358 -16834 -4342 -16800
rect -4298 -16834 -4282 -16800
rect -4180 -16834 -4164 -16800
rect -4120 -16834 -4104 -16800
rect -7605 -17459 -7505 -17268
rect 13619 -17459 13719 -17149
rect -7605 -17559 -7323 -17459
rect 13384 -17559 13719 -17459
<< viali >>
rect -7379 -1353 3329 -1260
rect -6218 -2073 -6174 -2039
rect -6040 -2073 -5996 -2039
rect -5862 -2073 -5818 -2039
rect -5684 -2073 -5640 -2039
rect -5506 -2073 -5462 -2039
rect -5328 -2073 -5284 -2039
rect -5150 -2073 -5106 -2039
rect -4972 -2073 -4928 -2039
rect -4794 -2073 -4750 -2039
rect -4616 -2073 -4572 -2039
rect -4438 -2073 -4394 -2039
rect -4260 -2073 -4216 -2039
rect -4082 -2073 -4038 -2039
rect -3904 -2073 -3860 -2039
rect -3726 -2073 -3682 -2039
rect -3548 -2073 -3504 -2039
rect -6302 -2388 -6268 -2132
rect -6124 -2388 -6090 -2132
rect -5946 -2388 -5912 -2132
rect -5768 -2388 -5734 -2132
rect -5590 -2388 -5556 -2132
rect -5412 -2388 -5378 -2132
rect -5234 -2388 -5200 -2132
rect -5056 -2388 -5022 -2132
rect -4878 -2388 -4844 -2132
rect -4700 -2388 -4666 -2132
rect -4522 -2388 -4488 -2132
rect -4344 -2388 -4310 -2132
rect -4166 -2388 -4132 -2132
rect -3988 -2388 -3954 -2132
rect -3810 -2388 -3776 -2132
rect -3632 -2388 -3598 -2132
rect -3454 -2388 -3420 -2132
rect -6218 -2481 -6174 -2447
rect -6040 -2481 -5996 -2447
rect -5862 -2481 -5818 -2447
rect -5684 -2481 -5640 -2447
rect -5506 -2481 -5462 -2447
rect -5328 -2481 -5284 -2447
rect -5150 -2481 -5106 -2447
rect -4972 -2481 -4928 -2447
rect -4794 -2481 -4750 -2447
rect -4616 -2481 -4572 -2447
rect -4438 -2481 -4394 -2447
rect -4260 -2481 -4216 -2447
rect -4082 -2481 -4038 -2447
rect -3904 -2481 -3860 -2447
rect -3726 -2481 -3682 -2447
rect -3548 -2481 -3504 -2447
rect -1370 -2825 -1326 -2791
rect -1192 -2825 -1148 -2791
rect -1014 -2825 -970 -2791
rect -836 -2825 -792 -2791
rect -658 -2825 -614 -2791
rect -480 -2825 -436 -2791
rect -302 -2825 -258 -2791
rect -124 -2825 -80 -2791
rect 54 -2825 98 -2791
rect 232 -2825 276 -2791
rect 410 -2825 454 -2791
rect 588 -2825 632 -2791
rect 766 -2825 810 -2791
rect 944 -2825 988 -2791
rect 1122 -2825 1166 -2791
rect 1300 -2825 1344 -2791
rect 1478 -2825 1522 -2791
rect 1656 -2825 1700 -2791
rect 1834 -2825 1878 -2791
rect 2012 -2825 2056 -2791
rect 2190 -2825 2234 -2791
rect 2368 -2825 2412 -2791
rect 2546 -2825 2590 -2791
rect -6218 -2943 -6174 -2909
rect -6040 -2943 -5996 -2909
rect -5862 -2943 -5818 -2909
rect -5684 -2943 -5640 -2909
rect -5506 -2943 -5462 -2909
rect -5328 -2943 -5284 -2909
rect -5150 -2943 -5106 -2909
rect -4972 -2943 -4928 -2909
rect -4794 -2943 -4750 -2909
rect -4616 -2943 -4572 -2909
rect -4438 -2943 -4394 -2909
rect -4260 -2943 -4216 -2909
rect -4082 -2943 -4038 -2909
rect -3904 -2943 -3860 -2909
rect -3726 -2943 -3682 -2909
rect -3548 -2943 -3504 -2909
rect -6302 -3258 -6268 -3002
rect -6124 -3258 -6090 -3002
rect -5946 -3258 -5912 -3002
rect -5768 -3258 -5734 -3002
rect -5590 -3258 -5556 -3002
rect -5412 -3258 -5378 -3002
rect -5234 -3258 -5200 -3002
rect -5056 -3258 -5022 -3002
rect -4878 -3258 -4844 -3002
rect -4700 -3258 -4666 -3002
rect -4522 -3258 -4488 -3002
rect -4344 -3258 -4310 -3002
rect -4166 -3258 -4132 -3002
rect -3988 -3258 -3954 -3002
rect -3810 -3258 -3776 -3002
rect -3632 -3258 -3598 -3002
rect -3454 -3258 -3420 -3002
rect -1454 -3140 -1420 -2884
rect -1276 -3140 -1242 -2884
rect -1098 -3140 -1064 -2884
rect -920 -3140 -886 -2884
rect -742 -3140 -708 -2884
rect -564 -3140 -530 -2884
rect -386 -3140 -352 -2884
rect -208 -3140 -174 -2884
rect -30 -3140 4 -2884
rect 148 -3140 182 -2884
rect 326 -3140 360 -2884
rect 504 -3140 538 -2884
rect 682 -3140 716 -2884
rect 860 -3140 894 -2884
rect 1038 -3140 1072 -2884
rect 1216 -3140 1250 -2884
rect 1394 -3140 1428 -2884
rect 1572 -3140 1606 -2884
rect 1750 -3140 1784 -2884
rect 1928 -3140 1962 -2884
rect 2106 -3140 2140 -2884
rect 2284 -3140 2318 -2884
rect 2462 -3140 2496 -2884
rect 2640 -3140 2674 -2884
rect -1370 -3233 -1326 -3199
rect -1192 -3233 -1148 -3199
rect -1014 -3233 -970 -3199
rect -836 -3233 -792 -3199
rect -658 -3233 -614 -3199
rect -480 -3233 -436 -3199
rect -302 -3233 -258 -3199
rect -124 -3233 -80 -3199
rect 54 -3233 98 -3199
rect 232 -3233 276 -3199
rect 410 -3233 454 -3199
rect 588 -3233 632 -3199
rect 766 -3233 810 -3199
rect 944 -3233 988 -3199
rect 1122 -3233 1166 -3199
rect 1300 -3233 1344 -3199
rect 1478 -3233 1522 -3199
rect 1656 -3233 1700 -3199
rect 1834 -3233 1878 -3199
rect 2012 -3233 2056 -3199
rect 2190 -3233 2234 -3199
rect 2368 -3233 2412 -3199
rect 2546 -3233 2590 -3199
rect -6218 -3351 -6174 -3317
rect -6040 -3351 -5996 -3317
rect -5862 -3351 -5818 -3317
rect -5684 -3351 -5640 -3317
rect -5506 -3351 -5462 -3317
rect -5328 -3351 -5284 -3317
rect -5150 -3351 -5106 -3317
rect -4972 -3351 -4928 -3317
rect -4794 -3351 -4750 -3317
rect -4616 -3351 -4572 -3317
rect -4438 -3351 -4394 -3317
rect -4260 -3351 -4216 -3317
rect -4082 -3351 -4038 -3317
rect -3904 -3351 -3860 -3317
rect -3726 -3351 -3682 -3317
rect -3548 -3351 -3504 -3317
rect -1370 -3725 -1326 -3691
rect -1192 -3725 -1148 -3691
rect -1014 -3725 -970 -3691
rect -836 -3725 -792 -3691
rect -658 -3725 -614 -3691
rect -480 -3725 -436 -3691
rect -302 -3725 -258 -3691
rect -124 -3725 -80 -3691
rect 54 -3725 98 -3691
rect 232 -3725 276 -3691
rect 410 -3725 454 -3691
rect 588 -3725 632 -3691
rect 766 -3725 810 -3691
rect 944 -3725 988 -3691
rect 1122 -3725 1166 -3691
rect 1300 -3725 1344 -3691
rect 1478 -3725 1522 -3691
rect 1656 -3725 1700 -3691
rect 1834 -3725 1878 -3691
rect 2012 -3725 2056 -3691
rect 2190 -3725 2234 -3691
rect 2368 -3725 2412 -3691
rect 2546 -3725 2590 -3691
rect -6218 -3813 -6174 -3779
rect -6040 -3813 -5996 -3779
rect -5862 -3813 -5818 -3779
rect -5684 -3813 -5640 -3779
rect -5506 -3813 -5462 -3779
rect -5328 -3813 -5284 -3779
rect -5150 -3813 -5106 -3779
rect -4972 -3813 -4928 -3779
rect -4794 -3813 -4750 -3779
rect -4616 -3813 -4572 -3779
rect -4438 -3813 -4394 -3779
rect -4260 -3813 -4216 -3779
rect -4082 -3813 -4038 -3779
rect -3904 -3813 -3860 -3779
rect -3726 -3813 -3682 -3779
rect -3548 -3813 -3504 -3779
rect -6302 -4128 -6268 -3872
rect -6124 -4128 -6090 -3872
rect -5946 -4128 -5912 -3872
rect -5768 -4128 -5734 -3872
rect -5590 -4128 -5556 -3872
rect -5412 -4128 -5378 -3872
rect -5234 -4128 -5200 -3872
rect -5056 -4128 -5022 -3872
rect -4878 -4128 -4844 -3872
rect -4700 -4128 -4666 -3872
rect -4522 -4128 -4488 -3872
rect -4344 -4128 -4310 -3872
rect -4166 -4128 -4132 -3872
rect -3988 -4128 -3954 -3872
rect -3810 -4128 -3776 -3872
rect -3632 -4128 -3598 -3872
rect -3454 -4128 -3420 -3872
rect -1454 -4040 -1420 -3784
rect -1276 -4040 -1242 -3784
rect -1098 -4040 -1064 -3784
rect -920 -4040 -886 -3784
rect -742 -4040 -708 -3784
rect -564 -4040 -530 -3784
rect -386 -4040 -352 -3784
rect -208 -4040 -174 -3784
rect -30 -4040 4 -3784
rect 148 -4040 182 -3784
rect 326 -4040 360 -3784
rect 504 -4040 538 -3784
rect 682 -4040 716 -3784
rect 860 -4040 894 -3784
rect 1038 -4040 1072 -3784
rect 1216 -4040 1250 -3784
rect 1394 -4040 1428 -3784
rect 1572 -4040 1606 -3784
rect 1750 -4040 1784 -3784
rect 1928 -4040 1962 -3784
rect 2106 -4040 2140 -3784
rect 2284 -4040 2318 -3784
rect 2462 -4040 2496 -3784
rect 2640 -4040 2674 -3784
rect -1370 -4133 -1326 -4099
rect -1192 -4133 -1148 -4099
rect -1014 -4133 -970 -4099
rect -836 -4133 -792 -4099
rect -658 -4133 -614 -4099
rect -480 -4133 -436 -4099
rect -302 -4133 -258 -4099
rect -124 -4133 -80 -4099
rect 54 -4133 98 -4099
rect 232 -4133 276 -4099
rect 410 -4133 454 -4099
rect 588 -4133 632 -4099
rect 766 -4133 810 -4099
rect 944 -4133 988 -4099
rect 1122 -4133 1166 -4099
rect 1300 -4133 1344 -4099
rect 1478 -4133 1522 -4099
rect 1656 -4133 1700 -4099
rect 1834 -4133 1878 -4099
rect 2012 -4133 2056 -4099
rect 2190 -4133 2234 -4099
rect 2368 -4133 2412 -4099
rect 2546 -4133 2590 -4099
rect -6218 -4221 -6174 -4187
rect -6040 -4221 -5996 -4187
rect -5862 -4221 -5818 -4187
rect -5684 -4221 -5640 -4187
rect -5506 -4221 -5462 -4187
rect -5328 -4221 -5284 -4187
rect -5150 -4221 -5106 -4187
rect -4972 -4221 -4928 -4187
rect -4794 -4221 -4750 -4187
rect -4616 -4221 -4572 -4187
rect -4438 -4221 -4394 -4187
rect -4260 -4221 -4216 -4187
rect -4082 -4221 -4038 -4187
rect -3904 -4221 -3860 -4187
rect -3726 -4221 -3682 -4187
rect -3548 -4221 -3504 -4187
rect -1370 -4625 -1326 -4591
rect -1192 -4625 -1148 -4591
rect -1014 -4625 -970 -4591
rect -836 -4625 -792 -4591
rect -658 -4625 -614 -4591
rect -480 -4625 -436 -4591
rect -302 -4625 -258 -4591
rect -124 -4625 -80 -4591
rect 54 -4625 98 -4591
rect 232 -4625 276 -4591
rect 410 -4625 454 -4591
rect 588 -4625 632 -4591
rect 766 -4625 810 -4591
rect 944 -4625 988 -4591
rect 1122 -4625 1166 -4591
rect 1300 -4625 1344 -4591
rect 1478 -4625 1522 -4591
rect 1656 -4625 1700 -4591
rect 1834 -4625 1878 -4591
rect 2012 -4625 2056 -4591
rect 2190 -4625 2234 -4591
rect 2368 -4625 2412 -4591
rect 2546 -4625 2590 -4591
rect -6218 -4683 -6174 -4649
rect -6040 -4683 -5996 -4649
rect -5862 -4683 -5818 -4649
rect -5684 -4683 -5640 -4649
rect -5506 -4683 -5462 -4649
rect -5328 -4683 -5284 -4649
rect -5150 -4683 -5106 -4649
rect -4972 -4683 -4928 -4649
rect -4794 -4683 -4750 -4649
rect -4616 -4683 -4572 -4649
rect -4438 -4683 -4394 -4649
rect -4260 -4683 -4216 -4649
rect -4082 -4683 -4038 -4649
rect -3904 -4683 -3860 -4649
rect -3726 -4683 -3682 -4649
rect -3548 -4683 -3504 -4649
rect -6302 -4998 -6268 -4742
rect -6124 -4998 -6090 -4742
rect -5946 -4998 -5912 -4742
rect -5768 -4998 -5734 -4742
rect -5590 -4998 -5556 -4742
rect -5412 -4998 -5378 -4742
rect -5234 -4998 -5200 -4742
rect -5056 -4998 -5022 -4742
rect -4878 -4998 -4844 -4742
rect -4700 -4998 -4666 -4742
rect -4522 -4998 -4488 -4742
rect -4344 -4998 -4310 -4742
rect -4166 -4998 -4132 -4742
rect -3988 -4998 -3954 -4742
rect -3810 -4998 -3776 -4742
rect -3632 -4998 -3598 -4742
rect -3454 -4998 -3420 -4742
rect -1454 -4940 -1420 -4684
rect -1276 -4940 -1242 -4684
rect -1098 -4940 -1064 -4684
rect -920 -4940 -886 -4684
rect -742 -4940 -708 -4684
rect -564 -4940 -530 -4684
rect -386 -4940 -352 -4684
rect -208 -4940 -174 -4684
rect -30 -4940 4 -4684
rect 148 -4940 182 -4684
rect 326 -4940 360 -4684
rect 504 -4940 538 -4684
rect 682 -4940 716 -4684
rect 860 -4940 894 -4684
rect 1038 -4940 1072 -4684
rect 1216 -4940 1250 -4684
rect 1394 -4940 1428 -4684
rect 1572 -4940 1606 -4684
rect 1750 -4940 1784 -4684
rect 1928 -4940 1962 -4684
rect 2106 -4940 2140 -4684
rect 2284 -4940 2318 -4684
rect 2462 -4940 2496 -4684
rect 2640 -4940 2674 -4684
rect -1370 -5033 -1326 -4999
rect -1192 -5033 -1148 -4999
rect -1014 -5033 -970 -4999
rect -836 -5033 -792 -4999
rect -658 -5033 -614 -4999
rect -480 -5033 -436 -4999
rect -302 -5033 -258 -4999
rect -124 -5033 -80 -4999
rect 54 -5033 98 -4999
rect 232 -5033 276 -4999
rect 410 -5033 454 -4999
rect 588 -5033 632 -4999
rect 766 -5033 810 -4999
rect 944 -5033 988 -4999
rect 1122 -5033 1166 -4999
rect 1300 -5033 1344 -4999
rect 1478 -5033 1522 -4999
rect 1656 -5033 1700 -4999
rect 1834 -5033 1878 -4999
rect 2012 -5033 2056 -4999
rect 2190 -5033 2234 -4999
rect 2368 -5033 2412 -4999
rect 2546 -5033 2590 -4999
rect -6218 -5091 -6174 -5057
rect -6040 -5091 -5996 -5057
rect -5862 -5091 -5818 -5057
rect -5684 -5091 -5640 -5057
rect -5506 -5091 -5462 -5057
rect -5328 -5091 -5284 -5057
rect -5150 -5091 -5106 -5057
rect -4972 -5091 -4928 -5057
rect -4794 -5091 -4750 -5057
rect -4616 -5091 -4572 -5057
rect -4438 -5091 -4394 -5057
rect -4260 -5091 -4216 -5057
rect -4082 -5091 -4038 -5057
rect -3904 -5091 -3860 -5057
rect -3726 -5091 -3682 -5057
rect -3548 -5091 -3504 -5057
rect -6218 -5553 -6174 -5519
rect -6040 -5553 -5996 -5519
rect -5862 -5553 -5818 -5519
rect -5684 -5553 -5640 -5519
rect -5506 -5553 -5462 -5519
rect -5328 -5553 -5284 -5519
rect -5150 -5553 -5106 -5519
rect -4972 -5553 -4928 -5519
rect -4794 -5553 -4750 -5519
rect -4616 -5553 -4572 -5519
rect -4438 -5553 -4394 -5519
rect -4260 -5553 -4216 -5519
rect -4082 -5553 -4038 -5519
rect -3904 -5553 -3860 -5519
rect -3726 -5553 -3682 -5519
rect -3548 -5553 -3504 -5519
rect -1370 -5525 -1326 -5491
rect -1192 -5525 -1148 -5491
rect -1014 -5525 -970 -5491
rect -836 -5525 -792 -5491
rect -658 -5525 -614 -5491
rect -480 -5525 -436 -5491
rect -302 -5525 -258 -5491
rect -124 -5525 -80 -5491
rect 54 -5525 98 -5491
rect 232 -5525 276 -5491
rect 410 -5525 454 -5491
rect 588 -5525 632 -5491
rect 766 -5525 810 -5491
rect 944 -5525 988 -5491
rect 1122 -5525 1166 -5491
rect 1300 -5525 1344 -5491
rect 1478 -5525 1522 -5491
rect 1656 -5525 1700 -5491
rect 1834 -5525 1878 -5491
rect 2012 -5525 2056 -5491
rect 2190 -5525 2234 -5491
rect 2368 -5525 2412 -5491
rect 2546 -5525 2590 -5491
rect -6302 -5868 -6268 -5612
rect -6124 -5868 -6090 -5612
rect -5946 -5868 -5912 -5612
rect -5768 -5868 -5734 -5612
rect -5590 -5868 -5556 -5612
rect -5412 -5868 -5378 -5612
rect -5234 -5868 -5200 -5612
rect -5056 -5868 -5022 -5612
rect -4878 -5868 -4844 -5612
rect -4700 -5868 -4666 -5612
rect -4522 -5868 -4488 -5612
rect -4344 -5868 -4310 -5612
rect -4166 -5868 -4132 -5612
rect -3988 -5868 -3954 -5612
rect -3810 -5868 -3776 -5612
rect -3632 -5868 -3598 -5612
rect -3454 -5868 -3420 -5612
rect -1454 -5840 -1420 -5584
rect -1276 -5840 -1242 -5584
rect -1098 -5840 -1064 -5584
rect -920 -5840 -886 -5584
rect -742 -5840 -708 -5584
rect -564 -5840 -530 -5584
rect -386 -5840 -352 -5584
rect -208 -5840 -174 -5584
rect -30 -5840 4 -5584
rect 148 -5840 182 -5584
rect 326 -5840 360 -5584
rect 504 -5840 538 -5584
rect 682 -5840 716 -5584
rect 860 -5840 894 -5584
rect 1038 -5840 1072 -5584
rect 1216 -5840 1250 -5584
rect 1394 -5840 1428 -5584
rect 1572 -5840 1606 -5584
rect 1750 -5840 1784 -5584
rect 1928 -5840 1962 -5584
rect 2106 -5840 2140 -5584
rect 2284 -5840 2318 -5584
rect 2462 -5840 2496 -5584
rect 2640 -5840 2674 -5584
rect -6218 -5961 -6174 -5927
rect -6040 -5961 -5996 -5927
rect -5862 -5961 -5818 -5927
rect -5684 -5961 -5640 -5927
rect -5506 -5961 -5462 -5927
rect -5328 -5961 -5284 -5927
rect -5150 -5961 -5106 -5927
rect -4972 -5961 -4928 -5927
rect -4794 -5961 -4750 -5927
rect -4616 -5961 -4572 -5927
rect -4438 -5961 -4394 -5927
rect -4260 -5961 -4216 -5927
rect -4082 -5961 -4038 -5927
rect -3904 -5961 -3860 -5927
rect -3726 -5961 -3682 -5927
rect -3548 -5961 -3504 -5927
rect -1370 -5933 -1326 -5899
rect -1192 -5933 -1148 -5899
rect -1014 -5933 -970 -5899
rect -836 -5933 -792 -5899
rect -658 -5933 -614 -5899
rect -480 -5933 -436 -5899
rect -302 -5933 -258 -5899
rect -124 -5933 -80 -5899
rect 54 -5933 98 -5899
rect 232 -5933 276 -5899
rect 410 -5933 454 -5899
rect 588 -5933 632 -5899
rect 766 -5933 810 -5899
rect 944 -5933 988 -5899
rect 1122 -5933 1166 -5899
rect 1300 -5933 1344 -5899
rect 1478 -5933 1522 -5899
rect 1656 -5933 1700 -5899
rect 1834 -5933 1878 -5899
rect 2012 -5933 2056 -5899
rect 2190 -5933 2234 -5899
rect 2368 -5933 2412 -5899
rect 2546 -5933 2590 -5899
rect -5544 -7824 -5500 -7790
rect -5366 -7824 -5322 -7790
rect -5188 -7824 -5144 -7790
rect -5010 -7824 -4966 -7790
rect -4832 -7824 -4788 -7790
rect -4654 -7824 -4610 -7790
rect -4476 -7824 -4432 -7790
rect -4298 -7824 -4254 -7790
rect -4120 -7824 -4076 -7790
rect -5628 -8130 -5594 -7874
rect -5450 -8130 -5416 -7874
rect -5272 -8130 -5238 -7874
rect -5094 -8130 -5060 -7874
rect -4916 -8130 -4882 -7874
rect -4738 -8130 -4704 -7874
rect -4560 -8130 -4526 -7874
rect -4382 -8130 -4348 -7874
rect -4204 -8130 -4170 -7874
rect -4026 -8130 -3992 -7874
rect -2089 -8082 -2045 -8048
rect -1911 -8082 -1867 -8048
rect -1733 -8082 -1689 -8048
rect -1555 -8082 -1511 -8048
rect -1377 -8082 -1333 -8048
rect -1199 -8082 -1155 -8048
rect -1021 -8082 -977 -8048
rect -843 -8082 -799 -8048
rect -665 -8082 -621 -8048
rect -487 -8082 -443 -8048
rect -309 -8082 -265 -8048
rect -131 -8082 -87 -8048
rect 47 -8082 91 -8048
rect 225 -8082 269 -8048
rect 403 -8082 447 -8048
rect 581 -8082 625 -8048
rect 759 -8082 803 -8048
rect 937 -8082 981 -8048
rect 1115 -8082 1159 -8048
rect 1293 -8082 1337 -8048
rect 1471 -8082 1515 -8048
rect 1649 -8082 1693 -8048
rect 1827 -8082 1871 -8048
rect 2005 -8082 2049 -8048
rect 2183 -8082 2227 -8048
rect 2361 -8082 2405 -8048
rect 2539 -8082 2583 -8048
rect 2717 -8082 2761 -8048
rect 2895 -8082 2939 -8048
rect 3073 -8082 3117 -8048
rect 3251 -8082 3295 -8048
rect 3429 -8082 3473 -8048
rect 3607 -8082 3651 -8048
rect 3785 -8082 3829 -8048
rect 3963 -8082 4007 -8048
rect -5544 -8214 -5500 -8180
rect -5366 -8214 -5322 -8180
rect -5188 -8214 -5144 -8180
rect -5010 -8214 -4966 -8180
rect -4832 -8214 -4788 -8180
rect -4654 -8214 -4610 -8180
rect -4476 -8214 -4432 -8180
rect -4298 -8214 -4254 -8180
rect -4120 -8214 -4076 -8180
rect -5544 -8374 -5500 -8340
rect -5366 -8374 -5322 -8340
rect -5188 -8374 -5144 -8340
rect -5010 -8374 -4966 -8340
rect -4832 -8374 -4788 -8340
rect -4654 -8374 -4610 -8340
rect -4476 -8374 -4432 -8340
rect -4298 -8374 -4254 -8340
rect -4120 -8374 -4076 -8340
rect -2173 -8388 -2139 -8132
rect -1995 -8388 -1961 -8132
rect -1817 -8388 -1783 -8132
rect -1639 -8388 -1605 -8132
rect -1461 -8388 -1427 -8132
rect -1283 -8388 -1249 -8132
rect -1105 -8388 -1071 -8132
rect -927 -8388 -893 -8132
rect -749 -8388 -715 -8132
rect -571 -8388 -537 -8132
rect -393 -8388 -359 -8132
rect -215 -8388 -181 -8132
rect -37 -8388 -3 -8132
rect 141 -8388 175 -8132
rect 319 -8388 353 -8132
rect 497 -8388 531 -8132
rect 675 -8388 709 -8132
rect 853 -8388 887 -8132
rect 1031 -8388 1065 -8132
rect 1209 -8388 1243 -8132
rect 1387 -8388 1421 -8132
rect 1565 -8388 1599 -8132
rect 1743 -8388 1777 -8132
rect 1921 -8388 1955 -8132
rect 2099 -8388 2133 -8132
rect 2277 -8388 2311 -8132
rect 2455 -8388 2489 -8132
rect 2633 -8388 2667 -8132
rect 2811 -8388 2845 -8132
rect 2989 -8388 3023 -8132
rect 3167 -8388 3201 -8132
rect 3345 -8388 3379 -8132
rect 3523 -8388 3557 -8132
rect 3701 -8388 3735 -8132
rect 3879 -8388 3913 -8132
rect 4057 -8388 4091 -8132
rect -5628 -8680 -5594 -8424
rect -5450 -8680 -5416 -8424
rect -5272 -8680 -5238 -8424
rect -5094 -8680 -5060 -8424
rect -4916 -8680 -4882 -8424
rect -4738 -8680 -4704 -8424
rect -4560 -8680 -4526 -8424
rect -4382 -8680 -4348 -8424
rect -4204 -8680 -4170 -8424
rect -4026 -8680 -3992 -8424
rect -2089 -8472 -2045 -8438
rect -1911 -8472 -1867 -8438
rect -1733 -8472 -1689 -8438
rect -1555 -8472 -1511 -8438
rect -1377 -8472 -1333 -8438
rect -1199 -8472 -1155 -8438
rect -1021 -8472 -977 -8438
rect -843 -8472 -799 -8438
rect -665 -8472 -621 -8438
rect -487 -8472 -443 -8438
rect -309 -8472 -265 -8438
rect -131 -8472 -87 -8438
rect 47 -8472 91 -8438
rect 225 -8472 269 -8438
rect 403 -8472 447 -8438
rect 581 -8472 625 -8438
rect 759 -8472 803 -8438
rect 937 -8472 981 -8438
rect 1115 -8472 1159 -8438
rect 1293 -8472 1337 -8438
rect 1471 -8472 1515 -8438
rect 1649 -8472 1693 -8438
rect 1827 -8472 1871 -8438
rect 2005 -8472 2049 -8438
rect 2183 -8472 2227 -8438
rect 2361 -8472 2405 -8438
rect 2539 -8472 2583 -8438
rect 2717 -8472 2761 -8438
rect 2895 -8472 2939 -8438
rect 3073 -8472 3117 -8438
rect 3251 -8472 3295 -8438
rect 3429 -8472 3473 -8438
rect 3607 -8472 3651 -8438
rect 3785 -8472 3829 -8438
rect 3963 -8472 4007 -8438
rect -5544 -8764 -5500 -8730
rect -5366 -8764 -5322 -8730
rect -5188 -8764 -5144 -8730
rect -5010 -8764 -4966 -8730
rect -4832 -8764 -4788 -8730
rect -4654 -8764 -4610 -8730
rect -4476 -8764 -4432 -8730
rect -4298 -8764 -4254 -8730
rect -4120 -8764 -4076 -8730
rect 6596 -8844 6640 -8810
rect 6774 -8844 6818 -8810
rect 6952 -8844 6996 -8810
rect 7130 -8844 7174 -8810
rect 7308 -8844 7352 -8810
rect 7486 -8844 7530 -8810
rect 7664 -8844 7708 -8810
rect 7842 -8844 7886 -8810
rect 8020 -8844 8064 -8810
rect 8198 -8844 8242 -8810
rect 8376 -8844 8420 -8810
rect 8554 -8844 8598 -8810
rect 8732 -8844 8776 -8810
rect 8910 -8844 8954 -8810
rect 9088 -8844 9132 -8810
rect 9266 -8844 9310 -8810
rect 10856 -8874 10900 -8840
rect 11148 -8874 11192 -8840
rect 11440 -8874 11484 -8840
rect 11732 -8874 11776 -8840
rect 12024 -8874 12068 -8840
rect 12316 -8874 12360 -8840
rect 12608 -8874 12652 -8840
rect -5544 -8924 -5500 -8890
rect -5366 -8924 -5322 -8890
rect -5188 -8924 -5144 -8890
rect -5010 -8924 -4966 -8890
rect -4832 -8924 -4788 -8890
rect -4654 -8924 -4610 -8890
rect -4476 -8924 -4432 -8890
rect -4298 -8924 -4254 -8890
rect -4120 -8924 -4076 -8890
rect -5628 -9230 -5594 -8974
rect -5450 -9230 -5416 -8974
rect -5272 -9230 -5238 -8974
rect -5094 -9230 -5060 -8974
rect -4916 -9230 -4882 -8974
rect -4738 -9230 -4704 -8974
rect -4560 -9230 -4526 -8974
rect -4382 -9230 -4348 -8974
rect -4204 -9230 -4170 -8974
rect -4026 -9230 -3992 -8974
rect -2089 -9082 -2045 -9048
rect -1911 -9082 -1867 -9048
rect -1733 -9082 -1689 -9048
rect -1555 -9082 -1511 -9048
rect -1377 -9082 -1333 -9048
rect -1199 -9082 -1155 -9048
rect -1021 -9082 -977 -9048
rect -843 -9082 -799 -9048
rect -665 -9082 -621 -9048
rect -487 -9082 -443 -9048
rect -309 -9082 -265 -9048
rect -131 -9082 -87 -9048
rect 47 -9082 91 -9048
rect 225 -9082 269 -9048
rect 403 -9082 447 -9048
rect 581 -9082 625 -9048
rect 759 -9082 803 -9048
rect 937 -9082 981 -9048
rect 1115 -9082 1159 -9048
rect 1293 -9082 1337 -9048
rect 1471 -9082 1515 -9048
rect 1649 -9082 1693 -9048
rect 1827 -9082 1871 -9048
rect 2005 -9082 2049 -9048
rect 2183 -9082 2227 -9048
rect 2361 -9082 2405 -9048
rect 2539 -9082 2583 -9048
rect 2717 -9082 2761 -9048
rect 2895 -9082 2939 -9048
rect 3073 -9082 3117 -9048
rect 3251 -9082 3295 -9048
rect 3429 -9082 3473 -9048
rect 3607 -9082 3651 -9048
rect 3785 -9082 3829 -9048
rect 3963 -9082 4007 -9048
rect -5544 -9314 -5500 -9280
rect -5366 -9314 -5322 -9280
rect -5188 -9314 -5144 -9280
rect -5010 -9314 -4966 -9280
rect -4832 -9314 -4788 -9280
rect -4654 -9314 -4610 -9280
rect -4476 -9314 -4432 -9280
rect -4298 -9314 -4254 -9280
rect -4120 -9314 -4076 -9280
rect -2173 -9388 -2139 -9132
rect -1995 -9388 -1961 -9132
rect -1817 -9388 -1783 -9132
rect -1639 -9388 -1605 -9132
rect -1461 -9388 -1427 -9132
rect -1283 -9388 -1249 -9132
rect -1105 -9388 -1071 -9132
rect -927 -9388 -893 -9132
rect -749 -9388 -715 -9132
rect -571 -9388 -537 -9132
rect -393 -9388 -359 -9132
rect -215 -9388 -181 -9132
rect -37 -9388 -3 -9132
rect 141 -9388 175 -9132
rect 319 -9388 353 -9132
rect 497 -9388 531 -9132
rect 675 -9388 709 -9132
rect 853 -9388 887 -9132
rect 1031 -9388 1065 -9132
rect 1209 -9388 1243 -9132
rect 1387 -9388 1421 -9132
rect 1565 -9388 1599 -9132
rect 1743 -9388 1777 -9132
rect 1921 -9388 1955 -9132
rect 2099 -9388 2133 -9132
rect 2277 -9388 2311 -9132
rect 2455 -9388 2489 -9132
rect 2633 -9388 2667 -9132
rect 2811 -9388 2845 -9132
rect 2989 -9388 3023 -9132
rect 3167 -9388 3201 -9132
rect 3345 -9388 3379 -9132
rect 3523 -9388 3557 -9132
rect 3701 -9388 3735 -9132
rect 3879 -9388 3913 -9132
rect 4057 -9388 4091 -9132
rect 6512 -9150 6546 -8894
rect 6690 -9150 6724 -8894
rect 6868 -9150 6902 -8894
rect 7046 -9150 7080 -8894
rect 7224 -9150 7258 -8894
rect 7402 -9150 7436 -8894
rect 7580 -9150 7614 -8894
rect 7758 -9150 7792 -8894
rect 7936 -9150 7970 -8894
rect 8114 -9150 8148 -8894
rect 8292 -9150 8326 -8894
rect 8470 -9150 8504 -8894
rect 8648 -9150 8682 -8894
rect 8826 -9150 8860 -8894
rect 9004 -9150 9038 -8894
rect 9182 -9150 9216 -8894
rect 9360 -9150 9394 -8894
rect 10772 -9180 10806 -8924
rect 10950 -9180 10984 -8924
rect 11064 -9180 11098 -8924
rect 11242 -9180 11276 -8924
rect 11356 -9180 11390 -8924
rect 11534 -9180 11568 -8924
rect 11648 -9180 11682 -8924
rect 11826 -9180 11860 -8924
rect 11940 -9180 11974 -8924
rect 12118 -9180 12152 -8924
rect 12232 -9180 12266 -8924
rect 12410 -9180 12444 -8924
rect 12524 -9180 12558 -8924
rect 12702 -9180 12736 -8924
rect 6596 -9234 6640 -9200
rect 6774 -9234 6818 -9200
rect 6952 -9234 6996 -9200
rect 7130 -9234 7174 -9200
rect 7308 -9234 7352 -9200
rect 7486 -9234 7530 -9200
rect 7664 -9234 7708 -9200
rect 7842 -9234 7886 -9200
rect 8020 -9234 8064 -9200
rect 8198 -9234 8242 -9200
rect 8376 -9234 8420 -9200
rect 8554 -9234 8598 -9200
rect 8732 -9234 8776 -9200
rect 8910 -9234 8954 -9200
rect 9088 -9234 9132 -9200
rect 9266 -9234 9310 -9200
rect 10856 -9264 10900 -9230
rect 11148 -9264 11192 -9230
rect 11440 -9264 11484 -9230
rect 11732 -9264 11776 -9230
rect 12024 -9264 12068 -9230
rect 12316 -9264 12360 -9230
rect 12608 -9264 12652 -9230
rect -5544 -9474 -5500 -9440
rect -5366 -9474 -5322 -9440
rect -5188 -9474 -5144 -9440
rect -5010 -9474 -4966 -9440
rect -4832 -9474 -4788 -9440
rect -4654 -9474 -4610 -9440
rect -4476 -9474 -4432 -9440
rect -4298 -9474 -4254 -9440
rect -4120 -9474 -4076 -9440
rect -2089 -9472 -2045 -9438
rect -1911 -9472 -1867 -9438
rect -1733 -9472 -1689 -9438
rect -1555 -9472 -1511 -9438
rect -1377 -9472 -1333 -9438
rect -1199 -9472 -1155 -9438
rect -1021 -9472 -977 -9438
rect -843 -9472 -799 -9438
rect -665 -9472 -621 -9438
rect -487 -9472 -443 -9438
rect -309 -9472 -265 -9438
rect -131 -9472 -87 -9438
rect 47 -9472 91 -9438
rect 225 -9472 269 -9438
rect 403 -9472 447 -9438
rect 581 -9472 625 -9438
rect 759 -9472 803 -9438
rect 937 -9472 981 -9438
rect 1115 -9472 1159 -9438
rect 1293 -9472 1337 -9438
rect 1471 -9472 1515 -9438
rect 1649 -9472 1693 -9438
rect 1827 -9472 1871 -9438
rect 2005 -9472 2049 -9438
rect 2183 -9472 2227 -9438
rect 2361 -9472 2405 -9438
rect 2539 -9472 2583 -9438
rect 2717 -9472 2761 -9438
rect 2895 -9472 2939 -9438
rect 3073 -9472 3117 -9438
rect 3251 -9472 3295 -9438
rect 3429 -9472 3473 -9438
rect 3607 -9472 3651 -9438
rect 3785 -9472 3829 -9438
rect 3963 -9472 4007 -9438
rect -5628 -9780 -5594 -9524
rect -5450 -9780 -5416 -9524
rect -5272 -9780 -5238 -9524
rect -5094 -9780 -5060 -9524
rect -4916 -9780 -4882 -9524
rect -4738 -9780 -4704 -9524
rect -4560 -9780 -4526 -9524
rect -4382 -9780 -4348 -9524
rect -4204 -9780 -4170 -9524
rect -4026 -9780 -3992 -9524
rect 10856 -9644 10900 -9610
rect 11148 -9644 11192 -9610
rect 11440 -9644 11484 -9610
rect 11732 -9644 11776 -9610
rect 12024 -9644 12068 -9610
rect 12316 -9644 12360 -9610
rect 12608 -9644 12652 -9610
rect 6596 -9744 6640 -9710
rect 6774 -9744 6818 -9710
rect 6952 -9744 6996 -9710
rect 7130 -9744 7174 -9710
rect 7308 -9744 7352 -9710
rect 7486 -9744 7530 -9710
rect 7664 -9744 7708 -9710
rect 7842 -9744 7886 -9710
rect 8020 -9744 8064 -9710
rect 8198 -9744 8242 -9710
rect 8376 -9744 8420 -9710
rect 8554 -9744 8598 -9710
rect 8732 -9744 8776 -9710
rect 8910 -9744 8954 -9710
rect 9088 -9744 9132 -9710
rect 9266 -9744 9310 -9710
rect -5544 -9864 -5500 -9830
rect -5366 -9864 -5322 -9830
rect -5188 -9864 -5144 -9830
rect -5010 -9864 -4966 -9830
rect -4832 -9864 -4788 -9830
rect -4654 -9864 -4610 -9830
rect -4476 -9864 -4432 -9830
rect -4298 -9864 -4254 -9830
rect -4120 -9864 -4076 -9830
rect -5544 -10024 -5500 -9990
rect -5366 -10024 -5322 -9990
rect -5188 -10024 -5144 -9990
rect -5010 -10024 -4966 -9990
rect -4832 -10024 -4788 -9990
rect -4654 -10024 -4610 -9990
rect -4476 -10024 -4432 -9990
rect -4298 -10024 -4254 -9990
rect -4120 -10024 -4076 -9990
rect -5628 -10330 -5594 -10074
rect -5450 -10330 -5416 -10074
rect -5272 -10330 -5238 -10074
rect -5094 -10330 -5060 -10074
rect -4916 -10330 -4882 -10074
rect -4738 -10330 -4704 -10074
rect -4560 -10330 -4526 -10074
rect -4382 -10330 -4348 -10074
rect -4204 -10330 -4170 -10074
rect -4026 -10330 -3992 -10074
rect -2089 -10082 -2045 -10048
rect -1911 -10082 -1867 -10048
rect -1733 -10082 -1689 -10048
rect -1555 -10082 -1511 -10048
rect -1377 -10082 -1333 -10048
rect -1199 -10082 -1155 -10048
rect -1021 -10082 -977 -10048
rect -843 -10082 -799 -10048
rect -665 -10082 -621 -10048
rect -487 -10082 -443 -10048
rect -309 -10082 -265 -10048
rect -131 -10082 -87 -10048
rect 47 -10082 91 -10048
rect 225 -10082 269 -10048
rect 403 -10082 447 -10048
rect 581 -10082 625 -10048
rect 759 -10082 803 -10048
rect 937 -10082 981 -10048
rect 1115 -10082 1159 -10048
rect 1293 -10082 1337 -10048
rect 1471 -10082 1515 -10048
rect 1649 -10082 1693 -10048
rect 1827 -10082 1871 -10048
rect 2005 -10082 2049 -10048
rect 2183 -10082 2227 -10048
rect 2361 -10082 2405 -10048
rect 2539 -10082 2583 -10048
rect 2717 -10082 2761 -10048
rect 2895 -10082 2939 -10048
rect 3073 -10082 3117 -10048
rect 3251 -10082 3295 -10048
rect 3429 -10082 3473 -10048
rect 3607 -10082 3651 -10048
rect 3785 -10082 3829 -10048
rect 3963 -10082 4007 -10048
rect 6512 -10050 6546 -9794
rect 6690 -10050 6724 -9794
rect 6868 -10050 6902 -9794
rect 7046 -10050 7080 -9794
rect 7224 -10050 7258 -9794
rect 7402 -10050 7436 -9794
rect 7580 -10050 7614 -9794
rect 7758 -10050 7792 -9794
rect 7936 -10050 7970 -9794
rect 8114 -10050 8148 -9794
rect 8292 -10050 8326 -9794
rect 8470 -10050 8504 -9794
rect 8648 -10050 8682 -9794
rect 8826 -10050 8860 -9794
rect 9004 -10050 9038 -9794
rect 9182 -10050 9216 -9794
rect 9360 -10050 9394 -9794
rect 10772 -9950 10806 -9694
rect 10950 -9950 10984 -9694
rect 11064 -9950 11098 -9694
rect 11242 -9950 11276 -9694
rect 11356 -9950 11390 -9694
rect 11534 -9950 11568 -9694
rect 11648 -9950 11682 -9694
rect 11826 -9950 11860 -9694
rect 11940 -9950 11974 -9694
rect 12118 -9950 12152 -9694
rect 12232 -9950 12266 -9694
rect 12410 -9950 12444 -9694
rect 12524 -9950 12558 -9694
rect 12702 -9950 12736 -9694
rect 10856 -10034 10900 -10000
rect 11148 -10034 11192 -10000
rect 11440 -10034 11484 -10000
rect 11732 -10034 11776 -10000
rect 12024 -10034 12068 -10000
rect 12316 -10034 12360 -10000
rect 12608 -10034 12652 -10000
rect -5544 -10414 -5500 -10380
rect -5366 -10414 -5322 -10380
rect -5188 -10414 -5144 -10380
rect -5010 -10414 -4966 -10380
rect -4832 -10414 -4788 -10380
rect -4654 -10414 -4610 -10380
rect -4476 -10414 -4432 -10380
rect -4298 -10414 -4254 -10380
rect -4120 -10414 -4076 -10380
rect -2173 -10388 -2139 -10132
rect -1995 -10388 -1961 -10132
rect -1817 -10388 -1783 -10132
rect -1639 -10388 -1605 -10132
rect -1461 -10388 -1427 -10132
rect -1283 -10388 -1249 -10132
rect -1105 -10388 -1071 -10132
rect -927 -10388 -893 -10132
rect -749 -10388 -715 -10132
rect -571 -10388 -537 -10132
rect -393 -10388 -359 -10132
rect -215 -10388 -181 -10132
rect -37 -10388 -3 -10132
rect 141 -10388 175 -10132
rect 319 -10388 353 -10132
rect 497 -10388 531 -10132
rect 675 -10388 709 -10132
rect 853 -10388 887 -10132
rect 1031 -10388 1065 -10132
rect 1209 -10388 1243 -10132
rect 1387 -10388 1421 -10132
rect 1565 -10388 1599 -10132
rect 1743 -10388 1777 -10132
rect 1921 -10388 1955 -10132
rect 2099 -10388 2133 -10132
rect 2277 -10388 2311 -10132
rect 2455 -10388 2489 -10132
rect 2633 -10388 2667 -10132
rect 2811 -10388 2845 -10132
rect 2989 -10388 3023 -10132
rect 3167 -10388 3201 -10132
rect 3345 -10388 3379 -10132
rect 3523 -10388 3557 -10132
rect 3701 -10388 3735 -10132
rect 3879 -10388 3913 -10132
rect 4057 -10388 4091 -10132
rect 6596 -10134 6640 -10100
rect 6774 -10134 6818 -10100
rect 6952 -10134 6996 -10100
rect 7130 -10134 7174 -10100
rect 7308 -10134 7352 -10100
rect 7486 -10134 7530 -10100
rect 7664 -10134 7708 -10100
rect 7842 -10134 7886 -10100
rect 8020 -10134 8064 -10100
rect 8198 -10134 8242 -10100
rect 8376 -10134 8420 -10100
rect 8554 -10134 8598 -10100
rect 8732 -10134 8776 -10100
rect 8910 -10134 8954 -10100
rect 9088 -10134 9132 -10100
rect 9266 -10134 9310 -10100
rect 10856 -10414 10900 -10380
rect 11148 -10414 11192 -10380
rect 11440 -10414 11484 -10380
rect 11732 -10414 11776 -10380
rect 12024 -10414 12068 -10380
rect 12316 -10414 12360 -10380
rect 12608 -10414 12652 -10380
rect -2089 -10472 -2045 -10438
rect -1911 -10472 -1867 -10438
rect -1733 -10472 -1689 -10438
rect -1555 -10472 -1511 -10438
rect -1377 -10472 -1333 -10438
rect -1199 -10472 -1155 -10438
rect -1021 -10472 -977 -10438
rect -843 -10472 -799 -10438
rect -665 -10472 -621 -10438
rect -487 -10472 -443 -10438
rect -309 -10472 -265 -10438
rect -131 -10472 -87 -10438
rect 47 -10472 91 -10438
rect 225 -10472 269 -10438
rect 403 -10472 447 -10438
rect 581 -10472 625 -10438
rect 759 -10472 803 -10438
rect 937 -10472 981 -10438
rect 1115 -10472 1159 -10438
rect 1293 -10472 1337 -10438
rect 1471 -10472 1515 -10438
rect 1649 -10472 1693 -10438
rect 1827 -10472 1871 -10438
rect 2005 -10472 2049 -10438
rect 2183 -10472 2227 -10438
rect 2361 -10472 2405 -10438
rect 2539 -10472 2583 -10438
rect 2717 -10472 2761 -10438
rect 2895 -10472 2939 -10438
rect 3073 -10472 3117 -10438
rect 3251 -10472 3295 -10438
rect 3429 -10472 3473 -10438
rect 3607 -10472 3651 -10438
rect 3785 -10472 3829 -10438
rect 3963 -10472 4007 -10438
rect -5544 -10574 -5500 -10540
rect -5366 -10574 -5322 -10540
rect -5188 -10574 -5144 -10540
rect -5010 -10574 -4966 -10540
rect -4832 -10574 -4788 -10540
rect -4654 -10574 -4610 -10540
rect -4476 -10574 -4432 -10540
rect -4298 -10574 -4254 -10540
rect -4120 -10574 -4076 -10540
rect -5628 -10880 -5594 -10624
rect -5450 -10880 -5416 -10624
rect -5272 -10880 -5238 -10624
rect -5094 -10880 -5060 -10624
rect -4916 -10880 -4882 -10624
rect -4738 -10880 -4704 -10624
rect -4560 -10880 -4526 -10624
rect -4382 -10880 -4348 -10624
rect -4204 -10880 -4170 -10624
rect -4026 -10880 -3992 -10624
rect 6596 -10644 6640 -10610
rect 6774 -10644 6818 -10610
rect 6952 -10644 6996 -10610
rect 7130 -10644 7174 -10610
rect 7308 -10644 7352 -10610
rect 7486 -10644 7530 -10610
rect 7664 -10644 7708 -10610
rect 7842 -10644 7886 -10610
rect 8020 -10644 8064 -10610
rect 8198 -10644 8242 -10610
rect 8376 -10644 8420 -10610
rect 8554 -10644 8598 -10610
rect 8732 -10644 8776 -10610
rect 8910 -10644 8954 -10610
rect 9088 -10644 9132 -10610
rect 9266 -10644 9310 -10610
rect -5544 -10964 -5500 -10930
rect -5366 -10964 -5322 -10930
rect -5188 -10964 -5144 -10930
rect -5010 -10964 -4966 -10930
rect -4832 -10964 -4788 -10930
rect -4654 -10964 -4610 -10930
rect -4476 -10964 -4432 -10930
rect -4298 -10964 -4254 -10930
rect -4120 -10964 -4076 -10930
rect 6512 -10950 6546 -10694
rect 6690 -10950 6724 -10694
rect 6868 -10950 6902 -10694
rect 7046 -10950 7080 -10694
rect 7224 -10950 7258 -10694
rect 7402 -10950 7436 -10694
rect 7580 -10950 7614 -10694
rect 7758 -10950 7792 -10694
rect 7936 -10950 7970 -10694
rect 8114 -10950 8148 -10694
rect 8292 -10950 8326 -10694
rect 8470 -10950 8504 -10694
rect 8648 -10950 8682 -10694
rect 8826 -10950 8860 -10694
rect 9004 -10950 9038 -10694
rect 9182 -10950 9216 -10694
rect 9360 -10950 9394 -10694
rect 10772 -10720 10806 -10464
rect 10950 -10720 10984 -10464
rect 11064 -10720 11098 -10464
rect 11242 -10720 11276 -10464
rect 11356 -10720 11390 -10464
rect 11534 -10720 11568 -10464
rect 11648 -10720 11682 -10464
rect 11826 -10720 11860 -10464
rect 11940 -10720 11974 -10464
rect 12118 -10720 12152 -10464
rect 12232 -10720 12266 -10464
rect 12410 -10720 12444 -10464
rect 12524 -10720 12558 -10464
rect 12702 -10720 12736 -10464
rect 10856 -10804 10900 -10770
rect 11148 -10804 11192 -10770
rect 11440 -10804 11484 -10770
rect 11732 -10804 11776 -10770
rect 12024 -10804 12068 -10770
rect 12316 -10804 12360 -10770
rect 12608 -10804 12652 -10770
rect 6596 -11034 6640 -11000
rect 6774 -11034 6818 -11000
rect 6952 -11034 6996 -11000
rect 7130 -11034 7174 -11000
rect 7308 -11034 7352 -11000
rect 7486 -11034 7530 -11000
rect 7664 -11034 7708 -11000
rect 7842 -11034 7886 -11000
rect 8020 -11034 8064 -11000
rect 8198 -11034 8242 -11000
rect 8376 -11034 8420 -11000
rect 8554 -11034 8598 -11000
rect 8732 -11034 8776 -11000
rect 8910 -11034 8954 -11000
rect 9088 -11034 9132 -11000
rect 9266 -11034 9310 -11000
rect -2089 -11082 -2045 -11048
rect -1911 -11082 -1867 -11048
rect -1733 -11082 -1689 -11048
rect -1555 -11082 -1511 -11048
rect -1377 -11082 -1333 -11048
rect -1199 -11082 -1155 -11048
rect -1021 -11082 -977 -11048
rect -843 -11082 -799 -11048
rect -665 -11082 -621 -11048
rect -487 -11082 -443 -11048
rect -309 -11082 -265 -11048
rect -131 -11082 -87 -11048
rect 47 -11082 91 -11048
rect 225 -11082 269 -11048
rect 403 -11082 447 -11048
rect 581 -11082 625 -11048
rect 759 -11082 803 -11048
rect 937 -11082 981 -11048
rect 1115 -11082 1159 -11048
rect 1293 -11082 1337 -11048
rect 1471 -11082 1515 -11048
rect 1649 -11082 1693 -11048
rect 1827 -11082 1871 -11048
rect 2005 -11082 2049 -11048
rect 2183 -11082 2227 -11048
rect 2361 -11082 2405 -11048
rect 2539 -11082 2583 -11048
rect 2717 -11082 2761 -11048
rect 2895 -11082 2939 -11048
rect 3073 -11082 3117 -11048
rect 3251 -11082 3295 -11048
rect 3429 -11082 3473 -11048
rect 3607 -11082 3651 -11048
rect 3785 -11082 3829 -11048
rect 3963 -11082 4007 -11048
rect -5544 -11124 -5500 -11090
rect -5366 -11124 -5322 -11090
rect -5188 -11124 -5144 -11090
rect -5010 -11124 -4966 -11090
rect -4832 -11124 -4788 -11090
rect -4654 -11124 -4610 -11090
rect -4476 -11124 -4432 -11090
rect -4298 -11124 -4254 -11090
rect -4120 -11124 -4076 -11090
rect -5628 -11430 -5594 -11174
rect -5450 -11430 -5416 -11174
rect -5272 -11430 -5238 -11174
rect -5094 -11430 -5060 -11174
rect -4916 -11430 -4882 -11174
rect -4738 -11430 -4704 -11174
rect -4560 -11430 -4526 -11174
rect -4382 -11430 -4348 -11174
rect -4204 -11430 -4170 -11174
rect -4026 -11430 -3992 -11174
rect -2173 -11388 -2139 -11132
rect -1995 -11388 -1961 -11132
rect -1817 -11388 -1783 -11132
rect -1639 -11388 -1605 -11132
rect -1461 -11388 -1427 -11132
rect -1283 -11388 -1249 -11132
rect -1105 -11388 -1071 -11132
rect -927 -11388 -893 -11132
rect -749 -11388 -715 -11132
rect -571 -11388 -537 -11132
rect -393 -11388 -359 -11132
rect -215 -11388 -181 -11132
rect -37 -11388 -3 -11132
rect 141 -11388 175 -11132
rect 319 -11388 353 -11132
rect 497 -11388 531 -11132
rect 675 -11388 709 -11132
rect 853 -11388 887 -11132
rect 1031 -11388 1065 -11132
rect 1209 -11388 1243 -11132
rect 1387 -11388 1421 -11132
rect 1565 -11388 1599 -11132
rect 1743 -11388 1777 -11132
rect 1921 -11388 1955 -11132
rect 2099 -11388 2133 -11132
rect 2277 -11388 2311 -11132
rect 2455 -11388 2489 -11132
rect 2633 -11388 2667 -11132
rect 2811 -11388 2845 -11132
rect 2989 -11388 3023 -11132
rect 3167 -11388 3201 -11132
rect 3345 -11388 3379 -11132
rect 3523 -11388 3557 -11132
rect 3701 -11388 3735 -11132
rect 3879 -11388 3913 -11132
rect 4057 -11388 4091 -11132
rect 10856 -11184 10900 -11150
rect 11148 -11184 11192 -11150
rect 11440 -11184 11484 -11150
rect 11732 -11184 11776 -11150
rect 12024 -11184 12068 -11150
rect 12316 -11184 12360 -11150
rect 12608 -11184 12652 -11150
rect -2089 -11472 -2045 -11438
rect -1911 -11472 -1867 -11438
rect -1733 -11472 -1689 -11438
rect -1555 -11472 -1511 -11438
rect -1377 -11472 -1333 -11438
rect -1199 -11472 -1155 -11438
rect -1021 -11472 -977 -11438
rect -843 -11472 -799 -11438
rect -665 -11472 -621 -11438
rect -487 -11472 -443 -11438
rect -309 -11472 -265 -11438
rect -131 -11472 -87 -11438
rect 47 -11472 91 -11438
rect 225 -11472 269 -11438
rect 403 -11472 447 -11438
rect 581 -11472 625 -11438
rect 759 -11472 803 -11438
rect 937 -11472 981 -11438
rect 1115 -11472 1159 -11438
rect 1293 -11472 1337 -11438
rect 1471 -11472 1515 -11438
rect 1649 -11472 1693 -11438
rect 1827 -11472 1871 -11438
rect 2005 -11472 2049 -11438
rect 2183 -11472 2227 -11438
rect 2361 -11472 2405 -11438
rect 2539 -11472 2583 -11438
rect 2717 -11472 2761 -11438
rect 2895 -11472 2939 -11438
rect 3073 -11472 3117 -11438
rect 3251 -11472 3295 -11438
rect 3429 -11472 3473 -11438
rect 3607 -11472 3651 -11438
rect 3785 -11472 3829 -11438
rect 3963 -11472 4007 -11438
rect -5544 -11514 -5500 -11480
rect -5366 -11514 -5322 -11480
rect -5188 -11514 -5144 -11480
rect -5010 -11514 -4966 -11480
rect -4832 -11514 -4788 -11480
rect -4654 -11514 -4610 -11480
rect -4476 -11514 -4432 -11480
rect -4298 -11514 -4254 -11480
rect -4120 -11514 -4076 -11480
rect 10772 -11490 10806 -11234
rect 10950 -11490 10984 -11234
rect 11064 -11490 11098 -11234
rect 11242 -11490 11276 -11234
rect 11356 -11490 11390 -11234
rect 11534 -11490 11568 -11234
rect 11648 -11490 11682 -11234
rect 11826 -11490 11860 -11234
rect 11940 -11490 11974 -11234
rect 12118 -11490 12152 -11234
rect 12232 -11490 12266 -11234
rect 12410 -11490 12444 -11234
rect 12524 -11490 12558 -11234
rect 12702 -11490 12736 -11234
rect 6596 -11544 6640 -11510
rect 6774 -11544 6818 -11510
rect 6952 -11544 6996 -11510
rect 7130 -11544 7174 -11510
rect 7308 -11544 7352 -11510
rect 7486 -11544 7530 -11510
rect 7664 -11544 7708 -11510
rect 7842 -11544 7886 -11510
rect 8020 -11544 8064 -11510
rect 8198 -11544 8242 -11510
rect 8376 -11544 8420 -11510
rect 8554 -11544 8598 -11510
rect 8732 -11544 8776 -11510
rect 8910 -11544 8954 -11510
rect 9088 -11544 9132 -11510
rect 9266 -11544 9310 -11510
rect 10856 -11574 10900 -11540
rect 11148 -11574 11192 -11540
rect 11440 -11574 11484 -11540
rect 11732 -11574 11776 -11540
rect 12024 -11574 12068 -11540
rect 12316 -11574 12360 -11540
rect 12608 -11574 12652 -11540
rect -5544 -11674 -5500 -11640
rect -5366 -11674 -5322 -11640
rect -5188 -11674 -5144 -11640
rect -5010 -11674 -4966 -11640
rect -4832 -11674 -4788 -11640
rect -4654 -11674 -4610 -11640
rect -4476 -11674 -4432 -11640
rect -4298 -11674 -4254 -11640
rect -4120 -11674 -4076 -11640
rect -5628 -11980 -5594 -11724
rect -5450 -11980 -5416 -11724
rect -5272 -11980 -5238 -11724
rect -5094 -11980 -5060 -11724
rect -4916 -11980 -4882 -11724
rect -4738 -11980 -4704 -11724
rect -4560 -11980 -4526 -11724
rect -4382 -11980 -4348 -11724
rect -4204 -11980 -4170 -11724
rect -4026 -11980 -3992 -11724
rect 6512 -11850 6546 -11594
rect 6690 -11850 6724 -11594
rect 6868 -11850 6902 -11594
rect 7046 -11850 7080 -11594
rect 7224 -11850 7258 -11594
rect 7402 -11850 7436 -11594
rect 7580 -11850 7614 -11594
rect 7758 -11850 7792 -11594
rect 7936 -11850 7970 -11594
rect 8114 -11850 8148 -11594
rect 8292 -11850 8326 -11594
rect 8470 -11850 8504 -11594
rect 8648 -11850 8682 -11594
rect 8826 -11850 8860 -11594
rect 9004 -11850 9038 -11594
rect 9182 -11850 9216 -11594
rect 9360 -11850 9394 -11594
rect 6596 -11934 6640 -11900
rect 6774 -11934 6818 -11900
rect 6952 -11934 6996 -11900
rect 7130 -11934 7174 -11900
rect 7308 -11934 7352 -11900
rect 7486 -11934 7530 -11900
rect 7664 -11934 7708 -11900
rect 7842 -11934 7886 -11900
rect 8020 -11934 8064 -11900
rect 8198 -11934 8242 -11900
rect 8376 -11934 8420 -11900
rect 8554 -11934 8598 -11900
rect 8732 -11934 8776 -11900
rect 8910 -11934 8954 -11900
rect 9088 -11934 9132 -11900
rect 9266 -11934 9310 -11900
rect -5544 -12064 -5500 -12030
rect -5366 -12064 -5322 -12030
rect -5188 -12064 -5144 -12030
rect -5010 -12064 -4966 -12030
rect -4832 -12064 -4788 -12030
rect -4654 -12064 -4610 -12030
rect -4476 -12064 -4432 -12030
rect -4298 -12064 -4254 -12030
rect -4120 -12064 -4076 -12030
rect -2089 -12082 -2045 -12048
rect -1911 -12082 -1867 -12048
rect -1733 -12082 -1689 -12048
rect -1555 -12082 -1511 -12048
rect -1377 -12082 -1333 -12048
rect -1199 -12082 -1155 -12048
rect -1021 -12082 -977 -12048
rect -843 -12082 -799 -12048
rect -665 -12082 -621 -12048
rect -487 -12082 -443 -12048
rect -309 -12082 -265 -12048
rect -131 -12082 -87 -12048
rect 47 -12082 91 -12048
rect 225 -12082 269 -12048
rect 403 -12082 447 -12048
rect 581 -12082 625 -12048
rect 759 -12082 803 -12048
rect 937 -12082 981 -12048
rect 1115 -12082 1159 -12048
rect 1293 -12082 1337 -12048
rect 1471 -12082 1515 -12048
rect 1649 -12082 1693 -12048
rect 1827 -12082 1871 -12048
rect 2005 -12082 2049 -12048
rect 2183 -12082 2227 -12048
rect 2361 -12082 2405 -12048
rect 2539 -12082 2583 -12048
rect 2717 -12082 2761 -12048
rect 2895 -12082 2939 -12048
rect 3073 -12082 3117 -12048
rect 3251 -12082 3295 -12048
rect 3429 -12082 3473 -12048
rect 3607 -12082 3651 -12048
rect 3785 -12082 3829 -12048
rect 3963 -12082 4007 -12048
rect -2173 -12388 -2139 -12132
rect -1995 -12388 -1961 -12132
rect -1817 -12388 -1783 -12132
rect -1639 -12388 -1605 -12132
rect -1461 -12388 -1427 -12132
rect -1283 -12388 -1249 -12132
rect -1105 -12388 -1071 -12132
rect -927 -12388 -893 -12132
rect -749 -12388 -715 -12132
rect -571 -12388 -537 -12132
rect -393 -12388 -359 -12132
rect -215 -12388 -181 -12132
rect -37 -12388 -3 -12132
rect 141 -12388 175 -12132
rect 319 -12388 353 -12132
rect 497 -12388 531 -12132
rect 675 -12388 709 -12132
rect 853 -12388 887 -12132
rect 1031 -12388 1065 -12132
rect 1209 -12388 1243 -12132
rect 1387 -12388 1421 -12132
rect 1565 -12388 1599 -12132
rect 1743 -12388 1777 -12132
rect 1921 -12388 1955 -12132
rect 2099 -12388 2133 -12132
rect 2277 -12388 2311 -12132
rect 2455 -12388 2489 -12132
rect 2633 -12388 2667 -12132
rect 2811 -12388 2845 -12132
rect 2989 -12388 3023 -12132
rect 3167 -12388 3201 -12132
rect 3345 -12388 3379 -12132
rect 3523 -12388 3557 -12132
rect 3701 -12388 3735 -12132
rect 3879 -12388 3913 -12132
rect 4057 -12388 4091 -12132
rect -2089 -12472 -2045 -12438
rect -1911 -12472 -1867 -12438
rect -1733 -12472 -1689 -12438
rect -1555 -12472 -1511 -12438
rect -1377 -12472 -1333 -12438
rect -1199 -12472 -1155 -12438
rect -1021 -12472 -977 -12438
rect -843 -12472 -799 -12438
rect -665 -12472 -621 -12438
rect -487 -12472 -443 -12438
rect -309 -12472 -265 -12438
rect -131 -12472 -87 -12438
rect 47 -12472 91 -12438
rect 225 -12472 269 -12438
rect 403 -12472 447 -12438
rect 581 -12472 625 -12438
rect 759 -12472 803 -12438
rect 937 -12472 981 -12438
rect 1115 -12472 1159 -12438
rect 1293 -12472 1337 -12438
rect 1471 -12472 1515 -12438
rect 1649 -12472 1693 -12438
rect 1827 -12472 1871 -12438
rect 2005 -12472 2049 -12438
rect 2183 -12472 2227 -12438
rect 2361 -12472 2405 -12438
rect 2539 -12472 2583 -12438
rect 2717 -12472 2761 -12438
rect 2895 -12472 2939 -12438
rect 3073 -12472 3117 -12438
rect 3251 -12472 3295 -12438
rect 3429 -12472 3473 -12438
rect 3607 -12472 3651 -12438
rect 3785 -12472 3829 -12438
rect 3963 -12472 4007 -12438
rect -5867 -12662 -5833 -12628
rect -5617 -12662 -5583 -12628
rect -5367 -12662 -5333 -12628
rect -5117 -12662 -5083 -12628
rect -4867 -12662 -4833 -12628
rect -4617 -12662 -4583 -12628
rect -4367 -12662 -4333 -12628
rect -4117 -12662 -4083 -12628
rect -5916 -12928 -5882 -12712
rect -5818 -12928 -5784 -12712
rect -5666 -12928 -5632 -12712
rect -5568 -12928 -5534 -12712
rect -5416 -12928 -5382 -12712
rect -5318 -12928 -5284 -12712
rect -5166 -12928 -5132 -12712
rect -5068 -12928 -5034 -12712
rect -4916 -12928 -4882 -12712
rect -4818 -12928 -4784 -12712
rect -4666 -12928 -4632 -12712
rect -4568 -12928 -4534 -12712
rect -4416 -12928 -4382 -12712
rect -4318 -12928 -4284 -12712
rect -4166 -12928 -4132 -12712
rect -4068 -12928 -4034 -12712
rect -5867 -13012 -5833 -12978
rect -5617 -13012 -5583 -12978
rect -5367 -13012 -5333 -12978
rect -5117 -13012 -5083 -12978
rect -4867 -13012 -4833 -12978
rect -4617 -13012 -4583 -12978
rect -4367 -13012 -4333 -12978
rect -4117 -13012 -4083 -12978
rect -2089 -13082 -2045 -13048
rect -1911 -13082 -1867 -13048
rect -1733 -13082 -1689 -13048
rect -1555 -13082 -1511 -13048
rect -1377 -13082 -1333 -13048
rect -1199 -13082 -1155 -13048
rect -1021 -13082 -977 -13048
rect -843 -13082 -799 -13048
rect -665 -13082 -621 -13048
rect -487 -13082 -443 -13048
rect -309 -13082 -265 -13048
rect -131 -13082 -87 -13048
rect 47 -13082 91 -13048
rect 225 -13082 269 -13048
rect 403 -13082 447 -13048
rect 581 -13082 625 -13048
rect 759 -13082 803 -13048
rect 937 -13082 981 -13048
rect 1115 -13082 1159 -13048
rect 1293 -13082 1337 -13048
rect 1471 -13082 1515 -13048
rect 1649 -13082 1693 -13048
rect 1827 -13082 1871 -13048
rect 2005 -13082 2049 -13048
rect 2183 -13082 2227 -13048
rect 2361 -13082 2405 -13048
rect 2539 -13082 2583 -13048
rect 2717 -13082 2761 -13048
rect 2895 -13082 2939 -13048
rect 3073 -13082 3117 -13048
rect 3251 -13082 3295 -13048
rect 3429 -13082 3473 -13048
rect 3607 -13082 3651 -13048
rect 3785 -13082 3829 -13048
rect 3963 -13082 4007 -13048
rect -5867 -13342 -5833 -13308
rect -5617 -13342 -5583 -13308
rect -5367 -13342 -5333 -13308
rect -5117 -13342 -5083 -13308
rect -4867 -13342 -4833 -13308
rect -4617 -13342 -4583 -13308
rect -4367 -13342 -4333 -13308
rect -4117 -13342 -4083 -13308
rect -5916 -13608 -5882 -13392
rect -5818 -13608 -5784 -13392
rect -5666 -13608 -5632 -13392
rect -5568 -13608 -5534 -13392
rect -5416 -13608 -5382 -13392
rect -5318 -13608 -5284 -13392
rect -5166 -13608 -5132 -13392
rect -5068 -13608 -5034 -13392
rect -4916 -13608 -4882 -13392
rect -4818 -13608 -4784 -13392
rect -4666 -13608 -4632 -13392
rect -4568 -13608 -4534 -13392
rect -4416 -13608 -4382 -13392
rect -4318 -13608 -4284 -13392
rect -4166 -13608 -4132 -13392
rect -4068 -13608 -4034 -13392
rect -2173 -13388 -2139 -13132
rect -1995 -13388 -1961 -13132
rect -1817 -13388 -1783 -13132
rect -1639 -13388 -1605 -13132
rect -1461 -13388 -1427 -13132
rect -1283 -13388 -1249 -13132
rect -1105 -13388 -1071 -13132
rect -927 -13388 -893 -13132
rect -749 -13388 -715 -13132
rect -571 -13388 -537 -13132
rect -393 -13388 -359 -13132
rect -215 -13388 -181 -13132
rect -37 -13388 -3 -13132
rect 141 -13388 175 -13132
rect 319 -13388 353 -13132
rect 497 -13388 531 -13132
rect 675 -13388 709 -13132
rect 853 -13388 887 -13132
rect 1031 -13388 1065 -13132
rect 1209 -13388 1243 -13132
rect 1387 -13388 1421 -13132
rect 1565 -13388 1599 -13132
rect 1743 -13388 1777 -13132
rect 1921 -13388 1955 -13132
rect 2099 -13388 2133 -13132
rect 2277 -13388 2311 -13132
rect 2455 -13388 2489 -13132
rect 2633 -13388 2667 -13132
rect 2811 -13388 2845 -13132
rect 2989 -13388 3023 -13132
rect 3167 -13388 3201 -13132
rect 3345 -13388 3379 -13132
rect 3523 -13388 3557 -13132
rect 3701 -13388 3735 -13132
rect 3879 -13388 3913 -13132
rect 4057 -13388 4091 -13132
rect -2089 -13472 -2045 -13438
rect -1911 -13472 -1867 -13438
rect -1733 -13472 -1689 -13438
rect -1555 -13472 -1511 -13438
rect -1377 -13472 -1333 -13438
rect -1199 -13472 -1155 -13438
rect -1021 -13472 -977 -13438
rect -843 -13472 -799 -13438
rect -665 -13472 -621 -13438
rect -487 -13472 -443 -13438
rect -309 -13472 -265 -13438
rect -131 -13472 -87 -13438
rect 47 -13472 91 -13438
rect 225 -13472 269 -13438
rect 403 -13472 447 -13438
rect 581 -13472 625 -13438
rect 759 -13472 803 -13438
rect 937 -13472 981 -13438
rect 1115 -13472 1159 -13438
rect 1293 -13472 1337 -13438
rect 1471 -13472 1515 -13438
rect 1649 -13472 1693 -13438
rect 1827 -13472 1871 -13438
rect 2005 -13472 2049 -13438
rect 2183 -13472 2227 -13438
rect 2361 -13472 2405 -13438
rect 2539 -13472 2583 -13438
rect 2717 -13472 2761 -13438
rect 2895 -13472 2939 -13438
rect 3073 -13472 3117 -13438
rect 3251 -13472 3295 -13438
rect 3429 -13472 3473 -13438
rect 3607 -13472 3651 -13438
rect 3785 -13472 3829 -13438
rect 3963 -13472 4007 -13438
rect -5867 -13692 -5833 -13658
rect -5617 -13692 -5583 -13658
rect -5367 -13692 -5333 -13658
rect -5117 -13692 -5083 -13658
rect -4867 -13692 -4833 -13658
rect -4617 -13692 -4583 -13658
rect -4367 -13692 -4333 -13658
rect -4117 -13692 -4083 -13658
rect -2089 -14082 -2045 -14048
rect -1911 -14082 -1867 -14048
rect -1733 -14082 -1689 -14048
rect -1555 -14082 -1511 -14048
rect -1377 -14082 -1333 -14048
rect -1199 -14082 -1155 -14048
rect -1021 -14082 -977 -14048
rect -843 -14082 -799 -14048
rect -665 -14082 -621 -14048
rect -487 -14082 -443 -14048
rect -309 -14082 -265 -14048
rect -131 -14082 -87 -14048
rect 47 -14082 91 -14048
rect 225 -14082 269 -14048
rect 403 -14082 447 -14048
rect 581 -14082 625 -14048
rect 759 -14082 803 -14048
rect 937 -14082 981 -14048
rect 1115 -14082 1159 -14048
rect 1293 -14082 1337 -14048
rect 1471 -14082 1515 -14048
rect 1649 -14082 1693 -14048
rect 1827 -14082 1871 -14048
rect 2005 -14082 2049 -14048
rect 2183 -14082 2227 -14048
rect 2361 -14082 2405 -14048
rect 2539 -14082 2583 -14048
rect 2717 -14082 2761 -14048
rect 2895 -14082 2939 -14048
rect 3073 -14082 3117 -14048
rect 3251 -14082 3295 -14048
rect 3429 -14082 3473 -14048
rect 3607 -14082 3651 -14048
rect 3785 -14082 3829 -14048
rect 3963 -14082 4007 -14048
rect 5661 -14082 5705 -14048
rect 5839 -14082 5883 -14048
rect 6017 -14082 6061 -14048
rect 6195 -14082 6239 -14048
rect 6373 -14082 6417 -14048
rect 6551 -14082 6595 -14048
rect 6729 -14082 6773 -14048
rect 6907 -14082 6951 -14048
rect 7085 -14082 7129 -14048
rect 7263 -14082 7307 -14048
rect 7441 -14082 7485 -14048
rect 7619 -14082 7663 -14048
rect 7797 -14082 7841 -14048
rect 7975 -14082 8019 -14048
rect 8153 -14082 8197 -14048
rect 8331 -14082 8375 -14048
rect 8509 -14082 8553 -14048
rect 8687 -14082 8731 -14048
rect 8865 -14082 8909 -14048
rect 9043 -14082 9087 -14048
rect 9221 -14082 9265 -14048
rect 9399 -14082 9443 -14048
rect 9577 -14082 9621 -14048
rect 9755 -14082 9799 -14048
rect 9933 -14082 9977 -14048
rect 10111 -14082 10155 -14048
rect 10289 -14082 10333 -14048
rect 10467 -14082 10511 -14048
rect 10645 -14082 10689 -14048
rect 10823 -14082 10867 -14048
rect 11001 -14082 11045 -14048
rect 11179 -14082 11223 -14048
rect 11357 -14082 11401 -14048
rect 11535 -14082 11579 -14048
rect 11713 -14082 11757 -14048
rect 11891 -14082 11935 -14048
rect 12069 -14082 12113 -14048
rect 12247 -14082 12291 -14048
rect 12425 -14082 12469 -14048
rect 12603 -14082 12647 -14048
rect -5944 -14344 -5900 -14310
rect -5766 -14344 -5722 -14310
rect -5588 -14344 -5544 -14310
rect -5410 -14344 -5366 -14310
rect -5232 -14344 -5188 -14310
rect -5054 -14344 -5010 -14310
rect -4876 -14344 -4832 -14310
rect -4698 -14344 -4654 -14310
rect -4520 -14344 -4476 -14310
rect -4342 -14344 -4298 -14310
rect -4164 -14344 -4120 -14310
rect -6028 -14650 -5994 -14394
rect -5850 -14650 -5816 -14394
rect -5672 -14650 -5638 -14394
rect -5494 -14650 -5460 -14394
rect -5316 -14650 -5282 -14394
rect -5138 -14650 -5104 -14394
rect -4960 -14650 -4926 -14394
rect -4782 -14650 -4748 -14394
rect -4604 -14650 -4570 -14394
rect -4426 -14650 -4392 -14394
rect -4248 -14650 -4214 -14394
rect -4070 -14650 -4036 -14394
rect -2173 -14388 -2139 -14132
rect -1995 -14388 -1961 -14132
rect -1817 -14388 -1783 -14132
rect -1639 -14388 -1605 -14132
rect -1461 -14388 -1427 -14132
rect -1283 -14388 -1249 -14132
rect -1105 -14388 -1071 -14132
rect -927 -14388 -893 -14132
rect -749 -14388 -715 -14132
rect -571 -14388 -537 -14132
rect -393 -14388 -359 -14132
rect -215 -14388 -181 -14132
rect -37 -14388 -3 -14132
rect 141 -14388 175 -14132
rect 319 -14388 353 -14132
rect 497 -14388 531 -14132
rect 675 -14388 709 -14132
rect 853 -14388 887 -14132
rect 1031 -14388 1065 -14132
rect 1209 -14388 1243 -14132
rect 1387 -14388 1421 -14132
rect 1565 -14388 1599 -14132
rect 1743 -14388 1777 -14132
rect 1921 -14388 1955 -14132
rect 2099 -14388 2133 -14132
rect 2277 -14388 2311 -14132
rect 2455 -14388 2489 -14132
rect 2633 -14388 2667 -14132
rect 2811 -14388 2845 -14132
rect 2989 -14388 3023 -14132
rect 3167 -14388 3201 -14132
rect 3345 -14388 3379 -14132
rect 3523 -14388 3557 -14132
rect 3701 -14388 3735 -14132
rect 3879 -14388 3913 -14132
rect 4057 -14388 4091 -14132
rect 5577 -14388 5611 -14132
rect 5755 -14388 5789 -14132
rect 5933 -14388 5967 -14132
rect 6111 -14388 6145 -14132
rect 6289 -14388 6323 -14132
rect 6467 -14388 6501 -14132
rect 6645 -14388 6679 -14132
rect 6823 -14388 6857 -14132
rect 7001 -14388 7035 -14132
rect 7179 -14388 7213 -14132
rect 7357 -14388 7391 -14132
rect 7535 -14388 7569 -14132
rect 7713 -14388 7747 -14132
rect 7891 -14388 7925 -14132
rect 8069 -14388 8103 -14132
rect 8247 -14388 8281 -14132
rect 8425 -14388 8459 -14132
rect 8603 -14388 8637 -14132
rect 8781 -14388 8815 -14132
rect 8959 -14388 8993 -14132
rect 9137 -14388 9171 -14132
rect 9315 -14388 9349 -14132
rect 9493 -14388 9527 -14132
rect 9671 -14388 9705 -14132
rect 9849 -14388 9883 -14132
rect 10027 -14388 10061 -14132
rect 10205 -14388 10239 -14132
rect 10383 -14388 10417 -14132
rect 10561 -14388 10595 -14132
rect 10739 -14388 10773 -14132
rect 10917 -14388 10951 -14132
rect 11095 -14388 11129 -14132
rect 11273 -14388 11307 -14132
rect 11451 -14388 11485 -14132
rect 11629 -14388 11663 -14132
rect 11807 -14388 11841 -14132
rect 11985 -14388 12019 -14132
rect 12163 -14388 12197 -14132
rect 12341 -14388 12375 -14132
rect 12519 -14388 12553 -14132
rect 12697 -14388 12731 -14132
rect -2089 -14472 -2045 -14438
rect -1911 -14472 -1867 -14438
rect -1733 -14472 -1689 -14438
rect -1555 -14472 -1511 -14438
rect -1377 -14472 -1333 -14438
rect -1199 -14472 -1155 -14438
rect -1021 -14472 -977 -14438
rect -843 -14472 -799 -14438
rect -665 -14472 -621 -14438
rect -487 -14472 -443 -14438
rect -309 -14472 -265 -14438
rect -131 -14472 -87 -14438
rect 47 -14472 91 -14438
rect 225 -14472 269 -14438
rect 403 -14472 447 -14438
rect 581 -14472 625 -14438
rect 759 -14472 803 -14438
rect 937 -14472 981 -14438
rect 1115 -14472 1159 -14438
rect 1293 -14472 1337 -14438
rect 1471 -14472 1515 -14438
rect 1649 -14472 1693 -14438
rect 1827 -14472 1871 -14438
rect 2005 -14472 2049 -14438
rect 2183 -14472 2227 -14438
rect 2361 -14472 2405 -14438
rect 2539 -14472 2583 -14438
rect 2717 -14472 2761 -14438
rect 2895 -14472 2939 -14438
rect 3073 -14472 3117 -14438
rect 3251 -14472 3295 -14438
rect 3429 -14472 3473 -14438
rect 3607 -14472 3651 -14438
rect 3785 -14472 3829 -14438
rect 3963 -14472 4007 -14438
rect 5661 -14472 5705 -14438
rect 5839 -14472 5883 -14438
rect 6017 -14472 6061 -14438
rect 6195 -14472 6239 -14438
rect 6373 -14472 6417 -14438
rect 6551 -14472 6595 -14438
rect 6729 -14472 6773 -14438
rect 6907 -14472 6951 -14438
rect 7085 -14472 7129 -14438
rect 7263 -14472 7307 -14438
rect 7441 -14472 7485 -14438
rect 7619 -14472 7663 -14438
rect 7797 -14472 7841 -14438
rect 7975 -14472 8019 -14438
rect 8153 -14472 8197 -14438
rect 8331 -14472 8375 -14438
rect 8509 -14472 8553 -14438
rect 8687 -14472 8731 -14438
rect 8865 -14472 8909 -14438
rect 9043 -14472 9087 -14438
rect 9221 -14472 9265 -14438
rect 9399 -14472 9443 -14438
rect 9577 -14472 9621 -14438
rect 9755 -14472 9799 -14438
rect 9933 -14472 9977 -14438
rect 10111 -14472 10155 -14438
rect 10289 -14472 10333 -14438
rect 10467 -14472 10511 -14438
rect 10645 -14472 10689 -14438
rect 10823 -14472 10867 -14438
rect 11001 -14472 11045 -14438
rect 11179 -14472 11223 -14438
rect 11357 -14472 11401 -14438
rect 11535 -14472 11579 -14438
rect 11713 -14472 11757 -14438
rect 11891 -14472 11935 -14438
rect 12069 -14472 12113 -14438
rect 12247 -14472 12291 -14438
rect 12425 -14472 12469 -14438
rect 12603 -14472 12647 -14438
rect -5944 -14734 -5900 -14700
rect -5766 -14734 -5722 -14700
rect -5588 -14734 -5544 -14700
rect -5410 -14734 -5366 -14700
rect -5232 -14734 -5188 -14700
rect -5054 -14734 -5010 -14700
rect -4876 -14734 -4832 -14700
rect -4698 -14734 -4654 -14700
rect -4520 -14734 -4476 -14700
rect -4342 -14734 -4298 -14700
rect -4164 -14734 -4120 -14700
rect -5944 -15044 -5900 -15010
rect -5766 -15044 -5722 -15010
rect -5588 -15044 -5544 -15010
rect -5410 -15044 -5366 -15010
rect -5232 -15044 -5188 -15010
rect -5054 -15044 -5010 -15010
rect -4876 -15044 -4832 -15010
rect -4698 -15044 -4654 -15010
rect -4520 -15044 -4476 -15010
rect -4342 -15044 -4298 -15010
rect -4164 -15044 -4120 -15010
rect -6028 -15350 -5994 -15094
rect -5850 -15350 -5816 -15094
rect -5672 -15350 -5638 -15094
rect -5494 -15350 -5460 -15094
rect -5316 -15350 -5282 -15094
rect -5138 -15350 -5104 -15094
rect -4960 -15350 -4926 -15094
rect -4782 -15350 -4748 -15094
rect -4604 -15350 -4570 -15094
rect -4426 -15350 -4392 -15094
rect -4248 -15350 -4214 -15094
rect -2089 -15082 -2045 -15048
rect -1911 -15082 -1867 -15048
rect -1733 -15082 -1689 -15048
rect -1555 -15082 -1511 -15048
rect -1377 -15082 -1333 -15048
rect -1199 -15082 -1155 -15048
rect -1021 -15082 -977 -15048
rect -843 -15082 -799 -15048
rect -665 -15082 -621 -15048
rect -487 -15082 -443 -15048
rect -309 -15082 -265 -15048
rect -131 -15082 -87 -15048
rect 47 -15082 91 -15048
rect 225 -15082 269 -15048
rect 403 -15082 447 -15048
rect 581 -15082 625 -15048
rect 759 -15082 803 -15048
rect 937 -15082 981 -15048
rect 1115 -15082 1159 -15048
rect 1293 -15082 1337 -15048
rect 1471 -15082 1515 -15048
rect 1649 -15082 1693 -15048
rect 1827 -15082 1871 -15048
rect 2005 -15082 2049 -15048
rect 2183 -15082 2227 -15048
rect 2361 -15082 2405 -15048
rect 2539 -15082 2583 -15048
rect 2717 -15082 2761 -15048
rect 2895 -15082 2939 -15048
rect 3073 -15082 3117 -15048
rect 3251 -15082 3295 -15048
rect 3429 -15082 3473 -15048
rect 3607 -15082 3651 -15048
rect 3785 -15082 3829 -15048
rect 3963 -15082 4007 -15048
rect 5661 -15082 5705 -15048
rect 5839 -15082 5883 -15048
rect 6017 -15082 6061 -15048
rect 6195 -15082 6239 -15048
rect 6373 -15082 6417 -15048
rect 6551 -15082 6595 -15048
rect 6729 -15082 6773 -15048
rect 6907 -15082 6951 -15048
rect 7085 -15082 7129 -15048
rect 7263 -15082 7307 -15048
rect 7441 -15082 7485 -15048
rect 7619 -15082 7663 -15048
rect 7797 -15082 7841 -15048
rect 7975 -15082 8019 -15048
rect 8153 -15082 8197 -15048
rect 8331 -15082 8375 -15048
rect 8509 -15082 8553 -15048
rect 8687 -15082 8731 -15048
rect 8865 -15082 8909 -15048
rect 9043 -15082 9087 -15048
rect 9221 -15082 9265 -15048
rect 9399 -15082 9443 -15048
rect 9577 -15082 9621 -15048
rect 9755 -15082 9799 -15048
rect 9933 -15082 9977 -15048
rect 10111 -15082 10155 -15048
rect 10289 -15082 10333 -15048
rect 10467 -15082 10511 -15048
rect 10645 -15082 10689 -15048
rect 10823 -15082 10867 -15048
rect 11001 -15082 11045 -15048
rect 11179 -15082 11223 -15048
rect 11357 -15082 11401 -15048
rect 11535 -15082 11579 -15048
rect 11713 -15082 11757 -15048
rect 11891 -15082 11935 -15048
rect 12069 -15082 12113 -15048
rect 12247 -15082 12291 -15048
rect 12425 -15082 12469 -15048
rect 12603 -15082 12647 -15048
rect -4070 -15350 -4036 -15094
rect -2173 -15388 -2139 -15132
rect -5944 -15434 -5900 -15400
rect -5766 -15434 -5722 -15400
rect -5588 -15434 -5544 -15400
rect -5410 -15434 -5366 -15400
rect -5232 -15434 -5188 -15400
rect -5054 -15434 -5010 -15400
rect -4876 -15434 -4832 -15400
rect -4698 -15434 -4654 -15400
rect -4520 -15434 -4476 -15400
rect -4342 -15434 -4298 -15400
rect -4164 -15434 -4120 -15400
rect -1995 -15388 -1961 -15132
rect -1817 -15388 -1783 -15132
rect -1639 -15388 -1605 -15132
rect -1461 -15388 -1427 -15132
rect -1283 -15388 -1249 -15132
rect -1105 -15388 -1071 -15132
rect -927 -15388 -893 -15132
rect -749 -15388 -715 -15132
rect -571 -15388 -537 -15132
rect -393 -15388 -359 -15132
rect -215 -15388 -181 -15132
rect -37 -15388 -3 -15132
rect 141 -15388 175 -15132
rect 319 -15388 353 -15132
rect 497 -15388 531 -15132
rect 675 -15388 709 -15132
rect 853 -15388 887 -15132
rect 1031 -15388 1065 -15132
rect 1209 -15388 1243 -15132
rect 1387 -15388 1421 -15132
rect 1565 -15388 1599 -15132
rect 1743 -15388 1777 -15132
rect 1921 -15388 1955 -15132
rect 2099 -15388 2133 -15132
rect 2277 -15388 2311 -15132
rect 2455 -15388 2489 -15132
rect 2633 -15388 2667 -15132
rect 2811 -15388 2845 -15132
rect 2989 -15388 3023 -15132
rect 3167 -15388 3201 -15132
rect 3345 -15388 3379 -15132
rect 3523 -15388 3557 -15132
rect 3701 -15388 3735 -15132
rect 3879 -15388 3913 -15132
rect 4057 -15388 4091 -15132
rect 5577 -15388 5611 -15132
rect 5755 -15388 5789 -15132
rect 5933 -15388 5967 -15132
rect 6111 -15388 6145 -15132
rect 6289 -15388 6323 -15132
rect 6467 -15388 6501 -15132
rect 6645 -15388 6679 -15132
rect 6823 -15388 6857 -15132
rect 7001 -15388 7035 -15132
rect 7179 -15388 7213 -15132
rect 7357 -15388 7391 -15132
rect 7535 -15388 7569 -15132
rect 7713 -15388 7747 -15132
rect 7891 -15388 7925 -15132
rect 8069 -15388 8103 -15132
rect 8247 -15388 8281 -15132
rect 8425 -15388 8459 -15132
rect 8603 -15388 8637 -15132
rect 8781 -15388 8815 -15132
rect 8959 -15388 8993 -15132
rect 9137 -15388 9171 -15132
rect 9315 -15388 9349 -15132
rect 9493 -15388 9527 -15132
rect 9671 -15388 9705 -15132
rect 9849 -15388 9883 -15132
rect 10027 -15388 10061 -15132
rect 10205 -15388 10239 -15132
rect 10383 -15388 10417 -15132
rect 10561 -15388 10595 -15132
rect 10739 -15388 10773 -15132
rect 10917 -15388 10951 -15132
rect 11095 -15388 11129 -15132
rect 11273 -15388 11307 -15132
rect 11451 -15388 11485 -15132
rect 11629 -15388 11663 -15132
rect 11807 -15388 11841 -15132
rect 11985 -15388 12019 -15132
rect 12163 -15388 12197 -15132
rect 12341 -15388 12375 -15132
rect 12519 -15388 12553 -15132
rect 12697 -15388 12731 -15132
rect -2089 -15472 -2045 -15438
rect -1911 -15472 -1867 -15438
rect -1733 -15472 -1689 -15438
rect -1555 -15472 -1511 -15438
rect -1377 -15472 -1333 -15438
rect -1199 -15472 -1155 -15438
rect -1021 -15472 -977 -15438
rect -843 -15472 -799 -15438
rect -665 -15472 -621 -15438
rect -487 -15472 -443 -15438
rect -309 -15472 -265 -15438
rect -131 -15472 -87 -15438
rect 47 -15472 91 -15438
rect 225 -15472 269 -15438
rect 403 -15472 447 -15438
rect 581 -15472 625 -15438
rect 759 -15472 803 -15438
rect 937 -15472 981 -15438
rect 1115 -15472 1159 -15438
rect 1293 -15472 1337 -15438
rect 1471 -15472 1515 -15438
rect 1649 -15472 1693 -15438
rect 1827 -15472 1871 -15438
rect 2005 -15472 2049 -15438
rect 2183 -15472 2227 -15438
rect 2361 -15472 2405 -15438
rect 2539 -15472 2583 -15438
rect 2717 -15472 2761 -15438
rect 2895 -15472 2939 -15438
rect 3073 -15472 3117 -15438
rect 3251 -15472 3295 -15438
rect 3429 -15472 3473 -15438
rect 3607 -15472 3651 -15438
rect 3785 -15472 3829 -15438
rect 3963 -15472 4007 -15438
rect 5661 -15472 5705 -15438
rect 5839 -15472 5883 -15438
rect 6017 -15472 6061 -15438
rect 6195 -15472 6239 -15438
rect 6373 -15472 6417 -15438
rect 6551 -15472 6595 -15438
rect 6729 -15472 6773 -15438
rect 6907 -15472 6951 -15438
rect 7085 -15472 7129 -15438
rect 7263 -15472 7307 -15438
rect 7441 -15472 7485 -15438
rect 7619 -15472 7663 -15438
rect 7797 -15472 7841 -15438
rect 7975 -15472 8019 -15438
rect 8153 -15472 8197 -15438
rect 8331 -15472 8375 -15438
rect 8509 -15472 8553 -15438
rect 8687 -15472 8731 -15438
rect 8865 -15472 8909 -15438
rect 9043 -15472 9087 -15438
rect 9221 -15472 9265 -15438
rect 9399 -15472 9443 -15438
rect 9577 -15472 9621 -15438
rect 9755 -15472 9799 -15438
rect 9933 -15472 9977 -15438
rect 10111 -15472 10155 -15438
rect 10289 -15472 10333 -15438
rect 10467 -15472 10511 -15438
rect 10645 -15472 10689 -15438
rect 10823 -15472 10867 -15438
rect 11001 -15472 11045 -15438
rect 11179 -15472 11223 -15438
rect 11357 -15472 11401 -15438
rect 11535 -15472 11579 -15438
rect 11713 -15472 11757 -15438
rect 11891 -15472 11935 -15438
rect 12069 -15472 12113 -15438
rect 12247 -15472 12291 -15438
rect 12425 -15472 12469 -15438
rect 12603 -15472 12647 -15438
rect -5944 -15744 -5900 -15710
rect -5766 -15744 -5722 -15710
rect -5588 -15744 -5544 -15710
rect -5410 -15744 -5366 -15710
rect -5232 -15744 -5188 -15710
rect -5054 -15744 -5010 -15710
rect -4876 -15744 -4832 -15710
rect -4698 -15744 -4654 -15710
rect -4520 -15744 -4476 -15710
rect -4342 -15744 -4298 -15710
rect -4164 -15744 -4120 -15710
rect -6028 -16050 -5994 -15794
rect -5850 -16050 -5816 -15794
rect -5672 -16050 -5638 -15794
rect -5494 -16050 -5460 -15794
rect -5316 -16050 -5282 -15794
rect -5138 -16050 -5104 -15794
rect -4960 -16050 -4926 -15794
rect -4782 -16050 -4748 -15794
rect -4604 -16050 -4570 -15794
rect -4426 -16050 -4392 -15794
rect -4248 -16050 -4214 -15794
rect -4070 -16050 -4036 -15794
rect -2089 -16082 -2045 -16048
rect -1911 -16082 -1867 -16048
rect -1733 -16082 -1689 -16048
rect -1555 -16082 -1511 -16048
rect -1377 -16082 -1333 -16048
rect -1199 -16082 -1155 -16048
rect -1021 -16082 -977 -16048
rect -843 -16082 -799 -16048
rect -665 -16082 -621 -16048
rect -487 -16082 -443 -16048
rect -309 -16082 -265 -16048
rect -131 -16082 -87 -16048
rect 47 -16082 91 -16048
rect 225 -16082 269 -16048
rect 403 -16082 447 -16048
rect 581 -16082 625 -16048
rect 759 -16082 803 -16048
rect 937 -16082 981 -16048
rect 1115 -16082 1159 -16048
rect 1293 -16082 1337 -16048
rect 1471 -16082 1515 -16048
rect 1649 -16082 1693 -16048
rect 1827 -16082 1871 -16048
rect 2005 -16082 2049 -16048
rect 2183 -16082 2227 -16048
rect 2361 -16082 2405 -16048
rect 2539 -16082 2583 -16048
rect 2717 -16082 2761 -16048
rect 2895 -16082 2939 -16048
rect 3073 -16082 3117 -16048
rect 3251 -16082 3295 -16048
rect 3429 -16082 3473 -16048
rect 3607 -16082 3651 -16048
rect 3785 -16082 3829 -16048
rect 3963 -16082 4007 -16048
rect 5661 -16082 5705 -16048
rect 5839 -16082 5883 -16048
rect 6017 -16082 6061 -16048
rect 6195 -16082 6239 -16048
rect 6373 -16082 6417 -16048
rect 6551 -16082 6595 -16048
rect 6729 -16082 6773 -16048
rect 6907 -16082 6951 -16048
rect 7085 -16082 7129 -16048
rect 7263 -16082 7307 -16048
rect 7441 -16082 7485 -16048
rect 7619 -16082 7663 -16048
rect 7797 -16082 7841 -16048
rect 7975 -16082 8019 -16048
rect 8153 -16082 8197 -16048
rect 8331 -16082 8375 -16048
rect 8509 -16082 8553 -16048
rect 8687 -16082 8731 -16048
rect 8865 -16082 8909 -16048
rect 9043 -16082 9087 -16048
rect 9221 -16082 9265 -16048
rect 9399 -16082 9443 -16048
rect 9577 -16082 9621 -16048
rect 9755 -16082 9799 -16048
rect 9933 -16082 9977 -16048
rect 10111 -16082 10155 -16048
rect 10289 -16082 10333 -16048
rect 10467 -16082 10511 -16048
rect 10645 -16082 10689 -16048
rect 10823 -16082 10867 -16048
rect 11001 -16082 11045 -16048
rect 11179 -16082 11223 -16048
rect 11357 -16082 11401 -16048
rect 11535 -16082 11579 -16048
rect 11713 -16082 11757 -16048
rect 11891 -16082 11935 -16048
rect 12069 -16082 12113 -16048
rect 12247 -16082 12291 -16048
rect 12425 -16082 12469 -16048
rect 12603 -16082 12647 -16048
rect -5944 -16134 -5900 -16100
rect -5766 -16134 -5722 -16100
rect -5588 -16134 -5544 -16100
rect -5410 -16134 -5366 -16100
rect -5232 -16134 -5188 -16100
rect -5054 -16134 -5010 -16100
rect -4876 -16134 -4832 -16100
rect -4698 -16134 -4654 -16100
rect -4520 -16134 -4476 -16100
rect -4342 -16134 -4298 -16100
rect -4164 -16134 -4120 -16100
rect -2173 -16388 -2139 -16132
rect -1995 -16388 -1961 -16132
rect -1817 -16388 -1783 -16132
rect -1639 -16388 -1605 -16132
rect -1461 -16388 -1427 -16132
rect -1283 -16388 -1249 -16132
rect -1105 -16388 -1071 -16132
rect -927 -16388 -893 -16132
rect -749 -16388 -715 -16132
rect -571 -16388 -537 -16132
rect -393 -16388 -359 -16132
rect -215 -16388 -181 -16132
rect -37 -16388 -3 -16132
rect 141 -16388 175 -16132
rect 319 -16388 353 -16132
rect 497 -16388 531 -16132
rect 675 -16388 709 -16132
rect 853 -16388 887 -16132
rect 1031 -16388 1065 -16132
rect 1209 -16388 1243 -16132
rect 1387 -16388 1421 -16132
rect 1565 -16388 1599 -16132
rect 1743 -16388 1777 -16132
rect 1921 -16388 1955 -16132
rect 2099 -16388 2133 -16132
rect 2277 -16388 2311 -16132
rect 2455 -16388 2489 -16132
rect 2633 -16388 2667 -16132
rect 2811 -16388 2845 -16132
rect 2989 -16388 3023 -16132
rect 3167 -16388 3201 -16132
rect 3345 -16388 3379 -16132
rect 3523 -16388 3557 -16132
rect 3701 -16388 3735 -16132
rect 3879 -16388 3913 -16132
rect 4057 -16388 4091 -16132
rect 5577 -16388 5611 -16132
rect 5755 -16388 5789 -16132
rect 5933 -16388 5967 -16132
rect 6111 -16388 6145 -16132
rect 6289 -16388 6323 -16132
rect 6467 -16388 6501 -16132
rect 6645 -16388 6679 -16132
rect 6823 -16388 6857 -16132
rect 7001 -16388 7035 -16132
rect 7179 -16388 7213 -16132
rect 7357 -16388 7391 -16132
rect 7535 -16388 7569 -16132
rect 7713 -16388 7747 -16132
rect 7891 -16388 7925 -16132
rect 8069 -16388 8103 -16132
rect 8247 -16388 8281 -16132
rect 8425 -16388 8459 -16132
rect 8603 -16388 8637 -16132
rect 8781 -16388 8815 -16132
rect 8959 -16388 8993 -16132
rect 9137 -16388 9171 -16132
rect 9315 -16388 9349 -16132
rect 9493 -16388 9527 -16132
rect 9671 -16388 9705 -16132
rect 9849 -16388 9883 -16132
rect 10027 -16388 10061 -16132
rect 10205 -16388 10239 -16132
rect 10383 -16388 10417 -16132
rect 10561 -16388 10595 -16132
rect 10739 -16388 10773 -16132
rect 10917 -16388 10951 -16132
rect 11095 -16388 11129 -16132
rect 11273 -16388 11307 -16132
rect 11451 -16388 11485 -16132
rect 11629 -16388 11663 -16132
rect 11807 -16388 11841 -16132
rect 11985 -16388 12019 -16132
rect 12163 -16388 12197 -16132
rect 12341 -16388 12375 -16132
rect 12519 -16388 12553 -16132
rect 12697 -16388 12731 -16132
rect -5944 -16444 -5900 -16410
rect -5766 -16444 -5722 -16410
rect -5588 -16444 -5544 -16410
rect -5410 -16444 -5366 -16410
rect -5232 -16444 -5188 -16410
rect -5054 -16444 -5010 -16410
rect -4876 -16444 -4832 -16410
rect -4698 -16444 -4654 -16410
rect -4520 -16444 -4476 -16410
rect -4342 -16444 -4298 -16410
rect -4164 -16444 -4120 -16410
rect -2089 -16472 -2045 -16438
rect -1911 -16472 -1867 -16438
rect -1733 -16472 -1689 -16438
rect -1555 -16472 -1511 -16438
rect -1377 -16472 -1333 -16438
rect -1199 -16472 -1155 -16438
rect -1021 -16472 -977 -16438
rect -843 -16472 -799 -16438
rect -665 -16472 -621 -16438
rect -487 -16472 -443 -16438
rect -309 -16472 -265 -16438
rect -131 -16472 -87 -16438
rect 47 -16472 91 -16438
rect 225 -16472 269 -16438
rect 403 -16472 447 -16438
rect 581 -16472 625 -16438
rect 759 -16472 803 -16438
rect 937 -16472 981 -16438
rect 1115 -16472 1159 -16438
rect 1293 -16472 1337 -16438
rect 1471 -16472 1515 -16438
rect 1649 -16472 1693 -16438
rect 1827 -16472 1871 -16438
rect 2005 -16472 2049 -16438
rect 2183 -16472 2227 -16438
rect 2361 -16472 2405 -16438
rect 2539 -16472 2583 -16438
rect 2717 -16472 2761 -16438
rect 2895 -16472 2939 -16438
rect 3073 -16472 3117 -16438
rect 3251 -16472 3295 -16438
rect 3429 -16472 3473 -16438
rect 3607 -16472 3651 -16438
rect 3785 -16472 3829 -16438
rect 3963 -16472 4007 -16438
rect 5661 -16472 5705 -16438
rect 5839 -16472 5883 -16438
rect 6017 -16472 6061 -16438
rect 6195 -16472 6239 -16438
rect 6373 -16472 6417 -16438
rect 6551 -16472 6595 -16438
rect 6729 -16472 6773 -16438
rect 6907 -16472 6951 -16438
rect 7085 -16472 7129 -16438
rect 7263 -16472 7307 -16438
rect 7441 -16472 7485 -16438
rect 7619 -16472 7663 -16438
rect 7797 -16472 7841 -16438
rect 7975 -16472 8019 -16438
rect 8153 -16472 8197 -16438
rect 8331 -16472 8375 -16438
rect 8509 -16472 8553 -16438
rect 8687 -16472 8731 -16438
rect 8865 -16472 8909 -16438
rect 9043 -16472 9087 -16438
rect 9221 -16472 9265 -16438
rect 9399 -16472 9443 -16438
rect 9577 -16472 9621 -16438
rect 9755 -16472 9799 -16438
rect 9933 -16472 9977 -16438
rect 10111 -16472 10155 -16438
rect 10289 -16472 10333 -16438
rect 10467 -16472 10511 -16438
rect 10645 -16472 10689 -16438
rect 10823 -16472 10867 -16438
rect 11001 -16472 11045 -16438
rect 11179 -16472 11223 -16438
rect 11357 -16472 11401 -16438
rect 11535 -16472 11579 -16438
rect 11713 -16472 11757 -16438
rect 11891 -16472 11935 -16438
rect 12069 -16472 12113 -16438
rect 12247 -16472 12291 -16438
rect 12425 -16472 12469 -16438
rect 12603 -16472 12647 -16438
rect -6028 -16750 -5994 -16494
rect -5850 -16750 -5816 -16494
rect -5672 -16750 -5638 -16494
rect -5494 -16750 -5460 -16494
rect -5316 -16750 -5282 -16494
rect -5138 -16750 -5104 -16494
rect -4960 -16750 -4926 -16494
rect -4782 -16750 -4748 -16494
rect -4604 -16750 -4570 -16494
rect -4426 -16750 -4392 -16494
rect -4248 -16750 -4214 -16494
rect -4070 -16750 -4036 -16494
rect -5944 -16834 -5900 -16800
rect -5766 -16834 -5722 -16800
rect -5588 -16834 -5544 -16800
rect -5410 -16834 -5366 -16800
rect -5232 -16834 -5188 -16800
rect -5054 -16834 -5010 -16800
rect -4876 -16834 -4832 -16800
rect -4698 -16834 -4654 -16800
rect -4520 -16834 -4476 -16800
rect -4342 -16834 -4298 -16800
rect -4164 -16834 -4120 -16800
rect -7323 -17559 13384 -17459
<< metal1 >>
rect -7605 -1260 3704 -1200
rect -7605 -1353 -7379 -1260
rect 3329 -1353 3704 -1260
rect -7605 -1467 3704 -1353
rect -5059 -1807 -5025 -1467
rect -5945 -1808 -3809 -1807
rect -5945 -1841 -3776 -1808
rect -6234 -2039 -6158 -2023
rect -6056 -2039 -5980 -2023
rect -5945 -2039 -5911 -1841
rect -5877 -1963 -5867 -1910
rect -5814 -1963 -5804 -1910
rect -5699 -1963 -5689 -1910
rect -5636 -1963 -5626 -1910
rect -5520 -1963 -5510 -1910
rect -5457 -1963 -5447 -1910
rect -5343 -1963 -5333 -1910
rect -5280 -1963 -5270 -1910
rect -5165 -1963 -5155 -1910
rect -5102 -1963 -5092 -1910
rect -4986 -1963 -4976 -1910
rect -4923 -1963 -4913 -1910
rect -4809 -1963 -4799 -1910
rect -4746 -1963 -4736 -1910
rect -4631 -1963 -4621 -1910
rect -4568 -1963 -4558 -1910
rect -4453 -1963 -4443 -1910
rect -4390 -1963 -4380 -1910
rect -4275 -1963 -4265 -1910
rect -4212 -1963 -4202 -1910
rect -4096 -1963 -4086 -1910
rect -4033 -1963 -4023 -1910
rect -3919 -1963 -3909 -1910
rect -3856 -1963 -3846 -1910
rect -5857 -2023 -5823 -1963
rect -5679 -2023 -5645 -1963
rect -5501 -2023 -5467 -1963
rect -5322 -2023 -5288 -1963
rect -5145 -2023 -5111 -1963
rect -4967 -2023 -4933 -1963
rect -4789 -2023 -4755 -1963
rect -4611 -2023 -4577 -1963
rect -4433 -2023 -4399 -1963
rect -4255 -2023 -4221 -1963
rect -4077 -2023 -4043 -1963
rect -3898 -2023 -3864 -1963
rect -6302 -2073 -6218 -2039
rect -6174 -2073 -6040 -2039
rect -5996 -2073 -5911 -2039
rect -6302 -2120 -6268 -2073
rect -6234 -2079 -6158 -2073
rect -6126 -2120 -6092 -2073
rect -6056 -2079 -5980 -2073
rect -5945 -2120 -5911 -2073
rect -5878 -2039 -5802 -2023
rect -5878 -2073 -5862 -2039
rect -5818 -2073 -5802 -2039
rect -5878 -2079 -5802 -2073
rect -5700 -2039 -5624 -2023
rect -5700 -2073 -5684 -2039
rect -5640 -2073 -5624 -2039
rect -5700 -2079 -5624 -2073
rect -5522 -2039 -5446 -2023
rect -5522 -2073 -5506 -2039
rect -5462 -2073 -5446 -2039
rect -5522 -2079 -5446 -2073
rect -5344 -2039 -5268 -2023
rect -5344 -2073 -5328 -2039
rect -5284 -2073 -5268 -2039
rect -5344 -2079 -5268 -2073
rect -5166 -2039 -5090 -2023
rect -5166 -2073 -5150 -2039
rect -5106 -2073 -5090 -2039
rect -5166 -2079 -5090 -2073
rect -4988 -2039 -4912 -2023
rect -4988 -2073 -4972 -2039
rect -4928 -2073 -4912 -2039
rect -4988 -2079 -4912 -2073
rect -4810 -2039 -4734 -2023
rect -4810 -2073 -4794 -2039
rect -4750 -2073 -4734 -2039
rect -4810 -2079 -4734 -2073
rect -4632 -2039 -4556 -2023
rect -4632 -2073 -4616 -2039
rect -4572 -2073 -4556 -2039
rect -4632 -2079 -4556 -2073
rect -4454 -2039 -4378 -2023
rect -4454 -2073 -4438 -2039
rect -4394 -2073 -4378 -2039
rect -4454 -2079 -4378 -2073
rect -4276 -2039 -4200 -2023
rect -4276 -2073 -4260 -2039
rect -4216 -2073 -4200 -2039
rect -4276 -2079 -4200 -2073
rect -4098 -2039 -4022 -2023
rect -4098 -2073 -4082 -2039
rect -4038 -2073 -4022 -2039
rect -4098 -2079 -4022 -2073
rect -3920 -2039 -3844 -2023
rect -3920 -2073 -3904 -2039
rect -3860 -2073 -3844 -2039
rect -3920 -2079 -3844 -2073
rect -3810 -2120 -3776 -1841
rect -1119 -1963 -1109 -1910
rect -1056 -1963 -1046 -1910
rect -3742 -2039 -3666 -2023
rect -3742 -2073 -3726 -2039
rect -3682 -2073 -3666 -2039
rect -3742 -2079 -3666 -2073
rect -3564 -2039 -3488 -2023
rect -3564 -2073 -3548 -2039
rect -3504 -2073 -3488 -2039
rect -3564 -2079 -3488 -2073
rect -6308 -2132 -6262 -2120
rect -6308 -2388 -6302 -2132
rect -6268 -2388 -6262 -2132
rect -6308 -2400 -6262 -2388
rect -6130 -2132 -6084 -2120
rect -6130 -2388 -6124 -2132
rect -6090 -2388 -6084 -2132
rect -6130 -2400 -6084 -2388
rect -5952 -2132 -5906 -2120
rect -5952 -2388 -5946 -2132
rect -5912 -2388 -5906 -2132
rect -5952 -2400 -5906 -2388
rect -5774 -2132 -5728 -2120
rect -5774 -2388 -5768 -2132
rect -5734 -2388 -5728 -2132
rect -5774 -2400 -5728 -2388
rect -5596 -2132 -5550 -2120
rect -5596 -2388 -5590 -2132
rect -5556 -2388 -5550 -2132
rect -5596 -2400 -5550 -2388
rect -5418 -2132 -5372 -2120
rect -5418 -2388 -5412 -2132
rect -5378 -2388 -5372 -2132
rect -5418 -2400 -5372 -2388
rect -5240 -2132 -5194 -2120
rect -5240 -2388 -5234 -2132
rect -5200 -2388 -5194 -2132
rect -5240 -2400 -5194 -2388
rect -5062 -2132 -5016 -2120
rect -5062 -2388 -5056 -2132
rect -5022 -2388 -5016 -2132
rect -5062 -2400 -5016 -2388
rect -4884 -2132 -4838 -2120
rect -4884 -2388 -4878 -2132
rect -4844 -2388 -4838 -2132
rect -4884 -2400 -4838 -2388
rect -4706 -2132 -4660 -2120
rect -4706 -2388 -4700 -2132
rect -4666 -2388 -4660 -2132
rect -4706 -2400 -4660 -2388
rect -4528 -2132 -4482 -2120
rect -4528 -2388 -4522 -2132
rect -4488 -2388 -4482 -2132
rect -4528 -2400 -4482 -2388
rect -4350 -2132 -4304 -2120
rect -4350 -2388 -4344 -2132
rect -4310 -2388 -4304 -2132
rect -4350 -2400 -4304 -2388
rect -4172 -2132 -4126 -2120
rect -4172 -2388 -4166 -2132
rect -4132 -2388 -4126 -2132
rect -4172 -2400 -4126 -2388
rect -3994 -2132 -3948 -2120
rect -3994 -2388 -3988 -2132
rect -3954 -2388 -3948 -2132
rect -3994 -2400 -3948 -2388
rect -3816 -2132 -3770 -2120
rect -3816 -2388 -3810 -2132
rect -3776 -2388 -3770 -2132
rect -3816 -2400 -3770 -2388
rect -3638 -2132 -3592 -2120
rect -3638 -2388 -3632 -2132
rect -3598 -2388 -3592 -2132
rect -3638 -2400 -3592 -2388
rect -3460 -2132 -3414 -2120
rect -3460 -2388 -3454 -2132
rect -3420 -2388 -3414 -2132
rect -3460 -2400 -3414 -2388
rect -6234 -2447 -6158 -2441
rect -6234 -2481 -6218 -2447
rect -6174 -2481 -6158 -2447
rect -6234 -2497 -6158 -2481
rect -6056 -2447 -5980 -2441
rect -6056 -2481 -6040 -2447
rect -5996 -2481 -5980 -2447
rect -6056 -2497 -5980 -2481
rect -6508 -2582 -6498 -2529
rect -6445 -2582 -6435 -2529
rect -6635 -3454 -6625 -3401
rect -6572 -3454 -6562 -3401
rect -6625 -5322 -6572 -3454
rect -6498 -3640 -6445 -2582
rect -6054 -2833 -6044 -2780
rect -5991 -2833 -5981 -2780
rect -6035 -2893 -6001 -2833
rect -6234 -2909 -6158 -2893
rect -6234 -2911 -6218 -2909
rect -6302 -2943 -6218 -2911
rect -6174 -2911 -6158 -2909
rect -6056 -2909 -5980 -2893
rect -6174 -2943 -6090 -2911
rect -6302 -2945 -6090 -2943
rect -6302 -2990 -6268 -2945
rect -6234 -2949 -6158 -2945
rect -6124 -2990 -6090 -2945
rect -6056 -2943 -6040 -2909
rect -5996 -2943 -5980 -2909
rect -6056 -2949 -5980 -2943
rect -5946 -2990 -5912 -2400
rect -5878 -2447 -5802 -2441
rect -5878 -2481 -5862 -2447
rect -5818 -2481 -5802 -2447
rect -5878 -2497 -5802 -2481
rect -5856 -2780 -5822 -2497
rect -5768 -2530 -5734 -2400
rect -5700 -2447 -5624 -2441
rect -5700 -2481 -5684 -2447
rect -5640 -2481 -5624 -2447
rect -5700 -2497 -5624 -2481
rect -5787 -2583 -5777 -2530
rect -5724 -2583 -5714 -2530
rect -5876 -2833 -5866 -2780
rect -5813 -2833 -5803 -2780
rect -5856 -2893 -5822 -2833
rect -5679 -2893 -5645 -2497
rect -5878 -2909 -5802 -2893
rect -5878 -2943 -5862 -2909
rect -5818 -2943 -5802 -2909
rect -5878 -2949 -5802 -2943
rect -5700 -2909 -5624 -2893
rect -5700 -2943 -5684 -2909
rect -5640 -2943 -5624 -2909
rect -5700 -2949 -5624 -2943
rect -5590 -2990 -5556 -2400
rect -5522 -2447 -5446 -2441
rect -5522 -2481 -5506 -2447
rect -5462 -2481 -5446 -2447
rect -5522 -2497 -5446 -2481
rect -5501 -2893 -5467 -2497
rect -5412 -2668 -5378 -2400
rect -5344 -2447 -5268 -2441
rect -5344 -2481 -5328 -2447
rect -5284 -2481 -5268 -2447
rect -5344 -2497 -5268 -2481
rect -5431 -2721 -5421 -2668
rect -5368 -2721 -5358 -2668
rect -5323 -2893 -5289 -2497
rect -5522 -2909 -5446 -2893
rect -5522 -2943 -5506 -2909
rect -5462 -2943 -5446 -2909
rect -5522 -2949 -5446 -2943
rect -5344 -2909 -5268 -2893
rect -5344 -2943 -5328 -2909
rect -5284 -2943 -5268 -2909
rect -5344 -2949 -5268 -2943
rect -5234 -2990 -5200 -2400
rect -5166 -2447 -5090 -2441
rect -5166 -2481 -5150 -2447
rect -5106 -2481 -5090 -2447
rect -5166 -2497 -5090 -2481
rect -5145 -2893 -5111 -2497
rect -5056 -2530 -5022 -2400
rect -4988 -2447 -4912 -2441
rect -4988 -2481 -4972 -2447
rect -4928 -2481 -4912 -2447
rect -4988 -2497 -4912 -2481
rect -5076 -2583 -5066 -2530
rect -5013 -2583 -5003 -2530
rect -4967 -2893 -4933 -2497
rect -5166 -2909 -5090 -2893
rect -5166 -2943 -5150 -2909
rect -5106 -2943 -5090 -2909
rect -5166 -2949 -5090 -2943
rect -4988 -2909 -4912 -2893
rect -4988 -2943 -4972 -2909
rect -4928 -2943 -4912 -2909
rect -4988 -2949 -4912 -2943
rect -4878 -2990 -4844 -2400
rect -4810 -2447 -4734 -2441
rect -4810 -2481 -4794 -2447
rect -4750 -2481 -4734 -2447
rect -4810 -2497 -4734 -2481
rect -4789 -2893 -4755 -2497
rect -4700 -2668 -4666 -2400
rect -4632 -2447 -4556 -2441
rect -4632 -2481 -4616 -2447
rect -4572 -2481 -4556 -2447
rect -4632 -2497 -4556 -2481
rect -4720 -2721 -4710 -2668
rect -4657 -2721 -4647 -2668
rect -4611 -2893 -4577 -2497
rect -4810 -2909 -4734 -2893
rect -4810 -2943 -4794 -2909
rect -4750 -2943 -4734 -2909
rect -4810 -2949 -4734 -2943
rect -4632 -2909 -4556 -2893
rect -4632 -2943 -4616 -2909
rect -4572 -2943 -4556 -2909
rect -4632 -2949 -4556 -2943
rect -4522 -2990 -4488 -2400
rect -4454 -2447 -4378 -2441
rect -4454 -2481 -4438 -2447
rect -4394 -2481 -4378 -2447
rect -4454 -2497 -4378 -2481
rect -4433 -2893 -4399 -2497
rect -4344 -2530 -4310 -2400
rect -4276 -2447 -4200 -2441
rect -4276 -2481 -4260 -2447
rect -4216 -2481 -4200 -2447
rect -4276 -2497 -4200 -2481
rect -4364 -2583 -4354 -2530
rect -4301 -2583 -4291 -2530
rect -4255 -2893 -4221 -2497
rect -4454 -2909 -4378 -2893
rect -4454 -2943 -4438 -2909
rect -4394 -2943 -4378 -2909
rect -4454 -2949 -4378 -2943
rect -4276 -2909 -4200 -2893
rect -4276 -2943 -4260 -2909
rect -4216 -2943 -4200 -2909
rect -4276 -2949 -4200 -2943
rect -4166 -2990 -4132 -2400
rect -4098 -2447 -4022 -2441
rect -4098 -2481 -4082 -2447
rect -4038 -2481 -4022 -2447
rect -4098 -2497 -4022 -2481
rect -4077 -2893 -4043 -2497
rect -3988 -2668 -3954 -2400
rect -3920 -2447 -3844 -2441
rect -3920 -2481 -3904 -2447
rect -3860 -2481 -3844 -2447
rect -3920 -2497 -3844 -2481
rect -3810 -2446 -3776 -2400
rect -3742 -2446 -3666 -2441
rect -3633 -2446 -3599 -2400
rect -3564 -2446 -3488 -2441
rect -3454 -2446 -3420 -2400
rect -1099 -2425 -1065 -1963
rect -3810 -2447 -3420 -2446
rect -3810 -2480 -3726 -2447
rect -4008 -2721 -3998 -2668
rect -3945 -2721 -3935 -2668
rect -3899 -2780 -3865 -2497
rect -3918 -2833 -3908 -2780
rect -3855 -2833 -3845 -2780
rect -3899 -2893 -3865 -2833
rect -4098 -2909 -4022 -2893
rect -4098 -2943 -4082 -2909
rect -4038 -2943 -4022 -2909
rect -4098 -2949 -4022 -2943
rect -3920 -2909 -3844 -2893
rect -3920 -2943 -3904 -2909
rect -3860 -2943 -3844 -2909
rect -3920 -2949 -3844 -2943
rect -3810 -2990 -3776 -2480
rect -3742 -2481 -3726 -2480
rect -3682 -2480 -3548 -2447
rect -3682 -2481 -3666 -2480
rect -3742 -2497 -3666 -2481
rect -3564 -2481 -3548 -2480
rect -3504 -2480 -3420 -2447
rect -1119 -2478 -1109 -2425
rect -1056 -2478 -1046 -2425
rect -762 -2478 -752 -2425
rect -699 -2478 -689 -2425
rect -3504 -2481 -3488 -2480
rect -3564 -2497 -3488 -2481
rect -2634 -2611 -2624 -2558
rect -2571 -2611 -2561 -2558
rect -1295 -2611 -1285 -2558
rect -1232 -2611 -1222 -2558
rect -3308 -2721 -3298 -2668
rect -3245 -2721 -3235 -2668
rect -3741 -2833 -3731 -2780
rect -3678 -2833 -3668 -2780
rect -3721 -2893 -3687 -2833
rect -3742 -2909 -3666 -2893
rect -3742 -2943 -3726 -2909
rect -3682 -2943 -3666 -2909
rect -3742 -2949 -3666 -2943
rect -3564 -2909 -3488 -2893
rect -3564 -2943 -3548 -2909
rect -3504 -2943 -3488 -2909
rect -3564 -2949 -3488 -2943
rect -6308 -3002 -6262 -2990
rect -6308 -3258 -6302 -3002
rect -6268 -3258 -6262 -3002
rect -6308 -3270 -6262 -3258
rect -6130 -3002 -6084 -2990
rect -6130 -3258 -6124 -3002
rect -6090 -3258 -6084 -3002
rect -6130 -3270 -6084 -3258
rect -5952 -3002 -5906 -2990
rect -5952 -3258 -5946 -3002
rect -5912 -3258 -5906 -3002
rect -5952 -3270 -5906 -3258
rect -5774 -3002 -5728 -2990
rect -5774 -3258 -5768 -3002
rect -5734 -3258 -5728 -3002
rect -5774 -3270 -5728 -3258
rect -5596 -3002 -5550 -2990
rect -5596 -3258 -5590 -3002
rect -5556 -3258 -5550 -3002
rect -5596 -3270 -5550 -3258
rect -5418 -3002 -5372 -2990
rect -5418 -3258 -5412 -3002
rect -5378 -3258 -5372 -3002
rect -5418 -3270 -5372 -3258
rect -5240 -3002 -5194 -2990
rect -5240 -3258 -5234 -3002
rect -5200 -3258 -5194 -3002
rect -5240 -3270 -5194 -3258
rect -5062 -3002 -5016 -2990
rect -5062 -3258 -5056 -3002
rect -5022 -3258 -5016 -3002
rect -5062 -3270 -5016 -3258
rect -4884 -3002 -4838 -2990
rect -4884 -3258 -4878 -3002
rect -4844 -3258 -4838 -3002
rect -4884 -3270 -4838 -3258
rect -4706 -3002 -4660 -2990
rect -4706 -3258 -4700 -3002
rect -4666 -3258 -4660 -3002
rect -4706 -3270 -4660 -3258
rect -4528 -3002 -4482 -2990
rect -4528 -3258 -4522 -3002
rect -4488 -3258 -4482 -3002
rect -4528 -3270 -4482 -3258
rect -4350 -3002 -4304 -2990
rect -4350 -3258 -4344 -3002
rect -4310 -3258 -4304 -3002
rect -4350 -3270 -4304 -3258
rect -4172 -3002 -4126 -2990
rect -4172 -3258 -4166 -3002
rect -4132 -3258 -4126 -3002
rect -4172 -3270 -4126 -3258
rect -3994 -3002 -3948 -2990
rect -3994 -3258 -3988 -3002
rect -3954 -3258 -3948 -3002
rect -3994 -3270 -3948 -3258
rect -3816 -3002 -3770 -2990
rect -3816 -3258 -3810 -3002
rect -3776 -3258 -3770 -3002
rect -3816 -3270 -3770 -3258
rect -3638 -3002 -3592 -2990
rect -3638 -3258 -3632 -3002
rect -3598 -3258 -3592 -3002
rect -3638 -3270 -3592 -3258
rect -3460 -3002 -3414 -2990
rect -3460 -3258 -3454 -3002
rect -3420 -3258 -3414 -3002
rect -3460 -3270 -3414 -3258
rect -6234 -3317 -6158 -3311
rect -6234 -3351 -6218 -3317
rect -6174 -3351 -6158 -3317
rect -6234 -3367 -6158 -3351
rect -6124 -3401 -6090 -3270
rect -6056 -3317 -5980 -3311
rect -6056 -3351 -6040 -3317
rect -5996 -3351 -5980 -3317
rect -6056 -3367 -5980 -3351
rect -6144 -3454 -6134 -3401
rect -6081 -3454 -6071 -3401
rect -6508 -3693 -6498 -3640
rect -6445 -3693 -6435 -3640
rect -6498 -4271 -6445 -3693
rect -6035 -3763 -6001 -3367
rect -6234 -3778 -6158 -3763
rect -6302 -3779 -6090 -3778
rect -6302 -3812 -6218 -3779
rect -6302 -3860 -6268 -3812
rect -6234 -3813 -6218 -3812
rect -6174 -3812 -6090 -3779
rect -6174 -3813 -6158 -3812
rect -6234 -3819 -6158 -3813
rect -6124 -3860 -6090 -3812
rect -6056 -3779 -5980 -3763
rect -6056 -3813 -6040 -3779
rect -5996 -3813 -5980 -3779
rect -6056 -3819 -5980 -3813
rect -5946 -3860 -5912 -3270
rect -5878 -3317 -5802 -3311
rect -5878 -3351 -5862 -3317
rect -5818 -3351 -5802 -3317
rect -5878 -3367 -5802 -3351
rect -5857 -3763 -5823 -3367
rect -5768 -3516 -5734 -3270
rect -5700 -3317 -5624 -3311
rect -5700 -3351 -5684 -3317
rect -5640 -3351 -5624 -3317
rect -5700 -3367 -5624 -3351
rect -5787 -3569 -5777 -3516
rect -5724 -3569 -5714 -3516
rect -5679 -3763 -5645 -3367
rect -5878 -3779 -5802 -3763
rect -5878 -3813 -5862 -3779
rect -5818 -3813 -5802 -3779
rect -5878 -3819 -5802 -3813
rect -5700 -3779 -5624 -3763
rect -5700 -3813 -5684 -3779
rect -5640 -3813 -5624 -3779
rect -5700 -3819 -5624 -3813
rect -5590 -3860 -5556 -3270
rect -5522 -3317 -5446 -3311
rect -5522 -3351 -5506 -3317
rect -5462 -3351 -5446 -3317
rect -5522 -3367 -5446 -3351
rect -5501 -3763 -5467 -3367
rect -5412 -3640 -5378 -3270
rect -5344 -3317 -5268 -3311
rect -5344 -3351 -5328 -3317
rect -5284 -3351 -5268 -3317
rect -5344 -3367 -5268 -3351
rect -5432 -3693 -5422 -3640
rect -5369 -3693 -5359 -3640
rect -5323 -3763 -5289 -3367
rect -5522 -3779 -5446 -3763
rect -5522 -3813 -5506 -3779
rect -5462 -3813 -5446 -3779
rect -5522 -3819 -5446 -3813
rect -5344 -3779 -5268 -3763
rect -5344 -3813 -5328 -3779
rect -5284 -3813 -5268 -3779
rect -5344 -3819 -5268 -3813
rect -5234 -3860 -5200 -3270
rect -5166 -3317 -5090 -3311
rect -5166 -3351 -5150 -3317
rect -5106 -3351 -5090 -3317
rect -5166 -3367 -5090 -3351
rect -5145 -3763 -5111 -3367
rect -5056 -3401 -5022 -3270
rect -4988 -3317 -4912 -3311
rect -4988 -3351 -4972 -3317
rect -4928 -3351 -4912 -3317
rect -4988 -3367 -4912 -3351
rect -5076 -3454 -5066 -3401
rect -5013 -3454 -5003 -3401
rect -4967 -3763 -4933 -3367
rect -5166 -3779 -5090 -3763
rect -5166 -3813 -5150 -3779
rect -5106 -3813 -5090 -3779
rect -5166 -3819 -5090 -3813
rect -4988 -3779 -4912 -3763
rect -4988 -3813 -4972 -3779
rect -4928 -3813 -4912 -3779
rect -4988 -3819 -4912 -3813
rect -4878 -3860 -4844 -3270
rect -4810 -3317 -4734 -3311
rect -4810 -3351 -4794 -3317
rect -4750 -3351 -4734 -3317
rect -4810 -3367 -4734 -3351
rect -4789 -3763 -4755 -3367
rect -4700 -3401 -4666 -3270
rect -4632 -3317 -4556 -3311
rect -4632 -3351 -4616 -3317
rect -4572 -3351 -4556 -3317
rect -4632 -3367 -4556 -3351
rect -4720 -3454 -4710 -3401
rect -4657 -3454 -4647 -3401
rect -4611 -3763 -4577 -3367
rect -4810 -3779 -4734 -3763
rect -4810 -3813 -4794 -3779
rect -4750 -3813 -4734 -3779
rect -4810 -3819 -4734 -3813
rect -4632 -3779 -4556 -3763
rect -4632 -3813 -4616 -3779
rect -4572 -3813 -4556 -3779
rect -4632 -3819 -4556 -3813
rect -4522 -3860 -4488 -3270
rect -4454 -3317 -4378 -3311
rect -4454 -3351 -4438 -3317
rect -4394 -3351 -4378 -3317
rect -4454 -3367 -4378 -3351
rect -4433 -3763 -4399 -3367
rect -4344 -3640 -4310 -3270
rect -4276 -3317 -4200 -3311
rect -4276 -3351 -4260 -3317
rect -4216 -3351 -4200 -3317
rect -4276 -3367 -4200 -3351
rect -4363 -3693 -4353 -3640
rect -4300 -3693 -4290 -3640
rect -4254 -3763 -4220 -3367
rect -4454 -3779 -4378 -3763
rect -4454 -3813 -4438 -3779
rect -4394 -3813 -4378 -3779
rect -4454 -3819 -4378 -3813
rect -4276 -3779 -4200 -3763
rect -4276 -3813 -4260 -3779
rect -4216 -3813 -4200 -3779
rect -4276 -3819 -4200 -3813
rect -4166 -3860 -4132 -3270
rect -4098 -3317 -4022 -3311
rect -4098 -3351 -4082 -3317
rect -4038 -3351 -4022 -3317
rect -4098 -3367 -4022 -3351
rect -4077 -3763 -4043 -3367
rect -3988 -3516 -3954 -3270
rect -3920 -3317 -3844 -3311
rect -3920 -3351 -3904 -3317
rect -3860 -3351 -3844 -3317
rect -3920 -3367 -3844 -3351
rect -4008 -3569 -3998 -3516
rect -3945 -3569 -3935 -3516
rect -3899 -3763 -3865 -3367
rect -4098 -3779 -4022 -3763
rect -4098 -3813 -4082 -3779
rect -4038 -3813 -4022 -3779
rect -4098 -3819 -4022 -3813
rect -3920 -3779 -3844 -3763
rect -3920 -3813 -3904 -3779
rect -3860 -3813 -3844 -3779
rect -3920 -3819 -3844 -3813
rect -3810 -3860 -3776 -3270
rect -3742 -3317 -3666 -3311
rect -3742 -3351 -3726 -3317
rect -3682 -3351 -3666 -3317
rect -3742 -3367 -3666 -3351
rect -3632 -3316 -3598 -3270
rect -3564 -3316 -3488 -3311
rect -3454 -3316 -3420 -3270
rect -3632 -3317 -3420 -3316
rect -3632 -3350 -3548 -3317
rect -3721 -3763 -3687 -3367
rect -3632 -3401 -3598 -3350
rect -3564 -3351 -3548 -3350
rect -3504 -3350 -3420 -3317
rect -3504 -3351 -3488 -3350
rect -3564 -3367 -3488 -3351
rect -3652 -3454 -3642 -3401
rect -3589 -3454 -3579 -3401
rect -3298 -3516 -3245 -2721
rect -3141 -3454 -3131 -3401
rect -3078 -3454 -3068 -3401
rect -3308 -3569 -3298 -3516
rect -3245 -3569 -3235 -3516
rect -3742 -3779 -3666 -3763
rect -3742 -3813 -3726 -3779
rect -3682 -3813 -3666 -3779
rect -3742 -3819 -3666 -3813
rect -3564 -3779 -3488 -3763
rect -3564 -3813 -3548 -3779
rect -3504 -3813 -3488 -3779
rect -3564 -3819 -3488 -3813
rect -6308 -3872 -6262 -3860
rect -6308 -4128 -6302 -3872
rect -6268 -4128 -6262 -3872
rect -6308 -4140 -6262 -4128
rect -6130 -3872 -6084 -3860
rect -6130 -4128 -6124 -3872
rect -6090 -4128 -6084 -3872
rect -6130 -4140 -6084 -4128
rect -5952 -3872 -5906 -3860
rect -5952 -4128 -5946 -3872
rect -5912 -4128 -5906 -3872
rect -5952 -4140 -5906 -4128
rect -5774 -3872 -5728 -3860
rect -5774 -4128 -5768 -3872
rect -5734 -4128 -5728 -3872
rect -5774 -4140 -5728 -4128
rect -5596 -3872 -5550 -3860
rect -5596 -4128 -5590 -3872
rect -5556 -4128 -5550 -3872
rect -5596 -4140 -5550 -4128
rect -5418 -3872 -5372 -3860
rect -5418 -4128 -5412 -3872
rect -5378 -4128 -5372 -3872
rect -5418 -4140 -5372 -4128
rect -5240 -3872 -5194 -3860
rect -5240 -4128 -5234 -3872
rect -5200 -4128 -5194 -3872
rect -5240 -4140 -5194 -4128
rect -5062 -3872 -5016 -3860
rect -5062 -4128 -5056 -3872
rect -5022 -4128 -5016 -3872
rect -5062 -4140 -5016 -4128
rect -4884 -3872 -4838 -3860
rect -4884 -4128 -4878 -3872
rect -4844 -4128 -4838 -3872
rect -4884 -4140 -4838 -4128
rect -4706 -3872 -4660 -3860
rect -4706 -4128 -4700 -3872
rect -4666 -4128 -4660 -3872
rect -4706 -4140 -4660 -4128
rect -4528 -3872 -4482 -3860
rect -4528 -4128 -4522 -3872
rect -4488 -4128 -4482 -3872
rect -4528 -4140 -4482 -4128
rect -4350 -3872 -4304 -3860
rect -4350 -4128 -4344 -3872
rect -4310 -4128 -4304 -3872
rect -4350 -4140 -4304 -4128
rect -4172 -3872 -4126 -3860
rect -4172 -4128 -4166 -3872
rect -4132 -4128 -4126 -3872
rect -4172 -4140 -4126 -4128
rect -3994 -3872 -3948 -3860
rect -3994 -4128 -3988 -3872
rect -3954 -4128 -3948 -3872
rect -3994 -4140 -3948 -4128
rect -3816 -3872 -3770 -3860
rect -3816 -4128 -3810 -3872
rect -3776 -4128 -3770 -3872
rect -3816 -4140 -3770 -4128
rect -3638 -3872 -3592 -3860
rect -3638 -4128 -3632 -3872
rect -3598 -4128 -3592 -3872
rect -3638 -4140 -3592 -4128
rect -3460 -3872 -3414 -3860
rect -3460 -4128 -3454 -3872
rect -3420 -4128 -3414 -3872
rect -3460 -4140 -3414 -4128
rect -6234 -4187 -6158 -4181
rect -6234 -4221 -6218 -4187
rect -6174 -4221 -6158 -4187
rect -6234 -4237 -6158 -4221
rect -6508 -4324 -6498 -4271
rect -6445 -4324 -6435 -4271
rect -6498 -5141 -6445 -4324
rect -6124 -4390 -6090 -4140
rect -6056 -4187 -5980 -4181
rect -6056 -4221 -6040 -4187
rect -5996 -4221 -5980 -4187
rect -6056 -4237 -5980 -4221
rect -6144 -4443 -6134 -4390
rect -6081 -4443 -6071 -4390
rect -6035 -4633 -6001 -4237
rect -6234 -4649 -6158 -4633
rect -6056 -4649 -5980 -4633
rect -6302 -4683 -6218 -4649
rect -6174 -4683 -6090 -4649
rect -6302 -4730 -6268 -4683
rect -6234 -4689 -6158 -4683
rect -6124 -4730 -6090 -4683
rect -6056 -4683 -6040 -4649
rect -5996 -4683 -5980 -4649
rect -6056 -4689 -5980 -4683
rect -5946 -4730 -5912 -4140
rect -5878 -4187 -5802 -4181
rect -5878 -4221 -5862 -4187
rect -5818 -4221 -5802 -4187
rect -5878 -4237 -5802 -4221
rect -5857 -4633 -5823 -4237
rect -5768 -4271 -5734 -4140
rect -5700 -4187 -5624 -4181
rect -5700 -4221 -5684 -4187
rect -5640 -4221 -5624 -4187
rect -5700 -4237 -5624 -4221
rect -5788 -4324 -5778 -4271
rect -5725 -4324 -5715 -4271
rect -5679 -4633 -5645 -4237
rect -5878 -4649 -5802 -4633
rect -5878 -4683 -5862 -4649
rect -5818 -4683 -5802 -4649
rect -5878 -4689 -5802 -4683
rect -5700 -4649 -5624 -4633
rect -5700 -4683 -5684 -4649
rect -5640 -4683 -5624 -4649
rect -5700 -4689 -5624 -4683
rect -5590 -4730 -5556 -4140
rect -5522 -4187 -5446 -4181
rect -5522 -4221 -5506 -4187
rect -5462 -4221 -5446 -4187
rect -5522 -4237 -5446 -4221
rect -5501 -4633 -5467 -4237
rect -5412 -4506 -5378 -4140
rect -5344 -4187 -5268 -4181
rect -5344 -4221 -5328 -4187
rect -5284 -4221 -5268 -4187
rect -5344 -4237 -5268 -4221
rect -5432 -4559 -5422 -4506
rect -5369 -4559 -5359 -4506
rect -5323 -4633 -5289 -4237
rect -5522 -4649 -5446 -4633
rect -5522 -4683 -5506 -4649
rect -5462 -4683 -5446 -4649
rect -5522 -4689 -5446 -4683
rect -5344 -4649 -5268 -4633
rect -5344 -4683 -5328 -4649
rect -5284 -4683 -5268 -4649
rect -5344 -4689 -5268 -4683
rect -5234 -4730 -5200 -4140
rect -5166 -4187 -5090 -4181
rect -5166 -4221 -5150 -4187
rect -5106 -4221 -5090 -4187
rect -5166 -4237 -5090 -4221
rect -5145 -4633 -5111 -4237
rect -5056 -4390 -5022 -4140
rect -4988 -4187 -4912 -4181
rect -4988 -4221 -4972 -4187
rect -4928 -4221 -4912 -4187
rect -4988 -4237 -4912 -4221
rect -5076 -4443 -5066 -4390
rect -5013 -4443 -5003 -4390
rect -4967 -4633 -4933 -4237
rect -5166 -4649 -5090 -4633
rect -5166 -4683 -5150 -4649
rect -5106 -4683 -5090 -4649
rect -5166 -4689 -5090 -4683
rect -4988 -4649 -4912 -4633
rect -4988 -4683 -4972 -4649
rect -4928 -4683 -4912 -4649
rect -4988 -4689 -4912 -4683
rect -4878 -4730 -4844 -4140
rect -4810 -4187 -4734 -4181
rect -4810 -4221 -4794 -4187
rect -4750 -4221 -4734 -4187
rect -4810 -4237 -4734 -4221
rect -4789 -4633 -4755 -4237
rect -4700 -4390 -4666 -4140
rect -4632 -4187 -4556 -4181
rect -4632 -4221 -4616 -4187
rect -4572 -4221 -4556 -4187
rect -4632 -4237 -4556 -4221
rect -4719 -4443 -4709 -4390
rect -4656 -4443 -4646 -4390
rect -4611 -4633 -4577 -4237
rect -4810 -4649 -4734 -4633
rect -4810 -4683 -4794 -4649
rect -4750 -4683 -4734 -4649
rect -4810 -4689 -4734 -4683
rect -4632 -4649 -4556 -4633
rect -4632 -4683 -4616 -4649
rect -4572 -4683 -4556 -4649
rect -4632 -4689 -4556 -4683
rect -4522 -4730 -4488 -4140
rect -4454 -4187 -4378 -4181
rect -4454 -4221 -4438 -4187
rect -4394 -4221 -4378 -4187
rect -4454 -4237 -4378 -4221
rect -4433 -4633 -4399 -4237
rect -4344 -4506 -4310 -4140
rect -4276 -4187 -4200 -4181
rect -4276 -4221 -4260 -4187
rect -4216 -4221 -4200 -4187
rect -4276 -4237 -4200 -4221
rect -4363 -4559 -4353 -4506
rect -4300 -4559 -4290 -4506
rect -4255 -4633 -4221 -4237
rect -4454 -4649 -4378 -4633
rect -4454 -4683 -4438 -4649
rect -4394 -4683 -4378 -4649
rect -4454 -4689 -4378 -4683
rect -4276 -4649 -4200 -4633
rect -4276 -4683 -4260 -4649
rect -4216 -4683 -4200 -4649
rect -4276 -4689 -4200 -4683
rect -4166 -4730 -4132 -4140
rect -4098 -4187 -4022 -4181
rect -4098 -4221 -4082 -4187
rect -4038 -4221 -4022 -4187
rect -4098 -4237 -4022 -4221
rect -4077 -4633 -4043 -4237
rect -3988 -4271 -3954 -4140
rect -3920 -4187 -3844 -4181
rect -3920 -4221 -3904 -4187
rect -3860 -4221 -3844 -4187
rect -3920 -4237 -3844 -4221
rect -4008 -4324 -3998 -4271
rect -3945 -4324 -3935 -4271
rect -3899 -4633 -3865 -4237
rect -4098 -4649 -4022 -4633
rect -4098 -4683 -4082 -4649
rect -4038 -4683 -4022 -4649
rect -4098 -4689 -4022 -4683
rect -3920 -4649 -3844 -4633
rect -3920 -4683 -3904 -4649
rect -3860 -4683 -3844 -4649
rect -3920 -4689 -3844 -4683
rect -3810 -4730 -3776 -4140
rect -3742 -4187 -3666 -4181
rect -3742 -4221 -3726 -4187
rect -3682 -4221 -3666 -4187
rect -3742 -4237 -3666 -4221
rect -3632 -4186 -3598 -4140
rect -3564 -4186 -3488 -4181
rect -3453 -4186 -3419 -4140
rect -3632 -4187 -3419 -4186
rect -3632 -4220 -3548 -4187
rect -3721 -4633 -3687 -4237
rect -3632 -4390 -3598 -4220
rect -3564 -4221 -3548 -4220
rect -3504 -4220 -3419 -4187
rect -3504 -4221 -3488 -4220
rect -3564 -4237 -3488 -4221
rect -3652 -4443 -3642 -4390
rect -3589 -4443 -3579 -4390
rect -3298 -4506 -3245 -3569
rect -3308 -4559 -3298 -4506
rect -3245 -4559 -3235 -4506
rect -3742 -4649 -3666 -4633
rect -3742 -4683 -3726 -4649
rect -3682 -4683 -3666 -4649
rect -3742 -4689 -3666 -4683
rect -3564 -4649 -3488 -4633
rect -3564 -4683 -3548 -4649
rect -3504 -4683 -3488 -4649
rect -3564 -4689 -3488 -4683
rect -6308 -4742 -6262 -4730
rect -6308 -4998 -6302 -4742
rect -6268 -4998 -6262 -4742
rect -6308 -5010 -6262 -4998
rect -6130 -4742 -6084 -4730
rect -6130 -4998 -6124 -4742
rect -6090 -4998 -6084 -4742
rect -6130 -5010 -6084 -4998
rect -5952 -4742 -5906 -4730
rect -5952 -4998 -5946 -4742
rect -5912 -4998 -5906 -4742
rect -5952 -5010 -5906 -4998
rect -5774 -4742 -5728 -4730
rect -5774 -4998 -5768 -4742
rect -5734 -4998 -5728 -4742
rect -5774 -5010 -5728 -4998
rect -5596 -4742 -5550 -4730
rect -5596 -4998 -5590 -4742
rect -5556 -4998 -5550 -4742
rect -5596 -5010 -5550 -4998
rect -5418 -4742 -5372 -4730
rect -5418 -4998 -5412 -4742
rect -5378 -4998 -5372 -4742
rect -5418 -5010 -5372 -4998
rect -5240 -4742 -5194 -4730
rect -5240 -4998 -5234 -4742
rect -5200 -4998 -5194 -4742
rect -5240 -5010 -5194 -4998
rect -5062 -4742 -5016 -4730
rect -5062 -4998 -5056 -4742
rect -5022 -4998 -5016 -4742
rect -5062 -5010 -5016 -4998
rect -4884 -4742 -4838 -4730
rect -4884 -4998 -4878 -4742
rect -4844 -4998 -4838 -4742
rect -4884 -5010 -4838 -4998
rect -4706 -4742 -4660 -4730
rect -4706 -4998 -4700 -4742
rect -4666 -4998 -4660 -4742
rect -4706 -5010 -4660 -4998
rect -4528 -4742 -4482 -4730
rect -4528 -4998 -4522 -4742
rect -4488 -4998 -4482 -4742
rect -4528 -5010 -4482 -4998
rect -4350 -4742 -4304 -4730
rect -4350 -4998 -4344 -4742
rect -4310 -4998 -4304 -4742
rect -4350 -5010 -4304 -4998
rect -4172 -4742 -4126 -4730
rect -4172 -4998 -4166 -4742
rect -4132 -4998 -4126 -4742
rect -4172 -5010 -4126 -4998
rect -3994 -4742 -3948 -4730
rect -3994 -4998 -3988 -4742
rect -3954 -4998 -3948 -4742
rect -3994 -5010 -3948 -4998
rect -3816 -4742 -3770 -4730
rect -3816 -4998 -3810 -4742
rect -3776 -4998 -3770 -4742
rect -3816 -5010 -3770 -4998
rect -3638 -4742 -3592 -4730
rect -3638 -4998 -3632 -4742
rect -3598 -4998 -3592 -4742
rect -3638 -5010 -3592 -4998
rect -3460 -4742 -3414 -4730
rect -3460 -4998 -3454 -4742
rect -3420 -4998 -3414 -4742
rect -3460 -5010 -3414 -4998
rect -6234 -5057 -6158 -5051
rect -6234 -5091 -6218 -5057
rect -6174 -5091 -6158 -5057
rect -6234 -5107 -6158 -5091
rect -6508 -5194 -6498 -5141
rect -6445 -5194 -6435 -5141
rect -6635 -5375 -6625 -5322
rect -6572 -5375 -6562 -5322
rect -6498 -6248 -6445 -5194
rect -6124 -5232 -6090 -5010
rect -6056 -5057 -5980 -5051
rect -6056 -5091 -6040 -5057
rect -5996 -5091 -5980 -5057
rect -6056 -5107 -5980 -5091
rect -6144 -5285 -6134 -5232
rect -6081 -5285 -6071 -5232
rect -6234 -5518 -6158 -5503
rect -6301 -5519 -6091 -5518
rect -6056 -5519 -5980 -5503
rect -5946 -5519 -5912 -5010
rect -5878 -5057 -5802 -5051
rect -5878 -5091 -5862 -5057
rect -5818 -5091 -5802 -5057
rect -5878 -5107 -5802 -5091
rect -5857 -5503 -5823 -5107
rect -5768 -5415 -5734 -5010
rect -5700 -5057 -5624 -5051
rect -5700 -5091 -5684 -5057
rect -5640 -5091 -5624 -5057
rect -5700 -5107 -5624 -5091
rect -5787 -5468 -5777 -5415
rect -5724 -5468 -5714 -5415
rect -5679 -5503 -5645 -5107
rect -6301 -5552 -6218 -5519
rect -6301 -5600 -6267 -5552
rect -6234 -5553 -6218 -5552
rect -6174 -5552 -6040 -5519
rect -6174 -5553 -6158 -5552
rect -6234 -5559 -6158 -5553
rect -6125 -5553 -6040 -5552
rect -5996 -5553 -5912 -5519
rect -6125 -5600 -6091 -5553
rect -6056 -5559 -5980 -5553
rect -5946 -5600 -5912 -5553
rect -5878 -5519 -5802 -5503
rect -5878 -5553 -5862 -5519
rect -5818 -5553 -5802 -5519
rect -5878 -5559 -5802 -5553
rect -5700 -5519 -5624 -5503
rect -5700 -5553 -5684 -5519
rect -5640 -5553 -5624 -5519
rect -5700 -5559 -5624 -5553
rect -5590 -5600 -5556 -5010
rect -5522 -5057 -5446 -5051
rect -5522 -5091 -5506 -5057
rect -5462 -5091 -5446 -5057
rect -5522 -5107 -5446 -5091
rect -5501 -5503 -5467 -5107
rect -5412 -5141 -5378 -5010
rect -5344 -5057 -5268 -5051
rect -5344 -5091 -5328 -5057
rect -5284 -5091 -5268 -5057
rect -5344 -5107 -5268 -5091
rect -5432 -5194 -5422 -5141
rect -5369 -5194 -5359 -5141
rect -5323 -5503 -5289 -5107
rect -5522 -5519 -5446 -5503
rect -5522 -5553 -5506 -5519
rect -5462 -5553 -5446 -5519
rect -5522 -5559 -5446 -5553
rect -5344 -5519 -5268 -5503
rect -5344 -5553 -5328 -5519
rect -5284 -5553 -5268 -5519
rect -5344 -5559 -5268 -5553
rect -5234 -5600 -5200 -5010
rect -5166 -5057 -5090 -5051
rect -5166 -5091 -5150 -5057
rect -5106 -5091 -5090 -5057
rect -5166 -5107 -5090 -5091
rect -5145 -5503 -5111 -5107
rect -5056 -5233 -5022 -5010
rect -4988 -5057 -4912 -5051
rect -4988 -5091 -4972 -5057
rect -4928 -5091 -4912 -5057
rect -4988 -5107 -4912 -5091
rect -5076 -5286 -5066 -5233
rect -5013 -5286 -5003 -5233
rect -4967 -5503 -4933 -5107
rect -5166 -5519 -5090 -5503
rect -5166 -5553 -5150 -5519
rect -5106 -5553 -5090 -5519
rect -5166 -5559 -5090 -5553
rect -4988 -5519 -4912 -5503
rect -4988 -5553 -4972 -5519
rect -4928 -5553 -4912 -5519
rect -4988 -5559 -4912 -5553
rect -4878 -5600 -4844 -5010
rect -4810 -5057 -4734 -5051
rect -4810 -5091 -4794 -5057
rect -4750 -5091 -4734 -5057
rect -4810 -5107 -4734 -5091
rect -4789 -5503 -4755 -5107
rect -4700 -5322 -4666 -5010
rect -4632 -5057 -4556 -5051
rect -4632 -5091 -4616 -5057
rect -4572 -5091 -4556 -5057
rect -4632 -5107 -4556 -5091
rect -4720 -5375 -4710 -5322
rect -4657 -5375 -4647 -5322
rect -4611 -5503 -4577 -5107
rect -4810 -5519 -4734 -5503
rect -4810 -5553 -4794 -5519
rect -4750 -5553 -4734 -5519
rect -4810 -5559 -4734 -5553
rect -4632 -5519 -4556 -5503
rect -4632 -5553 -4616 -5519
rect -4572 -5553 -4556 -5519
rect -4632 -5559 -4556 -5553
rect -4522 -5600 -4488 -5010
rect -4454 -5057 -4378 -5051
rect -4454 -5091 -4438 -5057
rect -4394 -5091 -4378 -5057
rect -4454 -5107 -4378 -5091
rect -4433 -5503 -4399 -5107
rect -4344 -5141 -4310 -5010
rect -4276 -5057 -4200 -5051
rect -4276 -5091 -4260 -5057
rect -4216 -5091 -4200 -5057
rect -4276 -5107 -4200 -5091
rect -4363 -5194 -4353 -5141
rect -4300 -5194 -4290 -5141
rect -4255 -5503 -4221 -5107
rect -4454 -5519 -4378 -5503
rect -4454 -5553 -4438 -5519
rect -4394 -5553 -4378 -5519
rect -4454 -5559 -4378 -5553
rect -4276 -5519 -4200 -5503
rect -4276 -5553 -4260 -5519
rect -4216 -5553 -4200 -5519
rect -4276 -5559 -4200 -5553
rect -4166 -5600 -4132 -5010
rect -4098 -5057 -4022 -5051
rect -4098 -5091 -4082 -5057
rect -4038 -5091 -4022 -5057
rect -4098 -5107 -4022 -5091
rect -4077 -5503 -4043 -5107
rect -3988 -5415 -3954 -5010
rect -3920 -5057 -3844 -5051
rect -3920 -5091 -3904 -5057
rect -3860 -5091 -3844 -5057
rect -3920 -5107 -3844 -5091
rect -4007 -5468 -3997 -5415
rect -3944 -5468 -3934 -5415
rect -3899 -5503 -3865 -5107
rect -4098 -5519 -4022 -5503
rect -4098 -5553 -4082 -5519
rect -4038 -5553 -4022 -5519
rect -4098 -5559 -4022 -5553
rect -3920 -5519 -3844 -5503
rect -3920 -5553 -3904 -5519
rect -3860 -5553 -3844 -5519
rect -3920 -5559 -3844 -5553
rect -3810 -5600 -3776 -5010
rect -3742 -5057 -3666 -5051
rect -3742 -5091 -3726 -5057
rect -3682 -5091 -3666 -5057
rect -3742 -5107 -3666 -5091
rect -3632 -5056 -3598 -5010
rect -3564 -5056 -3488 -5051
rect -3453 -5056 -3419 -5010
rect -3632 -5057 -3419 -5056
rect -3632 -5090 -3548 -5057
rect -3632 -5319 -3598 -5090
rect -3564 -5091 -3548 -5090
rect -3504 -5090 -3419 -5057
rect -3504 -5091 -3488 -5090
rect -3564 -5107 -3488 -5091
rect -3652 -5372 -3642 -5319
rect -3589 -5372 -3579 -5319
rect -3298 -5416 -3245 -4559
rect -3130 -5233 -3077 -3454
rect -3140 -5286 -3130 -5233
rect -3077 -5286 -3067 -5233
rect -2624 -5324 -2571 -2611
rect -1386 -2791 -1310 -2775
rect -1386 -2825 -1370 -2791
rect -1326 -2825 -1310 -2791
rect -1386 -2831 -1310 -2825
rect -1276 -2872 -1242 -2611
rect -1207 -2718 -1197 -2665
rect -1144 -2718 -1134 -2665
rect -1187 -2775 -1153 -2718
rect -1208 -2791 -1132 -2775
rect -1208 -2825 -1192 -2791
rect -1148 -2825 -1132 -2791
rect -1208 -2831 -1132 -2825
rect -1099 -2872 -1065 -2478
rect -940 -2611 -930 -2558
rect -877 -2611 -867 -2558
rect -1029 -2718 -1019 -2665
rect -966 -2718 -956 -2665
rect -1009 -2775 -975 -2718
rect -1030 -2791 -954 -2775
rect -1030 -2825 -1014 -2791
rect -970 -2825 -954 -2791
rect -1030 -2831 -954 -2825
rect -920 -2872 -886 -2611
rect -851 -2718 -841 -2665
rect -788 -2718 -778 -2665
rect -831 -2775 -797 -2718
rect -852 -2791 -776 -2775
rect -852 -2825 -836 -2791
rect -792 -2825 -776 -2791
rect -852 -2831 -776 -2825
rect -742 -2872 -708 -2478
rect -208 -2605 182 -2571
rect -674 -2791 -598 -2775
rect -674 -2825 -658 -2791
rect -614 -2825 -598 -2791
rect -674 -2831 -598 -2825
rect -496 -2791 -420 -2775
rect -496 -2825 -480 -2791
rect -436 -2825 -420 -2791
rect -496 -2831 -420 -2825
rect -318 -2791 -242 -2775
rect -318 -2825 -302 -2791
rect -258 -2825 -242 -2791
rect -318 -2831 -242 -2825
rect -208 -2872 -174 -2605
rect -139 -2718 -129 -2665
rect -76 -2718 -66 -2665
rect 40 -2718 50 -2665
rect 103 -2718 113 -2665
rect -119 -2775 -85 -2718
rect 59 -2775 93 -2718
rect -140 -2791 -64 -2775
rect -140 -2825 -124 -2791
rect -80 -2825 -64 -2791
rect -140 -2831 -64 -2825
rect 38 -2791 114 -2775
rect 38 -2825 54 -2791
rect 98 -2825 114 -2791
rect 38 -2831 114 -2825
rect 148 -2872 182 -2605
rect 217 -2718 227 -2665
rect 280 -2718 290 -2665
rect 237 -2775 271 -2718
rect 594 -2775 628 -1467
rect 1909 -2479 1919 -2426
rect 1972 -2479 1982 -2426
rect 2265 -2479 2275 -2426
rect 2328 -2479 2338 -2426
rect 1038 -2611 1428 -2577
rect 930 -2718 940 -2665
rect 993 -2718 1003 -2665
rect 949 -2775 983 -2718
rect 216 -2791 292 -2775
rect 216 -2825 232 -2791
rect 276 -2825 292 -2791
rect 216 -2831 292 -2825
rect 394 -2791 470 -2775
rect 394 -2825 410 -2791
rect 454 -2825 470 -2791
rect 394 -2831 470 -2825
rect 572 -2791 648 -2775
rect 572 -2825 588 -2791
rect 632 -2825 648 -2791
rect 572 -2831 648 -2825
rect 750 -2791 826 -2775
rect 750 -2825 766 -2791
rect 810 -2825 826 -2791
rect 750 -2831 826 -2825
rect 928 -2791 1004 -2775
rect 928 -2825 944 -2791
rect 988 -2825 1004 -2791
rect 928 -2831 1004 -2825
rect 1038 -2872 1072 -2611
rect 1107 -2718 1117 -2665
rect 1170 -2718 1180 -2665
rect 1285 -2718 1295 -2665
rect 1348 -2718 1358 -2665
rect 1127 -2775 1161 -2718
rect 1305 -2775 1339 -2718
rect 1106 -2791 1182 -2775
rect 1106 -2825 1122 -2791
rect 1166 -2825 1182 -2791
rect 1106 -2831 1182 -2825
rect 1284 -2791 1360 -2775
rect 1284 -2825 1300 -2791
rect 1344 -2825 1360 -2791
rect 1284 -2831 1360 -2825
rect 1394 -2872 1428 -2611
rect 1462 -2791 1538 -2775
rect 1462 -2825 1478 -2791
rect 1522 -2825 1538 -2791
rect 1462 -2831 1538 -2825
rect 1640 -2791 1716 -2775
rect 1640 -2825 1656 -2791
rect 1700 -2825 1716 -2791
rect 1640 -2831 1716 -2825
rect 1818 -2791 1894 -2775
rect 1818 -2825 1834 -2791
rect 1878 -2825 1894 -2791
rect 1818 -2831 1894 -2825
rect 1928 -2872 1962 -2479
rect 2087 -2607 2097 -2554
rect 2150 -2607 2160 -2554
rect 1997 -2718 2007 -2665
rect 2060 -2718 2070 -2665
rect 2017 -2775 2051 -2718
rect 1996 -2791 2072 -2775
rect 1996 -2825 2012 -2791
rect 2056 -2825 2072 -2791
rect 1996 -2831 2072 -2825
rect 2105 -2872 2139 -2607
rect 2176 -2718 2186 -2665
rect 2239 -2718 2249 -2665
rect 2195 -2775 2229 -2718
rect 2174 -2791 2250 -2775
rect 2174 -2825 2190 -2791
rect 2234 -2825 2250 -2791
rect 2174 -2831 2250 -2825
rect 2285 -2872 2319 -2479
rect 3183 -2480 3193 -2427
rect 3246 -2480 3256 -2427
rect 2443 -2607 2453 -2554
rect 2506 -2606 2931 -2554
rect 2506 -2607 2516 -2606
rect 2353 -2718 2363 -2665
rect 2416 -2718 2426 -2665
rect 2373 -2775 2407 -2718
rect 2352 -2791 2428 -2775
rect 2352 -2825 2368 -2791
rect 2412 -2825 2428 -2791
rect 2352 -2831 2428 -2825
rect 2462 -2872 2496 -2607
rect 2530 -2791 2606 -2775
rect 2530 -2825 2546 -2791
rect 2590 -2825 2606 -2791
rect 2530 -2831 2606 -2825
rect -1460 -2884 -1414 -2872
rect -1460 -3140 -1454 -2884
rect -1420 -3140 -1414 -2884
rect -1460 -3152 -1414 -3140
rect -1282 -2884 -1236 -2872
rect -1282 -3140 -1276 -2884
rect -1242 -3140 -1236 -2884
rect -1282 -3152 -1236 -3140
rect -1104 -2884 -1058 -2872
rect -1104 -3140 -1098 -2884
rect -1064 -3140 -1058 -2884
rect -1104 -3152 -1058 -3140
rect -926 -2884 -880 -2872
rect -926 -3140 -920 -2884
rect -886 -3140 -880 -2884
rect -926 -3152 -880 -3140
rect -748 -2884 -702 -2872
rect -748 -3140 -742 -2884
rect -708 -3140 -702 -2884
rect -748 -3152 -702 -3140
rect -570 -2884 -524 -2872
rect -570 -3140 -564 -2884
rect -530 -3140 -524 -2884
rect -570 -3152 -524 -3140
rect -392 -2884 -346 -2872
rect -392 -3140 -386 -2884
rect -352 -3140 -346 -2884
rect -392 -3152 -346 -3140
rect -214 -2884 -168 -2872
rect -214 -3140 -208 -2884
rect -174 -3140 -168 -2884
rect -214 -3152 -168 -3140
rect -36 -2884 10 -2872
rect -36 -3140 -30 -2884
rect 4 -3140 10 -2884
rect -36 -3152 10 -3140
rect 142 -2884 188 -2872
rect 142 -3140 148 -2884
rect 182 -3140 188 -2884
rect 142 -3152 188 -3140
rect 320 -2884 366 -2872
rect 320 -3140 326 -2884
rect 360 -3140 366 -2884
rect 320 -3152 366 -3140
rect 498 -2884 544 -2872
rect 498 -3140 504 -2884
rect 538 -3140 544 -2884
rect 498 -3152 544 -3140
rect 676 -2884 722 -2872
rect 676 -3140 682 -2884
rect 716 -3140 722 -2884
rect 676 -3152 722 -3140
rect 854 -2884 900 -2872
rect 854 -3140 860 -2884
rect 894 -3140 900 -2884
rect 854 -3152 900 -3140
rect 1032 -2884 1078 -2872
rect 1032 -3140 1038 -2884
rect 1072 -3140 1078 -2884
rect 1032 -3152 1078 -3140
rect 1210 -2884 1256 -2872
rect 1210 -3140 1216 -2884
rect 1250 -3140 1256 -2884
rect 1210 -3152 1256 -3140
rect 1388 -2884 1434 -2872
rect 1388 -3140 1394 -2884
rect 1428 -3140 1434 -2884
rect 1388 -3152 1434 -3140
rect 1566 -2884 1612 -2872
rect 1566 -3140 1572 -2884
rect 1606 -3140 1612 -2884
rect 1566 -3152 1612 -3140
rect 1744 -2884 1790 -2872
rect 1744 -3140 1750 -2884
rect 1784 -3140 1790 -2884
rect 1744 -3152 1790 -3140
rect 1922 -2884 1968 -2872
rect 1922 -3140 1928 -2884
rect 1962 -3140 1968 -2884
rect 1922 -3152 1968 -3140
rect 2100 -2884 2146 -2872
rect 2100 -3140 2106 -2884
rect 2140 -3140 2146 -2884
rect 2100 -3152 2146 -3140
rect 2278 -2884 2324 -2872
rect 2278 -3140 2284 -2884
rect 2318 -3140 2324 -2884
rect 2278 -3152 2324 -3140
rect 2456 -2884 2502 -2872
rect 2456 -3140 2462 -2884
rect 2496 -3140 2502 -2884
rect 2456 -3152 2502 -3140
rect 2634 -2884 2680 -2872
rect 2634 -3140 2640 -2884
rect 2674 -3140 2680 -2884
rect 2634 -3152 2680 -3140
rect -1454 -3282 -1420 -3152
rect -1386 -3199 -1310 -3193
rect -1386 -3233 -1370 -3199
rect -1326 -3233 -1310 -3199
rect -1386 -3249 -1310 -3233
rect -1365 -3282 -1331 -3249
rect -1276 -3282 -1242 -3152
rect -1208 -3199 -1132 -3193
rect -1208 -3233 -1192 -3199
rect -1148 -3233 -1132 -3199
rect -1208 -3249 -1132 -3233
rect -1030 -3199 -954 -3193
rect -1030 -3233 -1014 -3199
rect -970 -3233 -954 -3199
rect -1030 -3249 -954 -3233
rect -852 -3199 -776 -3193
rect -852 -3233 -836 -3199
rect -792 -3233 -776 -3199
rect -852 -3249 -776 -3233
rect -674 -3199 -598 -3193
rect -674 -3233 -658 -3199
rect -614 -3233 -598 -3199
rect -674 -3249 -598 -3233
rect -1454 -3316 -1242 -3282
rect -1454 -3317 -1420 -3316
rect -1655 -3510 -1645 -3449
rect -1584 -3510 -1574 -3449
rect -2014 -4465 -2004 -4412
rect -1951 -4465 -1941 -4412
rect -2003 -4517 -1950 -4465
rect -2634 -5377 -2624 -5324
rect -2571 -5377 -2561 -5324
rect -3308 -5469 -3298 -5416
rect -3245 -5469 -3235 -5416
rect -3742 -5519 -3666 -5503
rect -3742 -5553 -3726 -5519
rect -3682 -5553 -3666 -5519
rect -3742 -5559 -3666 -5553
rect -3564 -5519 -3488 -5503
rect -3564 -5553 -3548 -5519
rect -3504 -5553 -3488 -5519
rect -3564 -5559 -3488 -5553
rect -6308 -5612 -6262 -5600
rect -6308 -5868 -6302 -5612
rect -6268 -5868 -6262 -5612
rect -6308 -5880 -6262 -5868
rect -6130 -5612 -6084 -5600
rect -6130 -5868 -6124 -5612
rect -6090 -5868 -6084 -5612
rect -6130 -5880 -6084 -5868
rect -5952 -5612 -5906 -5600
rect -5952 -5868 -5946 -5612
rect -5912 -5868 -5906 -5612
rect -5952 -5880 -5906 -5868
rect -5774 -5612 -5728 -5600
rect -5774 -5868 -5768 -5612
rect -5734 -5868 -5728 -5612
rect -5774 -5880 -5728 -5868
rect -5596 -5612 -5550 -5600
rect -5596 -5868 -5590 -5612
rect -5556 -5868 -5550 -5612
rect -5596 -5880 -5550 -5868
rect -5418 -5612 -5372 -5600
rect -5418 -5868 -5412 -5612
rect -5378 -5868 -5372 -5612
rect -5418 -5880 -5372 -5868
rect -5240 -5612 -5194 -5600
rect -5240 -5868 -5234 -5612
rect -5200 -5868 -5194 -5612
rect -5240 -5880 -5194 -5868
rect -5062 -5612 -5016 -5600
rect -5062 -5868 -5056 -5612
rect -5022 -5868 -5016 -5612
rect -5062 -5880 -5016 -5868
rect -4884 -5612 -4838 -5600
rect -4884 -5868 -4878 -5612
rect -4844 -5868 -4838 -5612
rect -4884 -5880 -4838 -5868
rect -4706 -5612 -4660 -5600
rect -4706 -5868 -4700 -5612
rect -4666 -5868 -4660 -5612
rect -4706 -5880 -4660 -5868
rect -4528 -5612 -4482 -5600
rect -4528 -5868 -4522 -5612
rect -4488 -5868 -4482 -5612
rect -4528 -5880 -4482 -5868
rect -4350 -5612 -4304 -5600
rect -4350 -5868 -4344 -5612
rect -4310 -5868 -4304 -5612
rect -4350 -5880 -4304 -5868
rect -4172 -5612 -4126 -5600
rect -4172 -5868 -4166 -5612
rect -4132 -5868 -4126 -5612
rect -4172 -5880 -4126 -5868
rect -3994 -5612 -3948 -5600
rect -3994 -5868 -3988 -5612
rect -3954 -5868 -3948 -5612
rect -3994 -5880 -3948 -5868
rect -3816 -5612 -3770 -5600
rect -3816 -5868 -3810 -5612
rect -3776 -5868 -3770 -5612
rect -3816 -5880 -3770 -5868
rect -3638 -5612 -3592 -5600
rect -3638 -5868 -3632 -5612
rect -3598 -5868 -3592 -5612
rect -3638 -5880 -3592 -5868
rect -3460 -5612 -3414 -5600
rect -3460 -5868 -3454 -5612
rect -3420 -5868 -3414 -5612
rect -3460 -5880 -3414 -5868
rect -6234 -5927 -6158 -5921
rect -6234 -5961 -6218 -5927
rect -6174 -5961 -6158 -5927
rect -6234 -5977 -6158 -5961
rect -6056 -5927 -5980 -5921
rect -6056 -5961 -6040 -5927
rect -5996 -5961 -5980 -5927
rect -6056 -5977 -5980 -5961
rect -5946 -6016 -5912 -5880
rect -5878 -5927 -5802 -5921
rect -5878 -5961 -5862 -5927
rect -5818 -5961 -5802 -5927
rect -5878 -5977 -5802 -5961
rect -5966 -6069 -5956 -6016
rect -5903 -6069 -5893 -6016
rect -5768 -6131 -5734 -5880
rect -5700 -5927 -5624 -5921
rect -5700 -5961 -5684 -5927
rect -5640 -5961 -5624 -5927
rect -5700 -5977 -5624 -5961
rect -5590 -6016 -5556 -5880
rect -5522 -5927 -5446 -5921
rect -5522 -5961 -5506 -5927
rect -5462 -5961 -5446 -5927
rect -5522 -5977 -5446 -5961
rect -5611 -6069 -5601 -6016
rect -5548 -6069 -5538 -6016
rect -5788 -6184 -5778 -6131
rect -5725 -6184 -5715 -6131
rect -5412 -6248 -5378 -5880
rect -5344 -5927 -5268 -5921
rect -5344 -5961 -5328 -5927
rect -5284 -5961 -5268 -5927
rect -5344 -5977 -5268 -5961
rect -5234 -6016 -5200 -5880
rect -5166 -5927 -5090 -5921
rect -5166 -5961 -5150 -5927
rect -5106 -5961 -5090 -5927
rect -5166 -5977 -5090 -5961
rect -5254 -6069 -5244 -6016
rect -5191 -6069 -5181 -6016
rect -5056 -6131 -5022 -5880
rect -4988 -5927 -4912 -5921
rect -4988 -5961 -4972 -5927
rect -4928 -5961 -4912 -5927
rect -4988 -5977 -4912 -5961
rect -5075 -6184 -5065 -6131
rect -5012 -6184 -5002 -6131
rect -6508 -6301 -6498 -6248
rect -6445 -6301 -6435 -6248
rect -5431 -6301 -5421 -6248
rect -5368 -6301 -5358 -6248
rect -4967 -6376 -4933 -5977
rect -4878 -6016 -4844 -5880
rect -4810 -5927 -4734 -5921
rect -4810 -5961 -4794 -5927
rect -4750 -5961 -4734 -5927
rect -4810 -5977 -4734 -5961
rect -4898 -6069 -4888 -6016
rect -4835 -6069 -4825 -6016
rect -4700 -6248 -4666 -5880
rect -4632 -5927 -4556 -5921
rect -4632 -5961 -4616 -5927
rect -4572 -5961 -4556 -5927
rect -4632 -5977 -4556 -5961
rect -4720 -6301 -4710 -6248
rect -4657 -6301 -4647 -6248
rect -4613 -6376 -4579 -5977
rect -4522 -6016 -4488 -5880
rect -4454 -5927 -4378 -5921
rect -4454 -5961 -4438 -5927
rect -4394 -5961 -4378 -5927
rect -4454 -5977 -4378 -5961
rect -4542 -6069 -4532 -6016
rect -4479 -6069 -4469 -6016
rect -4344 -6131 -4310 -5880
rect -4276 -5927 -4200 -5921
rect -4276 -5961 -4260 -5927
rect -4216 -5961 -4200 -5927
rect -4276 -5977 -4200 -5961
rect -4166 -6016 -4132 -5880
rect -4098 -5927 -4022 -5921
rect -4098 -5961 -4082 -5927
rect -4038 -5961 -4022 -5927
rect -4098 -5977 -4022 -5961
rect -4185 -6069 -4175 -6016
rect -4122 -6069 -4112 -6016
rect -4364 -6184 -4354 -6131
rect -4301 -6184 -4291 -6131
rect -3988 -6247 -3954 -5880
rect -3920 -5927 -3844 -5921
rect -3920 -5961 -3904 -5927
rect -3860 -5961 -3844 -5927
rect -3920 -5977 -3844 -5961
rect -3810 -5928 -3776 -5880
rect -3742 -5927 -3666 -5921
rect -3742 -5928 -3726 -5927
rect -3810 -5961 -3726 -5928
rect -3682 -5928 -3666 -5927
rect -3632 -5928 -3598 -5880
rect -3564 -5927 -3488 -5921
rect -3564 -5928 -3548 -5927
rect -3682 -5961 -3548 -5928
rect -3504 -5928 -3488 -5927
rect -3455 -5928 -3421 -5880
rect -3504 -5961 -3421 -5928
rect -3810 -5962 -3421 -5961
rect -3810 -6016 -3776 -5962
rect -3742 -5977 -3666 -5962
rect -3564 -5977 -3488 -5962
rect -3830 -6069 -3820 -6016
rect -3767 -6069 -3757 -6016
rect -3298 -6131 -3245 -5469
rect -2624 -6007 -2571 -5377
rect -2634 -6060 -2624 -6007
rect -2571 -6060 -2561 -6007
rect -3308 -6184 -3298 -6131
rect -3245 -6184 -3235 -6131
rect -4008 -6300 -3998 -6247
rect -3945 -6300 -3935 -6247
rect -3988 -6301 -3954 -6300
rect -4967 -6378 -4579 -6376
rect -4967 -6410 -4786 -6378
rect -4796 -6431 -4786 -6410
rect -4733 -6410 -4579 -6378
rect -4733 -6431 -4723 -6410
rect -2002 -6714 -1950 -4517
rect -1886 -5285 -1876 -5232
rect -1823 -5285 -1813 -5232
rect -1646 -5278 -1585 -3510
rect -1296 -3624 -1286 -3571
rect -1233 -3624 -1223 -3571
rect -1386 -3691 -1310 -3675
rect -1386 -3725 -1370 -3691
rect -1326 -3725 -1310 -3691
rect -1386 -3731 -1310 -3725
rect -1276 -3772 -1242 -3624
rect -1186 -3675 -1152 -3249
rect -1118 -3509 -1108 -3456
rect -1055 -3509 -1045 -3456
rect -1208 -3691 -1132 -3675
rect -1208 -3725 -1192 -3691
rect -1148 -3725 -1132 -3691
rect -1208 -3731 -1132 -3725
rect -1098 -3772 -1064 -3509
rect -1009 -3675 -975 -3249
rect -939 -3624 -929 -3571
rect -876 -3624 -866 -3571
rect -1030 -3691 -954 -3675
rect -1030 -3725 -1014 -3691
rect -970 -3725 -954 -3691
rect -1030 -3731 -954 -3725
rect -919 -3772 -885 -3624
rect -831 -3675 -797 -3249
rect -653 -3282 -619 -3249
rect -563 -3282 -529 -3152
rect -496 -3199 -420 -3193
rect -496 -3233 -480 -3199
rect -436 -3233 -420 -3199
rect -496 -3249 -420 -3233
rect -474 -3282 -440 -3249
rect -385 -3282 -351 -3152
rect -318 -3199 -242 -3193
rect -318 -3233 -302 -3199
rect -258 -3233 -242 -3199
rect -318 -3249 -242 -3233
rect -295 -3282 -261 -3249
rect -653 -3301 -261 -3282
rect -653 -3316 -484 -3301
rect -494 -3354 -484 -3316
rect -431 -3316 -261 -3301
rect -431 -3354 -421 -3316
rect -760 -3509 -750 -3456
rect -697 -3509 -687 -3456
rect -406 -3509 -396 -3456
rect -343 -3509 -333 -3456
rect -852 -3691 -776 -3675
rect -852 -3725 -836 -3691
rect -792 -3725 -776 -3691
rect -852 -3731 -776 -3725
rect -742 -3772 -708 -3509
rect -583 -3624 -573 -3571
rect -520 -3624 -510 -3571
rect -674 -3691 -598 -3675
rect -674 -3725 -658 -3691
rect -614 -3725 -598 -3691
rect -674 -3731 -598 -3725
rect -564 -3772 -530 -3624
rect -496 -3691 -420 -3675
rect -496 -3725 -480 -3691
rect -436 -3725 -420 -3691
rect -496 -3731 -420 -3725
rect -386 -3772 -352 -3509
rect -208 -3571 -174 -3152
rect -140 -3199 -64 -3193
rect -140 -3233 -124 -3199
rect -80 -3233 -64 -3199
rect -140 -3249 -64 -3233
rect -227 -3624 -217 -3571
rect -164 -3624 -154 -3571
rect -318 -3691 -242 -3675
rect -318 -3725 -302 -3691
rect -258 -3725 -242 -3691
rect -318 -3731 -242 -3725
rect -208 -3772 -174 -3624
rect -119 -3675 -85 -3249
rect -30 -3456 4 -3152
rect 38 -3199 114 -3193
rect 38 -3233 54 -3199
rect 98 -3233 114 -3199
rect 38 -3249 114 -3233
rect 216 -3199 292 -3193
rect 216 -3233 232 -3199
rect 276 -3233 292 -3199
rect 216 -3249 292 -3233
rect 327 -3456 361 -3152
rect 394 -3199 470 -3193
rect 394 -3233 410 -3199
rect 454 -3233 470 -3199
rect 394 -3249 470 -3233
rect 414 -3283 448 -3249
rect 504 -3283 538 -3152
rect 572 -3199 648 -3193
rect 572 -3233 588 -3199
rect 632 -3233 648 -3199
rect 572 -3249 648 -3233
rect 592 -3283 626 -3249
rect 682 -3283 716 -3152
rect 750 -3199 826 -3193
rect 750 -3233 766 -3199
rect 810 -3233 826 -3199
rect 750 -3249 826 -3233
rect 771 -3283 805 -3249
rect 414 -3301 805 -3283
rect 414 -3317 583 -3301
rect 573 -3354 583 -3317
rect 636 -3317 805 -3301
rect 636 -3354 646 -3317
rect -49 -3509 -39 -3456
rect 14 -3509 24 -3456
rect 307 -3509 317 -3456
rect 370 -3509 380 -3456
rect -140 -3691 -64 -3675
rect -140 -3725 -124 -3691
rect -80 -3725 -64 -3691
rect -140 -3731 -64 -3725
rect -30 -3772 4 -3509
rect 589 -3598 623 -3354
rect 860 -3456 894 -3152
rect 928 -3199 1004 -3193
rect 928 -3233 944 -3199
rect 988 -3233 1004 -3199
rect 928 -3249 1004 -3233
rect 1106 -3199 1182 -3193
rect 1106 -3233 1122 -3199
rect 1166 -3233 1182 -3199
rect 1106 -3249 1182 -3233
rect 1216 -3456 1250 -3152
rect 1284 -3199 1360 -3193
rect 1284 -3233 1300 -3199
rect 1344 -3233 1360 -3199
rect 1284 -3249 1360 -3233
rect 840 -3509 850 -3456
rect 903 -3509 913 -3456
rect 1196 -3509 1206 -3456
rect 1259 -3509 1269 -3456
rect 59 -3632 1160 -3598
rect 59 -3675 93 -3632
rect 149 -3633 271 -3632
rect 38 -3691 114 -3675
rect 38 -3725 54 -3691
rect 98 -3725 114 -3691
rect 38 -3731 114 -3725
rect 149 -3772 183 -3633
rect 237 -3675 271 -3633
rect 948 -3675 982 -3632
rect 216 -3691 292 -3675
rect 216 -3725 232 -3691
rect 276 -3725 292 -3691
rect 216 -3731 292 -3725
rect 394 -3691 470 -3675
rect 394 -3725 410 -3691
rect 454 -3725 470 -3691
rect 394 -3731 470 -3725
rect 572 -3691 648 -3675
rect 572 -3725 588 -3691
rect 632 -3725 648 -3691
rect 572 -3731 648 -3725
rect 750 -3691 826 -3675
rect 750 -3725 766 -3691
rect 810 -3725 826 -3691
rect 750 -3731 826 -3725
rect 928 -3691 1004 -3675
rect 928 -3725 944 -3691
rect 988 -3725 1004 -3691
rect 928 -3731 1004 -3725
rect 1038 -3772 1072 -3632
rect 1126 -3675 1160 -3632
rect 1106 -3691 1182 -3675
rect 1106 -3725 1122 -3691
rect 1166 -3725 1182 -3691
rect 1106 -3731 1182 -3725
rect 1216 -3772 1250 -3509
rect 1306 -3675 1340 -3249
rect 1394 -3564 1428 -3152
rect 1462 -3199 1538 -3193
rect 1462 -3233 1478 -3199
rect 1522 -3233 1538 -3199
rect 1462 -3249 1538 -3233
rect 1482 -3283 1516 -3249
rect 1572 -3283 1606 -3152
rect 1640 -3199 1716 -3193
rect 1640 -3233 1656 -3199
rect 1700 -3233 1716 -3199
rect 1640 -3249 1716 -3233
rect 1662 -3283 1696 -3249
rect 1750 -3283 1784 -3152
rect 1818 -3199 1894 -3193
rect 1818 -3233 1834 -3199
rect 1878 -3233 1894 -3199
rect 1818 -3249 1894 -3233
rect 1996 -3199 2072 -3193
rect 1996 -3233 2012 -3199
rect 2056 -3233 2072 -3199
rect 1996 -3249 2072 -3233
rect 2174 -3199 2250 -3193
rect 2174 -3233 2190 -3199
rect 2234 -3233 2250 -3199
rect 2174 -3249 2250 -3233
rect 2352 -3199 2428 -3193
rect 2352 -3233 2368 -3199
rect 2412 -3233 2428 -3199
rect 2352 -3249 2428 -3233
rect 1840 -3283 1874 -3249
rect 1482 -3301 1874 -3283
rect 1482 -3317 1654 -3301
rect 1644 -3354 1654 -3317
rect 1707 -3317 1874 -3301
rect 1707 -3354 1717 -3317
rect 1552 -3509 1562 -3456
rect 1615 -3509 1625 -3456
rect 1909 -3509 1919 -3456
rect 1972 -3509 1982 -3456
rect 1374 -3617 1384 -3564
rect 1437 -3617 1447 -3564
rect 1284 -3691 1360 -3675
rect 1284 -3725 1300 -3691
rect 1344 -3725 1360 -3691
rect 1284 -3731 1360 -3725
rect 1394 -3772 1428 -3617
rect 1462 -3691 1538 -3675
rect 1462 -3725 1478 -3691
rect 1522 -3725 1538 -3691
rect 1462 -3731 1538 -3725
rect 1572 -3772 1606 -3509
rect 1731 -3617 1741 -3564
rect 1794 -3617 1804 -3564
rect 1640 -3691 1716 -3675
rect 1640 -3725 1656 -3691
rect 1700 -3725 1716 -3691
rect 1640 -3731 1716 -3725
rect 1750 -3772 1784 -3617
rect 1818 -3691 1894 -3675
rect 1818 -3725 1834 -3691
rect 1878 -3725 1894 -3691
rect 1818 -3731 1894 -3725
rect 1929 -3772 1963 -3509
rect 2017 -3675 2051 -3249
rect 2087 -3617 2097 -3564
rect 2150 -3617 2160 -3564
rect 1996 -3691 2072 -3675
rect 1996 -3725 2012 -3691
rect 2056 -3725 2072 -3691
rect 1996 -3731 2072 -3725
rect 2106 -3772 2140 -3617
rect 2196 -3675 2230 -3249
rect 2265 -3509 2275 -3456
rect 2328 -3509 2338 -3456
rect 2174 -3691 2250 -3675
rect 2174 -3725 2190 -3691
rect 2234 -3725 2250 -3691
rect 2174 -3731 2250 -3725
rect 2284 -3772 2318 -3509
rect 2373 -3675 2407 -3249
rect 2462 -3284 2496 -3152
rect 2530 -3199 2606 -3193
rect 2530 -3233 2546 -3199
rect 2590 -3233 2606 -3199
rect 2530 -3249 2606 -3233
rect 2551 -3284 2585 -3249
rect 2641 -3284 2675 -3152
rect 2462 -3318 2675 -3284
rect 2441 -3617 2451 -3564
rect 2504 -3617 2514 -3564
rect 2352 -3691 2428 -3675
rect 2352 -3725 2368 -3691
rect 2412 -3725 2428 -3691
rect 2352 -3731 2428 -3725
rect 2462 -3772 2496 -3617
rect 2530 -3691 2606 -3675
rect 2530 -3725 2546 -3691
rect 2590 -3725 2606 -3691
rect 2530 -3731 2606 -3725
rect -1460 -3784 -1414 -3772
rect -1460 -4040 -1454 -3784
rect -1420 -4040 -1414 -3784
rect -1460 -4052 -1414 -4040
rect -1282 -3784 -1236 -3772
rect -1282 -4040 -1276 -3784
rect -1242 -4040 -1236 -3784
rect -1282 -4052 -1236 -4040
rect -1104 -3784 -1058 -3772
rect -1104 -4040 -1098 -3784
rect -1064 -4040 -1058 -3784
rect -1104 -4052 -1058 -4040
rect -926 -3784 -880 -3772
rect -926 -4040 -920 -3784
rect -886 -4040 -880 -3784
rect -926 -4052 -880 -4040
rect -748 -3784 -702 -3772
rect -748 -4040 -742 -3784
rect -708 -4040 -702 -3784
rect -748 -4052 -702 -4040
rect -570 -3784 -524 -3772
rect -570 -4040 -564 -3784
rect -530 -4040 -524 -3784
rect -570 -4052 -524 -4040
rect -392 -3784 -346 -3772
rect -392 -4040 -386 -3784
rect -352 -4040 -346 -3784
rect -392 -4052 -346 -4040
rect -214 -3784 -168 -3772
rect -214 -4040 -208 -3784
rect -174 -4040 -168 -3784
rect -214 -4052 -168 -4040
rect -36 -3784 10 -3772
rect -36 -4040 -30 -3784
rect 4 -4040 10 -3784
rect -36 -4052 10 -4040
rect 142 -3784 188 -3772
rect 142 -4040 148 -3784
rect 182 -4040 188 -3784
rect 142 -4052 188 -4040
rect 320 -3784 366 -3772
rect 320 -4040 326 -3784
rect 360 -4040 366 -3784
rect 320 -4052 366 -4040
rect 498 -3784 544 -3772
rect 498 -4040 504 -3784
rect 538 -4040 544 -3784
rect 498 -4052 544 -4040
rect 676 -3784 722 -3772
rect 676 -4040 682 -3784
rect 716 -4040 722 -3784
rect 676 -4052 722 -4040
rect 854 -3784 900 -3772
rect 854 -4040 860 -3784
rect 894 -4040 900 -3784
rect 854 -4052 900 -4040
rect 1032 -3784 1078 -3772
rect 1032 -4040 1038 -3784
rect 1072 -4040 1078 -3784
rect 1032 -4052 1078 -4040
rect 1210 -3784 1256 -3772
rect 1210 -4040 1216 -3784
rect 1250 -4040 1256 -3784
rect 1210 -4052 1256 -4040
rect 1388 -3784 1434 -3772
rect 1388 -4040 1394 -3784
rect 1428 -4040 1434 -3784
rect 1388 -4052 1434 -4040
rect 1566 -3784 1612 -3772
rect 1566 -4040 1572 -3784
rect 1606 -4040 1612 -3784
rect 1566 -4052 1612 -4040
rect 1744 -3784 1790 -3772
rect 1744 -4040 1750 -3784
rect 1784 -4040 1790 -3784
rect 1744 -4052 1790 -4040
rect 1922 -3784 1968 -3772
rect 1922 -4040 1928 -3784
rect 1962 -4040 1968 -3784
rect 1922 -4052 1968 -4040
rect 2100 -3784 2146 -3772
rect 2100 -4040 2106 -3784
rect 2140 -4040 2146 -3784
rect 2100 -4052 2146 -4040
rect 2278 -3784 2324 -3772
rect 2278 -4040 2284 -3784
rect 2318 -4040 2324 -3784
rect 2278 -4052 2324 -4040
rect 2456 -3784 2502 -3772
rect 2456 -4040 2462 -3784
rect 2496 -4040 2502 -3784
rect 2456 -4052 2502 -4040
rect 2634 -3784 2680 -3772
rect 2634 -4040 2640 -3784
rect 2674 -4040 2680 -3784
rect 2634 -4052 2680 -4040
rect -1454 -4184 -1420 -4052
rect -1386 -4099 -1310 -4093
rect -1386 -4133 -1370 -4099
rect -1326 -4133 -1310 -4099
rect -1386 -4149 -1310 -4133
rect -1366 -4184 -1332 -4149
rect -1276 -4184 -1242 -4052
rect -1208 -4099 -1132 -4093
rect -1208 -4133 -1192 -4099
rect -1148 -4133 -1132 -4099
rect -1208 -4149 -1132 -4133
rect -1030 -4099 -954 -4093
rect -1030 -4133 -1014 -4099
rect -970 -4133 -954 -4099
rect -1030 -4149 -954 -4133
rect -852 -4099 -776 -4093
rect -852 -4133 -836 -4099
rect -792 -4133 -776 -4099
rect -852 -4149 -776 -4133
rect -674 -4099 -598 -4093
rect -674 -4133 -658 -4099
rect -614 -4133 -598 -4099
rect -674 -4149 -598 -4133
rect -496 -4099 -420 -4093
rect -496 -4133 -480 -4099
rect -436 -4133 -420 -4099
rect -496 -4149 -420 -4133
rect -318 -4099 -242 -4093
rect -318 -4133 -302 -4099
rect -258 -4133 -242 -4099
rect -318 -4149 -242 -4133
rect -140 -4099 -64 -4093
rect -140 -4133 -124 -4099
rect -80 -4133 -64 -4099
rect -140 -4149 -64 -4133
rect 38 -4099 114 -4093
rect 38 -4133 54 -4099
rect 98 -4133 114 -4099
rect 38 -4149 114 -4133
rect -1454 -4218 -1242 -4184
rect -1454 -4541 -1242 -4507
rect -1454 -4672 -1420 -4541
rect -1365 -4575 -1331 -4541
rect -1386 -4591 -1310 -4575
rect -1386 -4625 -1370 -4591
rect -1326 -4625 -1310 -4591
rect -1386 -4631 -1310 -4625
rect -1276 -4672 -1242 -4541
rect -1187 -4575 -1153 -4149
rect -1009 -4575 -975 -4149
rect -831 -4192 -797 -4149
rect -653 -4192 -619 -4149
rect -474 -4192 -440 -4149
rect -297 -4192 -263 -4149
rect -851 -4245 -841 -4192
rect -788 -4245 -778 -4192
rect -672 -4245 -662 -4192
rect -609 -4245 -599 -4192
rect -493 -4245 -483 -4192
rect -430 -4245 -420 -4192
rect -316 -4245 -306 -4192
rect -253 -4245 -243 -4192
rect -831 -4575 -797 -4245
rect -653 -4575 -619 -4245
rect -474 -4575 -440 -4245
rect -297 -4575 -263 -4245
rect -119 -4575 -85 -4149
rect -1208 -4591 -1132 -4575
rect -1208 -4625 -1192 -4591
rect -1148 -4625 -1132 -4591
rect -1208 -4631 -1132 -4625
rect -1030 -4591 -954 -4575
rect -1030 -4625 -1014 -4591
rect -970 -4625 -954 -4591
rect -1030 -4631 -954 -4625
rect -852 -4591 -776 -4575
rect -852 -4625 -836 -4591
rect -792 -4625 -776 -4591
rect -852 -4631 -776 -4625
rect -674 -4591 -598 -4575
rect -674 -4625 -658 -4591
rect -614 -4625 -598 -4591
rect -674 -4631 -598 -4625
rect -496 -4591 -420 -4575
rect -496 -4625 -480 -4591
rect -436 -4625 -420 -4591
rect -496 -4631 -420 -4625
rect -318 -4591 -242 -4575
rect -318 -4625 -302 -4591
rect -258 -4625 -242 -4591
rect -318 -4631 -242 -4625
rect -140 -4591 -64 -4575
rect -140 -4625 -124 -4591
rect -80 -4625 -64 -4591
rect -140 -4631 -64 -4625
rect 38 -4591 114 -4575
rect 38 -4625 54 -4591
rect 98 -4625 114 -4591
rect 38 -4631 114 -4625
rect 148 -4672 182 -4052
rect 216 -4099 292 -4093
rect 216 -4133 232 -4099
rect 276 -4133 292 -4099
rect 216 -4149 292 -4133
rect 326 -4304 360 -4052
rect 394 -4099 470 -4093
rect 394 -4133 410 -4099
rect 454 -4133 470 -4099
rect 394 -4149 470 -4133
rect 416 -4192 450 -4149
rect 397 -4245 407 -4192
rect 460 -4245 470 -4192
rect 307 -4357 317 -4304
rect 370 -4357 380 -4304
rect 216 -4591 292 -4575
rect 216 -4625 232 -4591
rect 276 -4625 292 -4591
rect 216 -4631 292 -4625
rect 326 -4672 360 -4357
rect 416 -4575 450 -4245
rect 504 -4412 538 -4052
rect 572 -4099 648 -4093
rect 572 -4133 588 -4099
rect 632 -4133 648 -4099
rect 572 -4149 648 -4133
rect 593 -4192 627 -4149
rect 573 -4245 583 -4192
rect 636 -4245 646 -4192
rect 485 -4465 495 -4412
rect 548 -4465 558 -4412
rect 394 -4591 470 -4575
rect 394 -4625 410 -4591
rect 454 -4625 470 -4591
rect 394 -4631 470 -4625
rect 504 -4672 538 -4465
rect 593 -4575 627 -4245
rect 682 -4304 716 -4052
rect 750 -4099 826 -4093
rect 750 -4133 766 -4099
rect 810 -4133 826 -4099
rect 750 -4149 826 -4133
rect 771 -4192 805 -4149
rect 751 -4245 761 -4192
rect 814 -4245 824 -4192
rect 663 -4357 673 -4304
rect 726 -4357 736 -4304
rect 572 -4591 648 -4575
rect 572 -4625 588 -4591
rect 632 -4625 648 -4591
rect 572 -4631 648 -4625
rect 682 -4672 716 -4357
rect 771 -4575 805 -4245
rect 860 -4412 894 -4052
rect 928 -4099 1004 -4093
rect 928 -4133 944 -4099
rect 988 -4133 1004 -4099
rect 928 -4149 1004 -4133
rect 840 -4465 850 -4412
rect 903 -4465 913 -4412
rect 750 -4591 826 -4575
rect 750 -4625 766 -4591
rect 810 -4625 826 -4591
rect 750 -4631 826 -4625
rect 860 -4672 894 -4465
rect 928 -4591 1004 -4575
rect 928 -4625 944 -4591
rect 988 -4625 1004 -4591
rect 928 -4631 1004 -4625
rect 1039 -4672 1073 -4052
rect 1106 -4099 1182 -4093
rect 1106 -4133 1122 -4099
rect 1166 -4133 1182 -4099
rect 1106 -4149 1182 -4133
rect 1284 -4099 1360 -4093
rect 1284 -4133 1300 -4099
rect 1344 -4133 1360 -4099
rect 1284 -4149 1360 -4133
rect 1462 -4099 1538 -4093
rect 1462 -4133 1478 -4099
rect 1522 -4133 1538 -4099
rect 1462 -4149 1538 -4133
rect 1640 -4099 1716 -4093
rect 1640 -4133 1656 -4099
rect 1700 -4133 1716 -4099
rect 1640 -4149 1716 -4133
rect 1818 -4099 1894 -4093
rect 1818 -4133 1834 -4099
rect 1878 -4133 1894 -4099
rect 1818 -4149 1894 -4133
rect 1996 -4099 2072 -4093
rect 1996 -4133 2012 -4099
rect 2056 -4133 2072 -4099
rect 1996 -4149 2072 -4133
rect 2174 -4099 2250 -4093
rect 2174 -4133 2190 -4099
rect 2234 -4133 2250 -4099
rect 2174 -4149 2250 -4133
rect 2352 -4099 2428 -4093
rect 2352 -4133 2368 -4099
rect 2412 -4133 2428 -4099
rect 2352 -4149 2428 -4133
rect 1305 -4575 1339 -4149
rect 1484 -4192 1518 -4149
rect 1661 -4192 1695 -4149
rect 1839 -4192 1873 -4149
rect 2017 -4192 2051 -4149
rect 1464 -4245 1474 -4192
rect 1527 -4245 1537 -4192
rect 1642 -4245 1652 -4192
rect 1705 -4245 1715 -4192
rect 1820 -4245 1830 -4192
rect 1883 -4245 1893 -4192
rect 1998 -4245 2008 -4192
rect 2061 -4245 2071 -4192
rect 1484 -4575 1518 -4245
rect 1661 -4575 1695 -4245
rect 1839 -4575 1873 -4245
rect 2017 -4575 2051 -4245
rect 2195 -4575 2229 -4149
rect 2373 -4575 2407 -4149
rect 2463 -4182 2497 -4052
rect 2530 -4099 2606 -4093
rect 2530 -4133 2546 -4099
rect 2590 -4133 2606 -4099
rect 2530 -4149 2606 -4133
rect 2552 -4182 2586 -4149
rect 2640 -4180 2674 -4052
rect 2640 -4182 2792 -4180
rect 2463 -4214 2792 -4182
rect 2463 -4216 2674 -4214
rect 2528 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect 2550 -4506 2584 -4327
rect 2758 -4446 2792 -4214
rect 2462 -4540 2674 -4506
rect 2736 -4507 2746 -4446
rect 2807 -4507 2817 -4446
rect 2758 -4508 2792 -4507
rect 1106 -4591 1182 -4575
rect 1106 -4625 1122 -4591
rect 1166 -4625 1182 -4591
rect 1106 -4631 1182 -4625
rect 1284 -4591 1360 -4575
rect 1284 -4625 1300 -4591
rect 1344 -4625 1360 -4591
rect 1284 -4631 1360 -4625
rect 1462 -4591 1538 -4575
rect 1462 -4625 1478 -4591
rect 1522 -4625 1538 -4591
rect 1462 -4631 1538 -4625
rect 1640 -4591 1716 -4575
rect 1640 -4625 1656 -4591
rect 1700 -4625 1716 -4591
rect 1640 -4631 1716 -4625
rect 1818 -4591 1894 -4575
rect 1818 -4625 1834 -4591
rect 1878 -4625 1894 -4591
rect 1818 -4631 1894 -4625
rect 1996 -4591 2072 -4575
rect 1996 -4625 2012 -4591
rect 2056 -4625 2072 -4591
rect 1996 -4631 2072 -4625
rect 2174 -4591 2250 -4575
rect 2174 -4625 2190 -4591
rect 2234 -4625 2250 -4591
rect 2174 -4631 2250 -4625
rect 2352 -4591 2428 -4575
rect 2352 -4625 2368 -4591
rect 2412 -4625 2428 -4591
rect 2352 -4631 2428 -4625
rect 2462 -4672 2496 -4540
rect 2550 -4575 2584 -4540
rect 2530 -4591 2606 -4575
rect 2530 -4625 2546 -4591
rect 2590 -4625 2606 -4591
rect 2530 -4631 2606 -4625
rect 2640 -4672 2674 -4540
rect -1460 -4684 -1414 -4672
rect -1460 -4940 -1454 -4684
rect -1420 -4940 -1414 -4684
rect -1460 -4952 -1414 -4940
rect -1282 -4684 -1236 -4672
rect -1282 -4940 -1276 -4684
rect -1242 -4940 -1236 -4684
rect -1282 -4952 -1236 -4940
rect -1104 -4684 -1058 -4672
rect -1104 -4940 -1098 -4684
rect -1064 -4940 -1058 -4684
rect -1104 -4952 -1058 -4940
rect -926 -4684 -880 -4672
rect -926 -4940 -920 -4684
rect -886 -4940 -880 -4684
rect -926 -4952 -880 -4940
rect -748 -4684 -702 -4672
rect -748 -4940 -742 -4684
rect -708 -4940 -702 -4684
rect -748 -4952 -702 -4940
rect -570 -4684 -524 -4672
rect -570 -4940 -564 -4684
rect -530 -4940 -524 -4684
rect -570 -4952 -524 -4940
rect -392 -4684 -346 -4672
rect -392 -4940 -386 -4684
rect -352 -4940 -346 -4684
rect -392 -4952 -346 -4940
rect -214 -4684 -168 -4672
rect -214 -4940 -208 -4684
rect -174 -4940 -168 -4684
rect -214 -4952 -168 -4940
rect -36 -4684 10 -4672
rect -36 -4940 -30 -4684
rect 4 -4940 10 -4684
rect -36 -4952 10 -4940
rect 142 -4684 188 -4672
rect 142 -4940 148 -4684
rect 182 -4940 188 -4684
rect 142 -4952 188 -4940
rect 320 -4684 366 -4672
rect 320 -4940 326 -4684
rect 360 -4940 366 -4684
rect 320 -4952 366 -4940
rect 498 -4684 544 -4672
rect 498 -4940 504 -4684
rect 538 -4940 544 -4684
rect 498 -4952 544 -4940
rect 676 -4684 722 -4672
rect 676 -4940 682 -4684
rect 716 -4940 722 -4684
rect 676 -4952 722 -4940
rect 854 -4684 900 -4672
rect 854 -4940 860 -4684
rect 894 -4940 900 -4684
rect 854 -4952 900 -4940
rect 1032 -4684 1078 -4672
rect 1032 -4940 1038 -4684
rect 1072 -4940 1078 -4684
rect 1032 -4952 1078 -4940
rect 1210 -4684 1256 -4672
rect 1210 -4940 1216 -4684
rect 1250 -4940 1256 -4684
rect 1210 -4952 1256 -4940
rect 1388 -4684 1434 -4672
rect 1388 -4940 1394 -4684
rect 1428 -4940 1434 -4684
rect 1388 -4952 1434 -4940
rect 1566 -4684 1612 -4672
rect 1566 -4940 1572 -4684
rect 1606 -4940 1612 -4684
rect 1566 -4952 1612 -4940
rect 1744 -4684 1790 -4672
rect 1744 -4940 1750 -4684
rect 1784 -4940 1790 -4684
rect 1744 -4952 1790 -4940
rect 1922 -4684 1968 -4672
rect 1922 -4940 1928 -4684
rect 1962 -4940 1968 -4684
rect 1922 -4952 1968 -4940
rect 2100 -4684 2146 -4672
rect 2100 -4940 2106 -4684
rect 2140 -4940 2146 -4684
rect 2100 -4952 2146 -4940
rect 2278 -4684 2324 -4672
rect 2278 -4940 2284 -4684
rect 2318 -4940 2324 -4684
rect 2278 -4952 2324 -4940
rect 2456 -4684 2502 -4672
rect 2456 -4940 2462 -4684
rect 2496 -4940 2502 -4684
rect 2456 -4952 2502 -4940
rect 2634 -4684 2680 -4672
rect 2634 -4940 2640 -4684
rect 2674 -4940 2680 -4684
rect 2634 -4952 2680 -4940
rect -1386 -4999 -1310 -4993
rect -1386 -5033 -1370 -4999
rect -1326 -5033 -1310 -4999
rect -1386 -5049 -1310 -5033
rect -1277 -5097 -1243 -4952
rect -1208 -4999 -1132 -4993
rect -1208 -5033 -1192 -4999
rect -1148 -5033 -1132 -4999
rect -1208 -5049 -1132 -5033
rect -1297 -5150 -1287 -5097
rect -1234 -5150 -1224 -5097
rect -1876 -5337 -1823 -5285
rect -1875 -6364 -1823 -5337
rect -1656 -5339 -1646 -5278
rect -1585 -5339 -1575 -5278
rect -1454 -5442 -1242 -5408
rect -1454 -5572 -1420 -5442
rect -1363 -5475 -1329 -5442
rect -1386 -5491 -1310 -5475
rect -1386 -5525 -1370 -5491
rect -1326 -5525 -1310 -5491
rect -1386 -5531 -1310 -5525
rect -1276 -5572 -1242 -5442
rect -1187 -5475 -1153 -5049
rect -1097 -5213 -1063 -4952
rect -1030 -4999 -954 -4993
rect -1030 -5033 -1014 -4999
rect -970 -5033 -954 -4999
rect -1030 -5049 -954 -5033
rect -1115 -5266 -1105 -5213
rect -1052 -5266 -1042 -5213
rect -1009 -5475 -975 -5049
rect -919 -5097 -885 -4952
rect -852 -4999 -776 -4993
rect -852 -5033 -836 -4999
rect -792 -5033 -776 -4999
rect -852 -5049 -776 -5033
rect -939 -5150 -929 -5097
rect -876 -5150 -866 -5097
rect -830 -5475 -796 -5049
rect -741 -5213 -707 -4952
rect -674 -4999 -598 -4993
rect -674 -5033 -658 -4999
rect -614 -5033 -598 -4999
rect -674 -5049 -598 -5033
rect -563 -5097 -529 -4952
rect -496 -4999 -420 -4993
rect -496 -5033 -480 -4999
rect -436 -5033 -420 -4999
rect -496 -5049 -420 -5033
rect -582 -5150 -572 -5097
rect -519 -5150 -509 -5097
rect -386 -5213 -352 -4952
rect -318 -4999 -242 -4993
rect -318 -5033 -302 -4999
rect -258 -5033 -242 -4999
rect -318 -5049 -242 -5033
rect -208 -5097 -174 -4952
rect -140 -4999 -64 -4993
rect -140 -5033 -124 -4999
rect -80 -5033 -64 -4999
rect -140 -5049 -64 -5033
rect -228 -5150 -218 -5097
rect -165 -5150 -155 -5097
rect -761 -5266 -751 -5213
rect -698 -5266 -688 -5213
rect -406 -5266 -396 -5213
rect -343 -5266 -333 -5213
rect -654 -5434 -262 -5400
rect -654 -5475 -620 -5434
rect -1208 -5491 -1132 -5475
rect -1208 -5525 -1192 -5491
rect -1148 -5525 -1132 -5491
rect -1208 -5531 -1132 -5525
rect -1030 -5491 -954 -5475
rect -1030 -5525 -1014 -5491
rect -970 -5525 -954 -5491
rect -1030 -5531 -954 -5525
rect -852 -5491 -776 -5475
rect -852 -5525 -836 -5491
rect -792 -5525 -776 -5491
rect -852 -5531 -776 -5525
rect -674 -5491 -598 -5475
rect -674 -5525 -658 -5491
rect -614 -5525 -598 -5491
rect -674 -5531 -598 -5525
rect -563 -5572 -529 -5434
rect -474 -5475 -440 -5434
rect -496 -5491 -420 -5475
rect -496 -5525 -480 -5491
rect -436 -5525 -420 -5491
rect -496 -5531 -420 -5525
rect -385 -5572 -351 -5434
rect -296 -5475 -262 -5434
rect -318 -5491 -242 -5475
rect -318 -5525 -302 -5491
rect -258 -5525 -242 -5491
rect -318 -5531 -242 -5525
rect -208 -5572 -174 -5150
rect -119 -5380 -85 -5049
rect -30 -5213 4 -4952
rect 59 -4993 93 -4992
rect 38 -4999 114 -4993
rect 38 -5033 54 -4999
rect 98 -5033 114 -4999
rect 38 -5049 114 -5033
rect 59 -5091 93 -5049
rect 148 -5091 182 -4952
rect 216 -4999 292 -4993
rect 216 -5033 232 -4999
rect 276 -5033 292 -4999
rect 216 -5049 292 -5033
rect 394 -4999 470 -4993
rect 394 -5033 410 -4999
rect 454 -5033 470 -4999
rect 394 -5049 470 -5033
rect 572 -4999 648 -4993
rect 572 -5033 588 -4999
rect 632 -5033 648 -4999
rect 572 -5049 648 -5033
rect 750 -4999 826 -4993
rect 750 -5033 766 -4999
rect 810 -5033 826 -4999
rect 750 -5049 826 -5033
rect 928 -4999 1004 -4993
rect 928 -5033 944 -4999
rect 988 -5033 1004 -4999
rect 928 -5049 1004 -5033
rect 236 -5091 270 -5049
rect 948 -5091 982 -5049
rect 1039 -5091 1073 -4952
rect 1106 -4999 1182 -4993
rect 1106 -5033 1122 -4999
rect 1166 -5033 1182 -4999
rect 1106 -5049 1182 -5033
rect 1128 -5091 1162 -5049
rect 59 -5125 1162 -5091
rect -51 -5266 -41 -5213
rect 12 -5266 22 -5213
rect 306 -5266 316 -5213
rect 369 -5266 379 -5213
rect -138 -5433 -128 -5380
rect -75 -5433 -65 -5380
rect -119 -5475 -85 -5433
rect -140 -5491 -64 -5475
rect -140 -5525 -124 -5491
rect -80 -5525 -64 -5491
rect -140 -5531 -64 -5525
rect -30 -5572 4 -5266
rect 40 -5433 50 -5380
rect 103 -5433 113 -5380
rect 218 -5433 228 -5380
rect 281 -5433 291 -5380
rect 59 -5475 93 -5433
rect 238 -5475 272 -5433
rect 38 -5491 114 -5475
rect 38 -5525 54 -5491
rect 98 -5525 114 -5491
rect 38 -5531 114 -5525
rect 216 -5491 292 -5475
rect 216 -5525 232 -5491
rect 276 -5525 292 -5491
rect 216 -5531 292 -5525
rect 326 -5572 360 -5266
rect 593 -5315 627 -5125
rect 1216 -5213 1250 -4952
rect 1284 -4999 1360 -4993
rect 1284 -5033 1300 -4999
rect 1344 -5033 1360 -4999
rect 1284 -5049 1360 -5033
rect 840 -5266 850 -5213
rect 903 -5266 913 -5213
rect 1197 -5266 1207 -5213
rect 1260 -5266 1270 -5213
rect 415 -5349 804 -5315
rect 415 -5475 449 -5349
rect 394 -5491 470 -5475
rect 394 -5525 410 -5491
rect 454 -5525 470 -5491
rect 394 -5531 470 -5525
rect 505 -5572 539 -5349
rect 592 -5475 626 -5349
rect 572 -5491 648 -5475
rect 572 -5525 588 -5491
rect 632 -5525 648 -5491
rect 572 -5531 648 -5525
rect 681 -5572 715 -5349
rect 770 -5475 804 -5349
rect 750 -5491 826 -5475
rect 750 -5525 766 -5491
rect 810 -5525 826 -5491
rect 750 -5531 826 -5525
rect 860 -5572 894 -5266
rect 930 -5434 940 -5381
rect 993 -5434 1003 -5381
rect 1109 -5433 1119 -5380
rect 1172 -5433 1182 -5380
rect 949 -5475 983 -5434
rect 1128 -5475 1162 -5433
rect 928 -5491 1004 -5475
rect 928 -5525 944 -5491
rect 988 -5525 1004 -5491
rect 928 -5531 1004 -5525
rect 1106 -5491 1182 -5475
rect 1106 -5525 1122 -5491
rect 1166 -5525 1182 -5491
rect 1106 -5531 1182 -5525
rect 1216 -5572 1250 -5266
rect 1306 -5380 1340 -5049
rect 1394 -5093 1428 -4952
rect 1462 -4999 1538 -4993
rect 1462 -5033 1478 -4999
rect 1522 -5033 1538 -4999
rect 1462 -5049 1538 -5033
rect 1375 -5146 1385 -5093
rect 1438 -5146 1448 -5093
rect 1286 -5433 1296 -5380
rect 1349 -5433 1359 -5380
rect 1306 -5475 1340 -5433
rect 1284 -5491 1360 -5475
rect 1284 -5525 1300 -5491
rect 1344 -5525 1360 -5491
rect 1284 -5531 1360 -5525
rect 1394 -5572 1428 -5146
rect 1572 -5213 1606 -4952
rect 1640 -4999 1716 -4993
rect 1640 -5033 1656 -4999
rect 1700 -5033 1716 -4999
rect 1640 -5049 1716 -5033
rect 1750 -5093 1784 -4952
rect 1818 -4999 1894 -4993
rect 1818 -5033 1834 -4999
rect 1878 -5033 1894 -4999
rect 1818 -5049 1894 -5033
rect 1730 -5146 1740 -5093
rect 1793 -5146 1803 -5093
rect 1927 -5213 1961 -4952
rect 1996 -4999 2072 -4993
rect 1996 -5033 2012 -4999
rect 2056 -5033 2072 -4999
rect 1996 -5049 2072 -5033
rect 1553 -5266 1563 -5213
rect 1616 -5266 1626 -5213
rect 1907 -5266 1917 -5213
rect 1970 -5266 1980 -5213
rect 1482 -5433 1874 -5399
rect 1482 -5475 1516 -5433
rect 1462 -5491 1538 -5475
rect 1462 -5525 1478 -5491
rect 1522 -5525 1538 -5491
rect 1462 -5531 1538 -5525
rect 1573 -5572 1607 -5433
rect 1661 -5475 1695 -5433
rect 1640 -5491 1716 -5475
rect 1640 -5525 1656 -5491
rect 1700 -5525 1716 -5491
rect 1640 -5531 1716 -5525
rect 1749 -5572 1783 -5433
rect 1840 -5475 1874 -5433
rect 2018 -5475 2052 -5049
rect 2106 -5093 2140 -4952
rect 2174 -4999 2250 -4993
rect 2174 -5033 2190 -4999
rect 2234 -5033 2250 -4999
rect 2174 -5049 2250 -5033
rect 2086 -5146 2096 -5093
rect 2149 -5146 2159 -5093
rect 2195 -5475 2229 -5049
rect 2284 -5213 2318 -4952
rect 2352 -4999 2428 -4993
rect 2352 -5033 2368 -4999
rect 2412 -5033 2428 -4999
rect 2352 -5049 2428 -5033
rect 2264 -5266 2274 -5213
rect 2327 -5266 2337 -5213
rect 2373 -5475 2407 -5049
rect 2462 -5093 2496 -4952
rect 2530 -4999 2606 -4993
rect 2530 -5033 2546 -4999
rect 2590 -5033 2606 -4999
rect 2530 -5049 2606 -5033
rect 2443 -5146 2453 -5093
rect 2506 -5146 2516 -5093
rect 2463 -5442 2674 -5408
rect 1818 -5491 1894 -5475
rect 1818 -5525 1834 -5491
rect 1878 -5525 1894 -5491
rect 1818 -5531 1894 -5525
rect 1996 -5491 2072 -5475
rect 1996 -5525 2012 -5491
rect 2056 -5525 2072 -5491
rect 1996 -5531 2072 -5525
rect 2174 -5491 2250 -5475
rect 2174 -5525 2190 -5491
rect 2234 -5525 2250 -5491
rect 2174 -5531 2250 -5525
rect 2352 -5491 2428 -5475
rect 2352 -5525 2368 -5491
rect 2412 -5525 2428 -5491
rect 2352 -5531 2428 -5525
rect 2463 -5572 2497 -5442
rect 2550 -5475 2584 -5442
rect 2530 -5491 2606 -5475
rect 2530 -5525 2546 -5491
rect 2590 -5525 2606 -5491
rect 2530 -5531 2606 -5525
rect 2640 -5572 2674 -5442
rect -1460 -5584 -1414 -5572
rect -1460 -5840 -1454 -5584
rect -1420 -5840 -1414 -5584
rect -1460 -5852 -1414 -5840
rect -1282 -5584 -1236 -5572
rect -1282 -5840 -1276 -5584
rect -1242 -5840 -1236 -5584
rect -1282 -5852 -1236 -5840
rect -1104 -5584 -1058 -5572
rect -1104 -5840 -1098 -5584
rect -1064 -5840 -1058 -5584
rect -1104 -5852 -1058 -5840
rect -926 -5584 -880 -5572
rect -926 -5840 -920 -5584
rect -886 -5840 -880 -5584
rect -926 -5852 -880 -5840
rect -748 -5584 -702 -5572
rect -748 -5840 -742 -5584
rect -708 -5840 -702 -5584
rect -748 -5852 -702 -5840
rect -570 -5584 -524 -5572
rect -570 -5840 -564 -5584
rect -530 -5840 -524 -5584
rect -570 -5852 -524 -5840
rect -392 -5584 -346 -5572
rect -392 -5840 -386 -5584
rect -352 -5840 -346 -5584
rect -392 -5852 -346 -5840
rect -214 -5584 -168 -5572
rect -214 -5840 -208 -5584
rect -174 -5840 -168 -5584
rect -214 -5852 -168 -5840
rect -36 -5584 10 -5572
rect -36 -5840 -30 -5584
rect 4 -5840 10 -5584
rect -36 -5852 10 -5840
rect 142 -5584 188 -5572
rect 142 -5840 148 -5584
rect 182 -5840 188 -5584
rect 142 -5852 188 -5840
rect 320 -5584 366 -5572
rect 320 -5840 326 -5584
rect 360 -5840 366 -5584
rect 320 -5852 366 -5840
rect 498 -5584 544 -5572
rect 498 -5840 504 -5584
rect 538 -5840 544 -5584
rect 498 -5852 544 -5840
rect 676 -5584 722 -5572
rect 676 -5840 682 -5584
rect 716 -5840 722 -5584
rect 676 -5852 722 -5840
rect 854 -5584 900 -5572
rect 854 -5840 860 -5584
rect 894 -5840 900 -5584
rect 854 -5852 900 -5840
rect 1032 -5584 1078 -5572
rect 1032 -5840 1038 -5584
rect 1072 -5840 1078 -5584
rect 1032 -5852 1078 -5840
rect 1210 -5584 1256 -5572
rect 1210 -5840 1216 -5584
rect 1250 -5840 1256 -5584
rect 1210 -5852 1256 -5840
rect 1388 -5584 1434 -5572
rect 1388 -5840 1394 -5584
rect 1428 -5840 1434 -5584
rect 1388 -5852 1434 -5840
rect 1566 -5584 1612 -5572
rect 1566 -5840 1572 -5584
rect 1606 -5840 1612 -5584
rect 1566 -5852 1612 -5840
rect 1744 -5584 1790 -5572
rect 1744 -5840 1750 -5584
rect 1784 -5840 1790 -5584
rect 1744 -5852 1790 -5840
rect 1922 -5584 1968 -5572
rect 1922 -5840 1928 -5584
rect 1962 -5840 1968 -5584
rect 1922 -5852 1968 -5840
rect 2100 -5584 2146 -5572
rect 2100 -5840 2106 -5584
rect 2140 -5840 2146 -5584
rect 2100 -5852 2146 -5840
rect 2278 -5584 2324 -5572
rect 2278 -5840 2284 -5584
rect 2318 -5840 2324 -5584
rect 2278 -5852 2324 -5840
rect 2456 -5584 2502 -5572
rect 2456 -5840 2462 -5584
rect 2496 -5840 2502 -5584
rect 2456 -5852 2502 -5840
rect 2634 -5584 2680 -5572
rect 2634 -5840 2640 -5584
rect 2674 -5840 2680 -5584
rect 2634 -5852 2680 -5840
rect -1386 -5899 -1310 -5893
rect -1386 -5933 -1370 -5899
rect -1326 -5933 -1310 -5899
rect -1386 -5949 -1310 -5933
rect -1274 -6364 -1240 -5852
rect -1208 -5899 -1132 -5893
rect -1208 -5933 -1192 -5899
rect -1148 -5933 -1132 -5899
rect -1208 -5949 -1132 -5933
rect -1886 -6417 -1876 -6364
rect -1823 -6417 -1813 -6364
rect -1292 -6417 -1282 -6364
rect -1229 -6417 -1219 -6364
rect -1099 -6479 -1065 -5852
rect -1030 -5899 -954 -5893
rect -1030 -5933 -1014 -5899
rect -970 -5933 -954 -5899
rect -1030 -5949 -954 -5933
rect -919 -6365 -885 -5852
rect -852 -5899 -776 -5893
rect -852 -5933 -836 -5899
rect -792 -5933 -776 -5899
rect -852 -5949 -776 -5933
rect -938 -6417 -928 -6365
rect -876 -6417 -866 -6365
rect -742 -6479 -708 -5852
rect -674 -5899 -598 -5893
rect -674 -5933 -658 -5899
rect -614 -5933 -598 -5899
rect -674 -5949 -598 -5933
rect -496 -5899 -420 -5893
rect -496 -5933 -480 -5899
rect -436 -5933 -420 -5899
rect -496 -5949 -420 -5933
rect -318 -5899 -242 -5893
rect -318 -5933 -302 -5899
rect -258 -5933 -242 -5899
rect -318 -5949 -242 -5933
rect -1120 -6532 -1110 -6479
rect -1057 -6532 -1047 -6479
rect -762 -6532 -752 -6479
rect -699 -6532 -689 -6479
rect -476 -6493 -442 -5949
rect -208 -6077 -174 -5852
rect -140 -5899 -64 -5893
rect -140 -5933 -124 -5899
rect -80 -5933 -64 -5899
rect -140 -5949 -64 -5933
rect 38 -5899 114 -5893
rect 38 -5933 54 -5899
rect 98 -5933 114 -5899
rect 38 -5949 114 -5933
rect 149 -6077 183 -5852
rect 216 -5899 292 -5893
rect 216 -5933 232 -5899
rect 276 -5933 292 -5899
rect 216 -5949 292 -5933
rect 394 -5899 470 -5893
rect 394 -5933 410 -5899
rect 454 -5933 470 -5899
rect 394 -5949 470 -5933
rect 572 -5899 648 -5893
rect 572 -5933 588 -5899
rect 632 -5933 648 -5899
rect 572 -5949 648 -5933
rect 750 -5899 826 -5893
rect 750 -5933 766 -5899
rect 810 -5933 826 -5899
rect 750 -5949 826 -5933
rect 928 -5899 1004 -5893
rect 928 -5933 944 -5899
rect 988 -5933 1004 -5899
rect 928 -5949 1004 -5933
rect -208 -6111 183 -6077
rect 237 -6250 271 -5949
rect 217 -6303 227 -6250
rect 280 -6303 290 -6250
rect 594 -6493 628 -5949
rect 951 -6250 985 -5949
rect 1038 -6081 1072 -5852
rect 1106 -5899 1182 -5893
rect 1106 -5933 1122 -5899
rect 1166 -5933 1182 -5899
rect 1106 -5949 1182 -5933
rect 1284 -5899 1360 -5893
rect 1284 -5933 1300 -5899
rect 1344 -5933 1360 -5899
rect 1284 -5949 1360 -5933
rect 1394 -6081 1428 -5852
rect 1462 -5899 1538 -5893
rect 1462 -5933 1478 -5899
rect 1522 -5933 1538 -5899
rect 1462 -5949 1538 -5933
rect 1640 -5899 1716 -5893
rect 1640 -5933 1656 -5899
rect 1700 -5933 1716 -5899
rect 1640 -5949 1716 -5933
rect 1818 -5899 1894 -5893
rect 1818 -5933 1834 -5899
rect 1878 -5933 1894 -5899
rect 1818 -5949 1894 -5933
rect 1038 -6115 1428 -6081
rect 932 -6303 942 -6250
rect 995 -6303 1005 -6250
rect 1662 -6493 1696 -5949
rect 1928 -6124 1962 -5852
rect 1996 -5899 2072 -5893
rect 1996 -5933 2012 -5899
rect 2056 -5933 2072 -5899
rect 1996 -5949 2072 -5933
rect 2106 -6007 2140 -5852
rect 2174 -5899 2250 -5893
rect 2174 -5933 2190 -5899
rect 2234 -5933 2250 -5899
rect 2174 -5949 2250 -5933
rect 2086 -6060 2096 -6007
rect 2149 -6060 2159 -6007
rect 2284 -6124 2318 -5852
rect 2352 -5899 2428 -5893
rect 2352 -5933 2368 -5899
rect 2412 -5933 2428 -5899
rect 2352 -5949 2428 -5933
rect 2462 -6007 2496 -5852
rect 2530 -5899 2606 -5893
rect 2530 -5933 2546 -5899
rect 2590 -5933 2606 -5899
rect 2530 -5949 2606 -5933
rect 2442 -6060 2452 -6007
rect 2505 -6060 2515 -6007
rect 1908 -6177 1918 -6124
rect 1971 -6177 1981 -6124
rect 2265 -6177 2275 -6124
rect 2328 -6177 2338 -6124
rect 2879 -6365 2931 -2606
rect 3194 -4805 3246 -2480
rect 3184 -4857 3194 -4805
rect 3246 -4857 3256 -4805
rect 4761 -4857 4771 -4805
rect 4823 -4857 4833 -4805
rect 2869 -6417 2879 -6365
rect 2931 -6417 2941 -6365
rect -476 -6527 1696 -6493
rect -742 -6598 -708 -6532
rect 4771 -6597 4823 -4857
rect 5027 -5059 5037 -5006
rect 5090 -5059 5100 -5006
rect 4895 -5265 4905 -5212
rect 4958 -5265 4968 -5212
rect -763 -6651 -753 -6598
rect -700 -6651 -690 -6598
rect 4762 -6650 4772 -6597
rect 4825 -6650 4835 -6597
rect -2013 -6767 -2003 -6714
rect -1950 -6767 -1940 -6714
rect 4771 -6891 4823 -6650
rect 4905 -6889 4958 -5265
rect 5037 -6887 5090 -5059
rect 4760 -6944 4770 -6891
rect 4823 -6944 4833 -6891
rect 4896 -6942 4906 -6889
rect 4959 -6942 4969 -6889
rect 5028 -6940 5038 -6887
rect 5091 -6940 5101 -6887
rect -3883 -7697 -3873 -7691
rect -5629 -7731 -3873 -7697
rect -5628 -7862 -5594 -7731
rect -5544 -7774 -5500 -7731
rect -5560 -7790 -5484 -7774
rect -5560 -7824 -5544 -7790
rect -5500 -7824 -5484 -7790
rect -5560 -7830 -5484 -7824
rect -5450 -7862 -5416 -7731
rect -5366 -7774 -5322 -7731
rect -5188 -7774 -5144 -7731
rect -5382 -7790 -5306 -7774
rect -5382 -7824 -5366 -7790
rect -5322 -7824 -5306 -7790
rect -5382 -7830 -5306 -7824
rect -5204 -7790 -5128 -7774
rect -5204 -7824 -5188 -7790
rect -5144 -7824 -5128 -7790
rect -5204 -7830 -5128 -7824
rect -5094 -7862 -5060 -7731
rect -5010 -7774 -4966 -7731
rect -4832 -7774 -4788 -7731
rect -5026 -7790 -4950 -7774
rect -5026 -7824 -5010 -7790
rect -4966 -7824 -4950 -7790
rect -5026 -7830 -4950 -7824
rect -4848 -7790 -4772 -7774
rect -4848 -7824 -4832 -7790
rect -4788 -7824 -4772 -7790
rect -4848 -7830 -4772 -7824
rect -4738 -7862 -4704 -7731
rect -4654 -7774 -4610 -7731
rect -4476 -7774 -4432 -7731
rect -4670 -7790 -4594 -7774
rect -4670 -7824 -4654 -7790
rect -4610 -7824 -4594 -7790
rect -4670 -7830 -4594 -7824
rect -4492 -7790 -4416 -7774
rect -4492 -7824 -4476 -7790
rect -4432 -7824 -4416 -7790
rect -4492 -7830 -4416 -7824
rect -4382 -7862 -4348 -7731
rect -4298 -7774 -4254 -7731
rect -3883 -7743 -3873 -7731
rect -3821 -7743 -3811 -7691
rect -4314 -7790 -4238 -7774
rect -4314 -7824 -4298 -7790
rect -4254 -7824 -4238 -7790
rect -4314 -7830 -4238 -7824
rect -4136 -7790 -4060 -7774
rect -3741 -7790 -3731 -7785
rect -4136 -7824 -4120 -7790
rect -4076 -7824 -4060 -7790
rect -4136 -7830 -4060 -7824
rect -4026 -7824 -3731 -7790
rect -4026 -7862 -3992 -7824
rect -3741 -7837 -3731 -7824
rect -3679 -7837 -3669 -7785
rect -3551 -7840 -3541 -7788
rect -3489 -7840 -3479 -7788
rect -5634 -7874 -5588 -7862
rect -5634 -8130 -5628 -7874
rect -5594 -8130 -5588 -7874
rect -5634 -8142 -5588 -8130
rect -5456 -7874 -5410 -7862
rect -5456 -8130 -5450 -7874
rect -5416 -8130 -5410 -7874
rect -5456 -8142 -5410 -8130
rect -5278 -7874 -5232 -7862
rect -5278 -8130 -5272 -7874
rect -5238 -8130 -5232 -7874
rect -5278 -8142 -5232 -8130
rect -5100 -7874 -5054 -7862
rect -5100 -8130 -5094 -7874
rect -5060 -8130 -5054 -7874
rect -5100 -8142 -5054 -8130
rect -4922 -7874 -4876 -7862
rect -4922 -8130 -4916 -7874
rect -4882 -8130 -4876 -7874
rect -4922 -8142 -4876 -8130
rect -4744 -7874 -4698 -7862
rect -4744 -8130 -4738 -7874
rect -4704 -8130 -4698 -7874
rect -4744 -8142 -4698 -8130
rect -4566 -7874 -4520 -7862
rect -4566 -8130 -4560 -7874
rect -4526 -8130 -4520 -7874
rect -4566 -8142 -4520 -8130
rect -4388 -7874 -4342 -7862
rect -4388 -8130 -4382 -7874
rect -4348 -8130 -4342 -7874
rect -4388 -8142 -4342 -8130
rect -4210 -7874 -4164 -7862
rect -4210 -8130 -4204 -7874
rect -4170 -8130 -4164 -7874
rect -4210 -8142 -4164 -8130
rect -4032 -7874 -3986 -7862
rect -4032 -8130 -4026 -7874
rect -3992 -8130 -3986 -7874
rect -4032 -8142 -3986 -8130
rect -5628 -8412 -5594 -8142
rect -5560 -8180 -5484 -8174
rect -5560 -8214 -5544 -8180
rect -5500 -8214 -5484 -8180
rect -5560 -8230 -5484 -8214
rect -5544 -8324 -5500 -8230
rect -5560 -8340 -5484 -8324
rect -5560 -8374 -5544 -8340
rect -5500 -8374 -5484 -8340
rect -5560 -8380 -5484 -8374
rect -5450 -8412 -5416 -8142
rect -5382 -8180 -5306 -8174
rect -5382 -8214 -5366 -8180
rect -5322 -8214 -5306 -8180
rect -5382 -8230 -5306 -8214
rect -5366 -8324 -5322 -8230
rect -5382 -8340 -5306 -8324
rect -5382 -8374 -5366 -8340
rect -5322 -8374 -5306 -8340
rect -5382 -8380 -5306 -8374
rect -5272 -8412 -5238 -8142
rect -5204 -8180 -5128 -8174
rect -5204 -8214 -5188 -8180
rect -5144 -8214 -5128 -8180
rect -5204 -8230 -5128 -8214
rect -5188 -8324 -5144 -8230
rect -5204 -8340 -5128 -8324
rect -5204 -8374 -5188 -8340
rect -5144 -8374 -5128 -8340
rect -5204 -8380 -5128 -8374
rect -5094 -8412 -5060 -8142
rect -5026 -8180 -4950 -8174
rect -5026 -8214 -5010 -8180
rect -4966 -8214 -4950 -8180
rect -5026 -8230 -4950 -8214
rect -5010 -8324 -4966 -8230
rect -5026 -8340 -4950 -8324
rect -5026 -8374 -5010 -8340
rect -4966 -8374 -4950 -8340
rect -5026 -8380 -4950 -8374
rect -4916 -8412 -4882 -8142
rect -4848 -8180 -4772 -8174
rect -4848 -8214 -4832 -8180
rect -4788 -8214 -4772 -8180
rect -4848 -8230 -4772 -8214
rect -4832 -8324 -4788 -8230
rect -4848 -8340 -4772 -8324
rect -4848 -8374 -4832 -8340
rect -4788 -8374 -4772 -8340
rect -4848 -8380 -4772 -8374
rect -4738 -8412 -4704 -8142
rect -4670 -8180 -4594 -8174
rect -4670 -8214 -4654 -8180
rect -4610 -8214 -4594 -8180
rect -4670 -8230 -4594 -8214
rect -4654 -8324 -4610 -8230
rect -4670 -8340 -4594 -8324
rect -4670 -8374 -4654 -8340
rect -4610 -8374 -4594 -8340
rect -4670 -8380 -4594 -8374
rect -4560 -8412 -4526 -8142
rect -4492 -8180 -4416 -8174
rect -4492 -8214 -4476 -8180
rect -4432 -8214 -4416 -8180
rect -4492 -8230 -4416 -8214
rect -4476 -8324 -4432 -8230
rect -4492 -8340 -4416 -8324
rect -4492 -8374 -4476 -8340
rect -4432 -8374 -4416 -8340
rect -4492 -8380 -4416 -8374
rect -4382 -8412 -4348 -8142
rect -4314 -8180 -4238 -8174
rect -4314 -8214 -4298 -8180
rect -4254 -8214 -4238 -8180
rect -4314 -8230 -4238 -8214
rect -4298 -8324 -4254 -8230
rect -4314 -8340 -4238 -8324
rect -4314 -8374 -4298 -8340
rect -4254 -8374 -4238 -8340
rect -4314 -8380 -4238 -8374
rect -4204 -8412 -4170 -8142
rect -4136 -8180 -4060 -8174
rect -4136 -8214 -4120 -8180
rect -4076 -8214 -4060 -8180
rect -4136 -8230 -4060 -8214
rect -4120 -8324 -4076 -8230
rect -4136 -8340 -4060 -8324
rect -4136 -8374 -4120 -8340
rect -4076 -8374 -4060 -8340
rect -4136 -8380 -4060 -8374
rect -4026 -8412 -3992 -8142
rect -5634 -8424 -5588 -8412
rect -5634 -8680 -5628 -8424
rect -5594 -8680 -5588 -8424
rect -5634 -8692 -5588 -8680
rect -5456 -8424 -5410 -8412
rect -5456 -8680 -5450 -8424
rect -5416 -8680 -5410 -8424
rect -5456 -8692 -5410 -8680
rect -5278 -8424 -5232 -8412
rect -5278 -8680 -5272 -8424
rect -5238 -8680 -5232 -8424
rect -5278 -8692 -5232 -8680
rect -5100 -8424 -5054 -8412
rect -5100 -8680 -5094 -8424
rect -5060 -8680 -5054 -8424
rect -5100 -8692 -5054 -8680
rect -4922 -8424 -4876 -8412
rect -4922 -8680 -4916 -8424
rect -4882 -8680 -4876 -8424
rect -4922 -8692 -4876 -8680
rect -4744 -8424 -4698 -8412
rect -4744 -8680 -4738 -8424
rect -4704 -8680 -4698 -8424
rect -4744 -8692 -4698 -8680
rect -4566 -8424 -4520 -8412
rect -4566 -8680 -4560 -8424
rect -4526 -8680 -4520 -8424
rect -4566 -8692 -4520 -8680
rect -4388 -8424 -4342 -8412
rect -4388 -8680 -4382 -8424
rect -4348 -8680 -4342 -8424
rect -4388 -8692 -4342 -8680
rect -4210 -8424 -4164 -8412
rect -4210 -8680 -4204 -8424
rect -4170 -8680 -4164 -8424
rect -4210 -8692 -4164 -8680
rect -4032 -8424 -3986 -8412
rect -4032 -8680 -4026 -8424
rect -3992 -8680 -3986 -8424
rect -4032 -8692 -3986 -8680
rect -5628 -8962 -5594 -8692
rect -5560 -8730 -5484 -8724
rect -5560 -8764 -5544 -8730
rect -5500 -8764 -5484 -8730
rect -5560 -8780 -5484 -8764
rect -5544 -8874 -5500 -8780
rect -5560 -8890 -5484 -8874
rect -5560 -8924 -5544 -8890
rect -5500 -8924 -5484 -8890
rect -5560 -8930 -5484 -8924
rect -5450 -8962 -5416 -8692
rect -5382 -8730 -5306 -8724
rect -5382 -8764 -5366 -8730
rect -5322 -8764 -5306 -8730
rect -5382 -8780 -5306 -8764
rect -5366 -8874 -5322 -8780
rect -5382 -8890 -5306 -8874
rect -5382 -8924 -5366 -8890
rect -5322 -8924 -5306 -8890
rect -5382 -8930 -5306 -8924
rect -5272 -8962 -5238 -8692
rect -5204 -8730 -5128 -8724
rect -5204 -8764 -5188 -8730
rect -5144 -8764 -5128 -8730
rect -5204 -8780 -5128 -8764
rect -5188 -8874 -5144 -8780
rect -5204 -8890 -5128 -8874
rect -5204 -8924 -5188 -8890
rect -5144 -8924 -5128 -8890
rect -5204 -8930 -5128 -8924
rect -5094 -8962 -5060 -8692
rect -5026 -8730 -4950 -8724
rect -5026 -8764 -5010 -8730
rect -4966 -8764 -4950 -8730
rect -5026 -8780 -4950 -8764
rect -5010 -8874 -4966 -8780
rect -5026 -8890 -4950 -8874
rect -5026 -8924 -5010 -8890
rect -4966 -8924 -4950 -8890
rect -5026 -8930 -4950 -8924
rect -4916 -8962 -4882 -8692
rect -4848 -8730 -4772 -8724
rect -4848 -8764 -4832 -8730
rect -4788 -8764 -4772 -8730
rect -4848 -8780 -4772 -8764
rect -4832 -8874 -4788 -8780
rect -4848 -8890 -4772 -8874
rect -4848 -8924 -4832 -8890
rect -4788 -8924 -4772 -8890
rect -4848 -8930 -4772 -8924
rect -4738 -8962 -4704 -8692
rect -4670 -8730 -4594 -8724
rect -4670 -8764 -4654 -8730
rect -4610 -8764 -4594 -8730
rect -4670 -8780 -4594 -8764
rect -4654 -8874 -4610 -8780
rect -4670 -8890 -4594 -8874
rect -4670 -8924 -4654 -8890
rect -4610 -8924 -4594 -8890
rect -4670 -8930 -4594 -8924
rect -4560 -8962 -4526 -8692
rect -4492 -8730 -4416 -8724
rect -4492 -8764 -4476 -8730
rect -4432 -8764 -4416 -8730
rect -4492 -8780 -4416 -8764
rect -4476 -8874 -4432 -8780
rect -4492 -8890 -4416 -8874
rect -4492 -8924 -4476 -8890
rect -4432 -8924 -4416 -8890
rect -4492 -8930 -4416 -8924
rect -4382 -8962 -4348 -8692
rect -4314 -8730 -4238 -8724
rect -4314 -8764 -4298 -8730
rect -4254 -8764 -4238 -8730
rect -4314 -8780 -4238 -8764
rect -4298 -8874 -4254 -8780
rect -4314 -8890 -4238 -8874
rect -4314 -8924 -4298 -8890
rect -4254 -8924 -4238 -8890
rect -4314 -8930 -4238 -8924
rect -4204 -8962 -4170 -8692
rect -4136 -8730 -4060 -8724
rect -4136 -8764 -4120 -8730
rect -4076 -8764 -4060 -8730
rect -4136 -8780 -4060 -8764
rect -4120 -8874 -4076 -8780
rect -4136 -8890 -4060 -8874
rect -4136 -8924 -4120 -8890
rect -4076 -8924 -4060 -8890
rect -4136 -8930 -4060 -8924
rect -4026 -8962 -3992 -8692
rect -5634 -8974 -5588 -8962
rect -5634 -9230 -5628 -8974
rect -5594 -9230 -5588 -8974
rect -5634 -9242 -5588 -9230
rect -5456 -8974 -5410 -8962
rect -5456 -9230 -5450 -8974
rect -5416 -9230 -5410 -8974
rect -5456 -9242 -5410 -9230
rect -5278 -8974 -5232 -8962
rect -5278 -9230 -5272 -8974
rect -5238 -9230 -5232 -8974
rect -5278 -9242 -5232 -9230
rect -5100 -8974 -5054 -8962
rect -5100 -9230 -5094 -8974
rect -5060 -9230 -5054 -8974
rect -5100 -9242 -5054 -9230
rect -4922 -8974 -4876 -8962
rect -4922 -9230 -4916 -8974
rect -4882 -9230 -4876 -8974
rect -4922 -9242 -4876 -9230
rect -4744 -8974 -4698 -8962
rect -4744 -9230 -4738 -8974
rect -4704 -9230 -4698 -8974
rect -4744 -9242 -4698 -9230
rect -4566 -8974 -4520 -8962
rect -4566 -9230 -4560 -8974
rect -4526 -9230 -4520 -8974
rect -4566 -9242 -4520 -9230
rect -4388 -8974 -4342 -8962
rect -4388 -9230 -4382 -8974
rect -4348 -9230 -4342 -8974
rect -4388 -9242 -4342 -9230
rect -4210 -8974 -4164 -8962
rect -4210 -9230 -4204 -8974
rect -4170 -9230 -4164 -8974
rect -4210 -9242 -4164 -9230
rect -4032 -8974 -3986 -8962
rect -4032 -9230 -4026 -8974
rect -3992 -9230 -3986 -8974
rect -4032 -9242 -3986 -9230
rect -5628 -9512 -5594 -9242
rect -5560 -9280 -5484 -9274
rect -5560 -9314 -5544 -9280
rect -5500 -9314 -5484 -9280
rect -5560 -9330 -5484 -9314
rect -5544 -9424 -5500 -9330
rect -5560 -9440 -5484 -9424
rect -5560 -9474 -5544 -9440
rect -5500 -9474 -5484 -9440
rect -5560 -9480 -5484 -9474
rect -5450 -9512 -5416 -9242
rect -5382 -9280 -5306 -9274
rect -5382 -9314 -5366 -9280
rect -5322 -9314 -5306 -9280
rect -5382 -9330 -5306 -9314
rect -5366 -9424 -5322 -9330
rect -5382 -9440 -5306 -9424
rect -5382 -9474 -5366 -9440
rect -5322 -9474 -5306 -9440
rect -5382 -9480 -5306 -9474
rect -5272 -9512 -5238 -9242
rect -5204 -9280 -5128 -9274
rect -5204 -9314 -5188 -9280
rect -5144 -9314 -5128 -9280
rect -5204 -9330 -5128 -9314
rect -5188 -9424 -5144 -9330
rect -5204 -9440 -5128 -9424
rect -5204 -9474 -5188 -9440
rect -5144 -9474 -5128 -9440
rect -5204 -9480 -5128 -9474
rect -5094 -9512 -5060 -9242
rect -5026 -9280 -4950 -9274
rect -5026 -9314 -5010 -9280
rect -4966 -9314 -4950 -9280
rect -5026 -9330 -4950 -9314
rect -5010 -9424 -4966 -9330
rect -5026 -9440 -4950 -9424
rect -5026 -9474 -5010 -9440
rect -4966 -9474 -4950 -9440
rect -5026 -9480 -4950 -9474
rect -4916 -9512 -4882 -9242
rect -4848 -9280 -4772 -9274
rect -4848 -9314 -4832 -9280
rect -4788 -9314 -4772 -9280
rect -4848 -9330 -4772 -9314
rect -4832 -9424 -4788 -9330
rect -4848 -9440 -4772 -9424
rect -4848 -9474 -4832 -9440
rect -4788 -9474 -4772 -9440
rect -4848 -9480 -4772 -9474
rect -4738 -9512 -4704 -9242
rect -4670 -9280 -4594 -9274
rect -4670 -9314 -4654 -9280
rect -4610 -9314 -4594 -9280
rect -4670 -9330 -4594 -9314
rect -4654 -9424 -4610 -9330
rect -4670 -9440 -4594 -9424
rect -4670 -9474 -4654 -9440
rect -4610 -9474 -4594 -9440
rect -4670 -9480 -4594 -9474
rect -4560 -9512 -4526 -9242
rect -4492 -9280 -4416 -9274
rect -4492 -9314 -4476 -9280
rect -4432 -9314 -4416 -9280
rect -4492 -9330 -4416 -9314
rect -4476 -9424 -4432 -9330
rect -4492 -9440 -4416 -9424
rect -4492 -9474 -4476 -9440
rect -4432 -9474 -4416 -9440
rect -4492 -9480 -4416 -9474
rect -4382 -9512 -4348 -9242
rect -4314 -9280 -4238 -9274
rect -4314 -9314 -4298 -9280
rect -4254 -9314 -4238 -9280
rect -4314 -9330 -4238 -9314
rect -4298 -9424 -4254 -9330
rect -4314 -9440 -4238 -9424
rect -4314 -9474 -4298 -9440
rect -4254 -9474 -4238 -9440
rect -4314 -9480 -4238 -9474
rect -4204 -9512 -4170 -9242
rect -4136 -9280 -4060 -9274
rect -4136 -9314 -4120 -9280
rect -4076 -9314 -4060 -9280
rect -4136 -9330 -4060 -9314
rect -4120 -9424 -4076 -9330
rect -4136 -9440 -4060 -9424
rect -4136 -9474 -4120 -9440
rect -4076 -9474 -4060 -9440
rect -4136 -9480 -4060 -9474
rect -4026 -9512 -3992 -9242
rect -5634 -9524 -5588 -9512
rect -5634 -9780 -5628 -9524
rect -5594 -9780 -5588 -9524
rect -5634 -9792 -5588 -9780
rect -5456 -9524 -5410 -9512
rect -5456 -9780 -5450 -9524
rect -5416 -9780 -5410 -9524
rect -5456 -9792 -5410 -9780
rect -5278 -9524 -5232 -9512
rect -5278 -9780 -5272 -9524
rect -5238 -9780 -5232 -9524
rect -5278 -9792 -5232 -9780
rect -5100 -9524 -5054 -9512
rect -5100 -9780 -5094 -9524
rect -5060 -9780 -5054 -9524
rect -5100 -9792 -5054 -9780
rect -4922 -9524 -4876 -9512
rect -4922 -9780 -4916 -9524
rect -4882 -9780 -4876 -9524
rect -4922 -9792 -4876 -9780
rect -4744 -9524 -4698 -9512
rect -4744 -9780 -4738 -9524
rect -4704 -9780 -4698 -9524
rect -4744 -9792 -4698 -9780
rect -4566 -9524 -4520 -9512
rect -4566 -9780 -4560 -9524
rect -4526 -9780 -4520 -9524
rect -4566 -9792 -4520 -9780
rect -4388 -9524 -4342 -9512
rect -4388 -9780 -4382 -9524
rect -4348 -9780 -4342 -9524
rect -4388 -9792 -4342 -9780
rect -4210 -9524 -4164 -9512
rect -4210 -9780 -4204 -9524
rect -4170 -9780 -4164 -9524
rect -4210 -9792 -4164 -9780
rect -4032 -9524 -3986 -9512
rect -4032 -9780 -4026 -9524
rect -3992 -9780 -3986 -9524
rect -4032 -9792 -3986 -9780
rect -5628 -10062 -5594 -9792
rect -5560 -9830 -5484 -9824
rect -5560 -9864 -5544 -9830
rect -5500 -9864 -5484 -9830
rect -5560 -9880 -5484 -9864
rect -5544 -9974 -5500 -9880
rect -5560 -9990 -5484 -9974
rect -5560 -10024 -5544 -9990
rect -5500 -10024 -5484 -9990
rect -5560 -10030 -5484 -10024
rect -5450 -10062 -5416 -9792
rect -5382 -9830 -5306 -9824
rect -5382 -9864 -5366 -9830
rect -5322 -9864 -5306 -9830
rect -5382 -9880 -5306 -9864
rect -5366 -9974 -5322 -9880
rect -5382 -9990 -5306 -9974
rect -5382 -10024 -5366 -9990
rect -5322 -10024 -5306 -9990
rect -5382 -10030 -5306 -10024
rect -5272 -10062 -5238 -9792
rect -5204 -9830 -5128 -9824
rect -5204 -9864 -5188 -9830
rect -5144 -9864 -5128 -9830
rect -5204 -9880 -5128 -9864
rect -5188 -9974 -5144 -9880
rect -5204 -9990 -5128 -9974
rect -5204 -10024 -5188 -9990
rect -5144 -10024 -5128 -9990
rect -5204 -10030 -5128 -10024
rect -5094 -10062 -5060 -9792
rect -5026 -9830 -4950 -9824
rect -5026 -9864 -5010 -9830
rect -4966 -9864 -4950 -9830
rect -5026 -9880 -4950 -9864
rect -5010 -9974 -4966 -9880
rect -5026 -9990 -4950 -9974
rect -5026 -10024 -5010 -9990
rect -4966 -10024 -4950 -9990
rect -5026 -10030 -4950 -10024
rect -4916 -10062 -4882 -9792
rect -4848 -9830 -4772 -9824
rect -4848 -9864 -4832 -9830
rect -4788 -9864 -4772 -9830
rect -4848 -9880 -4772 -9864
rect -4832 -9974 -4788 -9880
rect -4848 -9990 -4772 -9974
rect -4848 -10024 -4832 -9990
rect -4788 -10024 -4772 -9990
rect -4848 -10030 -4772 -10024
rect -4738 -10062 -4704 -9792
rect -4670 -9830 -4594 -9824
rect -4670 -9864 -4654 -9830
rect -4610 -9864 -4594 -9830
rect -4670 -9880 -4594 -9864
rect -4654 -9974 -4610 -9880
rect -4670 -9990 -4594 -9974
rect -4670 -10024 -4654 -9990
rect -4610 -10024 -4594 -9990
rect -4670 -10030 -4594 -10024
rect -4560 -10062 -4526 -9792
rect -4492 -9830 -4416 -9824
rect -4492 -9864 -4476 -9830
rect -4432 -9864 -4416 -9830
rect -4492 -9880 -4416 -9864
rect -4476 -9974 -4432 -9880
rect -4492 -9990 -4416 -9974
rect -4492 -10024 -4476 -9990
rect -4432 -10024 -4416 -9990
rect -4492 -10030 -4416 -10024
rect -4382 -10062 -4348 -9792
rect -4314 -9830 -4238 -9824
rect -4314 -9864 -4298 -9830
rect -4254 -9864 -4238 -9830
rect -4314 -9880 -4238 -9864
rect -4298 -9974 -4254 -9880
rect -4314 -9990 -4238 -9974
rect -4314 -10024 -4298 -9990
rect -4254 -10024 -4238 -9990
rect -4314 -10030 -4238 -10024
rect -4204 -10062 -4170 -9792
rect -4136 -9830 -4060 -9824
rect -4136 -9864 -4120 -9830
rect -4076 -9864 -4060 -9830
rect -4136 -9880 -4060 -9864
rect -4120 -9974 -4076 -9880
rect -4136 -9990 -4060 -9974
rect -4136 -10024 -4120 -9990
rect -4076 -10024 -4060 -9990
rect -4136 -10030 -4060 -10024
rect -4026 -10062 -3992 -9792
rect -5634 -10074 -5588 -10062
rect -5634 -10330 -5628 -10074
rect -5594 -10330 -5588 -10074
rect -5634 -10342 -5588 -10330
rect -5456 -10074 -5410 -10062
rect -5456 -10330 -5450 -10074
rect -5416 -10330 -5410 -10074
rect -5456 -10342 -5410 -10330
rect -5278 -10074 -5232 -10062
rect -5278 -10330 -5272 -10074
rect -5238 -10330 -5232 -10074
rect -5278 -10342 -5232 -10330
rect -5100 -10074 -5054 -10062
rect -5100 -10330 -5094 -10074
rect -5060 -10330 -5054 -10074
rect -5100 -10342 -5054 -10330
rect -4922 -10074 -4876 -10062
rect -4922 -10330 -4916 -10074
rect -4882 -10330 -4876 -10074
rect -4922 -10342 -4876 -10330
rect -4744 -10074 -4698 -10062
rect -4744 -10330 -4738 -10074
rect -4704 -10330 -4698 -10074
rect -4744 -10342 -4698 -10330
rect -4566 -10074 -4520 -10062
rect -4566 -10330 -4560 -10074
rect -4526 -10330 -4520 -10074
rect -4566 -10342 -4520 -10330
rect -4388 -10074 -4342 -10062
rect -4388 -10330 -4382 -10074
rect -4348 -10330 -4342 -10074
rect -4388 -10342 -4342 -10330
rect -4210 -10074 -4164 -10062
rect -4210 -10330 -4204 -10074
rect -4170 -10330 -4164 -10074
rect -4210 -10342 -4164 -10330
rect -4032 -10074 -3986 -10062
rect -4032 -10330 -4026 -10074
rect -3992 -10330 -3986 -10074
rect -4032 -10342 -3986 -10330
rect -5628 -10612 -5594 -10342
rect -5560 -10380 -5484 -10374
rect -5560 -10414 -5544 -10380
rect -5500 -10414 -5484 -10380
rect -5560 -10430 -5484 -10414
rect -5544 -10524 -5500 -10430
rect -5560 -10540 -5484 -10524
rect -5560 -10574 -5544 -10540
rect -5500 -10574 -5484 -10540
rect -5560 -10580 -5484 -10574
rect -5450 -10612 -5416 -10342
rect -5382 -10380 -5306 -10374
rect -5382 -10414 -5366 -10380
rect -5322 -10414 -5306 -10380
rect -5382 -10430 -5306 -10414
rect -5366 -10524 -5322 -10430
rect -5382 -10540 -5306 -10524
rect -5382 -10574 -5366 -10540
rect -5322 -10574 -5306 -10540
rect -5382 -10580 -5306 -10574
rect -5272 -10612 -5238 -10342
rect -5204 -10380 -5128 -10374
rect -5204 -10414 -5188 -10380
rect -5144 -10414 -5128 -10380
rect -5204 -10430 -5128 -10414
rect -5188 -10524 -5144 -10430
rect -5204 -10540 -5128 -10524
rect -5204 -10574 -5188 -10540
rect -5144 -10574 -5128 -10540
rect -5204 -10580 -5128 -10574
rect -5094 -10612 -5060 -10342
rect -5026 -10380 -4950 -10374
rect -5026 -10414 -5010 -10380
rect -4966 -10414 -4950 -10380
rect -5026 -10430 -4950 -10414
rect -5010 -10524 -4966 -10430
rect -5026 -10540 -4950 -10524
rect -5026 -10574 -5010 -10540
rect -4966 -10574 -4950 -10540
rect -5026 -10580 -4950 -10574
rect -4916 -10612 -4882 -10342
rect -4848 -10380 -4772 -10374
rect -4848 -10414 -4832 -10380
rect -4788 -10414 -4772 -10380
rect -4848 -10430 -4772 -10414
rect -4832 -10524 -4788 -10430
rect -4848 -10540 -4772 -10524
rect -4848 -10574 -4832 -10540
rect -4788 -10574 -4772 -10540
rect -4848 -10580 -4772 -10574
rect -4738 -10612 -4704 -10342
rect -4670 -10380 -4594 -10374
rect -4670 -10414 -4654 -10380
rect -4610 -10414 -4594 -10380
rect -4670 -10430 -4594 -10414
rect -4654 -10524 -4610 -10430
rect -4670 -10540 -4594 -10524
rect -4670 -10574 -4654 -10540
rect -4610 -10574 -4594 -10540
rect -4670 -10580 -4594 -10574
rect -4560 -10612 -4526 -10342
rect -4492 -10380 -4416 -10374
rect -4492 -10414 -4476 -10380
rect -4432 -10414 -4416 -10380
rect -4492 -10430 -4416 -10414
rect -4476 -10524 -4432 -10430
rect -4492 -10540 -4416 -10524
rect -4492 -10574 -4476 -10540
rect -4432 -10574 -4416 -10540
rect -4492 -10580 -4416 -10574
rect -4382 -10612 -4348 -10342
rect -4314 -10380 -4238 -10374
rect -4314 -10414 -4298 -10380
rect -4254 -10414 -4238 -10380
rect -4314 -10430 -4238 -10414
rect -4298 -10524 -4254 -10430
rect -4314 -10540 -4238 -10524
rect -4314 -10574 -4298 -10540
rect -4254 -10574 -4238 -10540
rect -4314 -10580 -4238 -10574
rect -4204 -10612 -4170 -10342
rect -4136 -10380 -4060 -10374
rect -4136 -10414 -4120 -10380
rect -4076 -10414 -4060 -10380
rect -4136 -10430 -4060 -10414
rect -4120 -10524 -4076 -10430
rect -4136 -10540 -4060 -10524
rect -4136 -10574 -4120 -10540
rect -4076 -10574 -4060 -10540
rect -4136 -10580 -4060 -10574
rect -4026 -10612 -3992 -10342
rect -5634 -10624 -5588 -10612
rect -5634 -10880 -5628 -10624
rect -5594 -10880 -5588 -10624
rect -5634 -10892 -5588 -10880
rect -5456 -10624 -5410 -10612
rect -5456 -10880 -5450 -10624
rect -5416 -10880 -5410 -10624
rect -5456 -10892 -5410 -10880
rect -5278 -10624 -5232 -10612
rect -5278 -10880 -5272 -10624
rect -5238 -10880 -5232 -10624
rect -5278 -10892 -5232 -10880
rect -5100 -10624 -5054 -10612
rect -5100 -10880 -5094 -10624
rect -5060 -10880 -5054 -10624
rect -5100 -10892 -5054 -10880
rect -4922 -10624 -4876 -10612
rect -4922 -10880 -4916 -10624
rect -4882 -10880 -4876 -10624
rect -4922 -10892 -4876 -10880
rect -4744 -10624 -4698 -10612
rect -4744 -10880 -4738 -10624
rect -4704 -10880 -4698 -10624
rect -4744 -10892 -4698 -10880
rect -4566 -10624 -4520 -10612
rect -4566 -10880 -4560 -10624
rect -4526 -10880 -4520 -10624
rect -4566 -10892 -4520 -10880
rect -4388 -10624 -4342 -10612
rect -4388 -10880 -4382 -10624
rect -4348 -10880 -4342 -10624
rect -4388 -10892 -4342 -10880
rect -4210 -10624 -4164 -10612
rect -4210 -10880 -4204 -10624
rect -4170 -10880 -4164 -10624
rect -4210 -10892 -4164 -10880
rect -4032 -10624 -3986 -10612
rect -4032 -10880 -4026 -10624
rect -3992 -10880 -3986 -10624
rect -4032 -10892 -3986 -10880
rect -5628 -11162 -5594 -10892
rect -5560 -10930 -5484 -10924
rect -5560 -10964 -5544 -10930
rect -5500 -10964 -5484 -10930
rect -5560 -10980 -5484 -10964
rect -5544 -11074 -5500 -10980
rect -5560 -11090 -5484 -11074
rect -5560 -11124 -5544 -11090
rect -5500 -11124 -5484 -11090
rect -5560 -11130 -5484 -11124
rect -5450 -11162 -5416 -10892
rect -5382 -10930 -5306 -10924
rect -5382 -10964 -5366 -10930
rect -5322 -10964 -5306 -10930
rect -5382 -10980 -5306 -10964
rect -5366 -11074 -5322 -10980
rect -5382 -11090 -5306 -11074
rect -5382 -11124 -5366 -11090
rect -5322 -11124 -5306 -11090
rect -5382 -11130 -5306 -11124
rect -5272 -11162 -5238 -10892
rect -5204 -10930 -5128 -10924
rect -5204 -10964 -5188 -10930
rect -5144 -10964 -5128 -10930
rect -5204 -10980 -5128 -10964
rect -5188 -11074 -5144 -10980
rect -5204 -11090 -5128 -11074
rect -5204 -11124 -5188 -11090
rect -5144 -11124 -5128 -11090
rect -5204 -11130 -5128 -11124
rect -5094 -11162 -5060 -10892
rect -5026 -10930 -4950 -10924
rect -5026 -10964 -5010 -10930
rect -4966 -10964 -4950 -10930
rect -5026 -10980 -4950 -10964
rect -5010 -11074 -4966 -10980
rect -5026 -11090 -4950 -11074
rect -5026 -11124 -5010 -11090
rect -4966 -11124 -4950 -11090
rect -5026 -11130 -4950 -11124
rect -4916 -11162 -4882 -10892
rect -4848 -10930 -4772 -10924
rect -4848 -10964 -4832 -10930
rect -4788 -10964 -4772 -10930
rect -4848 -10980 -4772 -10964
rect -4832 -11074 -4788 -10980
rect -4848 -11090 -4772 -11074
rect -4848 -11124 -4832 -11090
rect -4788 -11124 -4772 -11090
rect -4848 -11130 -4772 -11124
rect -4738 -11162 -4704 -10892
rect -4670 -10930 -4594 -10924
rect -4670 -10964 -4654 -10930
rect -4610 -10964 -4594 -10930
rect -4670 -10980 -4594 -10964
rect -4654 -11074 -4610 -10980
rect -4670 -11090 -4594 -11074
rect -4670 -11124 -4654 -11090
rect -4610 -11124 -4594 -11090
rect -4670 -11130 -4594 -11124
rect -4560 -11162 -4526 -10892
rect -4492 -10930 -4416 -10924
rect -4492 -10964 -4476 -10930
rect -4432 -10964 -4416 -10930
rect -4492 -10980 -4416 -10964
rect -4476 -11074 -4432 -10980
rect -4492 -11090 -4416 -11074
rect -4492 -11124 -4476 -11090
rect -4432 -11124 -4416 -11090
rect -4492 -11130 -4416 -11124
rect -4382 -11162 -4348 -10892
rect -4314 -10930 -4238 -10924
rect -4314 -10964 -4298 -10930
rect -4254 -10964 -4238 -10930
rect -4314 -10980 -4238 -10964
rect -4298 -11074 -4254 -10980
rect -4314 -11090 -4238 -11074
rect -4314 -11124 -4298 -11090
rect -4254 -11124 -4238 -11090
rect -4314 -11130 -4238 -11124
rect -4204 -11162 -4170 -10892
rect -4136 -10930 -4060 -10924
rect -4136 -10964 -4120 -10930
rect -4076 -10964 -4060 -10930
rect -4136 -10980 -4060 -10964
rect -4120 -11074 -4076 -10980
rect -4136 -11090 -4060 -11074
rect -4136 -11124 -4120 -11090
rect -4076 -11124 -4060 -11090
rect -4136 -11130 -4060 -11124
rect -4026 -11162 -3992 -10892
rect -5634 -11174 -5588 -11162
rect -5634 -11430 -5628 -11174
rect -5594 -11430 -5588 -11174
rect -5634 -11442 -5588 -11430
rect -5456 -11174 -5410 -11162
rect -5456 -11430 -5450 -11174
rect -5416 -11430 -5410 -11174
rect -5456 -11442 -5410 -11430
rect -5278 -11174 -5232 -11162
rect -5278 -11430 -5272 -11174
rect -5238 -11430 -5232 -11174
rect -5278 -11442 -5232 -11430
rect -5100 -11174 -5054 -11162
rect -5100 -11430 -5094 -11174
rect -5060 -11430 -5054 -11174
rect -5100 -11442 -5054 -11430
rect -4922 -11174 -4876 -11162
rect -4922 -11430 -4916 -11174
rect -4882 -11430 -4876 -11174
rect -4922 -11442 -4876 -11430
rect -4744 -11174 -4698 -11162
rect -4744 -11430 -4738 -11174
rect -4704 -11430 -4698 -11174
rect -4744 -11442 -4698 -11430
rect -4566 -11174 -4520 -11162
rect -4566 -11430 -4560 -11174
rect -4526 -11430 -4520 -11174
rect -4566 -11442 -4520 -11430
rect -4388 -11174 -4342 -11162
rect -4388 -11430 -4382 -11174
rect -4348 -11430 -4342 -11174
rect -4388 -11442 -4342 -11430
rect -4210 -11174 -4164 -11162
rect -4210 -11430 -4204 -11174
rect -4170 -11430 -4164 -11174
rect -4210 -11442 -4164 -11430
rect -4032 -11174 -3986 -11162
rect -4032 -11430 -4026 -11174
rect -3992 -11430 -3986 -11174
rect -4032 -11442 -3986 -11430
rect -5628 -11712 -5594 -11442
rect -5560 -11480 -5484 -11474
rect -5560 -11514 -5544 -11480
rect -5500 -11514 -5484 -11480
rect -5560 -11530 -5484 -11514
rect -5544 -11624 -5500 -11530
rect -5560 -11640 -5484 -11624
rect -5560 -11674 -5544 -11640
rect -5500 -11674 -5484 -11640
rect -5560 -11680 -5484 -11674
rect -5450 -11712 -5416 -11442
rect -5382 -11480 -5306 -11474
rect -5382 -11514 -5366 -11480
rect -5322 -11514 -5306 -11480
rect -5382 -11530 -5306 -11514
rect -5364 -11624 -5320 -11530
rect -5382 -11640 -5306 -11624
rect -5382 -11674 -5366 -11640
rect -5322 -11674 -5306 -11640
rect -5382 -11680 -5306 -11674
rect -5272 -11712 -5238 -11442
rect -5204 -11480 -5128 -11474
rect -5204 -11514 -5188 -11480
rect -5144 -11514 -5128 -11480
rect -5204 -11530 -5128 -11514
rect -5188 -11624 -5144 -11530
rect -5204 -11640 -5128 -11624
rect -5204 -11674 -5188 -11640
rect -5144 -11674 -5128 -11640
rect -5204 -11680 -5128 -11674
rect -5094 -11712 -5060 -11442
rect -5026 -11480 -4950 -11474
rect -5026 -11514 -5010 -11480
rect -4966 -11514 -4950 -11480
rect -5026 -11530 -4950 -11514
rect -5010 -11624 -4966 -11530
rect -5026 -11640 -4950 -11624
rect -5026 -11674 -5010 -11640
rect -4966 -11674 -4950 -11640
rect -5026 -11680 -4950 -11674
rect -4916 -11712 -4882 -11442
rect -4848 -11480 -4772 -11474
rect -4848 -11514 -4832 -11480
rect -4788 -11514 -4772 -11480
rect -4848 -11530 -4772 -11514
rect -4832 -11624 -4788 -11530
rect -4848 -11640 -4772 -11624
rect -4848 -11674 -4832 -11640
rect -4788 -11674 -4772 -11640
rect -4848 -11680 -4772 -11674
rect -4738 -11712 -4704 -11442
rect -4670 -11480 -4594 -11474
rect -4670 -11514 -4654 -11480
rect -4610 -11514 -4594 -11480
rect -4670 -11530 -4594 -11514
rect -4654 -11624 -4610 -11530
rect -4670 -11640 -4594 -11624
rect -4670 -11674 -4654 -11640
rect -4610 -11674 -4594 -11640
rect -4670 -11680 -4594 -11674
rect -4560 -11712 -4526 -11442
rect -4492 -11480 -4416 -11474
rect -4492 -11514 -4476 -11480
rect -4432 -11514 -4416 -11480
rect -4492 -11530 -4416 -11514
rect -4476 -11624 -4432 -11530
rect -4492 -11640 -4416 -11624
rect -4492 -11674 -4476 -11640
rect -4432 -11674 -4416 -11640
rect -4492 -11680 -4416 -11674
rect -4382 -11712 -4348 -11442
rect -4314 -11480 -4238 -11474
rect -4314 -11514 -4298 -11480
rect -4254 -11514 -4238 -11480
rect -4314 -11530 -4238 -11514
rect -4298 -11624 -4254 -11530
rect -4314 -11640 -4238 -11624
rect -4314 -11674 -4298 -11640
rect -4254 -11674 -4238 -11640
rect -4314 -11680 -4238 -11674
rect -4204 -11712 -4170 -11442
rect -4136 -11480 -4060 -11474
rect -4136 -11514 -4120 -11480
rect -4076 -11514 -4060 -11480
rect -4136 -11530 -4060 -11514
rect -4120 -11624 -4076 -11530
rect -4136 -11640 -4060 -11624
rect -4136 -11674 -4120 -11640
rect -4076 -11674 -4060 -11640
rect -4136 -11680 -4060 -11674
rect -4026 -11712 -3992 -11442
rect -5634 -11724 -5588 -11712
rect -5634 -11980 -5628 -11724
rect -5594 -11980 -5588 -11724
rect -5634 -11992 -5588 -11980
rect -5456 -11724 -5410 -11712
rect -5456 -11980 -5450 -11724
rect -5416 -11980 -5410 -11724
rect -5456 -11992 -5410 -11980
rect -5278 -11724 -5232 -11712
rect -5278 -11980 -5272 -11724
rect -5238 -11980 -5232 -11724
rect -5278 -11992 -5232 -11980
rect -5100 -11724 -5054 -11712
rect -5100 -11980 -5094 -11724
rect -5060 -11980 -5054 -11724
rect -5100 -11992 -5054 -11980
rect -4922 -11724 -4876 -11712
rect -4922 -11980 -4916 -11724
rect -4882 -11980 -4876 -11724
rect -4922 -11992 -4876 -11980
rect -4744 -11724 -4698 -11712
rect -4744 -11980 -4738 -11724
rect -4704 -11980 -4698 -11724
rect -4744 -11992 -4698 -11980
rect -4566 -11724 -4520 -11712
rect -4566 -11980 -4560 -11724
rect -4526 -11980 -4520 -11724
rect -4566 -11992 -4520 -11980
rect -4388 -11724 -4342 -11712
rect -4388 -11980 -4382 -11724
rect -4348 -11980 -4342 -11724
rect -4388 -11992 -4342 -11980
rect -4210 -11724 -4164 -11712
rect -4210 -11980 -4204 -11724
rect -4170 -11980 -4164 -11724
rect -4210 -11992 -4164 -11980
rect -4032 -11724 -3986 -11712
rect -4032 -11980 -4026 -11724
rect -3992 -11980 -3986 -11724
rect -4032 -11992 -3986 -11980
rect -5560 -12030 -5484 -12024
rect -5560 -12064 -5544 -12030
rect -5500 -12064 -5484 -12030
rect -5560 -12080 -5484 -12064
rect -5382 -12030 -5306 -12024
rect -5382 -12064 -5366 -12030
rect -5322 -12064 -5306 -12030
rect -5382 -12080 -5306 -12064
rect -5272 -12119 -5238 -11992
rect -5204 -12030 -5128 -12024
rect -5204 -12064 -5188 -12030
rect -5144 -12064 -5128 -12030
rect -5204 -12080 -5128 -12064
rect -5026 -12030 -4950 -12024
rect -5026 -12064 -5010 -12030
rect -4966 -12064 -4950 -12030
rect -5026 -12080 -4950 -12064
rect -4916 -12119 -4882 -11992
rect -4848 -12030 -4772 -12024
rect -4848 -12064 -4832 -12030
rect -4788 -12064 -4772 -12030
rect -4848 -12080 -4772 -12064
rect -4670 -12030 -4594 -12024
rect -4670 -12064 -4654 -12030
rect -4610 -12064 -4594 -12030
rect -4670 -12080 -4594 -12064
rect -4560 -12119 -4526 -11992
rect -4492 -12030 -4416 -12024
rect -4492 -12064 -4476 -12030
rect -4432 -12064 -4416 -12030
rect -4492 -12080 -4416 -12064
rect -4314 -12030 -4238 -12024
rect -4314 -12064 -4298 -12030
rect -4254 -12064 -4238 -12030
rect -4314 -12080 -4238 -12064
rect -4204 -12119 -4170 -11992
rect -4136 -12030 -4060 -12024
rect -4136 -12064 -4120 -12030
rect -4076 -12064 -4060 -12030
rect -4136 -12080 -4060 -12064
rect -4113 -12119 -4079 -12080
rect -4026 -12119 -3992 -11992
rect -5272 -12153 -3611 -12119
rect -5512 -12324 -5502 -12271
rect -5449 -12324 -5439 -12271
rect -6976 -12565 -6077 -12512
rect -6024 -12565 -6014 -12512
rect -5636 -12565 -5626 -12512
rect -5573 -12565 -5563 -12512
rect -6233 -13115 -6223 -13062
rect -6170 -13115 -6160 -13062
rect -6976 -13905 -6426 -13852
rect -6373 -13905 -6363 -13852
rect -6223 -14055 -6170 -13115
rect -6077 -13745 -6024 -12565
rect -5617 -12612 -5583 -12565
rect -5922 -12628 -5778 -12612
rect -5922 -12662 -5867 -12628
rect -5833 -12662 -5778 -12628
rect -5922 -12668 -5778 -12662
rect -5633 -12628 -5567 -12612
rect -5633 -12662 -5617 -12628
rect -5583 -12662 -5567 -12628
rect -5633 -12668 -5567 -12662
rect -5922 -12712 -5876 -12668
rect -5922 -12928 -5916 -12712
rect -5882 -12928 -5876 -12712
rect -5922 -12940 -5876 -12928
rect -5824 -12700 -5778 -12668
rect -5492 -12700 -5458 -12324
rect -5010 -12325 -5000 -12272
rect -4947 -12325 -4937 -12272
rect -4512 -12324 -4502 -12271
rect -4449 -12324 -4439 -12271
rect -5386 -12441 -5376 -12388
rect -5323 -12441 -5313 -12388
rect -5137 -12441 -5127 -12388
rect -5074 -12441 -5064 -12388
rect -5367 -12612 -5333 -12441
rect -5117 -12612 -5083 -12441
rect -5383 -12628 -5317 -12612
rect -5383 -12662 -5367 -12628
rect -5333 -12662 -5317 -12628
rect -5383 -12668 -5317 -12662
rect -5133 -12628 -5067 -12612
rect -5133 -12662 -5117 -12628
rect -5083 -12662 -5067 -12628
rect -5133 -12668 -5067 -12662
rect -4992 -12700 -4958 -12325
rect -4887 -12565 -4877 -12512
rect -4824 -12565 -4814 -12512
rect -4637 -12565 -4627 -12512
rect -4574 -12565 -4564 -12512
rect -4867 -12612 -4833 -12565
rect -4617 -12612 -4583 -12565
rect -4883 -12628 -4817 -12612
rect -4883 -12662 -4867 -12628
rect -4833 -12662 -4817 -12628
rect -4883 -12668 -4817 -12662
rect -4633 -12628 -4567 -12612
rect -4633 -12662 -4617 -12628
rect -4583 -12662 -4567 -12628
rect -4633 -12668 -4567 -12662
rect -4492 -12700 -4458 -12324
rect -4387 -12441 -4377 -12388
rect -4324 -12441 -4314 -12388
rect -4367 -12612 -4333 -12441
rect -3938 -12442 -3928 -12389
rect -3875 -12442 -3865 -12389
rect -4383 -12628 -4317 -12612
rect -4383 -12662 -4367 -12628
rect -4333 -12662 -4317 -12628
rect -4383 -12668 -4317 -12662
rect -4172 -12628 -4028 -12612
rect -4172 -12662 -4117 -12628
rect -4083 -12662 -4028 -12628
rect -4172 -12668 -4028 -12662
rect -4172 -12700 -4126 -12668
rect -5824 -12712 -5626 -12700
rect -5824 -12928 -5818 -12712
rect -5784 -12740 -5666 -12712
rect -5784 -12900 -5778 -12740
rect -5672 -12900 -5666 -12740
rect -5784 -12928 -5666 -12900
rect -5632 -12928 -5626 -12712
rect -5824 -12940 -5626 -12928
rect -5574 -12712 -5376 -12700
rect -5574 -12928 -5568 -12712
rect -5534 -12740 -5416 -12712
rect -5534 -12900 -5528 -12740
rect -5422 -12900 -5416 -12740
rect -5534 -12928 -5416 -12900
rect -5382 -12928 -5376 -12712
rect -5574 -12940 -5376 -12928
rect -5324 -12712 -5126 -12700
rect -5324 -12928 -5318 -12712
rect -5284 -12740 -5166 -12712
rect -5284 -12900 -5278 -12740
rect -5172 -12900 -5166 -12740
rect -5284 -12928 -5166 -12900
rect -5132 -12928 -5126 -12712
rect -5324 -12940 -5126 -12928
rect -5074 -12712 -4876 -12700
rect -5074 -12928 -5068 -12712
rect -5034 -12740 -4916 -12712
rect -5034 -12900 -5028 -12740
rect -4922 -12900 -4916 -12740
rect -5034 -12928 -4916 -12900
rect -4882 -12928 -4876 -12712
rect -4824 -12712 -4625 -12700
rect -4824 -12900 -4818 -12712
rect -5074 -12940 -4876 -12928
rect -4825 -12928 -4818 -12900
rect -4784 -12740 -4666 -12712
rect -4784 -12900 -4778 -12740
rect -4672 -12900 -4666 -12740
rect -4784 -12928 -4666 -12900
rect -4632 -12740 -4625 -12712
rect -4574 -12712 -4376 -12700
rect -4632 -12928 -4626 -12740
rect -4825 -12940 -4626 -12928
rect -4574 -12928 -4568 -12712
rect -4534 -12740 -4416 -12712
rect -4534 -12900 -4528 -12740
rect -4422 -12900 -4416 -12740
rect -4534 -12928 -4416 -12900
rect -4382 -12928 -4376 -12712
rect -4574 -12940 -4376 -12928
rect -4324 -12712 -4126 -12700
rect -4324 -12928 -4318 -12712
rect -4284 -12740 -4166 -12712
rect -4284 -12900 -4278 -12740
rect -4172 -12900 -4166 -12740
rect -4284 -12928 -4166 -12900
rect -4132 -12928 -4126 -12712
rect -4324 -12940 -4126 -12928
rect -4074 -12712 -4028 -12668
rect -4074 -12928 -4068 -12712
rect -4034 -12928 -4028 -12712
rect -4074 -12940 -4028 -12928
rect -5883 -12978 -5817 -12972
rect -5883 -13012 -5867 -12978
rect -5833 -13012 -5817 -12978
rect -5883 -13028 -5817 -13012
rect -5744 -13062 -5704 -12940
rect -5633 -12978 -5567 -12972
rect -5633 -13012 -5617 -12978
rect -5583 -13012 -5567 -12978
rect -5633 -13028 -5567 -13012
rect -5761 -13115 -5751 -13062
rect -5698 -13115 -5688 -13062
rect -5883 -13308 -5817 -13292
rect -5883 -13342 -5867 -13308
rect -5833 -13342 -5817 -13308
rect -5883 -13348 -5817 -13342
rect -5633 -13308 -5567 -13292
rect -5633 -13342 -5617 -13308
rect -5583 -13342 -5567 -13308
rect -5633 -13348 -5567 -13342
rect -5495 -13380 -5455 -12940
rect -5383 -12978 -5317 -12972
rect -5383 -13012 -5367 -12978
rect -5333 -13012 -5317 -12978
rect -5383 -13028 -5317 -13012
rect -5245 -13189 -5205 -12940
rect -5133 -12978 -5067 -12972
rect -5133 -13012 -5117 -12978
rect -5083 -13012 -5067 -12978
rect -5133 -13028 -5067 -13012
rect -5261 -13242 -5251 -13189
rect -5198 -13242 -5188 -13189
rect -5383 -13308 -5317 -13292
rect -5383 -13342 -5367 -13308
rect -5333 -13342 -5317 -13308
rect -5383 -13348 -5317 -13342
rect -5133 -13308 -5067 -13292
rect -5133 -13342 -5117 -13308
rect -5083 -13342 -5067 -13308
rect -5133 -13348 -5067 -13342
rect -4995 -13380 -4955 -12940
rect -4883 -12978 -4817 -12972
rect -4883 -13012 -4867 -12978
rect -4833 -13012 -4817 -12978
rect -4883 -13028 -4817 -13012
rect -4746 -13062 -4706 -12940
rect -4633 -12978 -4567 -12972
rect -4633 -13012 -4617 -12978
rect -4583 -13012 -4567 -12978
rect -4633 -13028 -4567 -13012
rect -4762 -13115 -4752 -13062
rect -4699 -13115 -4689 -13062
rect -4883 -13308 -4817 -13292
rect -4883 -13342 -4867 -13308
rect -4833 -13342 -4817 -13308
rect -4883 -13348 -4817 -13342
rect -4633 -13308 -4567 -13292
rect -4633 -13342 -4617 -13308
rect -4583 -13342 -4567 -13308
rect -4633 -13348 -4567 -13342
rect -4495 -13380 -4455 -12940
rect -4383 -12978 -4317 -12972
rect -4383 -13012 -4367 -12978
rect -4333 -13012 -4317 -12978
rect -4383 -13028 -4317 -13012
rect -4244 -13189 -4204 -12940
rect -4133 -12978 -4067 -12972
rect -4133 -13012 -4117 -12978
rect -4083 -13012 -4067 -12978
rect -4133 -13028 -4067 -13012
rect -4261 -13242 -4251 -13189
rect -4198 -13242 -4188 -13189
rect -4383 -13308 -4317 -13292
rect -4383 -13342 -4367 -13308
rect -4333 -13342 -4317 -13308
rect -4383 -13348 -4317 -13342
rect -4133 -13308 -4067 -13292
rect -4133 -13342 -4117 -13308
rect -4083 -13342 -4067 -13308
rect -4133 -13348 -4067 -13342
rect -5922 -13392 -5876 -13380
rect -5922 -13608 -5916 -13392
rect -5882 -13608 -5876 -13392
rect -5922 -13652 -5876 -13608
rect -5824 -13392 -5626 -13380
rect -5824 -13608 -5818 -13392
rect -5784 -13420 -5666 -13392
rect -5784 -13580 -5778 -13420
rect -5672 -13580 -5666 -13420
rect -5784 -13608 -5666 -13580
rect -5632 -13608 -5626 -13392
rect -5824 -13620 -5626 -13608
rect -5574 -13392 -5376 -13380
rect -5574 -13608 -5568 -13392
rect -5534 -13420 -5416 -13392
rect -5534 -13580 -5528 -13420
rect -5422 -13580 -5416 -13420
rect -5534 -13608 -5416 -13580
rect -5382 -13608 -5376 -13392
rect -5574 -13620 -5376 -13608
rect -5324 -13392 -5126 -13380
rect -5324 -13608 -5318 -13392
rect -5284 -13420 -5166 -13392
rect -5284 -13580 -5278 -13420
rect -5172 -13580 -5166 -13420
rect -5284 -13608 -5166 -13580
rect -5132 -13608 -5126 -13392
rect -5324 -13620 -5126 -13608
rect -5074 -13392 -4876 -13380
rect -5074 -13608 -5068 -13392
rect -5034 -13420 -4916 -13392
rect -5034 -13580 -5028 -13420
rect -4922 -13580 -4916 -13420
rect -5034 -13608 -4916 -13580
rect -4882 -13608 -4876 -13392
rect -5074 -13620 -4876 -13608
rect -4824 -13392 -4626 -13380
rect -4824 -13608 -4818 -13392
rect -4784 -13420 -4666 -13392
rect -4784 -13580 -4778 -13420
rect -4672 -13580 -4666 -13420
rect -4784 -13608 -4666 -13580
rect -4632 -13608 -4626 -13392
rect -4824 -13620 -4626 -13608
rect -4574 -13392 -4376 -13380
rect -4574 -13608 -4568 -13392
rect -4534 -13420 -4416 -13392
rect -4534 -13580 -4528 -13420
rect -4422 -13580 -4416 -13420
rect -4534 -13608 -4416 -13580
rect -4382 -13608 -4376 -13392
rect -4574 -13620 -4376 -13608
rect -4324 -13392 -4126 -13380
rect -4324 -13608 -4318 -13392
rect -4284 -13420 -4166 -13392
rect -4284 -13580 -4278 -13420
rect -4172 -13580 -4166 -13420
rect -4284 -13608 -4166 -13580
rect -4132 -13608 -4126 -13392
rect -4324 -13620 -4126 -13608
rect -5824 -13652 -5778 -13620
rect -5922 -13658 -5778 -13652
rect -5922 -13692 -5867 -13658
rect -5833 -13692 -5778 -13658
rect -5922 -13708 -5778 -13692
rect -6087 -13798 -6077 -13745
rect -6024 -13798 -6014 -13745
rect -5720 -13957 -5686 -13620
rect -5633 -13658 -5567 -13652
rect -5633 -13692 -5617 -13658
rect -5583 -13692 -5567 -13658
rect -5633 -13708 -5567 -13692
rect -5383 -13658 -5317 -13652
rect -5383 -13692 -5367 -13658
rect -5333 -13692 -5317 -13658
rect -5383 -13708 -5317 -13692
rect -5617 -13852 -5583 -13708
rect -5367 -13745 -5333 -13708
rect -5386 -13798 -5376 -13745
rect -5323 -13798 -5313 -13745
rect -5636 -13905 -5626 -13852
rect -5573 -13905 -5563 -13852
rect -5740 -14010 -5730 -13957
rect -5677 -14010 -5667 -13957
rect -5240 -14055 -5206 -13620
rect -5133 -13658 -5067 -13652
rect -5133 -13692 -5117 -13658
rect -5083 -13692 -5067 -13658
rect -5133 -13708 -5067 -13692
rect -4883 -13658 -4817 -13652
rect -4883 -13692 -4867 -13658
rect -4833 -13692 -4817 -13658
rect -4883 -13708 -4817 -13692
rect -5117 -13745 -5083 -13708
rect -5136 -13798 -5126 -13745
rect -5073 -13798 -5063 -13745
rect -4867 -13852 -4833 -13708
rect -4887 -13905 -4877 -13852
rect -4824 -13905 -4814 -13852
rect -4742 -13957 -4708 -13620
rect -4633 -13658 -4567 -13652
rect -4633 -13692 -4617 -13658
rect -4583 -13692 -4567 -13658
rect -4633 -13708 -4567 -13692
rect -4383 -13658 -4317 -13652
rect -4383 -13692 -4367 -13658
rect -4333 -13692 -4317 -13658
rect -4383 -13708 -4317 -13692
rect -4617 -13852 -4583 -13708
rect -4367 -13745 -4333 -13708
rect -4386 -13798 -4376 -13745
rect -4323 -13798 -4313 -13745
rect -4637 -13905 -4627 -13852
rect -4574 -13905 -4564 -13852
rect -4762 -14010 -4752 -13957
rect -4699 -14010 -4689 -13957
rect -4240 -14055 -4206 -13620
rect -4172 -13652 -4126 -13620
rect -4074 -13392 -4028 -13380
rect -4074 -13608 -4068 -13392
rect -4034 -13608 -4028 -13392
rect -4074 -13652 -4028 -13608
rect -4172 -13658 -4028 -13652
rect -4172 -13692 -4117 -13658
rect -4083 -13692 -4028 -13658
rect -4172 -13708 -4028 -13692
rect -3928 -13852 -3875 -12442
rect -3798 -13242 -3788 -13189
rect -3735 -13242 -3725 -13189
rect -3938 -13905 -3928 -13852
rect -3875 -13905 -3865 -13852
rect -3928 -13906 -3875 -13905
rect -3788 -13957 -3735 -13242
rect -3798 -14010 -3788 -13957
rect -3735 -14010 -3725 -13957
rect -6233 -14108 -6223 -14055
rect -6170 -14108 -6160 -14055
rect -5260 -14108 -5250 -14055
rect -5197 -14108 -5187 -14055
rect -4260 -14108 -4250 -14055
rect -4197 -14108 -4187 -14055
rect -6965 -14260 -4303 -14226
rect -6028 -14382 -5994 -14260
rect -5939 -14294 -5905 -14260
rect -5960 -14310 -5884 -14294
rect -5960 -14344 -5944 -14310
rect -5900 -14344 -5884 -14310
rect -5960 -14350 -5884 -14344
rect -5850 -14382 -5816 -14260
rect -5761 -14294 -5727 -14260
rect -5583 -14294 -5549 -14260
rect -5405 -14294 -5371 -14260
rect -5227 -14294 -5193 -14260
rect -5049 -14294 -5015 -14260
rect -4871 -14294 -4837 -14260
rect -4693 -14294 -4659 -14260
rect -4515 -14294 -4481 -14260
rect -4337 -14294 -4303 -14260
rect -4248 -14260 -4036 -14226
rect -5782 -14310 -5706 -14294
rect -5782 -14344 -5766 -14310
rect -5722 -14344 -5706 -14310
rect -5782 -14350 -5706 -14344
rect -5604 -14310 -5528 -14294
rect -5604 -14344 -5588 -14310
rect -5544 -14344 -5528 -14310
rect -5604 -14350 -5528 -14344
rect -5426 -14310 -5350 -14294
rect -5426 -14344 -5410 -14310
rect -5366 -14344 -5350 -14310
rect -5426 -14350 -5350 -14344
rect -5248 -14310 -5172 -14294
rect -5248 -14344 -5232 -14310
rect -5188 -14344 -5172 -14310
rect -5248 -14350 -5172 -14344
rect -5070 -14310 -4994 -14294
rect -5070 -14344 -5054 -14310
rect -5010 -14344 -4994 -14310
rect -5070 -14350 -4994 -14344
rect -4892 -14310 -4816 -14294
rect -4892 -14344 -4876 -14310
rect -4832 -14344 -4816 -14310
rect -4892 -14350 -4816 -14344
rect -4714 -14310 -4638 -14294
rect -4714 -14344 -4698 -14310
rect -4654 -14344 -4638 -14310
rect -4714 -14350 -4638 -14344
rect -4536 -14310 -4460 -14294
rect -4536 -14344 -4520 -14310
rect -4476 -14344 -4460 -14310
rect -4536 -14350 -4460 -14344
rect -4358 -14310 -4282 -14294
rect -4358 -14344 -4342 -14310
rect -4298 -14344 -4282 -14310
rect -4358 -14350 -4282 -14344
rect -4248 -14382 -4214 -14260
rect -4159 -14294 -4125 -14260
rect -4180 -14310 -4104 -14294
rect -4180 -14344 -4164 -14310
rect -4120 -14344 -4104 -14310
rect -4180 -14350 -4104 -14344
rect -4070 -14382 -4036 -14260
rect -6034 -14394 -5988 -14382
rect -6034 -14650 -6028 -14394
rect -5994 -14650 -5988 -14394
rect -6034 -14662 -5988 -14650
rect -5856 -14394 -5810 -14382
rect -5856 -14650 -5850 -14394
rect -5816 -14650 -5810 -14394
rect -5856 -14662 -5810 -14650
rect -5678 -14394 -5632 -14382
rect -5678 -14650 -5672 -14394
rect -5638 -14650 -5632 -14394
rect -5678 -14662 -5632 -14650
rect -5500 -14394 -5454 -14382
rect -5500 -14650 -5494 -14394
rect -5460 -14650 -5454 -14394
rect -5500 -14662 -5454 -14650
rect -5322 -14394 -5276 -14382
rect -5322 -14650 -5316 -14394
rect -5282 -14650 -5276 -14394
rect -5322 -14662 -5276 -14650
rect -5144 -14394 -5098 -14382
rect -5144 -14650 -5138 -14394
rect -5104 -14650 -5098 -14394
rect -5144 -14662 -5098 -14650
rect -4966 -14394 -4920 -14382
rect -4966 -14650 -4960 -14394
rect -4926 -14650 -4920 -14394
rect -4966 -14662 -4920 -14650
rect -4788 -14394 -4742 -14382
rect -4788 -14650 -4782 -14394
rect -4748 -14650 -4742 -14394
rect -4788 -14662 -4742 -14650
rect -4610 -14394 -4564 -14382
rect -4610 -14650 -4604 -14394
rect -4570 -14650 -4564 -14394
rect -4610 -14662 -4564 -14650
rect -4432 -14394 -4386 -14382
rect -4432 -14650 -4426 -14394
rect -4392 -14650 -4386 -14394
rect -4432 -14662 -4386 -14650
rect -4254 -14394 -4208 -14382
rect -4254 -14650 -4248 -14394
rect -4214 -14650 -4208 -14394
rect -4254 -14662 -4208 -14650
rect -4076 -14394 -4030 -14382
rect -4076 -14650 -4070 -14394
rect -4036 -14650 -4030 -14394
rect -4076 -14662 -4030 -14650
rect -5960 -14700 -5884 -14694
rect -5960 -14734 -5944 -14700
rect -5900 -14734 -5884 -14700
rect -5960 -14750 -5884 -14734
rect -5850 -14795 -5816 -14662
rect -5782 -14700 -5706 -14694
rect -5782 -14734 -5766 -14700
rect -5722 -14734 -5706 -14700
rect -5782 -14750 -5706 -14734
rect -6169 -14848 -6159 -14795
rect -6106 -14848 -6096 -14795
rect -5870 -14848 -5860 -14795
rect -5807 -14848 -5797 -14795
rect -6159 -15482 -6106 -14848
rect -6028 -14959 -5816 -14925
rect -6027 -15082 -5993 -14959
rect -5939 -14994 -5905 -14959
rect -5960 -15010 -5884 -14994
rect -5960 -15044 -5944 -15010
rect -5900 -15044 -5884 -15010
rect -5960 -15050 -5884 -15044
rect -5850 -15082 -5816 -14959
rect -5761 -14994 -5727 -14750
rect -5782 -15010 -5706 -14994
rect -5782 -15044 -5766 -15010
rect -5722 -15044 -5706 -15010
rect -5782 -15050 -5706 -15044
rect -5672 -15082 -5638 -14662
rect -5604 -14700 -5528 -14694
rect -5604 -14734 -5588 -14700
rect -5544 -14734 -5528 -14700
rect -5604 -14750 -5528 -14734
rect -5583 -14994 -5549 -14750
rect -5494 -14901 -5460 -14662
rect -5426 -14700 -5350 -14694
rect -5426 -14734 -5410 -14700
rect -5366 -14734 -5350 -14700
rect -5426 -14750 -5350 -14734
rect -5514 -14954 -5504 -14901
rect -5451 -14954 -5441 -14901
rect -5405 -14994 -5371 -14750
rect -5604 -15010 -5528 -14994
rect -5604 -15044 -5588 -15010
rect -5544 -15044 -5528 -15010
rect -5604 -15050 -5528 -15044
rect -5426 -15010 -5350 -14994
rect -5426 -15044 -5410 -15010
rect -5366 -15044 -5350 -15010
rect -5426 -15050 -5350 -15044
rect -5316 -15082 -5282 -14662
rect -5248 -14700 -5172 -14694
rect -5248 -14734 -5232 -14700
rect -5188 -14734 -5172 -14700
rect -5248 -14750 -5172 -14734
rect -5227 -14994 -5193 -14750
rect -5138 -14795 -5104 -14662
rect -5070 -14700 -4994 -14694
rect -5070 -14734 -5054 -14700
rect -5010 -14734 -4994 -14700
rect -5070 -14750 -4994 -14734
rect -5157 -14848 -5147 -14795
rect -5094 -14848 -5084 -14795
rect -5049 -14994 -5015 -14750
rect -5248 -15010 -5172 -14994
rect -5248 -15044 -5232 -15010
rect -5188 -15044 -5172 -15010
rect -5248 -15050 -5172 -15044
rect -5070 -15010 -4994 -14994
rect -5070 -15044 -5054 -15010
rect -5010 -15044 -4994 -15010
rect -5070 -15050 -4994 -15044
rect -4960 -15082 -4926 -14662
rect -4892 -14700 -4816 -14694
rect -4892 -14734 -4876 -14700
rect -4832 -14734 -4816 -14700
rect -4892 -14750 -4816 -14734
rect -4871 -14994 -4837 -14750
rect -4782 -14901 -4748 -14662
rect -4714 -14700 -4638 -14694
rect -4714 -14734 -4698 -14700
rect -4654 -14734 -4638 -14700
rect -4714 -14750 -4638 -14734
rect -4801 -14954 -4791 -14901
rect -4738 -14954 -4728 -14901
rect -4693 -14994 -4659 -14750
rect -4892 -15010 -4816 -14994
rect -4892 -15044 -4876 -15010
rect -4832 -15044 -4816 -15010
rect -4892 -15050 -4816 -15044
rect -4714 -15010 -4638 -14994
rect -4714 -15044 -4698 -15010
rect -4654 -15044 -4638 -15010
rect -4714 -15050 -4638 -15044
rect -4604 -15082 -4570 -14662
rect -4536 -14700 -4460 -14694
rect -4536 -14734 -4520 -14700
rect -4476 -14734 -4460 -14700
rect -4536 -14750 -4460 -14734
rect -4515 -14994 -4481 -14750
rect -4426 -14795 -4392 -14662
rect -4358 -14700 -4282 -14694
rect -4358 -14734 -4342 -14700
rect -4298 -14734 -4282 -14700
rect -4358 -14750 -4282 -14734
rect -4446 -14848 -4436 -14795
rect -4383 -14848 -4373 -14795
rect -4337 -14994 -4303 -14750
rect -4248 -14925 -4214 -14662
rect -4180 -14700 -4104 -14694
rect -4180 -14734 -4164 -14700
rect -4120 -14734 -4104 -14700
rect -4180 -14750 -4104 -14734
rect -3664 -14901 -3611 -12153
rect -3541 -13137 -3489 -7840
rect 4761 -7907 4771 -7854
rect 4824 -7907 4834 -7854
rect 4896 -7905 4906 -7852
rect 4959 -7905 4969 -7852
rect 5027 -7903 5037 -7850
rect 5090 -7903 5100 -7850
rect -3392 -7986 -3382 -7933
rect -3329 -7986 -3319 -7933
rect -1392 -7975 -1382 -7922
rect -1329 -7975 -1319 -7922
rect -3542 -13189 -3489 -13137
rect -3552 -13242 -3542 -13189
rect -3489 -13242 -3479 -13189
rect -3382 -14055 -3329 -7986
rect -1372 -8032 -1338 -7975
rect -1213 -7976 -1203 -7923
rect -1150 -7976 -1140 -7923
rect -1035 -7975 -1025 -7922
rect -972 -7975 -962 -7922
rect -858 -7975 -848 -7922
rect -795 -7975 -785 -7922
rect -680 -7975 -670 -7922
rect -617 -7975 -607 -7922
rect -500 -7975 -490 -7922
rect -437 -7975 -427 -7922
rect 745 -7975 755 -7922
rect 808 -7975 818 -7922
rect 922 -7975 932 -7922
rect 985 -7975 995 -7922
rect 1102 -7975 1112 -7922
rect 1165 -7975 1175 -7922
rect -1194 -8032 -1160 -7976
rect -1016 -8032 -982 -7975
rect -838 -8032 -804 -7975
rect -660 -8032 -626 -7975
rect -481 -8032 -447 -7975
rect 765 -8032 799 -7975
rect 942 -8032 976 -7975
rect 1121 -8032 1155 -7975
rect 1279 -7976 1289 -7923
rect 1342 -7976 1352 -7923
rect 1457 -7975 1467 -7922
rect 1520 -7975 1530 -7922
rect 1634 -7975 1644 -7922
rect 1697 -7975 1707 -7922
rect 2880 -7975 2890 -7922
rect 2943 -7975 2953 -7922
rect 3059 -7975 3069 -7922
rect 3122 -7975 3132 -7922
rect 3237 -7975 3247 -7922
rect 3300 -7975 3310 -7922
rect 3414 -7975 3424 -7922
rect 3477 -7975 3487 -7922
rect 1298 -8032 1332 -7976
rect 1476 -8032 1510 -7975
rect 1654 -8032 1688 -7975
rect 2900 -8032 2934 -7975
rect 3078 -8032 3112 -7975
rect 3256 -8032 3290 -7975
rect 3434 -8032 3468 -7975
rect 3593 -7976 3603 -7923
rect 3656 -7976 3666 -7923
rect 3768 -7975 3778 -7922
rect 3831 -7975 3841 -7922
rect 3612 -8032 3646 -7976
rect 3790 -8032 3824 -7975
rect 4198 -7976 4208 -7923
rect 4261 -7976 4271 -7923
rect -2105 -8048 -2029 -8032
rect -2105 -8082 -2089 -8048
rect -2045 -8082 -2029 -8048
rect -2105 -8088 -2029 -8082
rect -1927 -8048 -1851 -8032
rect -1927 -8082 -1911 -8048
rect -1867 -8082 -1851 -8048
rect -1927 -8088 -1851 -8082
rect -1749 -8048 -1673 -8032
rect -1749 -8082 -1733 -8048
rect -1689 -8082 -1673 -8048
rect -1749 -8088 -1673 -8082
rect -1571 -8048 -1495 -8032
rect -1571 -8082 -1555 -8048
rect -1511 -8082 -1495 -8048
rect -1571 -8088 -1495 -8082
rect -1393 -8048 -1317 -8032
rect -1393 -8082 -1377 -8048
rect -1333 -8082 -1317 -8048
rect -1393 -8088 -1317 -8082
rect -1215 -8048 -1139 -8032
rect -1215 -8082 -1199 -8048
rect -1155 -8082 -1139 -8048
rect -1215 -8088 -1139 -8082
rect -1037 -8048 -961 -8032
rect -1037 -8082 -1021 -8048
rect -977 -8082 -961 -8048
rect -1037 -8088 -961 -8082
rect -859 -8048 -783 -8032
rect -859 -8082 -843 -8048
rect -799 -8082 -783 -8048
rect -859 -8088 -783 -8082
rect -681 -8048 -605 -8032
rect -681 -8082 -665 -8048
rect -621 -8082 -605 -8048
rect -681 -8088 -605 -8082
rect -503 -8048 -427 -8032
rect -503 -8082 -487 -8048
rect -443 -8082 -427 -8048
rect -503 -8088 -427 -8082
rect -325 -8048 -249 -8032
rect -325 -8082 -309 -8048
rect -265 -8082 -249 -8048
rect -325 -8088 -249 -8082
rect -147 -8048 -71 -8032
rect -147 -8082 -131 -8048
rect -87 -8082 -71 -8048
rect -147 -8088 -71 -8082
rect 31 -8048 107 -8032
rect 31 -8082 47 -8048
rect 91 -8082 107 -8048
rect 31 -8088 107 -8082
rect 209 -8048 285 -8032
rect 209 -8082 225 -8048
rect 269 -8082 285 -8048
rect 209 -8088 285 -8082
rect 387 -8048 463 -8032
rect 387 -8082 403 -8048
rect 447 -8082 463 -8048
rect 387 -8088 463 -8082
rect 565 -8048 641 -8032
rect 565 -8082 581 -8048
rect 625 -8082 641 -8048
rect 565 -8088 641 -8082
rect 743 -8048 819 -8032
rect 743 -8082 759 -8048
rect 803 -8082 819 -8048
rect 743 -8088 819 -8082
rect 921 -8048 997 -8032
rect 921 -8082 937 -8048
rect 981 -8082 997 -8048
rect 921 -8088 997 -8082
rect 1099 -8048 1175 -8032
rect 1099 -8082 1115 -8048
rect 1159 -8082 1175 -8048
rect 1099 -8088 1175 -8082
rect 1277 -8048 1353 -8032
rect 1277 -8082 1293 -8048
rect 1337 -8082 1353 -8048
rect 1277 -8088 1353 -8082
rect 1455 -8048 1531 -8032
rect 1455 -8082 1471 -8048
rect 1515 -8082 1531 -8048
rect 1455 -8088 1531 -8082
rect 1633 -8048 1709 -8032
rect 1633 -8082 1649 -8048
rect 1693 -8082 1709 -8048
rect 1633 -8088 1709 -8082
rect 1811 -8048 1887 -8032
rect 1811 -8082 1827 -8048
rect 1871 -8082 1887 -8048
rect 1811 -8088 1887 -8082
rect 1989 -8048 2065 -8032
rect 1989 -8082 2005 -8048
rect 2049 -8082 2065 -8048
rect 1989 -8088 2065 -8082
rect 2167 -8048 2243 -8032
rect 2167 -8082 2183 -8048
rect 2227 -8082 2243 -8048
rect 2167 -8088 2243 -8082
rect 2345 -8048 2421 -8032
rect 2345 -8082 2361 -8048
rect 2405 -8082 2421 -8048
rect 2345 -8088 2421 -8082
rect 2523 -8048 2599 -8032
rect 2523 -8082 2539 -8048
rect 2583 -8082 2599 -8048
rect 2523 -8088 2599 -8082
rect 2701 -8048 2777 -8032
rect 2701 -8082 2717 -8048
rect 2761 -8082 2777 -8048
rect 2701 -8088 2777 -8082
rect 2879 -8048 2955 -8032
rect 2879 -8082 2895 -8048
rect 2939 -8082 2955 -8048
rect 2879 -8088 2955 -8082
rect 3057 -8048 3133 -8032
rect 3057 -8082 3073 -8048
rect 3117 -8082 3133 -8048
rect 3057 -8088 3133 -8082
rect 3235 -8048 3311 -8032
rect 3235 -8082 3251 -8048
rect 3295 -8082 3311 -8048
rect 3235 -8088 3311 -8082
rect 3413 -8048 3489 -8032
rect 3413 -8082 3429 -8048
rect 3473 -8082 3489 -8048
rect 3413 -8088 3489 -8082
rect 3591 -8048 3667 -8032
rect 3591 -8082 3607 -8048
rect 3651 -8082 3667 -8048
rect 3591 -8088 3667 -8082
rect 3769 -8048 3845 -8032
rect 3769 -8082 3785 -8048
rect 3829 -8082 3845 -8048
rect 3769 -8088 3845 -8082
rect 3947 -8048 4023 -8032
rect 3947 -8082 3963 -8048
rect 4007 -8082 4023 -8048
rect 3947 -8088 4023 -8082
rect -2179 -8132 -2133 -8120
rect -2179 -8388 -2173 -8132
rect -2139 -8388 -2133 -8132
rect -2179 -8400 -2133 -8388
rect -2001 -8132 -1955 -8120
rect -2001 -8388 -1995 -8132
rect -1961 -8388 -1955 -8132
rect -2001 -8400 -1955 -8388
rect -1823 -8132 -1777 -8120
rect -1823 -8388 -1817 -8132
rect -1783 -8388 -1777 -8132
rect -1823 -8400 -1777 -8388
rect -1645 -8132 -1599 -8120
rect -1645 -8388 -1639 -8132
rect -1605 -8388 -1599 -8132
rect -1645 -8400 -1599 -8388
rect -1467 -8132 -1421 -8120
rect -1467 -8388 -1461 -8132
rect -1427 -8388 -1421 -8132
rect -1467 -8400 -1421 -8388
rect -1289 -8132 -1243 -8120
rect -1289 -8388 -1283 -8132
rect -1249 -8388 -1243 -8132
rect -1289 -8400 -1243 -8388
rect -1111 -8132 -1065 -8120
rect -1111 -8388 -1105 -8132
rect -1071 -8388 -1065 -8132
rect -1111 -8400 -1065 -8388
rect -933 -8132 -887 -8120
rect -933 -8388 -927 -8132
rect -893 -8388 -887 -8132
rect -933 -8400 -887 -8388
rect -755 -8132 -709 -8120
rect -755 -8388 -749 -8132
rect -715 -8388 -709 -8132
rect -755 -8400 -709 -8388
rect -577 -8132 -531 -8120
rect -577 -8388 -571 -8132
rect -537 -8388 -531 -8132
rect -577 -8400 -531 -8388
rect -399 -8132 -353 -8120
rect -399 -8388 -393 -8132
rect -359 -8388 -353 -8132
rect -399 -8400 -353 -8388
rect -221 -8132 -175 -8120
rect -221 -8388 -215 -8132
rect -181 -8388 -175 -8132
rect -221 -8400 -175 -8388
rect -43 -8132 3 -8120
rect -43 -8388 -37 -8132
rect -3 -8388 3 -8132
rect -43 -8400 3 -8388
rect 135 -8132 181 -8120
rect 135 -8388 141 -8132
rect 175 -8388 181 -8132
rect 135 -8400 181 -8388
rect 313 -8132 359 -8120
rect 313 -8388 319 -8132
rect 353 -8388 359 -8132
rect 313 -8400 359 -8388
rect 491 -8132 537 -8120
rect 491 -8388 497 -8132
rect 531 -8388 537 -8132
rect 491 -8400 537 -8388
rect 669 -8132 715 -8120
rect 669 -8388 675 -8132
rect 709 -8388 715 -8132
rect 669 -8400 715 -8388
rect 847 -8132 893 -8120
rect 847 -8388 853 -8132
rect 887 -8388 893 -8132
rect 847 -8400 893 -8388
rect 1025 -8132 1071 -8120
rect 1025 -8388 1031 -8132
rect 1065 -8388 1071 -8132
rect 1025 -8400 1071 -8388
rect 1203 -8132 1249 -8120
rect 1203 -8388 1209 -8132
rect 1243 -8388 1249 -8132
rect 1203 -8400 1249 -8388
rect 1381 -8132 1427 -8120
rect 1381 -8388 1387 -8132
rect 1421 -8388 1427 -8132
rect 1381 -8400 1427 -8388
rect 1559 -8132 1605 -8120
rect 1559 -8388 1565 -8132
rect 1599 -8388 1605 -8132
rect 1559 -8400 1605 -8388
rect 1737 -8132 1783 -8120
rect 1737 -8388 1743 -8132
rect 1777 -8388 1783 -8132
rect 1737 -8400 1783 -8388
rect 1915 -8132 1961 -8120
rect 1915 -8388 1921 -8132
rect 1955 -8388 1961 -8132
rect 1915 -8400 1961 -8388
rect 2093 -8132 2139 -8120
rect 2093 -8388 2099 -8132
rect 2133 -8388 2139 -8132
rect 2093 -8400 2139 -8388
rect 2271 -8132 2317 -8120
rect 2271 -8388 2277 -8132
rect 2311 -8388 2317 -8132
rect 2271 -8400 2317 -8388
rect 2449 -8132 2495 -8120
rect 2449 -8388 2455 -8132
rect 2489 -8388 2495 -8132
rect 2449 -8400 2495 -8388
rect 2627 -8132 2673 -8120
rect 2627 -8388 2633 -8132
rect 2667 -8388 2673 -8132
rect 2627 -8400 2673 -8388
rect 2805 -8132 2851 -8120
rect 2805 -8388 2811 -8132
rect 2845 -8388 2851 -8132
rect 2805 -8400 2851 -8388
rect 2983 -8132 3029 -8120
rect 2983 -8388 2989 -8132
rect 3023 -8388 3029 -8132
rect 2983 -8400 3029 -8388
rect 3161 -8132 3207 -8120
rect 3161 -8388 3167 -8132
rect 3201 -8388 3207 -8132
rect 3161 -8400 3207 -8388
rect 3339 -8132 3385 -8120
rect 3339 -8388 3345 -8132
rect 3379 -8388 3385 -8132
rect 3339 -8400 3385 -8388
rect 3517 -8132 3563 -8120
rect 3517 -8388 3523 -8132
rect 3557 -8388 3563 -8132
rect 3517 -8400 3563 -8388
rect 3695 -8132 3741 -8120
rect 3695 -8388 3701 -8132
rect 3735 -8388 3741 -8132
rect 3695 -8400 3741 -8388
rect 3873 -8132 3919 -8120
rect 3873 -8388 3879 -8132
rect 3913 -8388 3919 -8132
rect 3873 -8400 3919 -8388
rect 4051 -8132 4097 -8120
rect 4051 -8388 4057 -8132
rect 4091 -8388 4097 -8132
rect 4051 -8400 4097 -8388
rect -2171 -8440 -2137 -8400
rect -2105 -8438 -2029 -8432
rect -2105 -8440 -2089 -8438
rect -2171 -8472 -2089 -8440
rect -2045 -8440 -2029 -8438
rect -1995 -8440 -1961 -8400
rect -2045 -8472 -1961 -8440
rect -2171 -8474 -1961 -8472
rect -2105 -8488 -2029 -8474
rect -1995 -8767 -1961 -8474
rect -1927 -8438 -1851 -8432
rect -1927 -8472 -1911 -8438
rect -1867 -8472 -1851 -8438
rect -1927 -8488 -1851 -8472
rect -1906 -8534 -1872 -8488
rect -1926 -8587 -1916 -8534
rect -1863 -8587 -1853 -8534
rect -1817 -8653 -1783 -8400
rect -1749 -8438 -1673 -8432
rect -1749 -8472 -1733 -8438
rect -1689 -8472 -1673 -8438
rect -1749 -8488 -1673 -8472
rect -1729 -8534 -1695 -8488
rect -1749 -8587 -1739 -8534
rect -1686 -8587 -1676 -8534
rect -1836 -8706 -1826 -8653
rect -1773 -8706 -1763 -8653
rect -2457 -8820 -2447 -8767
rect -2394 -8820 -2384 -8767
rect -2015 -8820 -2005 -8767
rect -1952 -8820 -1942 -8767
rect -2447 -12272 -2394 -8820
rect -2105 -9048 -2029 -9032
rect -2105 -9082 -2089 -9048
rect -2045 -9082 -2029 -9048
rect -2105 -9088 -2029 -9082
rect -1995 -9120 -1961 -8820
rect -1927 -9048 -1851 -9032
rect -1927 -9082 -1911 -9048
rect -1867 -9082 -1851 -9048
rect -1927 -9088 -1851 -9082
rect -1817 -9120 -1783 -8706
rect -1639 -8767 -1605 -8400
rect -1571 -8438 -1495 -8432
rect -1571 -8472 -1555 -8438
rect -1511 -8472 -1495 -8438
rect -1571 -8488 -1495 -8472
rect -1549 -8534 -1515 -8488
rect -1568 -8587 -1558 -8534
rect -1505 -8587 -1495 -8534
rect -1461 -8653 -1427 -8400
rect -1393 -8438 -1317 -8432
rect -1393 -8472 -1377 -8438
rect -1333 -8472 -1317 -8438
rect -1393 -8488 -1317 -8472
rect -1392 -8587 -1382 -8534
rect -1329 -8587 -1319 -8534
rect -1480 -8706 -1470 -8653
rect -1417 -8706 -1407 -8653
rect -1658 -8820 -1648 -8767
rect -1595 -8820 -1585 -8767
rect -1749 -9048 -1673 -9032
rect -1749 -9082 -1733 -9048
rect -1689 -9082 -1673 -9048
rect -1749 -9088 -1673 -9082
rect -1639 -9120 -1605 -8820
rect -1571 -9048 -1495 -9032
rect -1571 -9082 -1555 -9048
rect -1511 -9082 -1495 -9048
rect -1571 -9088 -1495 -9082
rect -1461 -9120 -1427 -8706
rect -1372 -9032 -1338 -8587
rect -1283 -8767 -1249 -8400
rect -1215 -8438 -1139 -8432
rect -1215 -8472 -1199 -8438
rect -1155 -8472 -1139 -8438
rect -1215 -8488 -1139 -8472
rect -1213 -8587 -1203 -8534
rect -1150 -8587 -1140 -8534
rect -1303 -8820 -1293 -8767
rect -1240 -8820 -1230 -8767
rect -1393 -9048 -1317 -9032
rect -1393 -9082 -1377 -9048
rect -1333 -9082 -1317 -9048
rect -1393 -9088 -1317 -9082
rect -1283 -9120 -1249 -8820
rect -1193 -9032 -1159 -8587
rect -1105 -8653 -1071 -8400
rect -1037 -8438 -961 -8432
rect -1037 -8472 -1021 -8438
rect -977 -8472 -961 -8438
rect -1037 -8488 -961 -8472
rect -1036 -8587 -1026 -8534
rect -973 -8587 -963 -8534
rect -1125 -8706 -1115 -8653
rect -1062 -8706 -1052 -8653
rect -1215 -9048 -1139 -9032
rect -1215 -9082 -1199 -9048
rect -1155 -9082 -1139 -9048
rect -1215 -9088 -1139 -9082
rect -1105 -9120 -1071 -8706
rect -1016 -9032 -982 -8587
rect -927 -8767 -893 -8400
rect -859 -8438 -783 -8432
rect -859 -8472 -843 -8438
rect -799 -8472 -783 -8438
rect -859 -8488 -783 -8472
rect -858 -8587 -848 -8534
rect -795 -8587 -785 -8534
rect -946 -8820 -936 -8767
rect -883 -8820 -873 -8767
rect -1037 -9048 -961 -9032
rect -1037 -9082 -1021 -9048
rect -977 -9082 -961 -9048
rect -1037 -9088 -961 -9082
rect -927 -9120 -893 -8820
rect -838 -9032 -804 -8587
rect -749 -8653 -715 -8400
rect -681 -8438 -605 -8432
rect -681 -8472 -665 -8438
rect -621 -8472 -605 -8438
rect -681 -8488 -605 -8472
rect -680 -8587 -670 -8534
rect -617 -8587 -607 -8534
rect -768 -8706 -758 -8653
rect -705 -8706 -695 -8653
rect -859 -9048 -783 -9032
rect -859 -9082 -843 -9048
rect -799 -9082 -783 -9048
rect -859 -9088 -783 -9082
rect -749 -9120 -715 -8706
rect -660 -9032 -626 -8587
rect -571 -8766 -537 -8400
rect -503 -8438 -427 -8432
rect -503 -8472 -487 -8438
rect -443 -8472 -427 -8438
rect -503 -8488 -427 -8472
rect -501 -8587 -491 -8534
rect -438 -8587 -428 -8534
rect -590 -8819 -580 -8766
rect -527 -8819 -517 -8766
rect -681 -9048 -605 -9032
rect -681 -9082 -665 -9048
rect -621 -9082 -605 -9048
rect -681 -9088 -605 -9082
rect -571 -9120 -537 -8819
rect -482 -9032 -448 -8587
rect -393 -8653 -359 -8400
rect -325 -8438 -249 -8432
rect -325 -8472 -309 -8438
rect -265 -8472 -249 -8438
rect -325 -8488 -249 -8472
rect -304 -8534 -270 -8488
rect -324 -8587 -314 -8534
rect -261 -8587 -251 -8534
rect -412 -8706 -402 -8653
rect -349 -8706 -339 -8653
rect -503 -9048 -427 -9032
rect -503 -9082 -487 -9048
rect -443 -9082 -427 -9048
rect -503 -9088 -427 -9082
rect -393 -9120 -359 -8706
rect -215 -8767 -181 -8400
rect -147 -8438 -71 -8432
rect -147 -8472 -131 -8438
rect -87 -8472 -71 -8438
rect -147 -8488 -71 -8472
rect -126 -8534 -92 -8488
rect -146 -8587 -136 -8534
rect -83 -8587 -73 -8534
rect -37 -8653 -3 -8400
rect 31 -8438 107 -8432
rect 31 -8472 47 -8438
rect 91 -8472 107 -8438
rect 31 -8488 107 -8472
rect 52 -8534 86 -8488
rect 32 -8587 42 -8534
rect 95 -8587 105 -8534
rect -57 -8706 -47 -8653
rect 6 -8706 16 -8653
rect -235 -8820 -225 -8767
rect -172 -8820 -162 -8767
rect -325 -9048 -249 -9032
rect -325 -9082 -309 -9048
rect -265 -9082 -249 -9048
rect -325 -9088 -249 -9082
rect -215 -9120 -181 -8820
rect -147 -9048 -71 -9032
rect -147 -9082 -131 -9048
rect -87 -9082 -71 -9048
rect -147 -9088 -71 -9082
rect -37 -9120 -3 -8706
rect 141 -8768 175 -8400
rect 209 -8438 285 -8432
rect 209 -8472 225 -8438
rect 269 -8472 285 -8438
rect 209 -8488 285 -8472
rect 230 -8534 264 -8488
rect 211 -8587 221 -8534
rect 274 -8587 284 -8534
rect 319 -8653 353 -8400
rect 387 -8438 463 -8432
rect 387 -8472 403 -8438
rect 447 -8472 463 -8438
rect 387 -8488 463 -8472
rect 408 -8534 442 -8488
rect 388 -8587 398 -8534
rect 451 -8587 461 -8534
rect 300 -8706 310 -8653
rect 363 -8706 373 -8653
rect 122 -8821 132 -8768
rect 185 -8821 195 -8768
rect 31 -9048 107 -9032
rect 31 -9082 47 -9048
rect 91 -9082 107 -9048
rect 31 -9088 107 -9082
rect 141 -9120 175 -8821
rect 209 -9048 285 -9032
rect 209 -9082 225 -9048
rect 269 -9082 285 -9048
rect 209 -9088 285 -9082
rect 319 -9120 353 -8706
rect 497 -8766 531 -8400
rect 565 -8438 641 -8432
rect 565 -8472 581 -8438
rect 625 -8472 641 -8438
rect 565 -8488 641 -8472
rect 586 -8534 620 -8488
rect 567 -8587 577 -8534
rect 630 -8587 640 -8534
rect 675 -8653 709 -8400
rect 743 -8438 819 -8432
rect 743 -8472 759 -8438
rect 803 -8472 819 -8438
rect 743 -8488 819 -8472
rect 744 -8587 754 -8534
rect 807 -8587 817 -8534
rect 656 -8706 666 -8653
rect 719 -8706 729 -8653
rect 479 -8819 489 -8766
rect 542 -8819 552 -8766
rect 387 -9048 463 -9032
rect 387 -9082 403 -9048
rect 447 -9082 463 -9048
rect 387 -9088 463 -9082
rect 497 -9120 531 -8819
rect 565 -9048 641 -9032
rect 565 -9082 581 -9048
rect 625 -9082 641 -9048
rect 565 -9088 641 -9082
rect 675 -9120 709 -8706
rect 764 -9032 798 -8587
rect 853 -8766 887 -8400
rect 921 -8438 997 -8432
rect 921 -8472 937 -8438
rect 981 -8472 997 -8438
rect 921 -8488 997 -8472
rect 922 -8587 932 -8534
rect 985 -8587 995 -8534
rect 833 -8819 843 -8766
rect 896 -8819 906 -8766
rect 743 -9048 819 -9032
rect 743 -9082 759 -9048
rect 803 -9082 819 -9048
rect 743 -9088 819 -9082
rect 853 -9120 887 -8819
rect 942 -9032 976 -8587
rect 1031 -8653 1065 -8400
rect 1099 -8438 1175 -8432
rect 1099 -8472 1115 -8438
rect 1159 -8472 1175 -8438
rect 1099 -8488 1175 -8472
rect 1101 -8587 1111 -8534
rect 1164 -8587 1174 -8534
rect 1012 -8706 1022 -8653
rect 1075 -8706 1085 -8653
rect 921 -9048 997 -9032
rect 921 -9082 937 -9048
rect 981 -9082 997 -9048
rect 921 -9088 997 -9082
rect 1031 -9120 1065 -8706
rect 1120 -9032 1154 -8587
rect 1209 -8767 1243 -8400
rect 1277 -8438 1353 -8432
rect 1277 -8472 1293 -8438
rect 1337 -8472 1353 -8438
rect 1277 -8488 1353 -8472
rect 1279 -8587 1289 -8534
rect 1342 -8587 1352 -8534
rect 1191 -8820 1201 -8767
rect 1254 -8820 1264 -8767
rect 1099 -9048 1175 -9032
rect 1099 -9082 1115 -9048
rect 1159 -9082 1175 -9048
rect 1099 -9088 1175 -9082
rect 1209 -9120 1243 -8820
rect 1298 -9032 1332 -8587
rect 1387 -8653 1421 -8400
rect 1455 -8438 1531 -8432
rect 1455 -8472 1471 -8438
rect 1515 -8472 1531 -8438
rect 1455 -8488 1531 -8472
rect 1456 -8587 1466 -8534
rect 1519 -8587 1529 -8534
rect 1367 -8706 1377 -8653
rect 1430 -8706 1440 -8653
rect 1277 -9048 1353 -9032
rect 1277 -9082 1293 -9048
rect 1337 -9082 1353 -9048
rect 1277 -9088 1353 -9082
rect 1387 -9120 1421 -8706
rect 1476 -9032 1510 -8587
rect 1565 -8767 1599 -8400
rect 1633 -8438 1709 -8432
rect 1633 -8472 1649 -8438
rect 1693 -8472 1709 -8438
rect 1633 -8488 1709 -8472
rect 1634 -8587 1644 -8534
rect 1697 -8587 1707 -8534
rect 1546 -8820 1556 -8767
rect 1609 -8820 1619 -8767
rect 1455 -9048 1531 -9032
rect 1455 -9082 1471 -9048
rect 1515 -9082 1531 -9048
rect 1455 -9088 1531 -9082
rect 1565 -9120 1599 -8820
rect 1654 -9032 1688 -8587
rect 1743 -8653 1777 -8400
rect 1811 -8438 1887 -8432
rect 1811 -8472 1827 -8438
rect 1871 -8472 1887 -8438
rect 1811 -8488 1887 -8472
rect 1832 -8534 1866 -8488
rect 1812 -8587 1822 -8534
rect 1875 -8587 1885 -8534
rect 1723 -8706 1733 -8653
rect 1786 -8706 1796 -8653
rect 1633 -9048 1709 -9032
rect 1633 -9082 1649 -9048
rect 1693 -9082 1709 -9048
rect 1633 -9088 1709 -9082
rect 1743 -9120 1777 -8706
rect 1921 -8767 1955 -8400
rect 1989 -8438 2065 -8432
rect 1989 -8472 2005 -8438
rect 2049 -8472 2065 -8438
rect 1989 -8488 2065 -8472
rect 2010 -8534 2044 -8488
rect 1990 -8587 2000 -8534
rect 2053 -8587 2063 -8534
rect 2099 -8653 2133 -8400
rect 2167 -8438 2243 -8432
rect 2167 -8472 2183 -8438
rect 2227 -8472 2243 -8438
rect 2167 -8488 2243 -8472
rect 2188 -8534 2222 -8488
rect 2168 -8587 2178 -8534
rect 2231 -8587 2241 -8534
rect 2080 -8706 2090 -8653
rect 2143 -8706 2153 -8653
rect 1901 -8820 1911 -8767
rect 1964 -8820 1974 -8767
rect 1811 -9048 1887 -9032
rect 1811 -9082 1827 -9048
rect 1871 -9082 1887 -9048
rect 1811 -9088 1887 -9082
rect 1921 -9120 1955 -8820
rect 1989 -9048 2065 -9032
rect 1989 -9082 2005 -9048
rect 2049 -9082 2065 -9048
rect 1989 -9088 2065 -9082
rect 2099 -9120 2133 -8706
rect 2277 -8767 2311 -8400
rect 2345 -8438 2421 -8432
rect 2345 -8472 2361 -8438
rect 2405 -8472 2421 -8438
rect 2345 -8488 2421 -8472
rect 2367 -8534 2401 -8488
rect 2347 -8587 2357 -8534
rect 2410 -8587 2420 -8534
rect 2455 -8653 2489 -8400
rect 2523 -8438 2599 -8432
rect 2523 -8472 2539 -8438
rect 2583 -8472 2599 -8438
rect 2523 -8488 2599 -8472
rect 2544 -8534 2578 -8488
rect 2524 -8587 2534 -8534
rect 2587 -8587 2597 -8534
rect 2436 -8706 2446 -8653
rect 2499 -8706 2509 -8653
rect 2257 -8820 2267 -8767
rect 2320 -8820 2330 -8767
rect 2167 -9048 2243 -9032
rect 2167 -9082 2183 -9048
rect 2227 -9082 2243 -9048
rect 2167 -9088 2243 -9082
rect 2277 -9120 2311 -8820
rect 2345 -9048 2421 -9032
rect 2345 -9082 2361 -9048
rect 2405 -9082 2421 -9048
rect 2345 -9088 2421 -9082
rect 2455 -9120 2489 -8706
rect 2633 -8767 2667 -8400
rect 2701 -8438 2777 -8432
rect 2701 -8472 2717 -8438
rect 2761 -8472 2777 -8438
rect 2701 -8488 2777 -8472
rect 2722 -8534 2756 -8488
rect 2702 -8587 2712 -8534
rect 2765 -8587 2775 -8534
rect 2811 -8653 2845 -8400
rect 2879 -8438 2955 -8432
rect 2879 -8472 2895 -8438
rect 2939 -8472 2955 -8438
rect 2879 -8488 2955 -8472
rect 2880 -8587 2890 -8534
rect 2943 -8587 2953 -8534
rect 2792 -8706 2802 -8653
rect 2855 -8706 2865 -8653
rect 2614 -8820 2624 -8767
rect 2677 -8820 2687 -8767
rect 2523 -9048 2599 -9032
rect 2523 -9082 2539 -9048
rect 2583 -9082 2599 -9048
rect 2523 -9088 2599 -9082
rect 2633 -9120 2667 -8820
rect 2701 -9048 2777 -9032
rect 2701 -9082 2717 -9048
rect 2761 -9082 2777 -9048
rect 2701 -9088 2777 -9082
rect 2811 -9120 2845 -8706
rect 2900 -9032 2934 -8587
rect 2989 -8767 3023 -8400
rect 3057 -8438 3133 -8432
rect 3057 -8472 3073 -8438
rect 3117 -8472 3133 -8438
rect 3057 -8488 3133 -8472
rect 3058 -8587 3068 -8534
rect 3121 -8587 3131 -8534
rect 2970 -8820 2980 -8767
rect 3033 -8820 3043 -8767
rect 2879 -9048 2955 -9032
rect 2879 -9082 2895 -9048
rect 2939 -9082 2955 -9048
rect 2879 -9088 2955 -9082
rect 2989 -9120 3023 -8820
rect 3078 -9032 3112 -8587
rect 3167 -8653 3201 -8400
rect 3235 -8438 3311 -8432
rect 3235 -8472 3251 -8438
rect 3295 -8472 3311 -8438
rect 3235 -8488 3311 -8472
rect 3236 -8587 3246 -8534
rect 3299 -8587 3309 -8534
rect 3148 -8706 3158 -8653
rect 3211 -8706 3221 -8653
rect 3057 -9048 3133 -9032
rect 3057 -9082 3073 -9048
rect 3117 -9082 3133 -9048
rect 3057 -9088 3133 -9082
rect 3167 -9120 3201 -8706
rect 3256 -9032 3290 -8587
rect 3345 -8767 3379 -8400
rect 3413 -8438 3489 -8432
rect 3413 -8472 3429 -8438
rect 3473 -8472 3489 -8438
rect 3413 -8488 3489 -8472
rect 3414 -8587 3424 -8534
rect 3477 -8587 3487 -8534
rect 3326 -8820 3336 -8767
rect 3389 -8820 3399 -8767
rect 3235 -9048 3311 -9032
rect 3235 -9082 3251 -9048
rect 3295 -9082 3311 -9048
rect 3235 -9088 3311 -9082
rect 3345 -9120 3379 -8820
rect 3434 -9032 3468 -8587
rect 3523 -8653 3557 -8400
rect 3591 -8438 3667 -8432
rect 3591 -8472 3607 -8438
rect 3651 -8472 3667 -8438
rect 3591 -8488 3667 -8472
rect 3592 -8587 3602 -8534
rect 3655 -8587 3665 -8534
rect 3503 -8706 3513 -8653
rect 3566 -8706 3576 -8653
rect 3413 -9048 3489 -9032
rect 3413 -9082 3429 -9048
rect 3473 -9082 3489 -9048
rect 3413 -9088 3489 -9082
rect 3523 -9120 3557 -8706
rect 3612 -9032 3646 -8587
rect 3701 -8767 3735 -8400
rect 3769 -8438 3845 -8432
rect 3769 -8472 3785 -8438
rect 3829 -8472 3845 -8438
rect 3769 -8488 3845 -8472
rect 3879 -8440 3913 -8400
rect 3947 -8438 4023 -8432
rect 3947 -8440 3963 -8438
rect 3879 -8472 3963 -8440
rect 4007 -8440 4023 -8438
rect 4056 -8440 4090 -8400
rect 4007 -8472 4090 -8440
rect 3879 -8474 4090 -8472
rect 3771 -8587 3781 -8534
rect 3834 -8587 3844 -8534
rect 3682 -8820 3692 -8767
rect 3745 -8820 3755 -8767
rect 3591 -9048 3667 -9032
rect 3591 -9082 3607 -9048
rect 3651 -9082 3667 -9048
rect 3591 -9088 3667 -9082
rect 3701 -9120 3735 -8820
rect 3790 -9032 3824 -8587
rect 3879 -8653 3913 -8474
rect 3947 -8488 4023 -8474
rect 3859 -8706 3869 -8653
rect 3922 -8706 3932 -8653
rect 3769 -9048 3845 -9032
rect 3769 -9082 3785 -9048
rect 3829 -9082 3845 -9048
rect 3769 -9088 3845 -9082
rect 3879 -9120 3913 -8706
rect 3947 -9048 4023 -9032
rect 3947 -9082 3963 -9048
rect 4007 -9082 4023 -9048
rect 3947 -9088 4023 -9082
rect -2179 -9132 -2133 -9120
rect -2179 -9388 -2173 -9132
rect -2139 -9388 -2133 -9132
rect -2179 -9400 -2133 -9388
rect -2001 -9132 -1955 -9120
rect -2001 -9388 -1995 -9132
rect -1961 -9388 -1955 -9132
rect -2001 -9400 -1955 -9388
rect -1823 -9132 -1777 -9120
rect -1823 -9388 -1817 -9132
rect -1783 -9388 -1777 -9132
rect -1823 -9400 -1777 -9388
rect -1645 -9132 -1599 -9120
rect -1645 -9388 -1639 -9132
rect -1605 -9388 -1599 -9132
rect -1645 -9400 -1599 -9388
rect -1467 -9132 -1421 -9120
rect -1467 -9388 -1461 -9132
rect -1427 -9388 -1421 -9132
rect -1467 -9400 -1421 -9388
rect -1289 -9132 -1243 -9120
rect -1289 -9388 -1283 -9132
rect -1249 -9388 -1243 -9132
rect -1289 -9400 -1243 -9388
rect -1111 -9132 -1065 -9120
rect -1111 -9388 -1105 -9132
rect -1071 -9388 -1065 -9132
rect -1111 -9400 -1065 -9388
rect -933 -9132 -887 -9120
rect -933 -9388 -927 -9132
rect -893 -9388 -887 -9132
rect -933 -9400 -887 -9388
rect -755 -9132 -709 -9120
rect -755 -9388 -749 -9132
rect -715 -9388 -709 -9132
rect -755 -9400 -709 -9388
rect -577 -9132 -531 -9120
rect -577 -9388 -571 -9132
rect -537 -9388 -531 -9132
rect -577 -9400 -531 -9388
rect -399 -9132 -353 -9120
rect -399 -9388 -393 -9132
rect -359 -9388 -353 -9132
rect -399 -9400 -353 -9388
rect -221 -9132 -175 -9120
rect -221 -9388 -215 -9132
rect -181 -9388 -175 -9132
rect -221 -9400 -175 -9388
rect -43 -9132 3 -9120
rect -43 -9388 -37 -9132
rect -3 -9388 3 -9132
rect -43 -9400 3 -9388
rect 135 -9132 181 -9120
rect 135 -9388 141 -9132
rect 175 -9388 181 -9132
rect 135 -9400 181 -9388
rect 313 -9132 359 -9120
rect 313 -9388 319 -9132
rect 353 -9388 359 -9132
rect 313 -9400 359 -9388
rect 491 -9132 537 -9120
rect 491 -9388 497 -9132
rect 531 -9388 537 -9132
rect 491 -9400 537 -9388
rect 669 -9132 715 -9120
rect 669 -9388 675 -9132
rect 709 -9388 715 -9132
rect 669 -9400 715 -9388
rect 847 -9132 893 -9120
rect 847 -9388 853 -9132
rect 887 -9388 893 -9132
rect 847 -9400 893 -9388
rect 1025 -9132 1071 -9120
rect 1025 -9388 1031 -9132
rect 1065 -9388 1071 -9132
rect 1025 -9400 1071 -9388
rect 1203 -9132 1249 -9120
rect 1203 -9388 1209 -9132
rect 1243 -9388 1249 -9132
rect 1203 -9400 1249 -9388
rect 1381 -9132 1427 -9120
rect 1381 -9388 1387 -9132
rect 1421 -9388 1427 -9132
rect 1381 -9400 1427 -9388
rect 1559 -9132 1605 -9120
rect 1559 -9388 1565 -9132
rect 1599 -9388 1605 -9132
rect 1559 -9400 1605 -9388
rect 1737 -9132 1783 -9120
rect 1737 -9388 1743 -9132
rect 1777 -9388 1783 -9132
rect 1737 -9400 1783 -9388
rect 1915 -9132 1961 -9120
rect 1915 -9388 1921 -9132
rect 1955 -9388 1961 -9132
rect 1915 -9400 1961 -9388
rect 2093 -9132 2139 -9120
rect 2093 -9388 2099 -9132
rect 2133 -9388 2139 -9132
rect 2093 -9400 2139 -9388
rect 2271 -9132 2317 -9120
rect 2271 -9388 2277 -9132
rect 2311 -9388 2317 -9132
rect 2271 -9400 2317 -9388
rect 2449 -9132 2495 -9120
rect 2449 -9388 2455 -9132
rect 2489 -9388 2495 -9132
rect 2449 -9400 2495 -9388
rect 2627 -9132 2673 -9120
rect 2627 -9388 2633 -9132
rect 2667 -9388 2673 -9132
rect 2627 -9400 2673 -9388
rect 2805 -9132 2851 -9120
rect 2805 -9388 2811 -9132
rect 2845 -9388 2851 -9132
rect 2805 -9400 2851 -9388
rect 2983 -9132 3029 -9120
rect 2983 -9388 2989 -9132
rect 3023 -9388 3029 -9132
rect 2983 -9400 3029 -9388
rect 3161 -9132 3207 -9120
rect 3161 -9388 3167 -9132
rect 3201 -9388 3207 -9132
rect 3161 -9400 3207 -9388
rect 3339 -9132 3385 -9120
rect 3339 -9388 3345 -9132
rect 3379 -9388 3385 -9132
rect 3339 -9400 3385 -9388
rect 3517 -9132 3563 -9120
rect 3517 -9388 3523 -9132
rect 3557 -9388 3563 -9132
rect 3517 -9400 3563 -9388
rect 3695 -9132 3741 -9120
rect 3695 -9388 3701 -9132
rect 3735 -9388 3741 -9132
rect 3695 -9400 3741 -9388
rect 3873 -9132 3919 -9120
rect 3873 -9388 3879 -9132
rect 3913 -9388 3919 -9132
rect 3873 -9400 3919 -9388
rect 4051 -9132 4097 -9120
rect 4051 -9388 4057 -9132
rect 4091 -9388 4097 -9132
rect 4051 -9400 4097 -9388
rect -2174 -9439 -2140 -9400
rect -2105 -9438 -2029 -9432
rect -2105 -9439 -2089 -9438
rect -2174 -9472 -2089 -9439
rect -2045 -9439 -2029 -9438
rect -1995 -9439 -1961 -9400
rect -2045 -9472 -1961 -9439
rect -2174 -9473 -1961 -9472
rect -2105 -9488 -2029 -9473
rect -2325 -9978 -2315 -9925
rect -2262 -9978 -2252 -9925
rect -2457 -12325 -2447 -12272
rect -2394 -12325 -2384 -12272
rect -3392 -14108 -3382 -14055
rect -3329 -14108 -3319 -14055
rect -4248 -14959 -4036 -14925
rect -3946 -14954 -3936 -14901
rect -3883 -14954 -3611 -14901
rect -4536 -15010 -4460 -14994
rect -4536 -15044 -4520 -15010
rect -4476 -15044 -4460 -15010
rect -4536 -15050 -4460 -15044
rect -4358 -15010 -4282 -14994
rect -4358 -15044 -4342 -15010
rect -4298 -15044 -4282 -15010
rect -4358 -15050 -4282 -15044
rect -4248 -15082 -4214 -14959
rect -4159 -14994 -4125 -14959
rect -4180 -15010 -4104 -14994
rect -4180 -15044 -4164 -15010
rect -4120 -15044 -4104 -15010
rect -4180 -15050 -4104 -15044
rect -4070 -15082 -4036 -14959
rect -3936 -15006 -3883 -14954
rect -6034 -15094 -5988 -15082
rect -6034 -15350 -6028 -15094
rect -5994 -15350 -5988 -15094
rect -6034 -15362 -5988 -15350
rect -5856 -15094 -5810 -15082
rect -5856 -15350 -5850 -15094
rect -5816 -15350 -5810 -15094
rect -5856 -15362 -5810 -15350
rect -5678 -15094 -5632 -15082
rect -5678 -15350 -5672 -15094
rect -5638 -15350 -5632 -15094
rect -5678 -15362 -5632 -15350
rect -5500 -15094 -5454 -15082
rect -5500 -15350 -5494 -15094
rect -5460 -15350 -5454 -15094
rect -5500 -15362 -5454 -15350
rect -5322 -15094 -5276 -15082
rect -5322 -15350 -5316 -15094
rect -5282 -15350 -5276 -15094
rect -5322 -15362 -5276 -15350
rect -5144 -15094 -5098 -15082
rect -5144 -15350 -5138 -15094
rect -5104 -15350 -5098 -15094
rect -5144 -15362 -5098 -15350
rect -4966 -15094 -4920 -15082
rect -4966 -15350 -4960 -15094
rect -4926 -15350 -4920 -15094
rect -4966 -15362 -4920 -15350
rect -4788 -15094 -4742 -15082
rect -4788 -15350 -4782 -15094
rect -4748 -15350 -4742 -15094
rect -4788 -15362 -4742 -15350
rect -4610 -15094 -4564 -15082
rect -4610 -15350 -4604 -15094
rect -4570 -15350 -4564 -15094
rect -4610 -15362 -4564 -15350
rect -4432 -15094 -4386 -15082
rect -4432 -15350 -4426 -15094
rect -4392 -15350 -4386 -15094
rect -4432 -15362 -4386 -15350
rect -4254 -15094 -4208 -15082
rect -4254 -15350 -4248 -15094
rect -4214 -15350 -4208 -15094
rect -4254 -15362 -4208 -15350
rect -4076 -15094 -4030 -15082
rect -4076 -15350 -4070 -15094
rect -4036 -15350 -4030 -15094
rect -4076 -15362 -4030 -15350
rect -5960 -15400 -5884 -15394
rect -5960 -15434 -5944 -15400
rect -5900 -15434 -5884 -15400
rect -5960 -15450 -5884 -15434
rect -6169 -15535 -6159 -15482
rect -6106 -15535 -6096 -15482
rect -6159 -16193 -6106 -15535
rect -5850 -15588 -5816 -15362
rect -5782 -15400 -5706 -15394
rect -5782 -15434 -5766 -15400
rect -5722 -15434 -5706 -15400
rect -5782 -15450 -5706 -15434
rect -5870 -15641 -5860 -15588
rect -5807 -15641 -5797 -15588
rect -5761 -15694 -5727 -15450
rect -5960 -15710 -5884 -15694
rect -5960 -15744 -5944 -15710
rect -5900 -15744 -5884 -15710
rect -5960 -15750 -5884 -15744
rect -5782 -15710 -5706 -15694
rect -5782 -15744 -5766 -15710
rect -5722 -15744 -5706 -15710
rect -5782 -15750 -5706 -15744
rect -5672 -15782 -5638 -15362
rect -5604 -15400 -5528 -15394
rect -5604 -15434 -5588 -15400
rect -5544 -15434 -5528 -15400
rect -5604 -15450 -5528 -15434
rect -5583 -15694 -5549 -15450
rect -5494 -15481 -5460 -15362
rect -5426 -15400 -5350 -15394
rect -5426 -15434 -5410 -15400
rect -5366 -15434 -5350 -15400
rect -5426 -15450 -5350 -15434
rect -5514 -15534 -5504 -15481
rect -5451 -15534 -5441 -15481
rect -5405 -15694 -5371 -15450
rect -5604 -15710 -5528 -15694
rect -5604 -15744 -5588 -15710
rect -5544 -15744 -5528 -15710
rect -5604 -15750 -5528 -15744
rect -5426 -15710 -5350 -15694
rect -5426 -15744 -5410 -15710
rect -5366 -15744 -5350 -15710
rect -5426 -15750 -5350 -15744
rect -5316 -15782 -5282 -15362
rect -5248 -15400 -5172 -15394
rect -5248 -15434 -5232 -15400
rect -5188 -15434 -5172 -15400
rect -5248 -15450 -5172 -15434
rect -5227 -15694 -5193 -15450
rect -5138 -15589 -5104 -15362
rect -5070 -15400 -4994 -15394
rect -5070 -15434 -5054 -15400
rect -5010 -15434 -4994 -15400
rect -5070 -15450 -4994 -15434
rect -5158 -15642 -5148 -15589
rect -5095 -15642 -5085 -15589
rect -5049 -15694 -5015 -15450
rect -5248 -15710 -5172 -15694
rect -5248 -15744 -5232 -15710
rect -5188 -15744 -5172 -15710
rect -5248 -15750 -5172 -15744
rect -5070 -15710 -4994 -15694
rect -5070 -15744 -5054 -15710
rect -5010 -15744 -4994 -15710
rect -5070 -15750 -4994 -15744
rect -4960 -15782 -4926 -15362
rect -4892 -15400 -4816 -15394
rect -4892 -15434 -4876 -15400
rect -4832 -15434 -4816 -15400
rect -4892 -15450 -4816 -15434
rect -4871 -15694 -4837 -15450
rect -4782 -15481 -4748 -15362
rect -4714 -15400 -4638 -15394
rect -4714 -15434 -4698 -15400
rect -4654 -15434 -4638 -15400
rect -4714 -15450 -4638 -15434
rect -4802 -15534 -4792 -15481
rect -4739 -15534 -4729 -15481
rect -4693 -15694 -4659 -15450
rect -4892 -15710 -4816 -15694
rect -4892 -15744 -4876 -15710
rect -4832 -15744 -4816 -15710
rect -4892 -15750 -4816 -15744
rect -4714 -15710 -4638 -15694
rect -4714 -15744 -4698 -15710
rect -4654 -15744 -4638 -15710
rect -4714 -15750 -4638 -15744
rect -4604 -15782 -4570 -15362
rect -4536 -15400 -4460 -15394
rect -4536 -15434 -4520 -15400
rect -4476 -15434 -4460 -15400
rect -4536 -15450 -4460 -15434
rect -4515 -15694 -4481 -15450
rect -4426 -15589 -4392 -15362
rect -4358 -15400 -4282 -15394
rect -4358 -15434 -4342 -15400
rect -4298 -15434 -4282 -15400
rect -4358 -15450 -4282 -15434
rect -4445 -15641 -4435 -15589
rect -4383 -15641 -4373 -15589
rect -4337 -15694 -4303 -15450
rect -4536 -15710 -4460 -15694
rect -4536 -15744 -4520 -15710
rect -4476 -15744 -4460 -15710
rect -4536 -15750 -4460 -15744
rect -4358 -15710 -4282 -15694
rect -4358 -15744 -4342 -15710
rect -4298 -15744 -4282 -15710
rect -4358 -15750 -4282 -15744
rect -4248 -15782 -4214 -15362
rect -4180 -15400 -4104 -15394
rect -4180 -15434 -4164 -15400
rect -4120 -15434 -4104 -15400
rect -4180 -15450 -4104 -15434
rect -3935 -15589 -3883 -15006
rect -3945 -15641 -3935 -15589
rect -3883 -15641 -3873 -15589
rect -4180 -15710 -4104 -15694
rect -4180 -15744 -4164 -15710
rect -4120 -15744 -4104 -15710
rect -4180 -15750 -4104 -15744
rect -6034 -15794 -5988 -15782
rect -6034 -16050 -6028 -15794
rect -5994 -16050 -5988 -15794
rect -6034 -16062 -5988 -16050
rect -5856 -15794 -5810 -15782
rect -5856 -16050 -5850 -15794
rect -5816 -16050 -5810 -15794
rect -5856 -16062 -5810 -16050
rect -5678 -15794 -5632 -15782
rect -5678 -16050 -5672 -15794
rect -5638 -16050 -5632 -15794
rect -5678 -16062 -5632 -16050
rect -5500 -15794 -5454 -15782
rect -5500 -16050 -5494 -15794
rect -5460 -16050 -5454 -15794
rect -5500 -16062 -5454 -16050
rect -5322 -15794 -5276 -15782
rect -5322 -16050 -5316 -15794
rect -5282 -16050 -5276 -15794
rect -5322 -16062 -5276 -16050
rect -5144 -15794 -5098 -15782
rect -5144 -16050 -5138 -15794
rect -5104 -16050 -5098 -15794
rect -5144 -16062 -5098 -16050
rect -4966 -15794 -4920 -15782
rect -4966 -16050 -4960 -15794
rect -4926 -16050 -4920 -15794
rect -4966 -16062 -4920 -16050
rect -4788 -15794 -4742 -15782
rect -4788 -16050 -4782 -15794
rect -4748 -16050 -4742 -15794
rect -4788 -16062 -4742 -16050
rect -4610 -15794 -4564 -15782
rect -4610 -16050 -4604 -15794
rect -4570 -16050 -4564 -15794
rect -4610 -16062 -4564 -16050
rect -4432 -15794 -4386 -15782
rect -4432 -16050 -4426 -15794
rect -4392 -16050 -4386 -15794
rect -4432 -16062 -4386 -16050
rect -4254 -15794 -4208 -15782
rect -4254 -16050 -4248 -15794
rect -4214 -16050 -4208 -15794
rect -4254 -16062 -4208 -16050
rect -4076 -15794 -4030 -15782
rect -4076 -16050 -4070 -15794
rect -4036 -16050 -4030 -15794
rect -4076 -16062 -4030 -16050
rect -6028 -16185 -5994 -16062
rect -5960 -16100 -5884 -16094
rect -5960 -16134 -5944 -16100
rect -5900 -16134 -5884 -16100
rect -5960 -16150 -5884 -16134
rect -5939 -16185 -5905 -16150
rect -5850 -16185 -5816 -16062
rect -5782 -16100 -5706 -16094
rect -5782 -16134 -5766 -16100
rect -5722 -16134 -5706 -16100
rect -5782 -16150 -5706 -16134
rect -6169 -16246 -6159 -16193
rect -6106 -16246 -6096 -16193
rect -6028 -16219 -5816 -16185
rect -6159 -17007 -6106 -16246
rect -5850 -16294 -5816 -16219
rect -5870 -16347 -5860 -16294
rect -5807 -16347 -5797 -16294
rect -5761 -16394 -5727 -16150
rect -5960 -16410 -5884 -16394
rect -5960 -16444 -5944 -16410
rect -5900 -16444 -5884 -16410
rect -5960 -16450 -5884 -16444
rect -5782 -16410 -5706 -16394
rect -5782 -16444 -5766 -16410
rect -5722 -16444 -5706 -16410
rect -5782 -16450 -5706 -16444
rect -5672 -16482 -5638 -16062
rect -5604 -16100 -5528 -16094
rect -5604 -16134 -5588 -16100
rect -5544 -16134 -5528 -16100
rect -5604 -16150 -5528 -16134
rect -5583 -16394 -5549 -16150
rect -5494 -16193 -5460 -16062
rect -5426 -16100 -5350 -16094
rect -5426 -16134 -5410 -16100
rect -5366 -16134 -5350 -16100
rect -5426 -16150 -5350 -16134
rect -5514 -16246 -5504 -16193
rect -5451 -16246 -5441 -16193
rect -5405 -16394 -5371 -16150
rect -5604 -16410 -5528 -16394
rect -5604 -16444 -5588 -16410
rect -5544 -16444 -5528 -16410
rect -5604 -16450 -5528 -16444
rect -5426 -16410 -5350 -16394
rect -5426 -16444 -5410 -16410
rect -5366 -16444 -5350 -16410
rect -5426 -16450 -5350 -16444
rect -5316 -16482 -5282 -16062
rect -5248 -16100 -5172 -16094
rect -5248 -16134 -5232 -16100
rect -5188 -16134 -5172 -16100
rect -5248 -16150 -5172 -16134
rect -5227 -16394 -5193 -16150
rect -5138 -16294 -5104 -16062
rect -5070 -16100 -4994 -16094
rect -5070 -16134 -5054 -16100
rect -5010 -16134 -4994 -16100
rect -5070 -16150 -4994 -16134
rect -5158 -16347 -5148 -16294
rect -5095 -16347 -5085 -16294
rect -5049 -16394 -5015 -16150
rect -5248 -16410 -5172 -16394
rect -5248 -16444 -5232 -16410
rect -5188 -16444 -5172 -16410
rect -5248 -16450 -5172 -16444
rect -5070 -16410 -4994 -16394
rect -5070 -16444 -5054 -16410
rect -5010 -16444 -4994 -16410
rect -5070 -16450 -4994 -16444
rect -4960 -16482 -4926 -16062
rect -4892 -16100 -4816 -16094
rect -4892 -16134 -4876 -16100
rect -4832 -16134 -4816 -16100
rect -4892 -16150 -4816 -16134
rect -4871 -16394 -4837 -16150
rect -4782 -16193 -4748 -16062
rect -4714 -16100 -4638 -16094
rect -4714 -16134 -4698 -16100
rect -4654 -16134 -4638 -16100
rect -4714 -16150 -4638 -16134
rect -4802 -16246 -4792 -16193
rect -4739 -16246 -4729 -16193
rect -4693 -16394 -4659 -16150
rect -4892 -16410 -4816 -16394
rect -4892 -16444 -4876 -16410
rect -4832 -16444 -4816 -16410
rect -4892 -16450 -4816 -16444
rect -4714 -16410 -4638 -16394
rect -4714 -16444 -4698 -16410
rect -4654 -16444 -4638 -16410
rect -4714 -16450 -4638 -16444
rect -4604 -16482 -4570 -16062
rect -4536 -16100 -4460 -16094
rect -4536 -16134 -4520 -16100
rect -4476 -16134 -4460 -16100
rect -4536 -16150 -4460 -16134
rect -4515 -16394 -4481 -16150
rect -4426 -16294 -4392 -16062
rect -4358 -16100 -4282 -16094
rect -4358 -16134 -4342 -16100
rect -4298 -16134 -4282 -16100
rect -4358 -16150 -4282 -16134
rect -4446 -16347 -4436 -16294
rect -4383 -16347 -4373 -16294
rect -4337 -16394 -4303 -16150
rect -4248 -16185 -4214 -16062
rect -4180 -16100 -4104 -16094
rect -4180 -16134 -4164 -16100
rect -4120 -16134 -4104 -16100
rect -4180 -16150 -4104 -16134
rect -4159 -16185 -4125 -16150
rect -4070 -16185 -4036 -16062
rect -4248 -16219 -4036 -16185
rect -4536 -16410 -4460 -16394
rect -4536 -16444 -4520 -16410
rect -4476 -16444 -4460 -16410
rect -4536 -16450 -4460 -16444
rect -4358 -16410 -4282 -16394
rect -4358 -16444 -4342 -16410
rect -4298 -16444 -4282 -16410
rect -4358 -16450 -4282 -16444
rect -4248 -16482 -4214 -16219
rect -3935 -16295 -3883 -15641
rect -2447 -15821 -2394 -12325
rect -2315 -14543 -2262 -9978
rect -2105 -10048 -2029 -10032
rect -2105 -10049 -2089 -10048
rect -2175 -10082 -2089 -10049
rect -2045 -10049 -2029 -10048
rect -1995 -10049 -1961 -9473
rect -1927 -9438 -1851 -9432
rect -1927 -9472 -1911 -9438
rect -1867 -9472 -1851 -9438
rect -1927 -9488 -1851 -9472
rect -1906 -9546 -1872 -9488
rect -1926 -9599 -1916 -9546
rect -1863 -9599 -1853 -9546
rect -1926 -9978 -1916 -9925
rect -1863 -9978 -1853 -9925
rect -1906 -10032 -1872 -9978
rect -2045 -10082 -1961 -10049
rect -2175 -10083 -1961 -10082
rect -2175 -10120 -2141 -10083
rect -2105 -10088 -2029 -10083
rect -1995 -10120 -1961 -10083
rect -1927 -10048 -1851 -10032
rect -1927 -10082 -1911 -10048
rect -1867 -10082 -1851 -10048
rect -1927 -10088 -1851 -10082
rect -1817 -10120 -1783 -9400
rect -1749 -9438 -1673 -9432
rect -1749 -9472 -1733 -9438
rect -1689 -9472 -1673 -9438
rect -1749 -9488 -1673 -9472
rect -1728 -9546 -1694 -9488
rect -1748 -9599 -1738 -9546
rect -1685 -9599 -1675 -9546
rect -1748 -9979 -1738 -9926
rect -1685 -9979 -1675 -9926
rect -1728 -10032 -1694 -9979
rect -1749 -10048 -1673 -10032
rect -1749 -10082 -1733 -10048
rect -1689 -10082 -1673 -10048
rect -1749 -10088 -1673 -10082
rect -1639 -10120 -1605 -9400
rect -1571 -9438 -1495 -9432
rect -1571 -9472 -1555 -9438
rect -1511 -9472 -1495 -9438
rect -1571 -9488 -1495 -9472
rect -1549 -9546 -1515 -9488
rect -1568 -9599 -1558 -9546
rect -1505 -9599 -1495 -9546
rect -1570 -9978 -1560 -9925
rect -1507 -9978 -1497 -9925
rect -1550 -10032 -1516 -9978
rect -1571 -10048 -1495 -10032
rect -1571 -10082 -1555 -10048
rect -1511 -10082 -1495 -10048
rect -1571 -10088 -1495 -10082
rect -1461 -10120 -1427 -9400
rect -1393 -9438 -1317 -9432
rect -1393 -9472 -1377 -9438
rect -1333 -9472 -1317 -9438
rect -1393 -9488 -1317 -9472
rect -1372 -9924 -1338 -9488
rect -1392 -9977 -1382 -9924
rect -1329 -9977 -1319 -9924
rect -1393 -10048 -1317 -10032
rect -1393 -10082 -1377 -10048
rect -1333 -10082 -1317 -10048
rect -1393 -10088 -1317 -10082
rect -1283 -10120 -1249 -9400
rect -1215 -9438 -1139 -9432
rect -1215 -9472 -1199 -9438
rect -1155 -9472 -1139 -9438
rect -1215 -9488 -1139 -9472
rect -1215 -10048 -1139 -10032
rect -1215 -10082 -1199 -10048
rect -1155 -10082 -1139 -10048
rect -1215 -10088 -1139 -10082
rect -1105 -10120 -1071 -9400
rect -1037 -9438 -961 -9432
rect -1037 -9472 -1021 -9438
rect -977 -9472 -961 -9438
rect -1037 -9488 -961 -9472
rect -1037 -10048 -961 -10032
rect -1037 -10082 -1021 -10048
rect -977 -10082 -961 -10048
rect -1037 -10088 -961 -10082
rect -927 -10120 -893 -9400
rect -859 -9438 -783 -9432
rect -859 -9472 -843 -9438
rect -799 -9472 -783 -9438
rect -859 -9488 -783 -9472
rect -859 -10048 -783 -10032
rect -859 -10082 -843 -10048
rect -799 -10082 -783 -10048
rect -859 -10088 -783 -10082
rect -749 -10120 -715 -9400
rect -681 -9438 -605 -9432
rect -681 -9472 -665 -9438
rect -621 -9472 -605 -9438
rect -681 -9488 -605 -9472
rect -681 -10048 -605 -10032
rect -681 -10082 -665 -10048
rect -621 -10082 -605 -10048
rect -681 -10088 -605 -10082
rect -571 -10120 -537 -9400
rect -503 -9438 -427 -9432
rect -503 -9472 -487 -9438
rect -443 -9472 -427 -9438
rect -503 -9488 -427 -9472
rect -503 -10048 -427 -10032
rect -503 -10082 -487 -10048
rect -443 -10082 -427 -10048
rect -503 -10088 -427 -10082
rect -393 -10120 -359 -9400
rect -325 -9438 -249 -9432
rect -325 -9472 -309 -9438
rect -265 -9472 -249 -9438
rect -325 -9488 -249 -9472
rect -303 -9546 -269 -9488
rect -322 -9599 -312 -9546
rect -259 -9599 -249 -9546
rect -324 -9978 -314 -9925
rect -261 -9978 -251 -9925
rect -304 -10032 -270 -9978
rect -325 -10048 -249 -10032
rect -325 -10082 -309 -10048
rect -265 -10082 -249 -10048
rect -325 -10088 -249 -10082
rect -215 -10120 -181 -9400
rect -147 -9438 -71 -9432
rect -147 -9472 -131 -9438
rect -87 -9472 -71 -9438
rect -147 -9488 -71 -9472
rect -126 -9545 -92 -9488
rect -146 -9598 -136 -9545
rect -83 -9598 -73 -9545
rect -146 -9979 -136 -9926
rect -83 -9979 -73 -9926
rect -126 -10032 -92 -9979
rect -147 -10048 -71 -10032
rect -147 -10082 -131 -10048
rect -87 -10082 -71 -10048
rect -147 -10088 -71 -10082
rect -37 -10120 -3 -9400
rect 31 -9438 107 -9432
rect 31 -9472 47 -9438
rect 91 -9472 107 -9438
rect 31 -9488 107 -9472
rect 52 -9546 86 -9488
rect 32 -9599 42 -9546
rect 95 -9599 105 -9546
rect 33 -9978 43 -9925
rect 96 -9978 106 -9925
rect 52 -10032 86 -9978
rect 31 -10048 107 -10032
rect 31 -10082 47 -10048
rect 91 -10082 107 -10048
rect 31 -10088 107 -10082
rect 141 -10120 175 -9400
rect 209 -9438 285 -9432
rect 209 -9472 225 -9438
rect 269 -9472 285 -9438
rect 209 -9488 285 -9472
rect 231 -9545 265 -9488
rect 212 -9598 222 -9545
rect 275 -9598 285 -9545
rect 210 -9978 220 -9925
rect 273 -9978 283 -9925
rect 230 -10032 264 -9978
rect 209 -10048 285 -10032
rect 209 -10082 225 -10048
rect 269 -10082 285 -10048
rect 209 -10088 285 -10082
rect 319 -10120 353 -9400
rect 387 -9438 463 -9432
rect 387 -9472 403 -9438
rect 447 -9472 463 -9438
rect 387 -9488 463 -9472
rect 408 -9546 442 -9488
rect 389 -9599 399 -9546
rect 452 -9599 462 -9546
rect 388 -9978 398 -9925
rect 451 -9978 461 -9925
rect 408 -10032 442 -9978
rect 387 -10048 463 -10032
rect 387 -10082 403 -10048
rect 447 -10082 463 -10048
rect 387 -10088 463 -10082
rect 497 -10120 531 -9400
rect 565 -9438 641 -9432
rect 565 -9472 581 -9438
rect 625 -9472 641 -9438
rect 565 -9488 641 -9472
rect 587 -9546 621 -9488
rect 567 -9599 577 -9546
rect 630 -9599 640 -9546
rect 566 -9978 576 -9925
rect 629 -9978 639 -9925
rect 586 -10032 620 -9978
rect 565 -10048 641 -10032
rect 565 -10082 581 -10048
rect 625 -10082 641 -10048
rect 565 -10088 641 -10082
rect 675 -10120 709 -9400
rect 743 -9438 819 -9432
rect 743 -9472 759 -9438
rect 803 -9472 819 -9438
rect 743 -9488 819 -9472
rect 921 -9438 997 -9432
rect 921 -9472 937 -9438
rect 981 -9472 997 -9438
rect 921 -9488 997 -9472
rect 743 -10048 819 -10032
rect 743 -10082 759 -10048
rect 803 -10082 819 -10048
rect 743 -10088 819 -10082
rect 921 -10048 997 -10032
rect 921 -10082 937 -10048
rect 981 -10082 997 -10048
rect 921 -10088 997 -10082
rect 1031 -10120 1065 -9400
rect 1099 -9438 1175 -9432
rect 1099 -9472 1115 -9438
rect 1159 -9472 1175 -9438
rect 1099 -9488 1175 -9472
rect 1099 -10048 1175 -10032
rect 1099 -10082 1115 -10048
rect 1159 -10082 1175 -10048
rect 1099 -10088 1175 -10082
rect 1209 -10120 1243 -9400
rect 1277 -9438 1353 -9432
rect 1277 -9472 1293 -9438
rect 1337 -9472 1353 -9438
rect 1277 -9488 1353 -9472
rect 1277 -10048 1353 -10032
rect 1277 -10082 1293 -10048
rect 1337 -10082 1353 -10048
rect 1277 -10088 1353 -10082
rect 1387 -10120 1421 -9400
rect 1455 -9438 1531 -9432
rect 1455 -9472 1471 -9438
rect 1515 -9472 1531 -9438
rect 1455 -9488 1531 -9472
rect 1455 -10048 1531 -10032
rect 1455 -10082 1471 -10048
rect 1515 -10082 1531 -10048
rect 1455 -10088 1531 -10082
rect 1565 -10120 1599 -9400
rect 1633 -9438 1709 -9432
rect 1633 -9472 1649 -9438
rect 1693 -9472 1709 -9438
rect 1633 -9488 1709 -9472
rect 1633 -10048 1709 -10032
rect 1633 -10082 1649 -10048
rect 1693 -10082 1709 -10048
rect 1633 -10088 1709 -10082
rect 1743 -10120 1777 -9400
rect 1832 -9432 1866 -9426
rect 1811 -9438 1887 -9432
rect 1811 -9472 1827 -9438
rect 1871 -9472 1887 -9438
rect 1811 -9488 1887 -9472
rect 1832 -10032 1866 -9488
rect 1811 -10048 1887 -10032
rect 1811 -10082 1827 -10048
rect 1871 -10082 1887 -10048
rect 1811 -10088 1887 -10082
rect 1921 -10120 1955 -9400
rect 2010 -9432 2044 -9426
rect 1989 -9438 2065 -9432
rect 1989 -9472 2005 -9438
rect 2049 -9472 2065 -9438
rect 1989 -9488 2065 -9472
rect 2010 -10032 2044 -9488
rect 1989 -10048 2065 -10032
rect 1989 -10082 2005 -10048
rect 2049 -10082 2065 -10048
rect 1989 -10088 2065 -10082
rect 2099 -10120 2133 -9400
rect 2188 -9432 2222 -9426
rect 2167 -9438 2243 -9432
rect 2167 -9472 2183 -9438
rect 2227 -9472 2243 -9438
rect 2167 -9488 2243 -9472
rect 2188 -9547 2222 -9488
rect 2168 -9600 2178 -9547
rect 2231 -9600 2241 -9547
rect 2188 -10032 2222 -9600
rect 2167 -10048 2243 -10032
rect 2167 -10082 2183 -10048
rect 2227 -10082 2243 -10048
rect 2167 -10088 2243 -10082
rect 2277 -10120 2311 -9400
rect 2345 -9438 2421 -9432
rect 2345 -9472 2361 -9438
rect 2405 -9472 2421 -9438
rect 2345 -9488 2421 -9472
rect 2366 -9546 2400 -9488
rect 2347 -9599 2357 -9546
rect 2410 -9599 2420 -9546
rect 2346 -9978 2356 -9925
rect 2409 -9978 2419 -9925
rect 2366 -10032 2400 -9978
rect 2345 -10048 2421 -10032
rect 2345 -10082 2361 -10048
rect 2405 -10082 2421 -10048
rect 2345 -10088 2421 -10082
rect 2455 -10120 2489 -9400
rect 2523 -9438 2599 -9432
rect 2523 -9472 2539 -9438
rect 2583 -9472 2599 -9438
rect 2523 -9488 2599 -9472
rect 2544 -9546 2578 -9488
rect 2524 -9599 2534 -9546
rect 2587 -9599 2597 -9546
rect 2524 -9978 2534 -9925
rect 2587 -9978 2597 -9925
rect 2544 -10032 2578 -9978
rect 2523 -10048 2599 -10032
rect 2523 -10082 2539 -10048
rect 2583 -10082 2599 -10048
rect 2523 -10088 2599 -10082
rect 2633 -10120 2667 -9400
rect 2701 -9438 2777 -9432
rect 2701 -9472 2717 -9438
rect 2761 -9472 2777 -9438
rect 2701 -9488 2777 -9472
rect 2722 -9546 2756 -9488
rect 2703 -9599 2713 -9546
rect 2766 -9599 2776 -9546
rect 2702 -9979 2712 -9926
rect 2765 -9979 2775 -9926
rect 2722 -10032 2756 -9979
rect 2701 -10048 2777 -10032
rect 2701 -10082 2717 -10048
rect 2761 -10082 2777 -10048
rect 2701 -10088 2777 -10082
rect 2811 -10120 2845 -9400
rect 2879 -9438 2955 -9432
rect 2879 -9472 2895 -9438
rect 2939 -9472 2955 -9438
rect 2879 -9488 2955 -9472
rect 2881 -9978 2891 -9925
rect 2944 -9978 2954 -9925
rect 2900 -10032 2934 -9978
rect 2879 -10048 2955 -10032
rect 2879 -10082 2895 -10048
rect 2939 -10082 2955 -10048
rect 2879 -10088 2955 -10082
rect 2989 -10120 3023 -9400
rect 3057 -9438 3133 -9432
rect 3057 -9472 3073 -9438
rect 3117 -9472 3133 -9438
rect 3057 -9488 3133 -9472
rect 3059 -9978 3069 -9925
rect 3122 -9978 3132 -9925
rect 3078 -10032 3112 -9978
rect 3057 -10048 3133 -10032
rect 3057 -10082 3073 -10048
rect 3117 -10082 3133 -10048
rect 3057 -10088 3133 -10082
rect 3167 -10120 3201 -9400
rect 3235 -9438 3311 -9432
rect 3235 -9472 3251 -9438
rect 3295 -9472 3311 -9438
rect 3235 -9488 3311 -9472
rect 3256 -9925 3290 -9488
rect 3236 -9978 3246 -9925
rect 3299 -9978 3309 -9925
rect 3256 -10032 3290 -9978
rect 3235 -10048 3311 -10032
rect 3235 -10082 3251 -10048
rect 3295 -10082 3311 -10048
rect 3235 -10088 3311 -10082
rect 3345 -10120 3379 -9400
rect 3413 -9438 3489 -9432
rect 3413 -9472 3429 -9438
rect 3473 -9472 3489 -9438
rect 3413 -9488 3489 -9472
rect 3413 -10048 3489 -10032
rect 3413 -10082 3429 -10048
rect 3473 -10082 3489 -10048
rect 3413 -10088 3489 -10082
rect 3523 -10120 3557 -9400
rect 3591 -9438 3667 -9432
rect 3591 -9472 3607 -9438
rect 3651 -9472 3667 -9438
rect 3591 -9488 3667 -9472
rect 3591 -10048 3667 -10032
rect 3591 -10082 3607 -10048
rect 3651 -10082 3667 -10048
rect 3591 -10088 3667 -10082
rect 3701 -10120 3735 -9400
rect 3769 -9438 3845 -9432
rect 3769 -9472 3785 -9438
rect 3829 -9472 3845 -9438
rect 3769 -9488 3845 -9472
rect 3879 -9439 3913 -9400
rect 3947 -9438 4023 -9432
rect 3947 -9439 3963 -9438
rect 3879 -9472 3963 -9439
rect 4007 -9439 4023 -9438
rect 4056 -9439 4090 -9400
rect 4007 -9472 4090 -9439
rect 3879 -9473 4090 -9472
rect 3769 -10048 3845 -10032
rect 3769 -10082 3785 -10048
rect 3829 -10082 3845 -10048
rect 3769 -10088 3845 -10082
rect 3879 -10047 3913 -9473
rect 3947 -9488 4023 -9473
rect 4208 -9546 4261 -7976
rect 4771 -9262 4823 -7907
rect 4771 -9314 4824 -9262
rect 4761 -9367 4771 -9314
rect 4824 -9367 4834 -9314
rect 4198 -9599 4208 -9546
rect 4261 -9599 4271 -9546
rect 3947 -10047 4023 -10032
rect 3879 -10048 4092 -10047
rect 3879 -10081 3963 -10048
rect 3879 -10120 3913 -10081
rect 3947 -10082 3963 -10081
rect 4007 -10081 4092 -10048
rect 4007 -10082 4023 -10081
rect 3947 -10088 4023 -10082
rect 4058 -10120 4092 -10081
rect -2179 -10132 -2133 -10120
rect -2179 -10388 -2173 -10132
rect -2139 -10388 -2133 -10132
rect -2179 -10400 -2133 -10388
rect -2001 -10132 -1955 -10120
rect -2001 -10388 -1995 -10132
rect -1961 -10388 -1955 -10132
rect -2001 -10400 -1955 -10388
rect -1823 -10132 -1777 -10120
rect -1823 -10388 -1817 -10132
rect -1783 -10388 -1777 -10132
rect -1823 -10400 -1777 -10388
rect -1645 -10132 -1599 -10120
rect -1645 -10388 -1639 -10132
rect -1605 -10388 -1599 -10132
rect -1645 -10400 -1599 -10388
rect -1467 -10132 -1421 -10120
rect -1467 -10388 -1461 -10132
rect -1427 -10388 -1421 -10132
rect -1467 -10400 -1421 -10388
rect -1289 -10132 -1243 -10120
rect -1289 -10388 -1283 -10132
rect -1249 -10388 -1243 -10132
rect -1289 -10400 -1243 -10388
rect -1111 -10132 -1065 -10120
rect -1111 -10388 -1105 -10132
rect -1071 -10388 -1065 -10132
rect -1111 -10400 -1065 -10388
rect -933 -10132 -887 -10120
rect -933 -10388 -927 -10132
rect -893 -10388 -887 -10132
rect -933 -10400 -887 -10388
rect -755 -10132 -709 -10120
rect -755 -10388 -749 -10132
rect -715 -10388 -709 -10132
rect -755 -10400 -709 -10388
rect -577 -10132 -531 -10120
rect -577 -10388 -571 -10132
rect -537 -10388 -531 -10132
rect -577 -10400 -531 -10388
rect -399 -10132 -353 -10120
rect -399 -10388 -393 -10132
rect -359 -10388 -353 -10132
rect -399 -10400 -353 -10388
rect -221 -10132 -175 -10120
rect -221 -10388 -215 -10132
rect -181 -10388 -175 -10132
rect -221 -10400 -175 -10388
rect -43 -10132 3 -10120
rect -43 -10388 -37 -10132
rect -3 -10388 3 -10132
rect -43 -10400 3 -10388
rect 135 -10132 181 -10120
rect 135 -10388 141 -10132
rect 175 -10388 181 -10132
rect 135 -10400 181 -10388
rect 313 -10132 359 -10120
rect 313 -10388 319 -10132
rect 353 -10388 359 -10132
rect 313 -10400 359 -10388
rect 491 -10132 537 -10120
rect 491 -10388 497 -10132
rect 531 -10388 537 -10132
rect 491 -10400 537 -10388
rect 669 -10132 715 -10120
rect 669 -10388 675 -10132
rect 709 -10388 715 -10132
rect 669 -10400 715 -10388
rect 847 -10132 893 -10120
rect 847 -10388 853 -10132
rect 887 -10388 893 -10132
rect 847 -10400 893 -10388
rect 1025 -10132 1071 -10120
rect 1025 -10388 1031 -10132
rect 1065 -10388 1071 -10132
rect 1025 -10400 1071 -10388
rect 1203 -10132 1249 -10120
rect 1203 -10388 1209 -10132
rect 1243 -10388 1249 -10132
rect 1203 -10400 1249 -10388
rect 1381 -10132 1427 -10120
rect 1381 -10388 1387 -10132
rect 1421 -10388 1427 -10132
rect 1381 -10400 1427 -10388
rect 1559 -10132 1605 -10120
rect 1559 -10388 1565 -10132
rect 1599 -10388 1605 -10132
rect 1559 -10400 1605 -10388
rect 1737 -10132 1783 -10120
rect 1737 -10388 1743 -10132
rect 1777 -10388 1783 -10132
rect 1737 -10400 1783 -10388
rect 1915 -10132 1961 -10120
rect 1915 -10388 1921 -10132
rect 1955 -10388 1961 -10132
rect 1915 -10400 1961 -10388
rect 2093 -10132 2139 -10120
rect 2093 -10388 2099 -10132
rect 2133 -10388 2139 -10132
rect 2093 -10400 2139 -10388
rect 2271 -10132 2317 -10120
rect 2271 -10388 2277 -10132
rect 2311 -10388 2317 -10132
rect 2271 -10400 2317 -10388
rect 2449 -10132 2495 -10120
rect 2449 -10388 2455 -10132
rect 2489 -10388 2495 -10132
rect 2449 -10400 2495 -10388
rect 2627 -10132 2673 -10120
rect 2627 -10388 2633 -10132
rect 2667 -10388 2673 -10132
rect 2627 -10400 2673 -10388
rect 2805 -10132 2851 -10120
rect 2805 -10388 2811 -10132
rect 2845 -10388 2851 -10132
rect 2805 -10400 2851 -10388
rect 2983 -10132 3029 -10120
rect 2983 -10388 2989 -10132
rect 3023 -10388 3029 -10132
rect 2983 -10400 3029 -10388
rect 3161 -10132 3207 -10120
rect 3161 -10388 3167 -10132
rect 3201 -10388 3207 -10132
rect 3161 -10400 3207 -10388
rect 3339 -10132 3385 -10120
rect 3339 -10388 3345 -10132
rect 3379 -10388 3385 -10132
rect 3339 -10400 3385 -10388
rect 3517 -10132 3563 -10120
rect 3517 -10388 3523 -10132
rect 3557 -10388 3563 -10132
rect 3517 -10400 3563 -10388
rect 3695 -10132 3741 -10120
rect 3695 -10388 3701 -10132
rect 3735 -10388 3741 -10132
rect 3695 -10400 3741 -10388
rect 3873 -10132 3919 -10120
rect 3873 -10388 3879 -10132
rect 3913 -10388 3919 -10132
rect 3873 -10400 3919 -10388
rect 4051 -10132 4097 -10120
rect 4051 -10388 4057 -10132
rect 4091 -10388 4097 -10132
rect 4051 -10400 4097 -10388
rect -2105 -10438 -2029 -10432
rect -2105 -10472 -2089 -10438
rect -2045 -10472 -2029 -10438
rect -2105 -10488 -2029 -10472
rect -1927 -10438 -1851 -10432
rect -1927 -10472 -1911 -10438
rect -1867 -10472 -1851 -10438
rect -1927 -10488 -1851 -10472
rect -1749 -10438 -1673 -10432
rect -1749 -10472 -1733 -10438
rect -1689 -10472 -1673 -10438
rect -1749 -10488 -1673 -10472
rect -1571 -10438 -1495 -10432
rect -1571 -10472 -1555 -10438
rect -1511 -10472 -1495 -10438
rect -1571 -10488 -1495 -10472
rect -1393 -10438 -1317 -10432
rect -1393 -10472 -1377 -10438
rect -1333 -10472 -1317 -10438
rect -1393 -10488 -1317 -10472
rect -1215 -10438 -1139 -10432
rect -1215 -10472 -1199 -10438
rect -1155 -10472 -1139 -10438
rect -1215 -10488 -1139 -10472
rect -1037 -10438 -961 -10432
rect -1037 -10472 -1021 -10438
rect -977 -10472 -961 -10438
rect -1037 -10488 -961 -10472
rect -859 -10438 -783 -10432
rect -859 -10472 -843 -10438
rect -799 -10472 -783 -10438
rect -859 -10488 -783 -10472
rect -681 -10438 -605 -10432
rect -681 -10472 -665 -10438
rect -621 -10472 -605 -10438
rect -681 -10488 -605 -10472
rect -503 -10438 -427 -10432
rect -503 -10472 -487 -10438
rect -443 -10472 -427 -10438
rect -503 -10488 -427 -10472
rect -325 -10438 -249 -10432
rect -325 -10472 -309 -10438
rect -265 -10472 -249 -10438
rect -325 -10488 -249 -10472
rect -147 -10438 -71 -10432
rect -147 -10472 -131 -10438
rect -87 -10472 -71 -10438
rect -147 -10488 -71 -10472
rect 31 -10438 107 -10432
rect 31 -10472 47 -10438
rect 91 -10472 107 -10438
rect 31 -10488 107 -10472
rect 209 -10438 285 -10432
rect 209 -10472 225 -10438
rect 269 -10472 285 -10438
rect 209 -10488 285 -10472
rect 387 -10438 463 -10432
rect 387 -10472 403 -10438
rect 447 -10472 463 -10438
rect 387 -10488 463 -10472
rect 565 -10438 641 -10432
rect 565 -10472 581 -10438
rect 625 -10472 641 -10438
rect 565 -10488 641 -10472
rect 743 -10438 819 -10432
rect 853 -10438 887 -10400
rect 941 -10432 975 -10431
rect 921 -10438 997 -10432
rect 1031 -10438 1065 -10400
rect 1653 -10432 1687 -10431
rect 1099 -10438 1175 -10432
rect 743 -10472 759 -10438
rect 803 -10472 937 -10438
rect 981 -10472 1115 -10438
rect 1159 -10472 1175 -10438
rect 743 -10488 819 -10472
rect 921 -10488 997 -10472
rect 1099 -10488 1175 -10472
rect 1277 -10438 1353 -10432
rect 1277 -10472 1293 -10438
rect 1337 -10472 1353 -10438
rect 1277 -10488 1353 -10472
rect 1455 -10438 1531 -10432
rect 1455 -10472 1471 -10438
rect 1515 -10472 1531 -10438
rect 1455 -10488 1531 -10472
rect 1633 -10438 1709 -10432
rect 1633 -10472 1649 -10438
rect 1693 -10472 1709 -10438
rect 1633 -10488 1709 -10472
rect 1811 -10438 1887 -10432
rect 1811 -10472 1827 -10438
rect 1871 -10472 1887 -10438
rect 1811 -10488 1887 -10472
rect 1989 -10438 2065 -10432
rect 1989 -10472 2005 -10438
rect 2049 -10472 2065 -10438
rect 1989 -10488 2065 -10472
rect 2167 -10438 2243 -10432
rect 2167 -10472 2183 -10438
rect 2227 -10472 2243 -10438
rect 2167 -10488 2243 -10472
rect 2345 -10438 2421 -10432
rect 2345 -10472 2361 -10438
rect 2405 -10472 2421 -10438
rect 2345 -10488 2421 -10472
rect 2523 -10438 2599 -10432
rect 2523 -10472 2539 -10438
rect 2583 -10472 2599 -10438
rect 2523 -10488 2599 -10472
rect 2701 -10438 2777 -10432
rect 2701 -10472 2717 -10438
rect 2761 -10472 2777 -10438
rect 2701 -10488 2777 -10472
rect 2879 -10438 2955 -10432
rect 2879 -10472 2895 -10438
rect 2939 -10472 2955 -10438
rect 2879 -10488 2955 -10472
rect 3057 -10438 3133 -10432
rect 3057 -10472 3073 -10438
rect 3117 -10472 3133 -10438
rect 3057 -10488 3133 -10472
rect 3235 -10438 3311 -10432
rect 3235 -10472 3251 -10438
rect 3295 -10472 3311 -10438
rect 3235 -10488 3311 -10472
rect 3413 -10438 3489 -10432
rect 3413 -10472 3429 -10438
rect 3473 -10472 3489 -10438
rect 3413 -10488 3489 -10472
rect 3591 -10438 3667 -10432
rect 3591 -10472 3607 -10438
rect 3651 -10472 3667 -10438
rect 3591 -10488 3667 -10472
rect 3769 -10438 3845 -10432
rect 3769 -10472 3785 -10438
rect 3829 -10472 3845 -10438
rect 3769 -10488 3845 -10472
rect 3947 -10438 4023 -10432
rect 3947 -10472 3963 -10438
rect 4007 -10472 4023 -10438
rect 3947 -10488 4023 -10472
rect -1837 -10961 -1827 -10908
rect -1774 -10961 -1764 -10908
rect -1480 -10961 -1470 -10908
rect -1417 -10961 -1407 -10908
rect -2105 -11048 -2029 -11032
rect -2105 -11082 -2089 -11048
rect -2045 -11082 -2029 -11048
rect -2105 -11088 -2029 -11082
rect -1927 -11048 -1851 -11032
rect -1927 -11082 -1911 -11048
rect -1867 -11082 -1851 -11048
rect -1927 -11088 -1851 -11082
rect -1818 -11120 -1784 -10961
rect -1749 -11048 -1673 -11032
rect -1749 -11082 -1733 -11048
rect -1689 -11082 -1673 -11048
rect -1749 -11088 -1673 -11082
rect -1571 -11048 -1495 -11032
rect -1571 -11082 -1555 -11048
rect -1511 -11082 -1495 -11048
rect -1571 -11088 -1495 -11082
rect -1461 -11120 -1427 -10961
rect -1372 -11032 -1338 -10488
rect -1193 -11032 -1159 -10488
rect -1124 -10961 -1114 -10908
rect -1061 -10961 -1051 -10908
rect -1393 -11048 -1317 -11032
rect -1393 -11082 -1377 -11048
rect -1333 -11082 -1317 -11048
rect -1393 -11088 -1317 -11082
rect -1215 -11048 -1139 -11032
rect -1215 -11082 -1199 -11048
rect -1155 -11082 -1139 -11048
rect -1215 -11088 -1139 -11082
rect -1105 -11120 -1071 -10961
rect -1016 -11032 -982 -10488
rect -838 -11032 -804 -10488
rect -768 -10961 -758 -10908
rect -705 -10961 -695 -10908
rect -1037 -11048 -961 -11032
rect -1037 -11082 -1021 -11048
rect -977 -11082 -961 -11048
rect -1037 -11088 -961 -11082
rect -859 -11048 -783 -11032
rect -859 -11082 -843 -11048
rect -799 -11082 -783 -11048
rect -859 -11088 -783 -11082
rect -749 -11120 -715 -10961
rect -659 -11032 -625 -10488
rect -482 -11032 -448 -10488
rect 941 -10908 975 -10488
rect -412 -10961 -402 -10908
rect -349 -10961 -339 -10908
rect -56 -10961 -46 -10908
rect 7 -10961 17 -10908
rect 299 -10961 309 -10908
rect 362 -10961 372 -10908
rect 655 -10961 665 -10908
rect 718 -10961 728 -10908
rect 921 -10961 931 -10908
rect 984 -10961 994 -10908
rect 1189 -10961 1199 -10908
rect 1252 -10961 1262 -10908
rect -681 -11048 -605 -11032
rect -681 -11082 -665 -11048
rect -621 -11082 -605 -11048
rect -681 -11088 -605 -11082
rect -503 -11048 -427 -11032
rect -503 -11082 -487 -11048
rect -443 -11082 -427 -11048
rect -503 -11088 -427 -11082
rect -393 -11120 -359 -10961
rect -325 -11048 -249 -11032
rect -325 -11082 -309 -11048
rect -265 -11082 -249 -11048
rect -325 -11088 -249 -11082
rect -147 -11048 -71 -11032
rect -147 -11082 -131 -11048
rect -87 -11082 -71 -11048
rect -147 -11088 -71 -11082
rect -36 -11120 -2 -10961
rect 31 -11048 107 -11032
rect 31 -11082 47 -11048
rect 91 -11082 107 -11048
rect 31 -11088 107 -11082
rect 209 -11048 285 -11032
rect 209 -11082 225 -11048
rect 269 -11082 285 -11048
rect 209 -11088 285 -11082
rect 319 -11120 353 -10961
rect 387 -11048 463 -11032
rect 387 -11082 403 -11048
rect 447 -11082 463 -11048
rect 387 -11088 463 -11082
rect 565 -11048 641 -11032
rect 565 -11082 581 -11048
rect 625 -11082 641 -11048
rect 565 -11088 641 -11082
rect 675 -11120 709 -10961
rect 941 -11032 975 -10961
rect 743 -11048 819 -11032
rect 743 -11082 759 -11048
rect 803 -11082 819 -11048
rect 743 -11088 819 -11082
rect 921 -11048 997 -11032
rect 921 -11082 937 -11048
rect 981 -11082 997 -11048
rect 921 -11088 997 -11082
rect 1099 -11048 1175 -11032
rect 1099 -11082 1115 -11048
rect 1159 -11082 1175 -11048
rect 1099 -11088 1175 -11082
rect 1209 -11120 1243 -10961
rect 1299 -11032 1333 -10488
rect 1477 -11032 1511 -10488
rect 1546 -10961 1556 -10908
rect 1609 -10961 1619 -10908
rect 1277 -11048 1353 -11032
rect 1277 -11082 1293 -11048
rect 1337 -11082 1353 -11048
rect 1277 -11088 1353 -11082
rect 1455 -11048 1531 -11032
rect 1455 -11082 1471 -11048
rect 1515 -11082 1531 -11048
rect 1455 -11088 1531 -11082
rect 1566 -11120 1600 -10961
rect 1653 -11032 1687 -10488
rect 1832 -11032 1866 -10488
rect 1903 -10961 1913 -10908
rect 1966 -10961 1976 -10908
rect 1633 -11048 1709 -11032
rect 1633 -11082 1649 -11048
rect 1693 -11082 1709 -11048
rect 1633 -11088 1709 -11082
rect 1811 -11048 1887 -11032
rect 1811 -11082 1827 -11048
rect 1871 -11082 1887 -11048
rect 1811 -11088 1887 -11082
rect 1922 -11120 1956 -10961
rect 2010 -11032 2044 -10488
rect 2188 -11032 2222 -10488
rect 2258 -10961 2268 -10908
rect 2321 -10961 2331 -10908
rect 2613 -10961 2623 -10908
rect 2676 -10961 2686 -10908
rect 2970 -10961 2980 -10908
rect 3033 -10961 3043 -10908
rect 3325 -10961 3335 -10908
rect 3388 -10961 3398 -10908
rect 1989 -11048 2065 -11032
rect 1989 -11082 2005 -11048
rect 2049 -11082 2065 -11048
rect 1989 -11088 2065 -11082
rect 2167 -11048 2243 -11032
rect 2167 -11082 2183 -11048
rect 2227 -11082 2243 -11048
rect 2167 -11088 2243 -11082
rect 2277 -11120 2311 -10961
rect 2345 -11048 2421 -11032
rect 2345 -11082 2361 -11048
rect 2405 -11082 2421 -11048
rect 2345 -11088 2421 -11082
rect 2523 -11048 2599 -11032
rect 2523 -11082 2539 -11048
rect 2583 -11082 2599 -11048
rect 2523 -11088 2599 -11082
rect 2633 -11120 2667 -10961
rect 2701 -11048 2777 -11032
rect 2701 -11082 2717 -11048
rect 2761 -11082 2777 -11048
rect 2701 -11088 2777 -11082
rect 2879 -11048 2955 -11032
rect 2879 -11082 2895 -11048
rect 2939 -11082 2955 -11048
rect 2879 -11088 2955 -11082
rect 2989 -11120 3023 -10961
rect 3057 -11048 3133 -11032
rect 3057 -11082 3073 -11048
rect 3117 -11082 3133 -11048
rect 3057 -11088 3133 -11082
rect 3235 -11048 3311 -11032
rect 3235 -11082 3251 -11048
rect 3295 -11082 3311 -11048
rect 3235 -11088 3311 -11082
rect 3345 -11120 3379 -10961
rect 3434 -11032 3468 -10488
rect 3613 -11032 3647 -10488
rect 3682 -10961 3692 -10908
rect 3745 -10961 3755 -10908
rect 3413 -11048 3489 -11032
rect 3413 -11082 3429 -11048
rect 3473 -11082 3489 -11048
rect 3413 -11088 3489 -11082
rect 3591 -11048 3667 -11032
rect 3591 -11082 3607 -11048
rect 3651 -11082 3667 -11048
rect 3591 -11088 3667 -11082
rect 3701 -11120 3735 -10961
rect 3791 -11032 3825 -10488
rect 3769 -11048 3845 -11032
rect 3769 -11082 3785 -11048
rect 3829 -11082 3845 -11048
rect 3769 -11088 3845 -11082
rect 3947 -11048 4023 -11032
rect 3947 -11082 3963 -11048
rect 4007 -11082 4023 -11048
rect 3947 -11088 4023 -11082
rect -2179 -11132 -2133 -11120
rect -2179 -11388 -2173 -11132
rect -2139 -11388 -2133 -11132
rect -2179 -11400 -2133 -11388
rect -2001 -11132 -1955 -11120
rect -2001 -11388 -1995 -11132
rect -1961 -11388 -1955 -11132
rect -2001 -11400 -1955 -11388
rect -1823 -11132 -1777 -11120
rect -1823 -11388 -1817 -11132
rect -1783 -11388 -1777 -11132
rect -1823 -11400 -1777 -11388
rect -1645 -11132 -1599 -11120
rect -1645 -11388 -1639 -11132
rect -1605 -11388 -1599 -11132
rect -1645 -11400 -1599 -11388
rect -1467 -11132 -1421 -11120
rect -1467 -11388 -1461 -11132
rect -1427 -11388 -1421 -11132
rect -1467 -11400 -1421 -11388
rect -1289 -11132 -1243 -11120
rect -1289 -11388 -1283 -11132
rect -1249 -11388 -1243 -11132
rect -1289 -11400 -1243 -11388
rect -1111 -11132 -1065 -11120
rect -1111 -11388 -1105 -11132
rect -1071 -11388 -1065 -11132
rect -1111 -11400 -1065 -11388
rect -933 -11132 -887 -11120
rect -933 -11388 -927 -11132
rect -893 -11388 -887 -11132
rect -933 -11400 -887 -11388
rect -755 -11132 -709 -11120
rect -755 -11388 -749 -11132
rect -715 -11388 -709 -11132
rect -755 -11400 -709 -11388
rect -577 -11132 -531 -11120
rect -577 -11388 -571 -11132
rect -537 -11388 -531 -11132
rect -577 -11400 -531 -11388
rect -399 -11132 -353 -11120
rect -399 -11388 -393 -11132
rect -359 -11388 -353 -11132
rect -399 -11400 -353 -11388
rect -221 -11132 -175 -11120
rect -221 -11388 -215 -11132
rect -181 -11388 -175 -11132
rect -221 -11400 -175 -11388
rect -43 -11132 3 -11120
rect -43 -11388 -37 -11132
rect -3 -11388 3 -11132
rect -43 -11400 3 -11388
rect 135 -11132 181 -11120
rect 135 -11388 141 -11132
rect 175 -11388 181 -11132
rect 135 -11400 181 -11388
rect 313 -11132 359 -11120
rect 313 -11388 319 -11132
rect 353 -11388 359 -11132
rect 313 -11400 359 -11388
rect 491 -11132 537 -11120
rect 491 -11388 497 -11132
rect 531 -11388 537 -11132
rect 491 -11400 537 -11388
rect 669 -11132 715 -11120
rect 669 -11388 675 -11132
rect 709 -11388 715 -11132
rect 669 -11400 715 -11388
rect 847 -11132 893 -11120
rect 847 -11388 853 -11132
rect 887 -11388 893 -11132
rect 847 -11400 893 -11388
rect 1025 -11132 1071 -11120
rect 1025 -11388 1031 -11132
rect 1065 -11388 1071 -11132
rect 1025 -11400 1071 -11388
rect 1203 -11132 1249 -11120
rect 1203 -11388 1209 -11132
rect 1243 -11388 1249 -11132
rect 1203 -11400 1249 -11388
rect 1381 -11132 1427 -11120
rect 1381 -11388 1387 -11132
rect 1421 -11388 1427 -11132
rect 1381 -11400 1427 -11388
rect 1559 -11132 1605 -11120
rect 1559 -11388 1565 -11132
rect 1599 -11388 1605 -11132
rect 1559 -11400 1605 -11388
rect 1737 -11132 1783 -11120
rect 1737 -11388 1743 -11132
rect 1777 -11388 1783 -11132
rect 1737 -11400 1783 -11388
rect 1915 -11132 1961 -11120
rect 1915 -11388 1921 -11132
rect 1955 -11388 1961 -11132
rect 1915 -11400 1961 -11388
rect 2093 -11132 2139 -11120
rect 2093 -11388 2099 -11132
rect 2133 -11388 2139 -11132
rect 2093 -11400 2139 -11388
rect 2271 -11132 2317 -11120
rect 2271 -11388 2277 -11132
rect 2311 -11388 2317 -11132
rect 2271 -11400 2317 -11388
rect 2449 -11132 2495 -11120
rect 2449 -11388 2455 -11132
rect 2489 -11388 2495 -11132
rect 2449 -11400 2495 -11388
rect 2627 -11132 2673 -11120
rect 2627 -11388 2633 -11132
rect 2667 -11388 2673 -11132
rect 2627 -11400 2673 -11388
rect 2805 -11132 2851 -11120
rect 2805 -11388 2811 -11132
rect 2845 -11388 2851 -11132
rect 2805 -11400 2851 -11388
rect 2983 -11132 3029 -11120
rect 2983 -11388 2989 -11132
rect 3023 -11388 3029 -11132
rect 2983 -11400 3029 -11388
rect 3161 -11132 3207 -11120
rect 3161 -11388 3167 -11132
rect 3201 -11388 3207 -11132
rect 3161 -11400 3207 -11388
rect 3339 -11132 3385 -11120
rect 3339 -11388 3345 -11132
rect 3379 -11388 3385 -11132
rect 3339 -11400 3385 -11388
rect 3517 -11132 3563 -11120
rect 3517 -11388 3523 -11132
rect 3557 -11388 3563 -11132
rect 3517 -11400 3563 -11388
rect 3695 -11132 3741 -11120
rect 3695 -11388 3701 -11132
rect 3735 -11388 3741 -11132
rect 3695 -11400 3741 -11388
rect 3873 -11132 3919 -11120
rect 3873 -11388 3879 -11132
rect 3913 -11388 3919 -11132
rect 3873 -11400 3919 -11388
rect 4051 -11132 4097 -11120
rect 4051 -11388 4057 -11132
rect 4091 -11388 4097 -11132
rect 4051 -11400 4097 -11388
rect -2172 -11439 -2138 -11400
rect -2105 -11438 -2029 -11432
rect -2105 -11439 -2089 -11438
rect -2172 -11472 -2089 -11439
rect -2045 -11439 -2029 -11438
rect -1995 -11439 -1961 -11400
rect -2045 -11472 -1961 -11439
rect -2172 -11473 -1961 -11472
rect -2105 -11488 -2029 -11473
rect -1995 -11637 -1961 -11473
rect -1927 -11438 -1851 -11432
rect -1927 -11472 -1911 -11438
rect -1867 -11472 -1851 -11438
rect -1927 -11488 -1851 -11472
rect -2014 -11690 -2004 -11637
rect -1951 -11690 -1941 -11637
rect -2105 -12047 -2029 -12032
rect -1995 -12047 -1961 -11690
rect -1905 -11919 -1871 -11488
rect -1925 -11972 -1915 -11919
rect -1862 -11972 -1852 -11919
rect -1905 -12032 -1871 -11972
rect -2176 -12048 -1961 -12047
rect -2176 -12081 -2089 -12048
rect -2176 -12120 -2142 -12081
rect -2105 -12082 -2089 -12081
rect -2045 -12081 -1961 -12048
rect -2045 -12082 -2029 -12081
rect -2105 -12088 -2029 -12082
rect -1995 -12120 -1961 -12081
rect -1927 -12048 -1851 -12032
rect -1927 -12082 -1911 -12048
rect -1867 -12082 -1851 -12048
rect -1927 -12088 -1851 -12082
rect -1818 -12120 -1784 -11400
rect -1749 -11438 -1673 -11432
rect -1749 -11472 -1733 -11438
rect -1689 -11472 -1673 -11438
rect -1749 -11488 -1673 -11472
rect -1728 -11919 -1694 -11488
rect -1639 -11528 -1605 -11400
rect -1571 -11438 -1495 -11432
rect -1571 -11472 -1555 -11438
rect -1511 -11472 -1495 -11438
rect -1571 -11488 -1495 -11472
rect -1659 -11581 -1649 -11528
rect -1596 -11581 -1586 -11528
rect -1549 -11919 -1515 -11488
rect -1748 -11972 -1738 -11919
rect -1685 -11972 -1675 -11919
rect -1569 -11972 -1559 -11919
rect -1506 -11972 -1496 -11919
rect -1728 -12032 -1694 -11972
rect -1549 -12032 -1515 -11972
rect -1749 -12048 -1673 -12032
rect -1749 -12082 -1733 -12048
rect -1689 -12082 -1673 -12048
rect -1749 -12088 -1673 -12082
rect -1571 -12048 -1495 -12032
rect -1571 -12082 -1555 -12048
rect -1511 -12082 -1495 -12048
rect -1571 -12088 -1495 -12082
rect -1461 -12120 -1427 -11400
rect -1393 -11438 -1317 -11432
rect -1393 -11472 -1377 -11438
rect -1333 -11472 -1317 -11438
rect -1393 -11488 -1317 -11472
rect -1372 -11919 -1338 -11488
rect -1283 -11526 -1249 -11400
rect -1215 -11438 -1139 -11432
rect -1215 -11472 -1199 -11438
rect -1155 -11472 -1139 -11438
rect -1215 -11488 -1139 -11472
rect -1284 -11528 -1249 -11526
rect -1303 -11581 -1293 -11528
rect -1240 -11581 -1230 -11528
rect -1391 -11972 -1381 -11919
rect -1328 -11972 -1318 -11919
rect -1372 -12032 -1338 -11972
rect -1393 -12048 -1317 -12032
rect -1393 -12082 -1377 -12048
rect -1333 -12082 -1317 -12048
rect -1393 -12088 -1317 -12082
rect -1284 -12120 -1250 -11581
rect -1194 -11919 -1160 -11488
rect -1213 -11972 -1203 -11919
rect -1150 -11972 -1140 -11919
rect -1194 -12032 -1160 -11972
rect -1215 -12048 -1139 -12032
rect -1215 -12082 -1199 -12048
rect -1155 -12082 -1139 -12048
rect -1215 -12088 -1139 -12082
rect -1105 -12120 -1071 -11400
rect -1037 -11438 -961 -11432
rect -1037 -11472 -1021 -11438
rect -977 -11472 -961 -11438
rect -1037 -11488 -961 -11472
rect -1016 -11919 -982 -11488
rect -927 -11528 -893 -11400
rect -859 -11438 -783 -11432
rect -859 -11472 -843 -11438
rect -799 -11472 -783 -11438
rect -859 -11488 -783 -11472
rect -947 -11581 -937 -11528
rect -884 -11581 -874 -11528
rect -838 -11919 -804 -11488
rect -1035 -11972 -1025 -11919
rect -972 -11972 -962 -11919
rect -858 -11972 -848 -11919
rect -795 -11972 -785 -11919
rect -1016 -12032 -982 -11972
rect -838 -12032 -804 -11972
rect -1037 -12048 -961 -12032
rect -1037 -12082 -1021 -12048
rect -977 -12082 -961 -12048
rect -1037 -12088 -961 -12082
rect -859 -12048 -783 -12032
rect -859 -12082 -843 -12048
rect -799 -12082 -783 -12048
rect -859 -12088 -783 -12082
rect -749 -12120 -715 -11400
rect -681 -11438 -605 -11432
rect -681 -11472 -665 -11438
rect -621 -11472 -605 -11438
rect -681 -11488 -605 -11472
rect -660 -11919 -626 -11488
rect -571 -11637 -537 -11400
rect -503 -11438 -427 -11432
rect -503 -11472 -487 -11438
rect -443 -11472 -427 -11438
rect -503 -11488 -427 -11472
rect -590 -11690 -580 -11637
rect -527 -11690 -517 -11637
rect -482 -11919 -448 -11488
rect -680 -11972 -670 -11919
rect -617 -11972 -607 -11919
rect -502 -11972 -492 -11919
rect -439 -11972 -429 -11919
rect -660 -12032 -626 -11972
rect -482 -12032 -448 -11972
rect -681 -12048 -605 -12032
rect -681 -12082 -665 -12048
rect -621 -12082 -605 -12048
rect -681 -12088 -605 -12082
rect -503 -12048 -427 -12032
rect -503 -12082 -487 -12048
rect -443 -12082 -427 -12048
rect -503 -12088 -427 -12082
rect -393 -12120 -359 -11400
rect -325 -11438 -249 -11432
rect -325 -11472 -309 -11438
rect -265 -11472 -249 -11438
rect -325 -11488 -249 -11472
rect -304 -11919 -270 -11488
rect -215 -11757 -181 -11400
rect -147 -11438 -71 -11432
rect -147 -11472 -131 -11438
rect -87 -11472 -71 -11438
rect -147 -11488 -71 -11472
rect -234 -11810 -224 -11757
rect -171 -11810 -161 -11757
rect -324 -11972 -314 -11919
rect -261 -11972 -251 -11919
rect -304 -12032 -270 -11972
rect -325 -12048 -249 -12032
rect -325 -12082 -309 -12048
rect -265 -12082 -249 -12048
rect -325 -12088 -249 -12082
rect -215 -12120 -181 -11810
rect -126 -11919 -92 -11488
rect -146 -11972 -136 -11919
rect -83 -11972 -73 -11919
rect -126 -12032 -92 -11972
rect -147 -12048 -71 -12032
rect -147 -12082 -131 -12048
rect -87 -12082 -71 -12048
rect -147 -12088 -71 -12082
rect -36 -12120 -2 -11400
rect 31 -11438 107 -11432
rect 31 -11472 47 -11438
rect 91 -11472 107 -11438
rect 31 -11488 107 -11472
rect 52 -11919 86 -11488
rect 141 -11757 175 -11400
rect 209 -11438 285 -11432
rect 209 -11472 225 -11438
rect 269 -11472 285 -11438
rect 209 -11488 285 -11472
rect 121 -11810 131 -11757
rect 184 -11810 194 -11757
rect 141 -11811 175 -11810
rect 230 -11919 264 -11488
rect 32 -11972 42 -11919
rect 95 -11972 105 -11919
rect 210 -11972 220 -11919
rect 273 -11972 283 -11919
rect 52 -12032 86 -11972
rect 230 -12032 264 -11972
rect 31 -12048 107 -12032
rect 31 -12082 47 -12048
rect 91 -12082 107 -12048
rect 31 -12088 107 -12082
rect 209 -12048 285 -12032
rect 209 -12082 225 -12048
rect 269 -12082 285 -12048
rect 209 -12088 285 -12082
rect 319 -12120 353 -11400
rect 387 -11438 463 -11432
rect 387 -11472 403 -11438
rect 447 -11472 463 -11438
rect 387 -11488 463 -11472
rect 408 -11919 442 -11488
rect 497 -11757 531 -11400
rect 565 -11438 641 -11432
rect 565 -11472 581 -11438
rect 625 -11472 641 -11438
rect 565 -11488 641 -11472
rect 477 -11810 487 -11757
rect 540 -11810 550 -11757
rect 389 -11972 399 -11919
rect 452 -11972 462 -11919
rect 408 -12032 442 -11972
rect 387 -12048 463 -12032
rect 387 -12082 403 -12048
rect 447 -12082 463 -12048
rect 387 -12088 463 -12082
rect 496 -12120 530 -11810
rect 586 -11919 620 -11488
rect 567 -11972 577 -11919
rect 630 -11972 640 -11919
rect 586 -12032 620 -11972
rect 565 -12048 641 -12032
rect 565 -12082 581 -12048
rect 625 -12082 641 -12048
rect 565 -12088 641 -12082
rect 675 -12120 709 -11400
rect 743 -11438 819 -11432
rect 853 -11438 887 -11400
rect 921 -11438 997 -11432
rect 1031 -11438 1065 -11400
rect 1099 -11438 1175 -11432
rect 743 -11472 759 -11438
rect 803 -11472 937 -11438
rect 981 -11472 1115 -11438
rect 1159 -11472 1175 -11438
rect 743 -11488 819 -11472
rect 921 -11488 997 -11472
rect 1099 -11488 1175 -11472
rect 942 -12032 976 -11488
rect 743 -12048 819 -12032
rect 743 -12082 759 -12048
rect 803 -12082 819 -12048
rect 743 -12088 819 -12082
rect 921 -12048 997 -12032
rect 921 -12082 937 -12048
rect 981 -12082 997 -12048
rect 921 -12088 997 -12082
rect 1099 -12048 1175 -12032
rect 1099 -12082 1115 -12048
rect 1159 -12082 1175 -12048
rect 1099 -12088 1175 -12082
rect 1209 -12120 1243 -11400
rect 1277 -11438 1353 -11432
rect 1277 -11472 1293 -11438
rect 1337 -11472 1353 -11438
rect 1277 -11488 1353 -11472
rect 1298 -11919 1332 -11488
rect 1387 -11528 1421 -11400
rect 1455 -11438 1531 -11432
rect 1455 -11472 1471 -11438
rect 1515 -11472 1531 -11438
rect 1455 -11488 1531 -11472
rect 1367 -11581 1377 -11528
rect 1430 -11581 1440 -11528
rect 1477 -11919 1511 -11488
rect 1278 -11972 1288 -11919
rect 1341 -11972 1351 -11919
rect 1458 -11972 1468 -11919
rect 1521 -11972 1531 -11919
rect 1298 -12032 1332 -11972
rect 1477 -12032 1511 -11972
rect 1277 -12048 1353 -12032
rect 1277 -12082 1293 -12048
rect 1337 -12082 1353 -12048
rect 1277 -12088 1353 -12082
rect 1455 -12048 1531 -12032
rect 1455 -12082 1471 -12048
rect 1515 -12082 1531 -12048
rect 1455 -12088 1531 -12082
rect 1566 -12120 1600 -11400
rect 1633 -11438 1709 -11432
rect 1633 -11472 1649 -11438
rect 1693 -11472 1709 -11438
rect 1633 -11488 1709 -11472
rect 1654 -11920 1688 -11488
rect 1743 -11528 1777 -11400
rect 1811 -11438 1887 -11432
rect 1811 -11472 1827 -11438
rect 1871 -11472 1887 -11438
rect 1811 -11488 1887 -11472
rect 1723 -11581 1733 -11528
rect 1786 -11581 1796 -11528
rect 1634 -11973 1644 -11920
rect 1697 -11973 1707 -11920
rect 1654 -12032 1688 -11973
rect 1633 -12048 1709 -12032
rect 1633 -12082 1649 -12048
rect 1693 -12082 1709 -12048
rect 1633 -12088 1709 -12082
rect 1744 -12120 1778 -11581
rect 1832 -11919 1866 -11488
rect 1813 -11972 1823 -11919
rect 1876 -11972 1886 -11919
rect 1832 -12032 1866 -11972
rect 1811 -12048 1887 -12032
rect 1811 -12082 1827 -12048
rect 1871 -12082 1887 -12048
rect 1811 -12088 1887 -12082
rect 1922 -12120 1956 -11400
rect 1989 -11438 2065 -11432
rect 1989 -11472 2005 -11438
rect 2049 -11472 2065 -11438
rect 1989 -11488 2065 -11472
rect 2010 -11919 2044 -11488
rect 2099 -11528 2133 -11400
rect 2167 -11438 2243 -11432
rect 2167 -11472 2183 -11438
rect 2227 -11472 2243 -11438
rect 2167 -11488 2243 -11472
rect 2079 -11581 2089 -11528
rect 2142 -11581 2152 -11528
rect 2188 -11919 2222 -11488
rect 1990 -11972 2000 -11919
rect 2053 -11972 2063 -11919
rect 2168 -11972 2178 -11919
rect 2231 -11972 2241 -11919
rect 2010 -12032 2044 -11972
rect 2188 -12032 2222 -11972
rect 1989 -12048 2065 -12032
rect 1989 -12082 2005 -12048
rect 2049 -12082 2065 -12048
rect 1989 -12088 2065 -12082
rect 2167 -12048 2243 -12032
rect 2167 -12082 2183 -12048
rect 2227 -12082 2243 -12048
rect 2167 -12088 2243 -12082
rect 2277 -12120 2311 -11400
rect 2345 -11438 2421 -11432
rect 2345 -11472 2361 -11438
rect 2405 -11472 2421 -11438
rect 2345 -11488 2421 -11472
rect 2366 -11919 2400 -11488
rect 2456 -11637 2490 -11400
rect 2523 -11438 2599 -11432
rect 2523 -11472 2539 -11438
rect 2583 -11472 2599 -11438
rect 2523 -11488 2599 -11472
rect 2436 -11690 2446 -11637
rect 2499 -11690 2509 -11637
rect 2544 -11919 2578 -11488
rect 2347 -11972 2357 -11919
rect 2410 -11972 2420 -11919
rect 2524 -11972 2534 -11919
rect 2587 -11972 2597 -11919
rect 2366 -12032 2400 -11972
rect 2544 -12032 2578 -11972
rect 2345 -12048 2421 -12032
rect 2345 -12082 2361 -12048
rect 2405 -12082 2421 -12048
rect 2345 -12088 2421 -12082
rect 2523 -12048 2599 -12032
rect 2523 -12082 2539 -12048
rect 2583 -12082 2599 -12048
rect 2523 -12088 2599 -12082
rect 2633 -12120 2667 -11400
rect 2701 -11438 2777 -11432
rect 2701 -11472 2717 -11438
rect 2761 -11472 2777 -11438
rect 2701 -11488 2777 -11472
rect 2722 -11919 2756 -11488
rect 2810 -11757 2844 -11400
rect 2879 -11438 2955 -11432
rect 2879 -11472 2895 -11438
rect 2939 -11472 2955 -11438
rect 2879 -11488 2955 -11472
rect 2790 -11810 2800 -11757
rect 2853 -11810 2863 -11757
rect 2703 -11972 2713 -11919
rect 2766 -11972 2776 -11919
rect 2722 -12032 2756 -11972
rect 2701 -12048 2777 -12032
rect 2701 -12082 2717 -12048
rect 2761 -12082 2777 -12048
rect 2701 -12088 2777 -12082
rect 2811 -12120 2845 -11810
rect 2900 -11919 2934 -11488
rect 2880 -11972 2890 -11919
rect 2943 -11972 2953 -11919
rect 2900 -12032 2934 -11972
rect 2879 -12048 2955 -12032
rect 2879 -12082 2895 -12048
rect 2939 -12082 2955 -12048
rect 2879 -12088 2955 -12082
rect 2989 -12120 3023 -11400
rect 3057 -11438 3133 -11432
rect 3057 -11472 3073 -11438
rect 3117 -11472 3133 -11438
rect 3057 -11488 3133 -11472
rect 3078 -11919 3112 -11488
rect 3166 -11757 3200 -11400
rect 3235 -11438 3311 -11432
rect 3235 -11472 3251 -11438
rect 3295 -11472 3311 -11438
rect 3235 -11488 3311 -11472
rect 3147 -11810 3157 -11757
rect 3210 -11810 3220 -11757
rect 3256 -11919 3290 -11488
rect 3058 -11972 3068 -11919
rect 3121 -11972 3131 -11919
rect 3237 -11972 3247 -11919
rect 3300 -11972 3310 -11919
rect 3078 -12032 3112 -11972
rect 3256 -12032 3290 -11972
rect 3057 -12048 3133 -12032
rect 3057 -12082 3073 -12048
rect 3117 -12082 3133 -12048
rect 3057 -12088 3133 -12082
rect 3235 -12048 3311 -12032
rect 3235 -12082 3251 -12048
rect 3295 -12082 3311 -12048
rect 3235 -12088 3311 -12082
rect 3345 -12120 3379 -11400
rect 3413 -11438 3489 -11432
rect 3413 -11472 3429 -11438
rect 3473 -11472 3489 -11438
rect 3413 -11488 3489 -11472
rect 3434 -11919 3468 -11488
rect 3522 -11757 3556 -11400
rect 3591 -11438 3667 -11432
rect 3591 -11472 3607 -11438
rect 3651 -11472 3667 -11438
rect 3591 -11488 3667 -11472
rect 3503 -11810 3513 -11757
rect 3566 -11810 3576 -11757
rect 3612 -11919 3646 -11488
rect 3415 -11972 3425 -11919
rect 3478 -11972 3488 -11919
rect 3593 -11972 3603 -11919
rect 3656 -11972 3666 -11919
rect 3434 -12032 3468 -11972
rect 3612 -12032 3646 -11972
rect 3413 -12048 3489 -12032
rect 3413 -12082 3429 -12048
rect 3473 -12082 3489 -12048
rect 3413 -12088 3489 -12082
rect 3591 -12048 3667 -12032
rect 3591 -12082 3607 -12048
rect 3651 -12082 3667 -12048
rect 3591 -12088 3667 -12082
rect 3701 -12120 3735 -11400
rect 3769 -11438 3845 -11432
rect 3769 -11472 3785 -11438
rect 3829 -11472 3845 -11438
rect 3769 -11488 3845 -11472
rect 3881 -11437 3915 -11400
rect 3947 -11437 4023 -11432
rect 4056 -11437 4090 -11400
rect 3881 -11438 4090 -11437
rect 3881 -11471 3963 -11438
rect 3790 -11919 3824 -11488
rect 3881 -11638 3915 -11471
rect 3947 -11472 3963 -11471
rect 4007 -11471 4090 -11438
rect 4007 -11472 4023 -11471
rect 3947 -11488 4023 -11472
rect 3861 -11691 3871 -11638
rect 3924 -11691 3934 -11638
rect 3771 -11972 3781 -11919
rect 3834 -11972 3844 -11919
rect 3790 -12032 3824 -11972
rect 3769 -12048 3845 -12032
rect 3769 -12082 3785 -12048
rect 3829 -12082 3845 -12048
rect 3769 -12088 3845 -12082
rect 3881 -12120 3915 -11691
rect 3947 -12048 4023 -12032
rect 3947 -12082 3963 -12048
rect 4007 -12082 4023 -12048
rect 3947 -12088 4023 -12082
rect -2179 -12132 -2133 -12120
rect -2179 -12388 -2173 -12132
rect -2139 -12388 -2133 -12132
rect -2179 -12400 -2133 -12388
rect -2001 -12132 -1955 -12120
rect -2001 -12388 -1995 -12132
rect -1961 -12388 -1955 -12132
rect -2001 -12400 -1955 -12388
rect -1823 -12132 -1777 -12120
rect -1823 -12388 -1817 -12132
rect -1783 -12388 -1777 -12132
rect -1823 -12400 -1777 -12388
rect -1645 -12132 -1599 -12120
rect -1645 -12388 -1639 -12132
rect -1605 -12388 -1599 -12132
rect -1645 -12400 -1599 -12388
rect -1467 -12132 -1421 -12120
rect -1467 -12388 -1461 -12132
rect -1427 -12388 -1421 -12132
rect -1467 -12400 -1421 -12388
rect -1289 -12132 -1243 -12120
rect -1289 -12388 -1283 -12132
rect -1249 -12388 -1243 -12132
rect -1289 -12400 -1243 -12388
rect -1111 -12132 -1065 -12120
rect -1111 -12388 -1105 -12132
rect -1071 -12388 -1065 -12132
rect -1111 -12400 -1065 -12388
rect -933 -12132 -887 -12120
rect -933 -12388 -927 -12132
rect -893 -12388 -887 -12132
rect -933 -12400 -887 -12388
rect -755 -12132 -709 -12120
rect -755 -12388 -749 -12132
rect -715 -12388 -709 -12132
rect -755 -12400 -709 -12388
rect -577 -12132 -531 -12120
rect -577 -12388 -571 -12132
rect -537 -12388 -531 -12132
rect -577 -12400 -531 -12388
rect -399 -12132 -353 -12120
rect -399 -12388 -393 -12132
rect -359 -12388 -353 -12132
rect -399 -12400 -353 -12388
rect -221 -12132 -175 -12120
rect -221 -12388 -215 -12132
rect -181 -12388 -175 -12132
rect -221 -12400 -175 -12388
rect -43 -12132 3 -12120
rect -43 -12388 -37 -12132
rect -3 -12388 3 -12132
rect -43 -12400 3 -12388
rect 135 -12132 181 -12120
rect 135 -12388 141 -12132
rect 175 -12388 181 -12132
rect 135 -12400 181 -12388
rect 313 -12132 359 -12120
rect 313 -12388 319 -12132
rect 353 -12388 359 -12132
rect 313 -12400 359 -12388
rect 491 -12132 537 -12120
rect 491 -12388 497 -12132
rect 531 -12388 537 -12132
rect 491 -12400 537 -12388
rect 669 -12132 715 -12120
rect 669 -12388 675 -12132
rect 709 -12388 715 -12132
rect 669 -12400 715 -12388
rect 847 -12132 893 -12120
rect 847 -12388 853 -12132
rect 887 -12388 893 -12132
rect 847 -12400 893 -12388
rect 1025 -12132 1071 -12120
rect 1025 -12388 1031 -12132
rect 1065 -12388 1071 -12132
rect 1025 -12400 1071 -12388
rect 1203 -12132 1249 -12120
rect 1203 -12388 1209 -12132
rect 1243 -12388 1249 -12132
rect 1203 -12400 1249 -12388
rect 1381 -12132 1427 -12120
rect 1381 -12388 1387 -12132
rect 1421 -12388 1427 -12132
rect 1381 -12400 1427 -12388
rect 1559 -12132 1605 -12120
rect 1559 -12388 1565 -12132
rect 1599 -12388 1605 -12132
rect 1559 -12400 1605 -12388
rect 1737 -12132 1783 -12120
rect 1737 -12388 1743 -12132
rect 1777 -12388 1783 -12132
rect 1737 -12400 1783 -12388
rect 1915 -12132 1961 -12120
rect 1915 -12388 1921 -12132
rect 1955 -12388 1961 -12132
rect 1915 -12400 1961 -12388
rect 2093 -12132 2139 -12120
rect 2093 -12388 2099 -12132
rect 2133 -12388 2139 -12132
rect 2093 -12400 2139 -12388
rect 2271 -12132 2317 -12120
rect 2271 -12388 2277 -12132
rect 2311 -12388 2317 -12132
rect 2271 -12400 2317 -12388
rect 2449 -12132 2495 -12120
rect 2449 -12388 2455 -12132
rect 2489 -12388 2495 -12132
rect 2449 -12400 2495 -12388
rect 2627 -12132 2673 -12120
rect 2627 -12388 2633 -12132
rect 2667 -12388 2673 -12132
rect 2627 -12400 2673 -12388
rect 2805 -12132 2851 -12120
rect 2805 -12388 2811 -12132
rect 2845 -12388 2851 -12132
rect 2805 -12400 2851 -12388
rect 2983 -12132 3029 -12120
rect 2983 -12388 2989 -12132
rect 3023 -12388 3029 -12132
rect 2983 -12400 3029 -12388
rect 3161 -12132 3207 -12120
rect 3161 -12388 3167 -12132
rect 3201 -12388 3207 -12132
rect 3161 -12400 3207 -12388
rect 3339 -12132 3385 -12120
rect 3339 -12388 3345 -12132
rect 3379 -12388 3385 -12132
rect 3339 -12400 3385 -12388
rect 3517 -12132 3563 -12120
rect 3517 -12388 3523 -12132
rect 3557 -12388 3563 -12132
rect 3517 -12400 3563 -12388
rect 3695 -12132 3741 -12120
rect 3695 -12388 3701 -12132
rect 3735 -12388 3741 -12132
rect 3695 -12400 3741 -12388
rect 3873 -12132 3919 -12120
rect 3873 -12388 3879 -12132
rect 3913 -12388 3919 -12132
rect 3873 -12400 3919 -12388
rect 4051 -12132 4097 -12120
rect 4051 -12388 4057 -12132
rect 4091 -12388 4097 -12132
rect 4051 -12400 4097 -12388
rect -2105 -12438 -2029 -12432
rect -2105 -12472 -2089 -12438
rect -2045 -12472 -2029 -12438
rect -2105 -12488 -2029 -12472
rect -1995 -12542 -1961 -12400
rect -1927 -12438 -1851 -12432
rect -1927 -12472 -1911 -12438
rect -1867 -12472 -1851 -12438
rect -1927 -12488 -1851 -12472
rect -2015 -12595 -2005 -12542
rect -1952 -12595 -1942 -12542
rect -2105 -13046 -2029 -13032
rect -1995 -13046 -1961 -12595
rect -1906 -13032 -1872 -12488
rect -2174 -13048 -1961 -13046
rect -2174 -13080 -2089 -13048
rect -2174 -13120 -2140 -13080
rect -2105 -13082 -2089 -13080
rect -2045 -13080 -1961 -13048
rect -2045 -13082 -2029 -13080
rect -2105 -13088 -2029 -13082
rect -1995 -13120 -1961 -13080
rect -1927 -13048 -1851 -13032
rect -1927 -13082 -1911 -13048
rect -1867 -13082 -1851 -13048
rect -1927 -13088 -1851 -13082
rect -1818 -13120 -1784 -12400
rect -1749 -12438 -1673 -12432
rect -1749 -12472 -1733 -12438
rect -1689 -12472 -1673 -12438
rect -1749 -12488 -1673 -12472
rect -1728 -13032 -1694 -12488
rect -1639 -12542 -1605 -12400
rect -1571 -12438 -1495 -12432
rect -1571 -12472 -1555 -12438
rect -1511 -12472 -1495 -12438
rect -1571 -12488 -1495 -12472
rect -1659 -12595 -1649 -12542
rect -1596 -12595 -1586 -12542
rect -1549 -13032 -1515 -12488
rect -1749 -13048 -1673 -13032
rect -1749 -13082 -1733 -13048
rect -1689 -13082 -1673 -13048
rect -1749 -13088 -1673 -13082
rect -1571 -13048 -1495 -13032
rect -1571 -13082 -1555 -13048
rect -1511 -13082 -1495 -13048
rect -1571 -13088 -1495 -13082
rect -1461 -13120 -1427 -12400
rect -1393 -12438 -1317 -12432
rect -1393 -12472 -1377 -12438
rect -1333 -12472 -1317 -12438
rect -1393 -12488 -1317 -12472
rect -1372 -13032 -1338 -12488
rect -1284 -12654 -1250 -12400
rect -1215 -12438 -1139 -12432
rect -1215 -12472 -1199 -12438
rect -1155 -12472 -1139 -12438
rect -1215 -12488 -1139 -12472
rect -1304 -12707 -1294 -12654
rect -1241 -12707 -1231 -12654
rect -1194 -13032 -1160 -12488
rect -1393 -13048 -1317 -13032
rect -1393 -13082 -1377 -13048
rect -1333 -13082 -1317 -13048
rect -1393 -13088 -1317 -13082
rect -1215 -13048 -1139 -13032
rect -1215 -13082 -1199 -13048
rect -1155 -13082 -1139 -13048
rect -1215 -13088 -1139 -13082
rect -1105 -13120 -1071 -12400
rect -1037 -12438 -961 -12432
rect -1037 -12472 -1021 -12438
rect -977 -12472 -961 -12438
rect -1037 -12488 -961 -12472
rect -1016 -13032 -982 -12488
rect -927 -12783 -893 -12400
rect -859 -12438 -783 -12432
rect -859 -12472 -843 -12438
rect -799 -12472 -783 -12438
rect -859 -12488 -783 -12472
rect -947 -12836 -937 -12783
rect -884 -12836 -874 -12783
rect -1037 -13048 -961 -13032
rect -1037 -13082 -1021 -13048
rect -977 -13082 -961 -13048
rect -1037 -13088 -961 -13082
rect -927 -13120 -893 -12836
rect -838 -13032 -804 -12488
rect -859 -13048 -783 -13032
rect -859 -13082 -843 -13048
rect -799 -13082 -783 -13048
rect -859 -13088 -783 -13082
rect -749 -13120 -715 -12400
rect -681 -12438 -605 -12432
rect -681 -12472 -665 -12438
rect -621 -12472 -605 -12438
rect -681 -12488 -605 -12472
rect -660 -13032 -626 -12488
rect -571 -12653 -537 -12400
rect -503 -12438 -427 -12432
rect -503 -12472 -487 -12438
rect -443 -12472 -427 -12438
rect -503 -12488 -427 -12472
rect -592 -12706 -582 -12653
rect -529 -12706 -519 -12653
rect -482 -13032 -448 -12488
rect -681 -13048 -605 -13032
rect -681 -13082 -665 -13048
rect -621 -13082 -605 -13048
rect -681 -13088 -605 -13082
rect -503 -13048 -427 -13032
rect -503 -13082 -487 -13048
rect -443 -13082 -427 -13048
rect -503 -13088 -427 -13082
rect -393 -13120 -359 -12400
rect -325 -12438 -249 -12432
rect -325 -12472 -309 -12438
rect -265 -12472 -249 -12438
rect -325 -12488 -249 -12472
rect -304 -13032 -270 -12488
rect -215 -12783 -181 -12400
rect -147 -12438 -71 -12432
rect -147 -12472 -131 -12438
rect -87 -12472 -71 -12438
rect -147 -12488 -71 -12472
rect -234 -12836 -224 -12783
rect -171 -12836 -161 -12783
rect -126 -13032 -92 -12488
rect -325 -13048 -249 -13032
rect -325 -13082 -309 -13048
rect -265 -13082 -249 -13048
rect -325 -13088 -249 -13082
rect -147 -13048 -71 -13032
rect -147 -13082 -131 -13048
rect -87 -13082 -71 -13048
rect -147 -13088 -71 -13082
rect -36 -13120 -2 -12400
rect 31 -12438 107 -12432
rect 31 -12472 47 -12438
rect 91 -12472 107 -12438
rect 31 -12488 107 -12472
rect 52 -13032 86 -12488
rect 141 -12653 175 -12400
rect 209 -12438 285 -12432
rect 209 -12472 225 -12438
rect 269 -12472 285 -12438
rect 209 -12488 285 -12472
rect 120 -12706 130 -12653
rect 183 -12706 193 -12653
rect 31 -13048 107 -13032
rect 31 -13082 47 -13048
rect 91 -13082 107 -13048
rect 31 -13088 107 -13082
rect 141 -13120 175 -12706
rect 230 -13032 264 -12488
rect 209 -13048 285 -13032
rect 209 -13082 225 -13048
rect 269 -13082 285 -13048
rect 209 -13088 285 -13082
rect 319 -13120 353 -12400
rect 387 -12438 463 -12432
rect 387 -12472 403 -12438
rect 447 -12472 463 -12438
rect 387 -12488 463 -12472
rect 408 -13032 442 -12488
rect 496 -12784 530 -12400
rect 565 -12438 641 -12432
rect 565 -12472 581 -12438
rect 625 -12472 641 -12438
rect 565 -12488 641 -12472
rect 476 -12837 486 -12784
rect 539 -12837 549 -12784
rect 587 -13032 621 -12488
rect 387 -13048 463 -13032
rect 387 -13082 403 -13048
rect 447 -13082 463 -13048
rect 387 -13088 463 -13082
rect 565 -13048 641 -13032
rect 565 -13082 581 -13048
rect 625 -13082 641 -13048
rect 565 -13088 641 -13082
rect 675 -13120 709 -12400
rect 743 -12438 819 -12432
rect 852 -12438 886 -12400
rect 921 -12438 997 -12432
rect 1031 -12438 1065 -12400
rect 1099 -12438 1175 -12432
rect 743 -12472 759 -12438
rect 803 -12472 937 -12438
rect 981 -12472 1115 -12438
rect 1159 -12472 1175 -12438
rect 743 -12488 819 -12472
rect 921 -12488 997 -12472
rect 1099 -12488 1175 -12472
rect 942 -13032 976 -12488
rect 743 -13048 819 -13032
rect 921 -13048 997 -13032
rect 1099 -13048 1175 -13032
rect 743 -13082 759 -13048
rect 803 -13082 937 -13048
rect 981 -13082 1115 -13048
rect 1159 -13082 1175 -13048
rect 743 -13088 819 -13082
rect 852 -13120 886 -13082
rect 921 -13088 997 -13082
rect 1032 -13120 1066 -13082
rect 1099 -13088 1175 -13082
rect 1209 -13120 1243 -12400
rect 1277 -12438 1353 -12432
rect 1277 -12472 1293 -12438
rect 1337 -12472 1353 -12438
rect 1277 -12488 1353 -12472
rect 1299 -13032 1333 -12488
rect 1388 -12783 1422 -12400
rect 1455 -12438 1531 -12432
rect 1455 -12472 1471 -12438
rect 1515 -12472 1531 -12438
rect 1455 -12488 1531 -12472
rect 1368 -12836 1378 -12783
rect 1431 -12836 1441 -12783
rect 1277 -13048 1353 -13032
rect 1277 -13082 1293 -13048
rect 1337 -13082 1353 -13048
rect 1277 -13088 1353 -13082
rect 1388 -13120 1422 -12836
rect 1476 -13032 1510 -12488
rect 1455 -13048 1531 -13032
rect 1455 -13082 1471 -13048
rect 1515 -13082 1531 -13048
rect 1455 -13088 1531 -13082
rect 1566 -13120 1600 -12400
rect 1633 -12438 1709 -12432
rect 1633 -12472 1649 -12438
rect 1693 -12472 1709 -12438
rect 1633 -12488 1709 -12472
rect 1655 -13032 1689 -12488
rect 1744 -12654 1778 -12400
rect 1811 -12438 1887 -12432
rect 1811 -12472 1827 -12438
rect 1871 -12472 1887 -12438
rect 1811 -12488 1887 -12472
rect 1725 -12707 1735 -12654
rect 1788 -12707 1798 -12654
rect 1833 -13032 1867 -12488
rect 1633 -13048 1709 -13032
rect 1633 -13082 1649 -13048
rect 1693 -13082 1709 -13048
rect 1633 -13088 1709 -13082
rect 1811 -13048 1887 -13032
rect 1811 -13082 1827 -13048
rect 1871 -13082 1887 -13048
rect 1811 -13088 1887 -13082
rect 1922 -13120 1956 -12400
rect 1989 -12438 2065 -12432
rect 1989 -12472 2005 -12438
rect 2049 -12472 2065 -12438
rect 1989 -12488 2065 -12472
rect 2009 -13032 2043 -12488
rect 2098 -12782 2132 -12400
rect 2167 -12438 2243 -12432
rect 2167 -12472 2183 -12438
rect 2227 -12472 2243 -12438
rect 2167 -12488 2243 -12472
rect 2078 -12835 2088 -12782
rect 2141 -12835 2151 -12782
rect 1989 -13048 2065 -13032
rect 1989 -13082 2005 -13048
rect 2049 -13082 2065 -13048
rect 1989 -13088 2065 -13082
rect 2098 -13120 2132 -12835
rect 2188 -13032 2222 -12488
rect 2167 -13048 2243 -13032
rect 2167 -13082 2183 -13048
rect 2227 -13082 2243 -13048
rect 2167 -13088 2243 -13082
rect 2277 -13120 2311 -12400
rect 2345 -12438 2421 -12432
rect 2345 -12472 2361 -12438
rect 2405 -12472 2421 -12438
rect 2345 -12488 2421 -12472
rect 2366 -13032 2400 -12488
rect 2455 -12653 2489 -12400
rect 2523 -12438 2599 -12432
rect 2523 -12472 2539 -12438
rect 2583 -12472 2599 -12438
rect 2523 -12488 2599 -12472
rect 2435 -12706 2445 -12653
rect 2498 -12706 2508 -12653
rect 2544 -13032 2578 -12488
rect 2345 -13048 2421 -13032
rect 2345 -13082 2361 -13048
rect 2405 -13082 2421 -13048
rect 2345 -13088 2421 -13082
rect 2523 -13048 2599 -13032
rect 2523 -13082 2539 -13048
rect 2583 -13082 2599 -13048
rect 2523 -13088 2599 -13082
rect 2633 -13120 2667 -12400
rect 2701 -12438 2777 -12432
rect 2701 -12472 2717 -12438
rect 2761 -12472 2777 -12438
rect 2701 -12488 2777 -12472
rect 2722 -13032 2756 -12488
rect 2811 -12782 2845 -12400
rect 2879 -12438 2955 -12432
rect 2879 -12472 2895 -12438
rect 2939 -12472 2955 -12438
rect 2879 -12488 2955 -12472
rect 2791 -12835 2801 -12782
rect 2854 -12835 2864 -12782
rect 2900 -13032 2934 -12488
rect 2701 -13048 2777 -13032
rect 2701 -13082 2717 -13048
rect 2761 -13082 2777 -13048
rect 2701 -13088 2777 -13082
rect 2879 -13048 2955 -13032
rect 2879 -13082 2895 -13048
rect 2939 -13082 2955 -13048
rect 2879 -13088 2955 -13082
rect 2989 -13120 3023 -12400
rect 3057 -12438 3133 -12432
rect 3057 -12472 3073 -12438
rect 3117 -12472 3133 -12438
rect 3057 -12488 3133 -12472
rect 3078 -13032 3112 -12488
rect 3167 -12650 3201 -12400
rect 3235 -12438 3311 -12432
rect 3235 -12472 3251 -12438
rect 3295 -12472 3311 -12438
rect 3235 -12488 3311 -12472
rect 3166 -12652 3201 -12650
rect 3148 -12705 3158 -12652
rect 3211 -12705 3221 -12652
rect 3057 -13048 3133 -13032
rect 3057 -13082 3073 -13048
rect 3117 -13082 3133 -13048
rect 3057 -13088 3133 -13082
rect 3166 -13120 3200 -12705
rect 3256 -13032 3290 -12488
rect 3235 -13048 3311 -13032
rect 3235 -13082 3251 -13048
rect 3295 -13082 3311 -13048
rect 3235 -13088 3311 -13082
rect 3345 -13120 3379 -12400
rect 3413 -12438 3489 -12432
rect 3413 -12472 3429 -12438
rect 3473 -12472 3489 -12438
rect 3413 -12488 3489 -12472
rect 3434 -13032 3468 -12488
rect 3524 -12542 3558 -12400
rect 3591 -12438 3667 -12432
rect 3591 -12472 3607 -12438
rect 3651 -12472 3667 -12438
rect 3591 -12488 3667 -12472
rect 3504 -12595 3514 -12542
rect 3567 -12595 3577 -12542
rect 3613 -13032 3647 -12488
rect 3413 -13048 3489 -13032
rect 3413 -13082 3429 -13048
rect 3473 -13082 3489 -13048
rect 3413 -13088 3489 -13082
rect 3591 -13048 3667 -13032
rect 3591 -13082 3607 -13048
rect 3651 -13082 3667 -13048
rect 3591 -13088 3667 -13082
rect 3701 -13120 3735 -12400
rect 3769 -12438 3845 -12432
rect 3769 -12472 3785 -12438
rect 3829 -12472 3845 -12438
rect 3769 -12488 3845 -12472
rect 3881 -12436 3915 -12400
rect 3947 -12436 4023 -12432
rect 4058 -12436 4092 -12400
rect 3881 -12438 4092 -12436
rect 3881 -12470 3963 -12438
rect 3790 -13032 3824 -12488
rect 3881 -12542 3915 -12470
rect 3947 -12472 3963 -12470
rect 4007 -12470 4092 -12438
rect 4007 -12472 4023 -12470
rect 3947 -12488 4023 -12472
rect 3861 -12595 3871 -12542
rect 3924 -12595 3934 -12542
rect 3769 -13048 3845 -13032
rect 3769 -13082 3785 -13048
rect 3829 -13082 3845 -13048
rect 3769 -13088 3845 -13082
rect 3881 -13047 3915 -12595
rect 3947 -13047 4023 -13032
rect 3881 -13048 4090 -13047
rect 3881 -13081 3963 -13048
rect 3881 -13120 3915 -13081
rect 3947 -13082 3963 -13081
rect 4007 -13081 4090 -13048
rect 4007 -13082 4023 -13081
rect 3947 -13088 4023 -13082
rect 4056 -13120 4090 -13081
rect -2179 -13132 -2133 -13120
rect -2179 -13388 -2173 -13132
rect -2139 -13388 -2133 -13132
rect -2179 -13400 -2133 -13388
rect -2001 -13132 -1955 -13120
rect -2001 -13388 -1995 -13132
rect -1961 -13388 -1955 -13132
rect -2001 -13400 -1955 -13388
rect -1823 -13132 -1777 -13120
rect -1823 -13388 -1817 -13132
rect -1783 -13388 -1777 -13132
rect -1823 -13400 -1777 -13388
rect -1645 -13132 -1599 -13120
rect -1645 -13388 -1639 -13132
rect -1605 -13388 -1599 -13132
rect -1645 -13400 -1599 -13388
rect -1467 -13132 -1421 -13120
rect -1467 -13388 -1461 -13132
rect -1427 -13388 -1421 -13132
rect -1467 -13400 -1421 -13388
rect -1289 -13132 -1243 -13120
rect -1289 -13388 -1283 -13132
rect -1249 -13388 -1243 -13132
rect -1289 -13400 -1243 -13388
rect -1111 -13132 -1065 -13120
rect -1111 -13388 -1105 -13132
rect -1071 -13388 -1065 -13132
rect -1111 -13400 -1065 -13388
rect -933 -13132 -887 -13120
rect -933 -13388 -927 -13132
rect -893 -13388 -887 -13132
rect -933 -13400 -887 -13388
rect -755 -13132 -709 -13120
rect -755 -13388 -749 -13132
rect -715 -13388 -709 -13132
rect -755 -13400 -709 -13388
rect -577 -13132 -531 -13120
rect -577 -13388 -571 -13132
rect -537 -13388 -531 -13132
rect -577 -13400 -531 -13388
rect -399 -13132 -353 -13120
rect -399 -13388 -393 -13132
rect -359 -13388 -353 -13132
rect -399 -13400 -353 -13388
rect -221 -13132 -175 -13120
rect -221 -13388 -215 -13132
rect -181 -13388 -175 -13132
rect -221 -13400 -175 -13388
rect -43 -13132 3 -13120
rect -43 -13388 -37 -13132
rect -3 -13388 3 -13132
rect -43 -13400 3 -13388
rect 135 -13132 181 -13120
rect 135 -13388 141 -13132
rect 175 -13388 181 -13132
rect 135 -13400 181 -13388
rect 313 -13132 359 -13120
rect 313 -13388 319 -13132
rect 353 -13388 359 -13132
rect 313 -13400 359 -13388
rect 491 -13132 537 -13120
rect 491 -13388 497 -13132
rect 531 -13388 537 -13132
rect 491 -13400 537 -13388
rect 669 -13132 715 -13120
rect 669 -13388 675 -13132
rect 709 -13388 715 -13132
rect 669 -13400 715 -13388
rect 847 -13132 893 -13120
rect 847 -13388 853 -13132
rect 887 -13388 893 -13132
rect 847 -13400 893 -13388
rect 1025 -13132 1071 -13120
rect 1025 -13388 1031 -13132
rect 1065 -13388 1071 -13132
rect 1025 -13400 1071 -13388
rect 1203 -13132 1249 -13120
rect 1203 -13388 1209 -13132
rect 1243 -13388 1249 -13132
rect 1203 -13400 1249 -13388
rect 1381 -13132 1427 -13120
rect 1381 -13388 1387 -13132
rect 1421 -13388 1427 -13132
rect 1381 -13400 1427 -13388
rect 1559 -13132 1605 -13120
rect 1559 -13388 1565 -13132
rect 1599 -13388 1605 -13132
rect 1559 -13400 1605 -13388
rect 1737 -13132 1783 -13120
rect 1737 -13388 1743 -13132
rect 1777 -13388 1783 -13132
rect 1737 -13400 1783 -13388
rect 1915 -13132 1961 -13120
rect 1915 -13388 1921 -13132
rect 1955 -13388 1961 -13132
rect 1915 -13400 1961 -13388
rect 2093 -13132 2139 -13120
rect 2093 -13388 2099 -13132
rect 2133 -13388 2139 -13132
rect 2093 -13400 2139 -13388
rect 2271 -13132 2317 -13120
rect 2271 -13388 2277 -13132
rect 2311 -13388 2317 -13132
rect 2271 -13400 2317 -13388
rect 2449 -13132 2495 -13120
rect 2449 -13388 2455 -13132
rect 2489 -13388 2495 -13132
rect 2449 -13400 2495 -13388
rect 2627 -13132 2673 -13120
rect 2627 -13388 2633 -13132
rect 2667 -13388 2673 -13132
rect 2627 -13400 2673 -13388
rect 2805 -13132 2851 -13120
rect 2805 -13388 2811 -13132
rect 2845 -13388 2851 -13132
rect 2805 -13400 2851 -13388
rect 2983 -13132 3029 -13120
rect 2983 -13388 2989 -13132
rect 3023 -13388 3029 -13132
rect 2983 -13400 3029 -13388
rect 3161 -13132 3207 -13120
rect 3161 -13388 3167 -13132
rect 3201 -13388 3207 -13132
rect 3161 -13400 3207 -13388
rect 3339 -13132 3385 -13120
rect 3339 -13388 3345 -13132
rect 3379 -13388 3385 -13132
rect 3339 -13400 3385 -13388
rect 3517 -13132 3563 -13120
rect 3517 -13388 3523 -13132
rect 3557 -13388 3563 -13132
rect 3517 -13400 3563 -13388
rect 3695 -13132 3741 -13120
rect 3695 -13388 3701 -13132
rect 3735 -13388 3741 -13132
rect 3695 -13400 3741 -13388
rect 3873 -13132 3919 -13120
rect 3873 -13388 3879 -13132
rect 3913 -13388 3919 -13132
rect 3873 -13400 3919 -13388
rect 4051 -13132 4097 -13120
rect 4051 -13388 4057 -13132
rect 4091 -13388 4097 -13132
rect 4051 -13400 4097 -13388
rect -2105 -13438 -2029 -13432
rect -2105 -13472 -2089 -13438
rect -2045 -13472 -2029 -13438
rect -2105 -13488 -2029 -13472
rect -1995 -13545 -1961 -13400
rect -1927 -13438 -1851 -13432
rect -1927 -13472 -1911 -13438
rect -1867 -13472 -1851 -13438
rect -1927 -13488 -1851 -13472
rect -1749 -13438 -1673 -13432
rect -1749 -13472 -1733 -13438
rect -1689 -13472 -1673 -13438
rect -1749 -13488 -1673 -13472
rect -2014 -13598 -2004 -13545
rect -1951 -13598 -1941 -13545
rect -1905 -14032 -1871 -13488
rect -1728 -14032 -1694 -13488
rect -1638 -13672 -1604 -13400
rect -1571 -13438 -1495 -13432
rect -1571 -13472 -1555 -13438
rect -1511 -13472 -1495 -13438
rect -1571 -13488 -1495 -13472
rect -1393 -13438 -1317 -13432
rect -1393 -13472 -1377 -13438
rect -1333 -13472 -1317 -13438
rect -1393 -13488 -1317 -13472
rect -1658 -13725 -1648 -13672
rect -1595 -13725 -1585 -13672
rect -1550 -14032 -1516 -13488
rect -1282 -13672 -1248 -13400
rect -1215 -13438 -1139 -13432
rect -1215 -13472 -1199 -13438
rect -1155 -13472 -1139 -13438
rect -1215 -13488 -1139 -13472
rect -1037 -13438 -961 -13432
rect -1037 -13472 -1021 -13438
rect -977 -13472 -961 -13438
rect -1037 -13488 -961 -13472
rect -927 -13672 -893 -13400
rect -859 -13438 -783 -13432
rect -859 -13472 -843 -13438
rect -799 -13472 -783 -13438
rect -859 -13488 -783 -13472
rect -681 -13438 -605 -13432
rect -681 -13472 -665 -13438
rect -621 -13472 -605 -13438
rect -681 -13488 -605 -13472
rect -571 -13545 -537 -13400
rect -503 -13438 -427 -13432
rect -503 -13472 -487 -13438
rect -443 -13472 -427 -13438
rect -503 -13488 -427 -13472
rect -325 -13438 -249 -13432
rect -325 -13472 -309 -13438
rect -265 -13472 -249 -13438
rect -325 -13488 -249 -13472
rect -591 -13598 -581 -13545
rect -528 -13598 -518 -13545
rect -1301 -13725 -1291 -13672
rect -1238 -13725 -1228 -13672
rect -947 -13725 -937 -13672
rect -884 -13725 -874 -13672
rect -927 -13726 -893 -13725
rect -304 -14032 -270 -13488
rect -216 -13794 -182 -13400
rect -147 -13438 -71 -13432
rect -147 -13472 -131 -13438
rect -87 -13472 -71 -13438
rect -147 -13488 -71 -13472
rect 31 -13438 107 -13432
rect 31 -13472 47 -13438
rect 91 -13472 107 -13438
rect 31 -13488 107 -13472
rect -235 -13847 -225 -13794
rect -172 -13847 -162 -13794
rect -125 -14032 -91 -13488
rect 52 -14032 86 -13488
rect 141 -13794 175 -13400
rect 209 -13438 285 -13432
rect 209 -13472 225 -13438
rect 269 -13472 285 -13438
rect 209 -13488 285 -13472
rect 387 -13438 463 -13432
rect 387 -13472 403 -13438
rect 447 -13472 463 -13438
rect 387 -13488 463 -13472
rect 123 -13847 133 -13794
rect 186 -13847 196 -13794
rect 230 -14032 264 -13488
rect 408 -14032 442 -13488
rect 496 -13795 530 -13400
rect 942 -13432 976 -13430
rect 565 -13438 641 -13432
rect 565 -13472 581 -13438
rect 625 -13472 641 -13438
rect 565 -13488 641 -13472
rect 743 -13438 819 -13432
rect 743 -13472 759 -13438
rect 803 -13472 819 -13438
rect 743 -13488 819 -13472
rect 921 -13438 997 -13432
rect 921 -13472 937 -13438
rect 981 -13472 997 -13438
rect 921 -13488 997 -13472
rect 1099 -13438 1175 -13432
rect 1099 -13472 1115 -13438
rect 1159 -13472 1175 -13438
rect 1099 -13488 1175 -13472
rect 1277 -13438 1353 -13432
rect 1277 -13472 1293 -13438
rect 1337 -13472 1353 -13438
rect 1277 -13488 1353 -13472
rect 477 -13848 487 -13795
rect 540 -13848 550 -13795
rect 587 -14032 621 -13488
rect 942 -14032 976 -13488
rect 1388 -13672 1422 -13400
rect 1455 -13438 1531 -13432
rect 1455 -13472 1471 -13438
rect 1515 -13472 1531 -13438
rect 1455 -13488 1531 -13472
rect 1633 -13438 1709 -13432
rect 1633 -13472 1649 -13438
rect 1693 -13472 1709 -13438
rect 1633 -13488 1709 -13472
rect 1743 -13672 1777 -13400
rect 1811 -13438 1887 -13432
rect 1811 -13472 1827 -13438
rect 1871 -13472 1887 -13438
rect 1811 -13488 1887 -13472
rect 1989 -13438 2065 -13432
rect 1989 -13472 2005 -13438
rect 2049 -13472 2065 -13438
rect 1989 -13488 2065 -13472
rect 2100 -13672 2134 -13400
rect 2167 -13438 2243 -13432
rect 2167 -13472 2183 -13438
rect 2227 -13472 2243 -13438
rect 2167 -13488 2243 -13472
rect 2345 -13438 2421 -13432
rect 2345 -13472 2361 -13438
rect 2405 -13472 2421 -13438
rect 2345 -13488 2421 -13472
rect 1369 -13725 1379 -13672
rect 1432 -13725 1442 -13672
rect 1722 -13725 1732 -13672
rect 1785 -13725 1795 -13672
rect 2081 -13725 2091 -13672
rect 2144 -13725 2154 -13672
rect 2366 -14032 2400 -13488
rect 2455 -13545 2489 -13400
rect 2523 -13438 2599 -13432
rect 2523 -13472 2539 -13438
rect 2583 -13472 2599 -13438
rect 2523 -13488 2599 -13472
rect 2701 -13438 2777 -13432
rect 2701 -13472 2717 -13438
rect 2761 -13472 2777 -13438
rect 2701 -13488 2777 -13472
rect 2436 -13598 2446 -13545
rect 2499 -13598 2509 -13545
rect 2544 -14032 2578 -13488
rect 2723 -14032 2757 -13488
rect 2812 -13794 2846 -13400
rect 2879 -13438 2955 -13432
rect 2879 -13472 2895 -13438
rect 2939 -13472 2955 -13438
rect 2879 -13488 2955 -13472
rect 3057 -13438 3133 -13432
rect 3057 -13472 3073 -13438
rect 3117 -13472 3133 -13438
rect 3057 -13488 3133 -13472
rect 2792 -13847 2802 -13794
rect 2855 -13847 2865 -13794
rect 2901 -14032 2935 -13488
rect 3078 -14032 3112 -13488
rect 3166 -13795 3200 -13400
rect 3257 -13432 3291 -13431
rect 3235 -13438 3311 -13432
rect 3235 -13472 3251 -13438
rect 3295 -13472 3311 -13438
rect 3235 -13488 3311 -13472
rect 3413 -13438 3489 -13432
rect 3413 -13472 3429 -13438
rect 3473 -13472 3489 -13438
rect 3413 -13488 3489 -13472
rect 3147 -13848 3157 -13795
rect 3210 -13848 3220 -13795
rect 3257 -14032 3291 -13488
rect 3523 -13794 3557 -13400
rect 3591 -13438 3667 -13432
rect 3591 -13472 3607 -13438
rect 3651 -13472 3667 -13438
rect 3591 -13488 3667 -13472
rect 3769 -13438 3845 -13432
rect 3769 -13472 3785 -13438
rect 3829 -13472 3845 -13438
rect 3769 -13488 3845 -13472
rect 3879 -13545 3913 -13400
rect 3947 -13438 4023 -13432
rect 3947 -13472 3963 -13438
rect 4007 -13472 4023 -13438
rect 3947 -13488 4023 -13472
rect 3860 -13598 3870 -13545
rect 3923 -13598 3933 -13545
rect 3502 -13847 3512 -13794
rect 3565 -13847 3575 -13794
rect 3523 -13848 3557 -13847
rect -2105 -14048 -2029 -14032
rect -2105 -14082 -2089 -14048
rect -2045 -14082 -2029 -14048
rect -2105 -14088 -2029 -14082
rect -1927 -14048 -1851 -14032
rect -1927 -14082 -1911 -14048
rect -1867 -14082 -1851 -14048
rect -1927 -14088 -1851 -14082
rect -1749 -14048 -1673 -14032
rect -1749 -14082 -1733 -14048
rect -1689 -14082 -1673 -14048
rect -1749 -14088 -1673 -14082
rect -1571 -14048 -1495 -14032
rect -1571 -14082 -1555 -14048
rect -1511 -14082 -1495 -14048
rect -1571 -14088 -1495 -14082
rect -1393 -14048 -1317 -14032
rect -1393 -14082 -1377 -14048
rect -1333 -14082 -1317 -14048
rect -1393 -14088 -1317 -14082
rect -1215 -14048 -1139 -14032
rect -1215 -14082 -1199 -14048
rect -1155 -14082 -1139 -14048
rect -1215 -14088 -1139 -14082
rect -1037 -14048 -961 -14032
rect -1037 -14082 -1021 -14048
rect -977 -14082 -961 -14048
rect -1037 -14088 -961 -14082
rect -859 -14048 -783 -14032
rect -859 -14082 -843 -14048
rect -799 -14082 -783 -14048
rect -859 -14088 -783 -14082
rect -681 -14048 -605 -14032
rect -681 -14082 -665 -14048
rect -621 -14082 -605 -14048
rect -681 -14088 -605 -14082
rect -503 -14048 -427 -14032
rect -503 -14082 -487 -14048
rect -443 -14082 -427 -14048
rect -503 -14088 -427 -14082
rect -325 -14048 -249 -14032
rect -325 -14082 -309 -14048
rect -265 -14082 -249 -14048
rect -325 -14088 -249 -14082
rect -147 -14048 -71 -14032
rect -147 -14082 -131 -14048
rect -87 -14082 -71 -14048
rect -147 -14088 -71 -14082
rect 31 -14048 107 -14032
rect 31 -14082 47 -14048
rect 91 -14082 107 -14048
rect 31 -14088 107 -14082
rect 209 -14048 285 -14032
rect 209 -14082 225 -14048
rect 269 -14082 285 -14048
rect 209 -14088 285 -14082
rect 387 -14048 463 -14032
rect 387 -14082 403 -14048
rect 447 -14082 463 -14048
rect 387 -14088 463 -14082
rect 565 -14048 641 -14032
rect 565 -14082 581 -14048
rect 625 -14082 641 -14048
rect 565 -14088 641 -14082
rect 743 -14048 819 -14032
rect 921 -14048 997 -14032
rect 1099 -14048 1175 -14032
rect 743 -14082 759 -14048
rect 803 -14082 937 -14048
rect 981 -14082 1115 -14048
rect 1159 -14082 1175 -14048
rect 743 -14088 819 -14082
rect 853 -14120 887 -14082
rect 921 -14088 997 -14082
rect 1032 -14120 1066 -14082
rect 1099 -14088 1175 -14082
rect 1277 -14048 1353 -14032
rect 1277 -14082 1293 -14048
rect 1337 -14082 1353 -14048
rect 1277 -14088 1353 -14082
rect 1455 -14048 1531 -14032
rect 1455 -14082 1471 -14048
rect 1515 -14082 1531 -14048
rect 1455 -14088 1531 -14082
rect 1633 -14048 1709 -14032
rect 1633 -14082 1649 -14048
rect 1693 -14082 1709 -14048
rect 1633 -14088 1709 -14082
rect 1811 -14048 1887 -14032
rect 1811 -14082 1827 -14048
rect 1871 -14082 1887 -14048
rect 1811 -14088 1887 -14082
rect 1989 -14048 2065 -14032
rect 1989 -14082 2005 -14048
rect 2049 -14082 2065 -14048
rect 1989 -14088 2065 -14082
rect 2167 -14048 2243 -14032
rect 2167 -14082 2183 -14048
rect 2227 -14082 2243 -14048
rect 2167 -14088 2243 -14082
rect 2345 -14048 2421 -14032
rect 2345 -14082 2361 -14048
rect 2405 -14082 2421 -14048
rect 2345 -14088 2421 -14082
rect 2523 -14048 2599 -14032
rect 2523 -14082 2539 -14048
rect 2583 -14082 2599 -14048
rect 2523 -14088 2599 -14082
rect 2701 -14048 2777 -14032
rect 2701 -14082 2717 -14048
rect 2761 -14082 2777 -14048
rect 2701 -14088 2777 -14082
rect 2879 -14048 2955 -14032
rect 2879 -14082 2895 -14048
rect 2939 -14082 2955 -14048
rect 2879 -14088 2955 -14082
rect 3057 -14048 3133 -14032
rect 3057 -14082 3073 -14048
rect 3117 -14082 3133 -14048
rect 3057 -14088 3133 -14082
rect 3235 -14048 3311 -14032
rect 3235 -14082 3251 -14048
rect 3295 -14082 3311 -14048
rect 3235 -14088 3311 -14082
rect 3413 -14048 3489 -14032
rect 3413 -14082 3429 -14048
rect 3473 -14082 3489 -14048
rect 3413 -14088 3489 -14082
rect 3591 -14048 3667 -14032
rect 3591 -14082 3607 -14048
rect 3651 -14082 3667 -14048
rect 3591 -14088 3667 -14082
rect 3769 -14048 3845 -14032
rect 3769 -14082 3785 -14048
rect 3829 -14082 3845 -14048
rect 3769 -14088 3845 -14082
rect 3947 -14048 4023 -14032
rect 3947 -14082 3963 -14048
rect 4007 -14082 4023 -14048
rect 3947 -14088 4023 -14082
rect -2179 -14132 -2133 -14120
rect -2179 -14388 -2173 -14132
rect -2139 -14388 -2133 -14132
rect -2179 -14400 -2133 -14388
rect -2001 -14132 -1955 -14120
rect -2001 -14388 -1995 -14132
rect -1961 -14388 -1955 -14132
rect -2001 -14400 -1955 -14388
rect -1823 -14132 -1777 -14120
rect -1823 -14388 -1817 -14132
rect -1783 -14388 -1777 -14132
rect -1823 -14400 -1777 -14388
rect -1645 -14132 -1599 -14120
rect -1645 -14388 -1639 -14132
rect -1605 -14388 -1599 -14132
rect -1645 -14400 -1599 -14388
rect -1467 -14132 -1421 -14120
rect -1467 -14388 -1461 -14132
rect -1427 -14388 -1421 -14132
rect -1467 -14400 -1421 -14388
rect -1289 -14132 -1243 -14120
rect -1289 -14388 -1283 -14132
rect -1249 -14388 -1243 -14132
rect -1289 -14400 -1243 -14388
rect -1111 -14132 -1065 -14120
rect -1111 -14388 -1105 -14132
rect -1071 -14388 -1065 -14132
rect -1111 -14400 -1065 -14388
rect -933 -14132 -887 -14120
rect -933 -14388 -927 -14132
rect -893 -14388 -887 -14132
rect -933 -14400 -887 -14388
rect -755 -14132 -709 -14120
rect -755 -14388 -749 -14132
rect -715 -14388 -709 -14132
rect -755 -14400 -709 -14388
rect -577 -14132 -531 -14120
rect -577 -14388 -571 -14132
rect -537 -14388 -531 -14132
rect -577 -14400 -531 -14388
rect -399 -14132 -353 -14120
rect -399 -14388 -393 -14132
rect -359 -14388 -353 -14132
rect -399 -14400 -353 -14388
rect -221 -14132 -175 -14120
rect -221 -14388 -215 -14132
rect -181 -14388 -175 -14132
rect -221 -14400 -175 -14388
rect -43 -14132 3 -14120
rect -43 -14388 -37 -14132
rect -3 -14388 3 -14132
rect -43 -14400 3 -14388
rect 135 -14132 181 -14120
rect 135 -14388 141 -14132
rect 175 -14388 181 -14132
rect 135 -14400 181 -14388
rect 313 -14132 359 -14120
rect 313 -14388 319 -14132
rect 353 -14388 359 -14132
rect 313 -14400 359 -14388
rect 491 -14132 537 -14120
rect 491 -14388 497 -14132
rect 531 -14388 537 -14132
rect 491 -14400 537 -14388
rect 669 -14132 715 -14120
rect 669 -14388 675 -14132
rect 709 -14388 715 -14132
rect 669 -14400 715 -14388
rect 847 -14132 893 -14120
rect 847 -14388 853 -14132
rect 887 -14388 893 -14132
rect 847 -14400 893 -14388
rect 1025 -14132 1071 -14120
rect 1025 -14388 1031 -14132
rect 1065 -14388 1071 -14132
rect 1025 -14400 1071 -14388
rect 1203 -14132 1249 -14120
rect 1203 -14388 1209 -14132
rect 1243 -14388 1249 -14132
rect 1203 -14400 1249 -14388
rect 1381 -14132 1427 -14120
rect 1381 -14388 1387 -14132
rect 1421 -14388 1427 -14132
rect 1381 -14400 1427 -14388
rect 1559 -14132 1605 -14120
rect 1559 -14388 1565 -14132
rect 1599 -14388 1605 -14132
rect 1559 -14400 1605 -14388
rect 1737 -14132 1783 -14120
rect 1737 -14388 1743 -14132
rect 1777 -14388 1783 -14132
rect 1737 -14400 1783 -14388
rect 1915 -14132 1961 -14120
rect 1915 -14388 1921 -14132
rect 1955 -14388 1961 -14132
rect 1915 -14400 1961 -14388
rect 2093 -14132 2139 -14120
rect 2093 -14388 2099 -14132
rect 2133 -14388 2139 -14132
rect 2093 -14400 2139 -14388
rect 2271 -14132 2317 -14120
rect 2271 -14388 2277 -14132
rect 2311 -14388 2317 -14132
rect 2271 -14400 2317 -14388
rect 2449 -14132 2495 -14120
rect 2449 -14388 2455 -14132
rect 2489 -14388 2495 -14132
rect 2449 -14400 2495 -14388
rect 2627 -14132 2673 -14120
rect 2627 -14388 2633 -14132
rect 2667 -14388 2673 -14132
rect 2627 -14400 2673 -14388
rect 2805 -14132 2851 -14120
rect 2805 -14388 2811 -14132
rect 2845 -14388 2851 -14132
rect 2805 -14400 2851 -14388
rect 2983 -14132 3029 -14120
rect 2983 -14388 2989 -14132
rect 3023 -14388 3029 -14132
rect 2983 -14400 3029 -14388
rect 3161 -14132 3207 -14120
rect 3161 -14388 3167 -14132
rect 3201 -14388 3207 -14132
rect 3161 -14400 3207 -14388
rect 3339 -14132 3385 -14120
rect 3339 -14388 3345 -14132
rect 3379 -14388 3385 -14132
rect 3339 -14400 3385 -14388
rect 3517 -14132 3563 -14120
rect 3517 -14388 3523 -14132
rect 3557 -14388 3563 -14132
rect 3517 -14400 3563 -14388
rect 3695 -14132 3741 -14120
rect 3695 -14388 3701 -14132
rect 3735 -14388 3741 -14132
rect 3695 -14400 3741 -14388
rect 3873 -14132 3919 -14120
rect 3873 -14388 3879 -14132
rect 3913 -14388 3919 -14132
rect 3873 -14400 3919 -14388
rect 4051 -14132 4097 -14120
rect 4051 -14388 4057 -14132
rect 4091 -14388 4097 -14132
rect 4051 -14400 4097 -14388
rect -2173 -14441 -2139 -14400
rect -2105 -14438 -2029 -14432
rect -2105 -14441 -2089 -14438
rect -2173 -14472 -2089 -14441
rect -2045 -14441 -2029 -14438
rect -1995 -14441 -1961 -14400
rect -2045 -14472 -1961 -14441
rect -2173 -14475 -1961 -14472
rect -2105 -14488 -2029 -14475
rect -2325 -14596 -2315 -14543
rect -2262 -14596 -2252 -14543
rect -2105 -15045 -2029 -15032
rect -1995 -15045 -1961 -14475
rect -1927 -14438 -1851 -14432
rect -1927 -14472 -1911 -14438
rect -1867 -14472 -1851 -14438
rect -1927 -14488 -1851 -14472
rect -2176 -15048 -1961 -15045
rect -2176 -15079 -2089 -15048
rect -2176 -15120 -2142 -15079
rect -2105 -15082 -2089 -15079
rect -2045 -15079 -1961 -15048
rect -2045 -15082 -2029 -15079
rect -2105 -15088 -2029 -15082
rect -1995 -15120 -1961 -15079
rect -1927 -15048 -1851 -15032
rect -1927 -15082 -1911 -15048
rect -1867 -15082 -1851 -15048
rect -1927 -15088 -1851 -15082
rect -1817 -15120 -1783 -14400
rect -1749 -14438 -1673 -14432
rect -1749 -14472 -1733 -14438
rect -1689 -14472 -1673 -14438
rect -1749 -14488 -1673 -14472
rect -1749 -15048 -1673 -15032
rect -1749 -15082 -1733 -15048
rect -1689 -15082 -1673 -15048
rect -1749 -15088 -1673 -15082
rect -1639 -15120 -1605 -14400
rect -1571 -14438 -1495 -14432
rect -1571 -14472 -1555 -14438
rect -1511 -14472 -1495 -14438
rect -1571 -14488 -1495 -14472
rect -1571 -15048 -1495 -15032
rect -1571 -15082 -1555 -15048
rect -1511 -15082 -1495 -15048
rect -1571 -15088 -1495 -15082
rect -1461 -15120 -1427 -14400
rect -1393 -14438 -1317 -14432
rect -1393 -14472 -1377 -14438
rect -1333 -14472 -1317 -14438
rect -1393 -14488 -1317 -14472
rect -1371 -14543 -1337 -14488
rect -1391 -14596 -1381 -14543
rect -1328 -14596 -1318 -14543
rect -1371 -15032 -1337 -14596
rect -1393 -15048 -1317 -15032
rect -1393 -15082 -1377 -15048
rect -1333 -15082 -1317 -15048
rect -1393 -15088 -1317 -15082
rect -1283 -15120 -1249 -14400
rect -1215 -14438 -1139 -14432
rect -1215 -14472 -1199 -14438
rect -1155 -14472 -1139 -14438
rect -1215 -14488 -1139 -14472
rect -1194 -14543 -1160 -14488
rect -1214 -14596 -1204 -14543
rect -1151 -14596 -1141 -14543
rect -1215 -15048 -1139 -15032
rect -1215 -15082 -1199 -15048
rect -1155 -15082 -1139 -15048
rect -1215 -15088 -1139 -15082
rect -1104 -15120 -1070 -14400
rect -1037 -14438 -961 -14432
rect -1037 -14472 -1021 -14438
rect -977 -14472 -961 -14438
rect -1037 -14488 -961 -14472
rect -1016 -14543 -982 -14488
rect -1036 -14596 -1026 -14543
rect -973 -14596 -963 -14543
rect -1037 -15048 -961 -15032
rect -1037 -15082 -1021 -15048
rect -977 -15082 -961 -15048
rect -1037 -15088 -961 -15082
rect -927 -15120 -893 -14400
rect -859 -14438 -783 -14432
rect -859 -14472 -843 -14438
rect -799 -14472 -783 -14438
rect -859 -14488 -783 -14472
rect -838 -14543 -804 -14488
rect -858 -14596 -848 -14543
rect -795 -14596 -785 -14543
rect -857 -14979 -847 -14926
rect -794 -14979 -784 -14926
rect -838 -15032 -804 -14979
rect -859 -15048 -783 -15032
rect -859 -15082 -843 -15048
rect -799 -15082 -783 -15048
rect -859 -15088 -783 -15082
rect -749 -15120 -715 -14400
rect -681 -14438 -605 -14432
rect -681 -14472 -665 -14438
rect -621 -14472 -605 -14438
rect -681 -14488 -605 -14472
rect -659 -14543 -625 -14488
rect -679 -14596 -669 -14543
rect -616 -14596 -606 -14543
rect -679 -14979 -669 -14926
rect -616 -14979 -606 -14926
rect -660 -15032 -626 -14979
rect -681 -15048 -605 -15032
rect -681 -15082 -665 -15048
rect -621 -15082 -605 -15048
rect -681 -15088 -605 -15082
rect -571 -15120 -537 -14400
rect -503 -14438 -427 -14432
rect -503 -14472 -487 -14438
rect -443 -14472 -427 -14438
rect -503 -14488 -427 -14472
rect -482 -14543 -448 -14488
rect -501 -14596 -491 -14543
rect -438 -14596 -428 -14543
rect -501 -14979 -491 -14926
rect -438 -14979 -428 -14926
rect -481 -15032 -447 -14979
rect -503 -15048 -427 -15032
rect -503 -15082 -487 -15048
rect -443 -15082 -427 -15048
rect -503 -15088 -427 -15082
rect -393 -15120 -359 -14400
rect -325 -14438 -249 -14432
rect -325 -14472 -309 -14438
rect -265 -14472 -249 -14438
rect -325 -14488 -249 -14472
rect -304 -14927 -270 -14488
rect -324 -14980 -314 -14927
rect -261 -14980 -251 -14927
rect -304 -15032 -270 -14980
rect -325 -15048 -249 -15032
rect -325 -15082 -309 -15048
rect -265 -15082 -249 -15048
rect -325 -15088 -249 -15082
rect -215 -15120 -181 -14400
rect -147 -14438 -71 -14432
rect -147 -14472 -131 -14438
rect -87 -14472 -71 -14438
rect -147 -14488 -71 -14472
rect -126 -14926 -92 -14488
rect -147 -14979 -137 -14926
rect -84 -14979 -74 -14926
rect -126 -15032 -92 -14979
rect -147 -15048 -71 -15032
rect -147 -15082 -131 -15048
rect -87 -15082 -71 -15048
rect -147 -15088 -71 -15082
rect -37 -15120 -3 -14400
rect 31 -14438 107 -14432
rect 31 -14472 47 -14438
rect 91 -14472 107 -14438
rect 31 -14488 107 -14472
rect 52 -14926 86 -14488
rect 33 -14979 43 -14926
rect 96 -14979 106 -14926
rect 52 -15032 86 -14979
rect 31 -15048 107 -15032
rect 31 -15082 47 -15048
rect 91 -15082 107 -15048
rect 31 -15088 107 -15082
rect 141 -15120 175 -14400
rect 209 -14438 285 -14432
rect 209 -14472 225 -14438
rect 269 -14472 285 -14438
rect 209 -14488 285 -14472
rect 209 -15048 285 -15032
rect 209 -15082 225 -15048
rect 269 -15082 285 -15048
rect 209 -15088 285 -15082
rect 319 -15120 353 -14400
rect 387 -14438 463 -14432
rect 387 -14472 403 -14438
rect 447 -14472 463 -14438
rect 387 -14488 463 -14472
rect 387 -15048 463 -15032
rect 387 -15082 403 -15048
rect 447 -15082 463 -15048
rect 387 -15088 463 -15082
rect 497 -15120 531 -14400
rect 565 -14438 641 -14432
rect 565 -14472 581 -14438
rect 625 -14472 641 -14438
rect 565 -14488 641 -14472
rect 565 -15048 641 -15032
rect 565 -15082 581 -15048
rect 625 -15082 641 -15048
rect 565 -15088 641 -15082
rect 675 -15120 709 -14400
rect 743 -14438 819 -14432
rect 743 -14472 759 -14438
rect 803 -14472 819 -14438
rect 743 -14488 819 -14472
rect 921 -14438 997 -14432
rect 921 -14472 937 -14438
rect 981 -14472 997 -14438
rect 921 -14488 997 -14472
rect 743 -15048 819 -15032
rect 743 -15082 759 -15048
rect 803 -15082 819 -15048
rect 743 -15088 819 -15082
rect 921 -15048 997 -15032
rect 921 -15082 937 -15048
rect 981 -15082 997 -15048
rect 921 -15088 997 -15082
rect 1031 -15120 1065 -14400
rect 1099 -14438 1175 -14432
rect 1099 -14472 1115 -14438
rect 1159 -14472 1175 -14438
rect 1099 -14488 1175 -14472
rect 1099 -15048 1175 -15032
rect 1099 -15082 1115 -15048
rect 1159 -15082 1175 -15048
rect 1099 -15088 1175 -15082
rect 1209 -15120 1243 -14400
rect 1277 -14438 1353 -14432
rect 1277 -14472 1293 -14438
rect 1337 -14472 1353 -14438
rect 1277 -14488 1353 -14472
rect 1298 -14543 1332 -14488
rect 1278 -14596 1288 -14543
rect 1341 -14596 1351 -14543
rect 1279 -14980 1289 -14927
rect 1342 -14980 1352 -14927
rect 1298 -15032 1332 -14980
rect 1277 -15048 1353 -15032
rect 1277 -15082 1293 -15048
rect 1337 -15082 1353 -15048
rect 1277 -15088 1353 -15082
rect 1387 -15120 1421 -14400
rect 1455 -14438 1531 -14432
rect 1455 -14472 1471 -14438
rect 1515 -14472 1531 -14438
rect 1455 -14488 1531 -14472
rect 1477 -14543 1511 -14488
rect 1456 -14596 1466 -14543
rect 1519 -14596 1529 -14543
rect 1457 -14979 1467 -14926
rect 1520 -14979 1530 -14926
rect 1476 -15032 1510 -14979
rect 1455 -15048 1531 -15032
rect 1455 -15082 1471 -15048
rect 1515 -15082 1531 -15048
rect 1455 -15088 1531 -15082
rect 1565 -15120 1599 -14400
rect 1633 -14438 1709 -14432
rect 1633 -14472 1649 -14438
rect 1693 -14472 1709 -14438
rect 1633 -14488 1709 -14472
rect 1654 -14543 1688 -14488
rect 1634 -14596 1644 -14543
rect 1697 -14596 1707 -14543
rect 1634 -14979 1644 -14926
rect 1697 -14979 1707 -14926
rect 1654 -15032 1688 -14979
rect 1633 -15048 1709 -15032
rect 1633 -15082 1649 -15048
rect 1693 -15082 1709 -15048
rect 1633 -15088 1709 -15082
rect 1744 -15120 1778 -14400
rect 1811 -14438 1887 -14432
rect 1811 -14472 1827 -14438
rect 1871 -14472 1887 -14438
rect 1811 -14488 1887 -14472
rect 1832 -14542 1866 -14488
rect 1813 -14595 1823 -14542
rect 1876 -14595 1886 -14542
rect 1812 -14979 1822 -14926
rect 1875 -14979 1885 -14926
rect 1833 -15032 1867 -14979
rect 1811 -15048 1887 -15032
rect 1811 -15082 1827 -15048
rect 1871 -15082 1887 -15048
rect 1811 -15088 1887 -15082
rect 1921 -15120 1955 -14400
rect 1989 -14438 2065 -14432
rect 1989 -14472 2005 -14438
rect 2049 -14472 2065 -14438
rect 1989 -14488 2065 -14472
rect 2010 -14543 2044 -14488
rect 1990 -14596 2000 -14543
rect 2053 -14596 2063 -14543
rect 1989 -14979 1999 -14926
rect 2052 -14979 2062 -14926
rect 2010 -15032 2044 -14979
rect 1989 -15048 2065 -15032
rect 1989 -15082 2005 -15048
rect 2049 -15082 2065 -15048
rect 1989 -15088 2065 -15082
rect 2100 -15120 2134 -14400
rect 2167 -14438 2243 -14432
rect 2167 -14472 2183 -14438
rect 2227 -14472 2243 -14438
rect 2167 -14488 2243 -14472
rect 2188 -14543 2222 -14488
rect 2168 -14596 2178 -14543
rect 2231 -14596 2241 -14543
rect 2170 -14979 2180 -14926
rect 2233 -14979 2243 -14926
rect 2189 -15032 2223 -14979
rect 2167 -15048 2243 -15032
rect 2167 -15082 2183 -15048
rect 2227 -15082 2243 -15048
rect 2167 -15088 2243 -15082
rect 2277 -15120 2311 -14400
rect 2345 -14438 2421 -14432
rect 2345 -14472 2361 -14438
rect 2405 -14472 2421 -14438
rect 2345 -14488 2421 -14472
rect 2345 -15048 2421 -15032
rect 2345 -15082 2361 -15048
rect 2405 -15082 2421 -15048
rect 2345 -15088 2421 -15082
rect 2455 -15120 2489 -14400
rect 2523 -14438 2599 -14432
rect 2523 -14472 2539 -14438
rect 2583 -14472 2599 -14438
rect 2523 -14488 2599 -14472
rect 2523 -15048 2599 -15032
rect 2523 -15082 2539 -15048
rect 2583 -15082 2599 -15048
rect 2523 -15088 2599 -15082
rect 2633 -15120 2667 -14400
rect 2701 -14438 2777 -14432
rect 2701 -14472 2717 -14438
rect 2761 -14472 2777 -14438
rect 2701 -14488 2777 -14472
rect 2701 -15048 2777 -15032
rect 2701 -15082 2717 -15048
rect 2761 -15082 2777 -15048
rect 2701 -15088 2777 -15082
rect 2811 -15120 2845 -14400
rect 2879 -14438 2955 -14432
rect 2879 -14472 2895 -14438
rect 2939 -14472 2955 -14438
rect 2879 -14488 2955 -14472
rect 2879 -15048 2955 -15032
rect 2879 -15082 2895 -15048
rect 2939 -15082 2955 -15048
rect 2879 -15088 2955 -15082
rect 2989 -15120 3023 -14400
rect 3057 -14438 3133 -14432
rect 3057 -14472 3073 -14438
rect 3117 -14472 3133 -14438
rect 3057 -14488 3133 -14472
rect 3057 -15048 3133 -15032
rect 3057 -15082 3073 -15048
rect 3117 -15082 3133 -15048
rect 3057 -15088 3133 -15082
rect 3167 -15120 3201 -14400
rect 3235 -14438 3311 -14432
rect 3235 -14472 3251 -14438
rect 3295 -14472 3311 -14438
rect 3235 -14488 3311 -14472
rect 3236 -14597 3246 -14544
rect 3299 -14597 3309 -14544
rect 3256 -15032 3290 -14597
rect 3235 -15048 3311 -15032
rect 3235 -15082 3251 -15048
rect 3295 -15082 3311 -15048
rect 3235 -15088 3311 -15082
rect 3345 -15120 3379 -14400
rect 3413 -14438 3489 -14432
rect 3413 -14472 3429 -14438
rect 3473 -14472 3489 -14438
rect 3413 -14488 3489 -14472
rect 3434 -14543 3468 -14488
rect 3414 -14596 3424 -14543
rect 3477 -14596 3487 -14543
rect 3415 -14979 3425 -14926
rect 3478 -14979 3488 -14926
rect 3434 -15032 3468 -14979
rect 3413 -15048 3489 -15032
rect 3413 -15082 3429 -15048
rect 3473 -15082 3489 -15048
rect 3413 -15088 3489 -15082
rect 3524 -15120 3558 -14400
rect 3591 -14438 3667 -14432
rect 3591 -14472 3607 -14438
rect 3651 -14472 3667 -14438
rect 3591 -14488 3667 -14472
rect 3612 -14543 3646 -14488
rect 3592 -14596 3602 -14543
rect 3655 -14596 3665 -14543
rect 3593 -14979 3603 -14926
rect 3656 -14979 3666 -14926
rect 3612 -15032 3646 -14979
rect 3591 -15048 3667 -15032
rect 3591 -15082 3607 -15048
rect 3651 -15082 3667 -15048
rect 3591 -15088 3667 -15082
rect 3701 -15120 3735 -14400
rect 3769 -14438 3845 -14432
rect 3769 -14472 3785 -14438
rect 3829 -14472 3845 -14438
rect 3769 -14488 3845 -14472
rect 3879 -14439 3913 -14400
rect 3947 -14438 4023 -14432
rect 3947 -14439 3963 -14438
rect 3879 -14472 3963 -14439
rect 4007 -14439 4023 -14438
rect 4057 -14439 4091 -14400
rect 4007 -14472 4091 -14439
rect 3879 -14473 4091 -14472
rect 3791 -14543 3825 -14488
rect 3771 -14596 3781 -14543
rect 3834 -14596 3844 -14543
rect 3770 -14979 3780 -14926
rect 3833 -14979 3843 -14926
rect 3790 -15032 3824 -14979
rect 3769 -15048 3845 -15032
rect 3769 -15082 3785 -15048
rect 3829 -15082 3845 -15048
rect 3769 -15088 3845 -15082
rect 3879 -15047 3913 -14473
rect 3947 -14488 4023 -14473
rect 4905 -14545 4958 -7905
rect 5037 -13296 5090 -7903
rect 5174 -7908 5184 -7855
rect 5237 -7908 5247 -7855
rect 5327 -7903 5337 -7850
rect 5390 -7903 5400 -7850
rect 5185 -8635 5237 -7908
rect 5175 -8687 5185 -8635
rect 5237 -8687 5247 -8635
rect 5337 -9925 5390 -7903
rect 11647 -8716 11681 -8715
rect 6690 -8760 6815 -8726
rect 6580 -8810 6656 -8794
rect 6580 -8844 6596 -8810
rect 6640 -8844 6656 -8810
rect 6580 -8850 6656 -8844
rect 6690 -8882 6724 -8760
rect 6781 -8794 6815 -8760
rect 11044 -8769 11054 -8716
rect 11107 -8769 11117 -8716
rect 11335 -8769 11345 -8716
rect 11398 -8769 11408 -8716
rect 11628 -8769 11638 -8716
rect 11691 -8769 11701 -8716
rect 11922 -8769 11932 -8716
rect 11985 -8769 11995 -8716
rect 12212 -8769 12222 -8716
rect 12275 -8769 12285 -8716
rect 6758 -8810 6834 -8794
rect 6758 -8844 6774 -8810
rect 6818 -8844 6834 -8810
rect 6758 -8850 6834 -8844
rect 6936 -8810 7012 -8794
rect 6936 -8844 6952 -8810
rect 6996 -8844 7012 -8810
rect 6936 -8850 7012 -8844
rect 7114 -8810 7190 -8794
rect 7114 -8844 7130 -8810
rect 7174 -8844 7190 -8810
rect 7114 -8850 7190 -8844
rect 7292 -8810 7368 -8794
rect 7292 -8844 7308 -8810
rect 7352 -8844 7368 -8810
rect 7292 -8850 7368 -8844
rect 7470 -8810 7546 -8794
rect 7470 -8844 7486 -8810
rect 7530 -8844 7546 -8810
rect 7470 -8850 7546 -8844
rect 7648 -8810 7724 -8794
rect 7648 -8844 7664 -8810
rect 7708 -8844 7724 -8810
rect 7648 -8850 7724 -8844
rect 7826 -8810 7902 -8794
rect 7826 -8844 7842 -8810
rect 7886 -8844 7902 -8810
rect 7826 -8850 7902 -8844
rect 8004 -8810 8080 -8794
rect 8004 -8844 8020 -8810
rect 8064 -8844 8080 -8810
rect 8004 -8850 8080 -8844
rect 8182 -8810 8258 -8794
rect 8182 -8844 8198 -8810
rect 8242 -8844 8258 -8810
rect 8182 -8850 8258 -8844
rect 8360 -8810 8436 -8794
rect 8360 -8844 8376 -8810
rect 8420 -8844 8436 -8810
rect 8360 -8850 8436 -8844
rect 8538 -8810 8614 -8794
rect 8538 -8844 8554 -8810
rect 8598 -8844 8614 -8810
rect 8538 -8850 8614 -8844
rect 8716 -8810 8792 -8794
rect 8716 -8844 8732 -8810
rect 8776 -8844 8792 -8810
rect 8716 -8850 8792 -8844
rect 8894 -8810 8970 -8794
rect 9072 -8808 9148 -8794
rect 9250 -8808 9326 -8794
rect 8894 -8844 8910 -8810
rect 8954 -8844 8970 -8810
rect 8894 -8850 8970 -8844
rect 9004 -8810 9395 -8808
rect 9004 -8842 9088 -8810
rect 9004 -8882 9038 -8842
rect 9072 -8844 9088 -8842
rect 9132 -8842 9266 -8810
rect 9132 -8844 9148 -8842
rect 9072 -8850 9148 -8844
rect 9183 -8882 9217 -8842
rect 9250 -8844 9266 -8842
rect 9310 -8842 9395 -8810
rect 9310 -8844 9326 -8842
rect 9250 -8850 9326 -8844
rect 9361 -8882 9395 -8842
rect 10840 -8840 10916 -8824
rect 10840 -8874 10856 -8840
rect 10900 -8874 10916 -8840
rect 10840 -8880 10916 -8874
rect 6506 -8894 6552 -8882
rect 6506 -9150 6512 -8894
rect 6546 -9150 6552 -8894
rect 6506 -9162 6552 -9150
rect 6684 -8894 6730 -8882
rect 6684 -9150 6690 -8894
rect 6724 -9150 6730 -8894
rect 6684 -9162 6730 -9150
rect 6862 -8894 6908 -8882
rect 6862 -9150 6868 -8894
rect 6902 -9150 6908 -8894
rect 6862 -9162 6908 -9150
rect 7040 -8894 7086 -8882
rect 7040 -9150 7046 -8894
rect 7080 -9150 7086 -8894
rect 7040 -9162 7086 -9150
rect 7218 -8894 7264 -8882
rect 7218 -9150 7224 -8894
rect 7258 -9150 7264 -8894
rect 7218 -9162 7264 -9150
rect 7396 -8894 7442 -8882
rect 7396 -9150 7402 -8894
rect 7436 -9150 7442 -8894
rect 7396 -9162 7442 -9150
rect 7574 -8894 7620 -8882
rect 7574 -9150 7580 -8894
rect 7614 -9150 7620 -8894
rect 7574 -9162 7620 -9150
rect 7752 -8894 7798 -8882
rect 7752 -9150 7758 -8894
rect 7792 -9150 7798 -8894
rect 7752 -9162 7798 -9150
rect 7930 -8894 7976 -8882
rect 7930 -9150 7936 -8894
rect 7970 -9150 7976 -8894
rect 7930 -9162 7976 -9150
rect 8108 -8894 8154 -8882
rect 8108 -9150 8114 -8894
rect 8148 -9150 8154 -8894
rect 8108 -9162 8154 -9150
rect 8286 -8894 8332 -8882
rect 8286 -9150 8292 -8894
rect 8326 -9150 8332 -8894
rect 8286 -9162 8332 -9150
rect 8464 -8894 8510 -8882
rect 8464 -9150 8470 -8894
rect 8504 -9150 8510 -8894
rect 8464 -9162 8510 -9150
rect 8642 -8894 8688 -8882
rect 8642 -9150 8648 -8894
rect 8682 -9150 8688 -8894
rect 8642 -9162 8688 -9150
rect 8820 -8894 8866 -8882
rect 8820 -9150 8826 -8894
rect 8860 -9150 8866 -8894
rect 8820 -9162 8866 -9150
rect 8998 -8894 9044 -8882
rect 8998 -9150 9004 -8894
rect 9038 -9150 9044 -8894
rect 8998 -9162 9044 -9150
rect 9176 -8894 9222 -8882
rect 9176 -9150 9182 -8894
rect 9216 -9150 9222 -8894
rect 9176 -9162 9222 -9150
rect 9354 -8894 9400 -8882
rect 9354 -9150 9360 -8894
rect 9394 -9150 9400 -8894
rect 11063 -8912 11097 -8769
rect 11132 -8840 11208 -8824
rect 11132 -8874 11148 -8840
rect 11192 -8874 11208 -8840
rect 11132 -8880 11208 -8874
rect 11354 -8912 11388 -8769
rect 11424 -8840 11500 -8824
rect 11424 -8874 11440 -8840
rect 11484 -8874 11500 -8840
rect 11424 -8880 11500 -8874
rect 11647 -8912 11681 -8769
rect 11716 -8840 11792 -8824
rect 11716 -8874 11732 -8840
rect 11776 -8874 11792 -8840
rect 11716 -8880 11792 -8874
rect 11941 -8912 11975 -8769
rect 12008 -8840 12084 -8824
rect 12008 -8874 12024 -8840
rect 12068 -8874 12084 -8840
rect 12008 -8880 12084 -8874
rect 12231 -8840 12265 -8769
rect 12300 -8840 12376 -8824
rect 12592 -8840 12668 -8824
rect 12231 -8874 12316 -8840
rect 12360 -8874 12608 -8840
rect 12652 -8874 12738 -8840
rect 12231 -8912 12265 -8874
rect 12300 -8880 12376 -8874
rect 12522 -8912 12556 -8874
rect 12592 -8880 12668 -8874
rect 12704 -8912 12738 -8874
rect 9354 -9162 9400 -9150
rect 10766 -8924 10812 -8912
rect 6513 -9201 6547 -9162
rect 6580 -9200 6656 -9194
rect 6580 -9201 6596 -9200
rect 6513 -9234 6596 -9201
rect 6640 -9201 6656 -9200
rect 6689 -9201 6723 -9162
rect 6640 -9234 6723 -9201
rect 6513 -9235 6723 -9234
rect 6758 -9200 6834 -9194
rect 6758 -9234 6774 -9200
rect 6818 -9234 6834 -9200
rect 6580 -9250 6656 -9235
rect 6758 -9250 6834 -9234
rect 6779 -9314 6813 -9250
rect 6759 -9367 6769 -9314
rect 6822 -9367 6832 -9314
rect 6669 -9598 6679 -9545
rect 6732 -9598 6742 -9545
rect 6580 -9710 6656 -9694
rect 6580 -9744 6596 -9710
rect 6640 -9744 6656 -9710
rect 6580 -9750 6656 -9744
rect 6690 -9782 6724 -9598
rect 6779 -9694 6813 -9367
rect 6758 -9710 6834 -9694
rect 6758 -9744 6774 -9710
rect 6818 -9744 6834 -9710
rect 6758 -9750 6834 -9744
rect 6868 -9782 6902 -9162
rect 6936 -9200 7012 -9194
rect 6936 -9234 6952 -9200
rect 6996 -9234 7012 -9200
rect 6936 -9250 7012 -9234
rect 6957 -9315 6991 -9250
rect 6937 -9368 6947 -9315
rect 7000 -9368 7010 -9315
rect 6957 -9621 6991 -9368
rect 7046 -9621 7080 -9162
rect 7114 -9200 7190 -9194
rect 7114 -9234 7130 -9200
rect 7174 -9234 7190 -9200
rect 7114 -9250 7190 -9234
rect 7135 -9315 7169 -9250
rect 7116 -9368 7126 -9315
rect 7179 -9368 7189 -9315
rect 6957 -9655 7080 -9621
rect 6957 -9694 6991 -9655
rect 6936 -9710 7012 -9694
rect 6936 -9744 6952 -9710
rect 6996 -9744 7012 -9710
rect 6936 -9750 7012 -9744
rect 7046 -9782 7080 -9655
rect 7135 -9694 7169 -9368
rect 7114 -9710 7190 -9694
rect 7114 -9744 7130 -9710
rect 7174 -9744 7190 -9710
rect 7114 -9750 7190 -9744
rect 7224 -9782 7258 -9162
rect 7292 -9200 7368 -9194
rect 7292 -9234 7308 -9200
rect 7352 -9234 7368 -9200
rect 7292 -9250 7368 -9234
rect 7313 -9313 7347 -9250
rect 7293 -9366 7303 -9313
rect 7356 -9366 7366 -9313
rect 7313 -9694 7347 -9366
rect 7292 -9710 7368 -9694
rect 7292 -9744 7308 -9710
rect 7352 -9744 7368 -9710
rect 7292 -9750 7368 -9744
rect 7402 -9782 7436 -9162
rect 7470 -9200 7546 -9194
rect 7470 -9234 7486 -9200
rect 7530 -9234 7546 -9200
rect 7470 -9250 7546 -9234
rect 7491 -9313 7525 -9250
rect 7472 -9366 7482 -9313
rect 7535 -9366 7545 -9313
rect 7491 -9694 7525 -9366
rect 7470 -9710 7546 -9694
rect 7470 -9744 7486 -9710
rect 7530 -9744 7546 -9710
rect 7470 -9750 7546 -9744
rect 7580 -9782 7614 -9162
rect 7648 -9200 7724 -9194
rect 7648 -9234 7664 -9200
rect 7708 -9234 7724 -9200
rect 7648 -9250 7724 -9234
rect 7669 -9315 7703 -9250
rect 7649 -9368 7659 -9315
rect 7712 -9368 7722 -9315
rect 7669 -9694 7703 -9368
rect 7648 -9710 7724 -9694
rect 7648 -9744 7664 -9710
rect 7708 -9744 7724 -9710
rect 7648 -9750 7724 -9744
rect 7758 -9782 7792 -9162
rect 7826 -9200 7902 -9194
rect 7826 -9234 7842 -9200
rect 7886 -9234 7902 -9200
rect 7826 -9250 7902 -9234
rect 7847 -9314 7881 -9250
rect 7827 -9367 7837 -9314
rect 7890 -9367 7900 -9314
rect 7847 -9694 7881 -9367
rect 7826 -9710 7902 -9694
rect 7826 -9744 7842 -9710
rect 7886 -9744 7902 -9710
rect 7826 -9750 7902 -9744
rect 7936 -9782 7970 -9162
rect 8004 -9200 8080 -9194
rect 8004 -9234 8020 -9200
rect 8064 -9234 8080 -9200
rect 8004 -9250 8080 -9234
rect 8025 -9315 8059 -9250
rect 8005 -9368 8015 -9315
rect 8068 -9368 8078 -9315
rect 8025 -9694 8059 -9368
rect 8004 -9710 8080 -9694
rect 8004 -9744 8020 -9710
rect 8064 -9744 8080 -9710
rect 8004 -9750 8080 -9744
rect 8113 -9782 8147 -9162
rect 8182 -9200 8258 -9194
rect 8182 -9234 8198 -9200
rect 8242 -9234 8258 -9200
rect 8182 -9250 8258 -9234
rect 8203 -9314 8237 -9250
rect 8184 -9367 8194 -9314
rect 8247 -9367 8257 -9314
rect 8203 -9694 8237 -9367
rect 8182 -9710 8258 -9694
rect 8182 -9744 8198 -9710
rect 8242 -9744 8258 -9710
rect 8182 -9750 8258 -9744
rect 8292 -9782 8326 -9162
rect 8360 -9200 8436 -9194
rect 8360 -9234 8376 -9200
rect 8420 -9234 8436 -9200
rect 8360 -9250 8436 -9234
rect 8381 -9314 8415 -9250
rect 8361 -9367 8371 -9314
rect 8424 -9367 8434 -9314
rect 8381 -9694 8415 -9367
rect 8360 -9710 8436 -9694
rect 8360 -9744 8376 -9710
rect 8420 -9744 8436 -9710
rect 8360 -9750 8436 -9744
rect 8470 -9782 8504 -9162
rect 8538 -9200 8614 -9194
rect 8538 -9234 8554 -9200
rect 8598 -9234 8614 -9200
rect 8538 -9250 8614 -9234
rect 8559 -9314 8593 -9250
rect 8539 -9367 8549 -9314
rect 8602 -9367 8612 -9314
rect 8559 -9694 8593 -9367
rect 8538 -9710 8614 -9694
rect 8538 -9744 8554 -9710
rect 8598 -9744 8614 -9710
rect 8538 -9750 8614 -9744
rect 8648 -9782 8682 -9162
rect 8716 -9200 8792 -9194
rect 8716 -9234 8732 -9200
rect 8776 -9234 8792 -9200
rect 8716 -9250 8792 -9234
rect 8737 -9315 8771 -9250
rect 8717 -9368 8727 -9315
rect 8780 -9368 8790 -9315
rect 8737 -9694 8771 -9368
rect 8716 -9710 8792 -9694
rect 8716 -9744 8732 -9710
rect 8776 -9744 8792 -9710
rect 8716 -9750 8792 -9744
rect 8826 -9782 8860 -9162
rect 8894 -9200 8970 -9194
rect 8894 -9234 8910 -9200
rect 8954 -9234 8970 -9200
rect 8894 -9250 8970 -9234
rect 8915 -9314 8949 -9250
rect 8896 -9367 8906 -9314
rect 8959 -9367 8969 -9314
rect 8915 -9694 8949 -9367
rect 8894 -9710 8970 -9694
rect 8894 -9744 8910 -9710
rect 8954 -9744 8970 -9710
rect 8894 -9750 8970 -9744
rect 9004 -9709 9038 -9162
rect 10766 -9180 10772 -8924
rect 10806 -9180 10812 -8924
rect 10766 -9192 10812 -9180
rect 10944 -8924 10990 -8912
rect 10944 -9180 10950 -8924
rect 10984 -9145 10990 -8924
rect 11058 -8924 11104 -8912
rect 11058 -9145 11064 -8924
rect 10984 -9179 11064 -9145
rect 10984 -9180 10990 -9179
rect 10944 -9192 10990 -9180
rect 11058 -9180 11064 -9179
rect 11098 -9180 11104 -8924
rect 11058 -9192 11104 -9180
rect 11236 -8924 11282 -8912
rect 11236 -9180 11242 -8924
rect 11276 -9180 11282 -8924
rect 11236 -9192 11282 -9180
rect 11350 -8924 11396 -8912
rect 11350 -9180 11356 -8924
rect 11390 -9180 11396 -8924
rect 11350 -9192 11396 -9180
rect 11528 -8924 11574 -8912
rect 11528 -9180 11534 -8924
rect 11568 -9180 11574 -8924
rect 11528 -9192 11574 -9180
rect 11642 -8924 11688 -8912
rect 11642 -9180 11648 -8924
rect 11682 -9180 11688 -8924
rect 11642 -9192 11688 -9180
rect 11820 -8924 11866 -8912
rect 11820 -9180 11826 -8924
rect 11860 -9180 11866 -8924
rect 11820 -9192 11866 -9180
rect 11934 -8924 11980 -8912
rect 11934 -9180 11940 -8924
rect 11974 -9180 11980 -8924
rect 11934 -9192 11980 -9180
rect 12112 -8924 12158 -8912
rect 12112 -9180 12118 -8924
rect 12152 -9180 12158 -8924
rect 12112 -9192 12158 -9180
rect 12226 -8924 12272 -8912
rect 12226 -9180 12232 -8924
rect 12266 -9180 12272 -8924
rect 12226 -9192 12272 -9180
rect 12404 -8924 12450 -8912
rect 12404 -9180 12410 -8924
rect 12444 -9180 12450 -8924
rect 12404 -9192 12450 -9180
rect 12518 -8924 12564 -8912
rect 12518 -9180 12524 -8924
rect 12558 -9180 12564 -8924
rect 12518 -9192 12564 -9180
rect 12696 -8924 12742 -8912
rect 12696 -9180 12702 -8924
rect 12736 -9180 12742 -8924
rect 12696 -9192 12742 -9180
rect 9072 -9200 9148 -9194
rect 9072 -9234 9088 -9200
rect 9132 -9234 9148 -9200
rect 9072 -9250 9148 -9234
rect 9250 -9200 9326 -9194
rect 9250 -9234 9266 -9200
rect 9310 -9234 9326 -9200
rect 9250 -9250 9326 -9234
rect 10772 -9230 10806 -9192
rect 10840 -9230 10916 -9224
rect 10950 -9230 10984 -9192
rect 10772 -9264 10856 -9230
rect 10900 -9264 10984 -9230
rect 10840 -9280 10916 -9264
rect 10861 -9594 10895 -9280
rect 11063 -9387 11097 -9192
rect 11132 -9230 11208 -9224
rect 11132 -9264 11148 -9230
rect 11192 -9264 11208 -9230
rect 11132 -9280 11208 -9264
rect 11154 -9374 11188 -9280
rect 11134 -9387 11144 -9374
rect 11063 -9421 11144 -9387
rect 11134 -9427 11144 -9421
rect 11197 -9427 11207 -9374
rect 11154 -9594 11188 -9427
rect 10840 -9610 10916 -9594
rect 10840 -9644 10856 -9610
rect 10900 -9644 10916 -9610
rect 10840 -9650 10916 -9644
rect 11132 -9610 11208 -9594
rect 11132 -9644 11148 -9610
rect 11192 -9644 11208 -9610
rect 11132 -9650 11208 -9644
rect 11242 -9682 11276 -9192
rect 11424 -9230 11500 -9224
rect 11424 -9264 11440 -9230
rect 11484 -9264 11500 -9230
rect 11424 -9280 11500 -9264
rect 11445 -9375 11479 -9280
rect 11426 -9428 11436 -9375
rect 11489 -9428 11499 -9375
rect 11445 -9594 11479 -9428
rect 11424 -9610 11500 -9594
rect 11424 -9644 11440 -9610
rect 11484 -9644 11500 -9610
rect 11424 -9650 11500 -9644
rect 11534 -9682 11568 -9192
rect 11716 -9230 11792 -9224
rect 11716 -9264 11732 -9230
rect 11776 -9264 11792 -9230
rect 11716 -9280 11792 -9264
rect 11738 -9375 11772 -9280
rect 11718 -9428 11728 -9375
rect 11781 -9428 11791 -9375
rect 11738 -9594 11772 -9428
rect 11716 -9610 11792 -9594
rect 11716 -9644 11732 -9610
rect 11776 -9644 11792 -9610
rect 11716 -9650 11792 -9644
rect 11825 -9682 11859 -9192
rect 12008 -9230 12084 -9224
rect 12008 -9264 12024 -9230
rect 12068 -9264 12084 -9230
rect 12008 -9280 12084 -9264
rect 12030 -9376 12064 -9280
rect 12010 -9429 12020 -9376
rect 12073 -9429 12083 -9376
rect 12030 -9594 12064 -9429
rect 12008 -9610 12084 -9594
rect 12008 -9644 12024 -9610
rect 12068 -9644 12084 -9610
rect 12008 -9650 12084 -9644
rect 12118 -9682 12152 -9192
rect 12300 -9230 12376 -9224
rect 12300 -9264 12316 -9230
rect 12360 -9264 12376 -9230
rect 12300 -9280 12376 -9264
rect 12321 -9375 12355 -9280
rect 12302 -9428 12312 -9375
rect 12365 -9428 12375 -9375
rect 12321 -9594 12355 -9428
rect 12300 -9610 12376 -9594
rect 12300 -9644 12316 -9610
rect 12360 -9644 12376 -9610
rect 12300 -9650 12376 -9644
rect 12410 -9682 12444 -9192
rect 12592 -9230 12668 -9224
rect 12592 -9264 12608 -9230
rect 12652 -9264 12668 -9230
rect 12592 -9280 12668 -9264
rect 12613 -9594 12647 -9280
rect 12592 -9610 12668 -9594
rect 12525 -9644 12608 -9610
rect 12652 -9644 12736 -9610
rect 12525 -9682 12559 -9644
rect 12592 -9650 12668 -9644
rect 12702 -9682 12736 -9644
rect 10766 -9694 10812 -9682
rect 9072 -9709 9148 -9694
rect 9250 -9709 9326 -9694
rect 9004 -9710 9394 -9709
rect 9004 -9743 9088 -9710
rect 9004 -9782 9038 -9743
rect 9072 -9744 9088 -9743
rect 9132 -9743 9266 -9710
rect 9132 -9744 9148 -9743
rect 9072 -9750 9148 -9744
rect 9182 -9782 9216 -9743
rect 9250 -9744 9266 -9743
rect 9310 -9743 9394 -9710
rect 9310 -9744 9326 -9743
rect 9250 -9750 9326 -9744
rect 9360 -9782 9394 -9743
rect 6506 -9794 6552 -9782
rect 5327 -9978 5337 -9925
rect 5390 -9978 5400 -9925
rect 6506 -10050 6512 -9794
rect 6546 -10050 6552 -9794
rect 6506 -10062 6552 -10050
rect 6684 -9794 6730 -9782
rect 6684 -10050 6690 -9794
rect 6724 -10050 6730 -9794
rect 6684 -10062 6730 -10050
rect 6862 -9794 6908 -9782
rect 6862 -10050 6868 -9794
rect 6902 -10050 6908 -9794
rect 6862 -10062 6908 -10050
rect 7040 -9794 7086 -9782
rect 7040 -10050 7046 -9794
rect 7080 -10050 7086 -9794
rect 7040 -10062 7086 -10050
rect 7218 -9794 7264 -9782
rect 7218 -10050 7224 -9794
rect 7258 -10050 7264 -9794
rect 7218 -10062 7264 -10050
rect 7396 -9794 7442 -9782
rect 7396 -10050 7402 -9794
rect 7436 -10050 7442 -9794
rect 7396 -10062 7442 -10050
rect 7574 -9794 7620 -9782
rect 7574 -10050 7580 -9794
rect 7614 -10050 7620 -9794
rect 7574 -10062 7620 -10050
rect 7752 -9794 7798 -9782
rect 7752 -10050 7758 -9794
rect 7792 -10050 7798 -9794
rect 7752 -10062 7798 -10050
rect 7930 -9794 7976 -9782
rect 7930 -10050 7936 -9794
rect 7970 -10050 7976 -9794
rect 7930 -10062 7976 -10050
rect 8108 -9794 8154 -9782
rect 8108 -10050 8114 -9794
rect 8148 -10050 8154 -9794
rect 8108 -10062 8154 -10050
rect 8286 -9794 8332 -9782
rect 8286 -10050 8292 -9794
rect 8326 -10050 8332 -9794
rect 8286 -10062 8332 -10050
rect 8464 -9794 8510 -9782
rect 8464 -10050 8470 -9794
rect 8504 -10050 8510 -9794
rect 8464 -10062 8510 -10050
rect 8642 -9794 8688 -9782
rect 8642 -10050 8648 -9794
rect 8682 -10050 8688 -9794
rect 8642 -10062 8688 -10050
rect 8820 -9794 8866 -9782
rect 8820 -10050 8826 -9794
rect 8860 -10050 8866 -9794
rect 8820 -10062 8866 -10050
rect 8998 -9794 9044 -9782
rect 8998 -10050 9004 -9794
rect 9038 -10050 9044 -9794
rect 8998 -10062 9044 -10050
rect 9176 -9794 9222 -9782
rect 9176 -10050 9182 -9794
rect 9216 -10050 9222 -9794
rect 9176 -10062 9222 -10050
rect 9354 -9794 9400 -9782
rect 9354 -10050 9360 -9794
rect 9394 -10050 9400 -9794
rect 10766 -9950 10772 -9694
rect 10806 -9950 10812 -9694
rect 10766 -9962 10812 -9950
rect 10944 -9694 10990 -9682
rect 10944 -9950 10950 -9694
rect 10984 -9950 10990 -9694
rect 10944 -9962 10990 -9950
rect 11058 -9694 11104 -9682
rect 11058 -9950 11064 -9694
rect 11098 -9950 11104 -9694
rect 11058 -9962 11104 -9950
rect 11236 -9694 11282 -9682
rect 11236 -9950 11242 -9694
rect 11276 -9950 11282 -9694
rect 11236 -9962 11282 -9950
rect 11350 -9694 11396 -9682
rect 11350 -9950 11356 -9694
rect 11390 -9950 11396 -9694
rect 11350 -9962 11396 -9950
rect 11528 -9694 11574 -9682
rect 11528 -9950 11534 -9694
rect 11568 -9950 11574 -9694
rect 11528 -9962 11574 -9950
rect 11642 -9694 11688 -9682
rect 11642 -9950 11648 -9694
rect 11682 -9950 11688 -9694
rect 11642 -9962 11688 -9950
rect 11820 -9694 11866 -9682
rect 11820 -9950 11826 -9694
rect 11860 -9950 11866 -9694
rect 11820 -9962 11866 -9950
rect 11934 -9694 11980 -9682
rect 11934 -9950 11940 -9694
rect 11974 -9950 11980 -9694
rect 11934 -9962 11980 -9950
rect 12112 -9694 12158 -9682
rect 12112 -9950 12118 -9694
rect 12152 -9950 12158 -9694
rect 12112 -9962 12158 -9950
rect 12226 -9694 12272 -9682
rect 12226 -9950 12232 -9694
rect 12266 -9950 12272 -9694
rect 12226 -9962 12272 -9950
rect 12404 -9694 12450 -9682
rect 12404 -9950 12410 -9694
rect 12444 -9950 12450 -9694
rect 12404 -9962 12450 -9950
rect 12518 -9694 12564 -9682
rect 12518 -9950 12524 -9694
rect 12558 -9950 12564 -9694
rect 12518 -9962 12564 -9950
rect 12696 -9694 12742 -9682
rect 12696 -9950 12702 -9694
rect 12736 -9950 12742 -9694
rect 12696 -9962 12742 -9950
rect 10773 -10001 10807 -9962
rect 10840 -10000 10916 -9994
rect 10840 -10001 10856 -10000
rect 10773 -10034 10856 -10001
rect 10900 -10001 10916 -10000
rect 10951 -10001 10985 -9962
rect 10900 -10034 10985 -10001
rect 10773 -10035 10985 -10034
rect 10840 -10050 10916 -10035
rect 9354 -10062 9400 -10050
rect 6513 -10099 6547 -10062
rect 6580 -10099 6656 -10094
rect 6690 -10099 6724 -10062
rect 6513 -10100 6724 -10099
rect 6513 -10133 6596 -10100
rect 6580 -10134 6596 -10133
rect 6640 -10133 6724 -10100
rect 6640 -10134 6656 -10133
rect 6580 -10150 6656 -10134
rect 6690 -10313 6724 -10133
rect 6758 -10100 6834 -10094
rect 6758 -10134 6774 -10100
rect 6818 -10134 6834 -10100
rect 6758 -10150 6834 -10134
rect 6670 -10366 6680 -10313
rect 6733 -10366 6743 -10313
rect 6868 -10467 6902 -10062
rect 6936 -10100 7012 -10094
rect 6936 -10134 6952 -10100
rect 6996 -10134 7012 -10100
rect 6936 -10150 7012 -10134
rect 6848 -10520 6858 -10467
rect 6911 -10520 6921 -10467
rect 6580 -10610 6656 -10594
rect 6580 -10644 6596 -10610
rect 6640 -10644 6656 -10610
rect 6580 -10650 6656 -10644
rect 6758 -10610 6834 -10594
rect 6758 -10644 6774 -10610
rect 6818 -10644 6834 -10610
rect 6758 -10650 6834 -10644
rect 6868 -10682 6902 -10520
rect 6958 -10594 6992 -10150
rect 6936 -10610 7012 -10594
rect 6936 -10644 6952 -10610
rect 6996 -10644 7012 -10610
rect 6936 -10650 7012 -10644
rect 7046 -10682 7080 -10062
rect 7114 -10100 7190 -10094
rect 7114 -10134 7130 -10100
rect 7174 -10134 7190 -10100
rect 7114 -10150 7190 -10134
rect 7136 -10594 7170 -10150
rect 7224 -10466 7258 -10062
rect 7292 -10100 7368 -10094
rect 7292 -10134 7308 -10100
rect 7352 -10134 7368 -10100
rect 7292 -10150 7368 -10134
rect 7204 -10519 7214 -10466
rect 7267 -10519 7277 -10466
rect 7114 -10610 7190 -10594
rect 7114 -10644 7130 -10610
rect 7174 -10644 7190 -10610
rect 7114 -10650 7190 -10644
rect 7224 -10682 7258 -10519
rect 7313 -10594 7347 -10150
rect 7292 -10610 7368 -10594
rect 7292 -10644 7308 -10610
rect 7352 -10644 7368 -10610
rect 7292 -10650 7368 -10644
rect 7402 -10682 7436 -10062
rect 7470 -10100 7546 -10094
rect 7470 -10134 7486 -10100
rect 7530 -10134 7546 -10100
rect 7470 -10150 7546 -10134
rect 7492 -10594 7526 -10150
rect 7580 -10466 7614 -10062
rect 7648 -10100 7724 -10094
rect 7648 -10134 7664 -10100
rect 7708 -10134 7724 -10100
rect 7648 -10150 7724 -10134
rect 7561 -10519 7571 -10466
rect 7624 -10519 7634 -10466
rect 7470 -10610 7546 -10594
rect 7470 -10644 7486 -10610
rect 7530 -10644 7546 -10610
rect 7470 -10650 7546 -10644
rect 7580 -10682 7614 -10519
rect 7669 -10594 7703 -10150
rect 7648 -10610 7724 -10594
rect 7648 -10644 7664 -10610
rect 7708 -10644 7724 -10610
rect 7648 -10650 7724 -10644
rect 7758 -10682 7792 -10062
rect 7826 -10100 7902 -10094
rect 7826 -10134 7842 -10100
rect 7886 -10134 7902 -10100
rect 7826 -10150 7902 -10134
rect 7847 -10594 7881 -10150
rect 7936 -10466 7970 -10062
rect 8004 -10100 8080 -10094
rect 8004 -10134 8020 -10100
rect 8064 -10134 8080 -10100
rect 8004 -10150 8080 -10134
rect 7917 -10519 7927 -10466
rect 7980 -10519 7990 -10466
rect 7826 -10610 7902 -10594
rect 7826 -10644 7842 -10610
rect 7886 -10644 7902 -10610
rect 7826 -10650 7902 -10644
rect 7936 -10682 7970 -10519
rect 8025 -10594 8059 -10150
rect 8004 -10610 8080 -10594
rect 8004 -10644 8020 -10610
rect 8064 -10644 8080 -10610
rect 8004 -10650 8080 -10644
rect 8113 -10682 8147 -10062
rect 8182 -10100 8258 -10094
rect 8182 -10134 8198 -10100
rect 8242 -10134 8258 -10100
rect 8182 -10150 8258 -10134
rect 8203 -10594 8237 -10150
rect 8292 -10467 8326 -10062
rect 8360 -10100 8436 -10094
rect 8360 -10134 8376 -10100
rect 8420 -10134 8436 -10100
rect 8360 -10150 8436 -10134
rect 8273 -10520 8283 -10467
rect 8336 -10520 8346 -10467
rect 8182 -10610 8258 -10594
rect 8182 -10644 8198 -10610
rect 8242 -10644 8258 -10610
rect 8182 -10650 8258 -10644
rect 8292 -10682 8326 -10520
rect 8382 -10594 8416 -10150
rect 8360 -10610 8436 -10594
rect 8360 -10644 8376 -10610
rect 8420 -10644 8436 -10610
rect 8360 -10650 8436 -10644
rect 8470 -10682 8504 -10062
rect 8538 -10100 8614 -10094
rect 8538 -10134 8554 -10100
rect 8598 -10134 8614 -10100
rect 8538 -10150 8614 -10134
rect 8559 -10594 8593 -10150
rect 8648 -10466 8682 -10062
rect 8716 -10100 8792 -10094
rect 8716 -10134 8732 -10100
rect 8776 -10134 8792 -10100
rect 8716 -10150 8792 -10134
rect 8628 -10519 8638 -10466
rect 8691 -10519 8701 -10466
rect 8538 -10610 8614 -10594
rect 8538 -10644 8554 -10610
rect 8598 -10644 8614 -10610
rect 8538 -10650 8614 -10644
rect 8648 -10682 8682 -10519
rect 8737 -10594 8771 -10150
rect 8716 -10610 8792 -10594
rect 8716 -10644 8732 -10610
rect 8776 -10644 8792 -10610
rect 8716 -10650 8792 -10644
rect 8826 -10682 8860 -10062
rect 8894 -10100 8970 -10094
rect 8894 -10134 8910 -10100
rect 8954 -10134 8970 -10100
rect 8894 -10150 8970 -10134
rect 8915 -10594 8949 -10150
rect 9004 -10467 9038 -10062
rect 9072 -10100 9148 -10094
rect 9072 -10134 9088 -10100
rect 9132 -10134 9148 -10100
rect 9072 -10150 9148 -10134
rect 9250 -10100 9326 -10094
rect 9250 -10134 9266 -10100
rect 9310 -10134 9326 -10100
rect 9250 -10150 9326 -10134
rect 9161 -10367 9171 -10314
rect 9224 -10367 9234 -10314
rect 10862 -10364 10896 -10050
rect 8985 -10520 8995 -10467
rect 9048 -10520 9058 -10467
rect 8894 -10610 8970 -10594
rect 8894 -10644 8910 -10610
rect 8954 -10644 8970 -10610
rect 8894 -10650 8970 -10644
rect 9004 -10682 9038 -10520
rect 9072 -10610 9148 -10594
rect 9072 -10644 9088 -10610
rect 9132 -10644 9148 -10610
rect 9072 -10650 9148 -10644
rect 9181 -10614 9215 -10367
rect 10840 -10380 10916 -10364
rect 10772 -10414 10856 -10380
rect 10900 -10414 10986 -10380
rect 10772 -10452 10806 -10414
rect 10840 -10420 10916 -10414
rect 10952 -10452 10986 -10414
rect 11063 -10452 11097 -9962
rect 11132 -10000 11208 -9994
rect 11132 -10034 11148 -10000
rect 11192 -10034 11208 -10000
rect 11132 -10050 11208 -10034
rect 11153 -10364 11187 -10050
rect 11132 -10380 11208 -10364
rect 11132 -10414 11148 -10380
rect 11192 -10414 11208 -10380
rect 11132 -10420 11208 -10414
rect 11356 -10452 11390 -9962
rect 11424 -10000 11500 -9994
rect 11424 -10034 11440 -10000
rect 11484 -10034 11500 -10000
rect 11424 -10050 11500 -10034
rect 11446 -10364 11480 -10050
rect 11424 -10380 11500 -10364
rect 11424 -10414 11440 -10380
rect 11484 -10414 11500 -10380
rect 11424 -10420 11500 -10414
rect 11648 -10452 11682 -9962
rect 11716 -10000 11792 -9994
rect 11716 -10034 11732 -10000
rect 11776 -10034 11792 -10000
rect 11716 -10050 11792 -10034
rect 11737 -10364 11771 -10050
rect 11716 -10380 11792 -10364
rect 11716 -10414 11732 -10380
rect 11776 -10414 11792 -10380
rect 11716 -10420 11792 -10414
rect 11940 -10452 11974 -9962
rect 12008 -10000 12084 -9994
rect 12008 -10034 12024 -10000
rect 12068 -10034 12084 -10000
rect 12008 -10050 12084 -10034
rect 12028 -10364 12062 -10050
rect 12008 -10380 12084 -10364
rect 12008 -10414 12024 -10380
rect 12068 -10414 12084 -10380
rect 12008 -10420 12084 -10414
rect 12232 -10452 12266 -9962
rect 12300 -10000 12376 -9994
rect 12300 -10034 12316 -10000
rect 12360 -10034 12376 -10000
rect 12300 -10050 12376 -10034
rect 12592 -10000 12668 -9994
rect 12592 -10034 12608 -10000
rect 12652 -10034 12668 -10000
rect 12592 -10050 12668 -10034
rect 12320 -10364 12354 -10050
rect 12613 -10364 12647 -10050
rect 12300 -10380 12376 -10364
rect 12300 -10414 12316 -10380
rect 12360 -10414 12376 -10380
rect 12300 -10420 12376 -10414
rect 12592 -10380 12668 -10364
rect 12592 -10414 12608 -10380
rect 12652 -10414 12668 -10380
rect 12592 -10420 12668 -10414
rect 10766 -10464 10812 -10452
rect 9250 -10610 9326 -10594
rect 9250 -10614 9266 -10610
rect 9181 -10644 9266 -10614
rect 9310 -10614 9326 -10610
rect 9310 -10644 9393 -10614
rect 9181 -10648 9393 -10644
rect 9181 -10682 9215 -10648
rect 9250 -10650 9326 -10648
rect 9359 -10682 9393 -10648
rect 6506 -10694 6552 -10682
rect 6506 -10950 6512 -10694
rect 6546 -10950 6552 -10694
rect 6506 -10962 6552 -10950
rect 6684 -10694 6730 -10682
rect 6684 -10950 6690 -10694
rect 6724 -10950 6730 -10694
rect 6684 -10962 6730 -10950
rect 6862 -10694 6908 -10682
rect 6862 -10950 6868 -10694
rect 6902 -10950 6908 -10694
rect 6862 -10962 6908 -10950
rect 7040 -10694 7086 -10682
rect 7040 -10950 7046 -10694
rect 7080 -10950 7086 -10694
rect 7040 -10962 7086 -10950
rect 7218 -10694 7264 -10682
rect 7218 -10950 7224 -10694
rect 7258 -10950 7264 -10694
rect 7218 -10962 7264 -10950
rect 7396 -10694 7442 -10682
rect 7396 -10950 7402 -10694
rect 7436 -10950 7442 -10694
rect 7396 -10962 7442 -10950
rect 7574 -10694 7620 -10682
rect 7574 -10950 7580 -10694
rect 7614 -10950 7620 -10694
rect 7574 -10962 7620 -10950
rect 7752 -10694 7798 -10682
rect 7752 -10950 7758 -10694
rect 7792 -10950 7798 -10694
rect 7752 -10962 7798 -10950
rect 7930 -10694 7976 -10682
rect 7930 -10950 7936 -10694
rect 7970 -10950 7976 -10694
rect 7930 -10962 7976 -10950
rect 8108 -10694 8154 -10682
rect 8108 -10950 8114 -10694
rect 8148 -10950 8154 -10694
rect 8108 -10962 8154 -10950
rect 8286 -10694 8332 -10682
rect 8286 -10950 8292 -10694
rect 8326 -10950 8332 -10694
rect 8286 -10962 8332 -10950
rect 8464 -10694 8510 -10682
rect 8464 -10950 8470 -10694
rect 8504 -10950 8510 -10694
rect 8464 -10962 8510 -10950
rect 8642 -10694 8688 -10682
rect 8642 -10950 8648 -10694
rect 8682 -10950 8688 -10694
rect 8642 -10962 8688 -10950
rect 8820 -10694 8866 -10682
rect 8820 -10950 8826 -10694
rect 8860 -10950 8866 -10694
rect 8820 -10962 8866 -10950
rect 8998 -10694 9044 -10682
rect 8998 -10950 9004 -10694
rect 9038 -10950 9044 -10694
rect 8998 -10962 9044 -10950
rect 9176 -10694 9222 -10682
rect 9176 -10950 9182 -10694
rect 9216 -10950 9222 -10694
rect 9176 -10962 9222 -10950
rect 9354 -10694 9400 -10682
rect 9354 -10950 9360 -10694
rect 9394 -10950 9400 -10694
rect 10766 -10720 10772 -10464
rect 10806 -10720 10812 -10464
rect 10766 -10732 10812 -10720
rect 10944 -10464 10990 -10452
rect 10944 -10720 10950 -10464
rect 10984 -10720 10990 -10464
rect 10944 -10732 10990 -10720
rect 11058 -10464 11104 -10452
rect 11058 -10720 11064 -10464
rect 11098 -10720 11104 -10464
rect 11058 -10732 11104 -10720
rect 11236 -10464 11282 -10452
rect 11236 -10720 11242 -10464
rect 11276 -10720 11282 -10464
rect 11236 -10732 11282 -10720
rect 11350 -10464 11396 -10452
rect 11350 -10720 11356 -10464
rect 11390 -10720 11396 -10464
rect 11350 -10732 11396 -10720
rect 11528 -10464 11574 -10452
rect 11528 -10720 11534 -10464
rect 11568 -10720 11574 -10464
rect 11528 -10732 11574 -10720
rect 11642 -10464 11688 -10452
rect 11642 -10720 11648 -10464
rect 11682 -10720 11688 -10464
rect 11642 -10732 11688 -10720
rect 11820 -10464 11866 -10452
rect 11820 -10720 11826 -10464
rect 11860 -10720 11866 -10464
rect 11820 -10732 11866 -10720
rect 11934 -10464 11980 -10452
rect 11934 -10720 11940 -10464
rect 11974 -10720 11980 -10464
rect 11934 -10732 11980 -10720
rect 12112 -10464 12158 -10452
rect 12112 -10720 12118 -10464
rect 12152 -10720 12158 -10464
rect 12112 -10732 12158 -10720
rect 12226 -10464 12272 -10452
rect 12226 -10720 12232 -10464
rect 12266 -10720 12272 -10464
rect 12226 -10732 12272 -10720
rect 12404 -10464 12450 -10452
rect 12404 -10720 12410 -10464
rect 12444 -10720 12450 -10464
rect 12404 -10732 12450 -10720
rect 12518 -10464 12564 -10452
rect 12518 -10720 12524 -10464
rect 12558 -10720 12564 -10464
rect 12518 -10732 12564 -10720
rect 12696 -10464 12742 -10452
rect 12696 -10720 12702 -10464
rect 12736 -10720 12742 -10464
rect 12696 -10732 12742 -10720
rect 10840 -10770 10916 -10764
rect 10840 -10804 10856 -10770
rect 10900 -10804 10916 -10770
rect 10840 -10820 10916 -10804
rect 11132 -10770 11208 -10764
rect 11132 -10804 11148 -10770
rect 11192 -10804 11208 -10770
rect 11132 -10820 11208 -10804
rect 9354 -10962 9400 -10950
rect 6510 -11003 6544 -10962
rect 6580 -11000 6656 -10994
rect 6580 -11003 6596 -11000
rect 6510 -11034 6596 -11003
rect 6640 -11003 6656 -11000
rect 6688 -11003 6722 -10962
rect 6758 -11000 6834 -10994
rect 6758 -11003 6774 -11000
rect 6640 -11034 6774 -11003
rect 6818 -11003 6834 -11000
rect 6868 -11003 6902 -10962
rect 6818 -11034 6902 -11003
rect 6510 -11037 6902 -11034
rect 6580 -11050 6656 -11037
rect 6758 -11050 6834 -11037
rect 6580 -11510 6656 -11494
rect 6580 -11544 6596 -11510
rect 6640 -11544 6656 -11510
rect 6580 -11550 6656 -11544
rect 6758 -11510 6834 -11494
rect 6758 -11544 6774 -11510
rect 6818 -11544 6834 -11510
rect 6758 -11550 6834 -11544
rect 6868 -11582 6902 -11037
rect 6936 -11000 7012 -10994
rect 6936 -11034 6952 -11000
rect 6996 -11034 7012 -11000
rect 6936 -11050 7012 -11034
rect 6958 -11494 6992 -11050
rect 7046 -11366 7080 -10962
rect 7114 -11000 7190 -10994
rect 7114 -11034 7130 -11000
rect 7174 -11034 7190 -11000
rect 7114 -11050 7190 -11034
rect 7027 -11419 7037 -11366
rect 7090 -11419 7100 -11366
rect 6936 -11510 7012 -11494
rect 6936 -11544 6952 -11510
rect 6996 -11544 7012 -11510
rect 6936 -11550 7012 -11544
rect 7046 -11582 7080 -11419
rect 7135 -11494 7169 -11050
rect 7114 -11510 7190 -11494
rect 7114 -11544 7130 -11510
rect 7174 -11544 7190 -11510
rect 7114 -11550 7190 -11544
rect 7224 -11582 7258 -10962
rect 7313 -10994 7347 -10993
rect 7292 -11000 7368 -10994
rect 7292 -11034 7308 -11000
rect 7352 -11034 7368 -11000
rect 7292 -11050 7368 -11034
rect 7313 -11494 7347 -11050
rect 7402 -11366 7436 -10962
rect 7491 -10994 7525 -10993
rect 7470 -11000 7546 -10994
rect 7470 -11034 7486 -11000
rect 7530 -11034 7546 -11000
rect 7470 -11050 7546 -11034
rect 7383 -11419 7393 -11366
rect 7446 -11419 7456 -11366
rect 7292 -11510 7368 -11494
rect 7292 -11544 7308 -11510
rect 7352 -11544 7368 -11510
rect 7292 -11550 7368 -11544
rect 7402 -11582 7436 -11419
rect 7491 -11494 7525 -11050
rect 7470 -11510 7546 -11494
rect 7470 -11544 7486 -11510
rect 7530 -11544 7546 -11510
rect 7470 -11550 7546 -11544
rect 7580 -11582 7614 -10962
rect 7669 -10994 7703 -10993
rect 7648 -11000 7724 -10994
rect 7648 -11034 7664 -11000
rect 7708 -11034 7724 -11000
rect 7648 -11050 7724 -11034
rect 7669 -11494 7703 -11050
rect 7758 -11367 7792 -10962
rect 7848 -10994 7882 -10993
rect 7826 -11000 7902 -10994
rect 7826 -11034 7842 -11000
rect 7886 -11034 7902 -11000
rect 7826 -11050 7902 -11034
rect 7738 -11420 7748 -11367
rect 7801 -11420 7811 -11367
rect 7648 -11510 7724 -11494
rect 7648 -11544 7664 -11510
rect 7708 -11544 7724 -11510
rect 7648 -11550 7724 -11544
rect 7758 -11582 7792 -11420
rect 7848 -11494 7882 -11050
rect 7826 -11510 7902 -11494
rect 7826 -11544 7842 -11510
rect 7886 -11544 7902 -11510
rect 7826 -11550 7902 -11544
rect 7936 -11582 7970 -10962
rect 8004 -11000 8080 -10994
rect 8004 -11034 8020 -11000
rect 8064 -11034 8080 -11000
rect 8004 -11050 8080 -11034
rect 8024 -11494 8058 -11050
rect 8113 -11366 8147 -10962
rect 8182 -11000 8258 -10994
rect 8182 -11034 8198 -11000
rect 8242 -11034 8258 -11000
rect 8182 -11050 8258 -11034
rect 8093 -11419 8103 -11366
rect 8156 -11419 8166 -11366
rect 8004 -11510 8080 -11494
rect 8004 -11544 8020 -11510
rect 8064 -11544 8080 -11510
rect 8004 -11550 8080 -11544
rect 8113 -11582 8147 -11419
rect 8203 -11494 8237 -11050
rect 8182 -11510 8258 -11494
rect 8182 -11544 8198 -11510
rect 8242 -11544 8258 -11510
rect 8182 -11550 8258 -11544
rect 8292 -11582 8326 -10962
rect 8360 -11000 8436 -10994
rect 8360 -11034 8376 -11000
rect 8420 -11034 8436 -11000
rect 8360 -11050 8436 -11034
rect 8381 -11494 8415 -11050
rect 8470 -11366 8504 -10962
rect 8538 -11000 8614 -10994
rect 8538 -11034 8554 -11000
rect 8598 -11034 8614 -11000
rect 8538 -11050 8614 -11034
rect 8451 -11419 8461 -11366
rect 8514 -11419 8524 -11366
rect 8360 -11510 8436 -11494
rect 8360 -11544 8376 -11510
rect 8420 -11544 8436 -11510
rect 8360 -11550 8436 -11544
rect 8470 -11582 8504 -11419
rect 8559 -11494 8593 -11050
rect 8538 -11510 8614 -11494
rect 8538 -11544 8554 -11510
rect 8598 -11544 8614 -11510
rect 8538 -11550 8614 -11544
rect 8648 -11582 8682 -10962
rect 8716 -11000 8792 -10994
rect 8716 -11034 8732 -11000
rect 8776 -11034 8792 -11000
rect 8716 -11050 8792 -11034
rect 8737 -11494 8771 -11050
rect 8826 -11366 8860 -10962
rect 8894 -11000 8970 -10994
rect 8894 -11034 8910 -11000
rect 8954 -11034 8970 -11000
rect 8894 -11050 8970 -11034
rect 8807 -11419 8817 -11366
rect 8870 -11419 8880 -11366
rect 8716 -11510 8792 -11494
rect 8716 -11544 8732 -11510
rect 8776 -11544 8792 -11510
rect 8716 -11550 8792 -11544
rect 8826 -11582 8860 -11419
rect 8915 -11494 8949 -11050
rect 8894 -11510 8970 -11494
rect 8894 -11544 8910 -11510
rect 8954 -11544 8970 -11510
rect 8894 -11550 8970 -11544
rect 9004 -11582 9038 -10962
rect 9072 -11000 9148 -10994
rect 9072 -11034 9088 -11000
rect 9132 -11034 9148 -11000
rect 9072 -11050 9148 -11034
rect 9250 -11000 9326 -10994
rect 9250 -11034 9266 -11000
rect 9310 -11034 9326 -11000
rect 9250 -11050 9326 -11034
rect 9093 -11494 9127 -11050
rect 10860 -11134 10894 -10820
rect 11152 -11134 11186 -10820
rect 10772 -11149 10806 -11148
rect 10840 -11149 10916 -11134
rect 10772 -11150 10986 -11149
rect 10772 -11183 10856 -11150
rect 10772 -11222 10806 -11183
rect 10840 -11184 10856 -11183
rect 10900 -11183 10986 -11150
rect 10900 -11184 10916 -11183
rect 10840 -11190 10916 -11184
rect 10952 -11222 10986 -11183
rect 11132 -11150 11208 -11134
rect 11132 -11184 11148 -11150
rect 11192 -11184 11208 -11150
rect 11132 -11190 11208 -11184
rect 11244 -11222 11278 -10732
rect 11424 -10770 11500 -10764
rect 11424 -10804 11440 -10770
rect 11484 -10804 11500 -10770
rect 11424 -10820 11500 -10804
rect 11446 -11134 11480 -10820
rect 11424 -11150 11500 -11134
rect 11424 -11184 11440 -11150
rect 11484 -11184 11500 -11150
rect 11424 -11190 11500 -11184
rect 11534 -11222 11568 -10732
rect 11716 -10770 11792 -10764
rect 11716 -10804 11732 -10770
rect 11776 -10804 11792 -10770
rect 11716 -10820 11792 -10804
rect 11737 -11134 11771 -10820
rect 11716 -11150 11792 -11134
rect 11716 -11184 11732 -11150
rect 11776 -11184 11792 -11150
rect 11716 -11190 11792 -11184
rect 11826 -11222 11860 -10732
rect 12008 -10770 12084 -10764
rect 12008 -10804 12024 -10770
rect 12068 -10804 12084 -10770
rect 12008 -10820 12084 -10804
rect 12029 -11134 12063 -10820
rect 12008 -11150 12084 -11134
rect 12008 -11184 12024 -11150
rect 12068 -11184 12084 -11150
rect 12008 -11190 12084 -11184
rect 12118 -11222 12152 -10732
rect 12300 -10770 12376 -10764
rect 12300 -10804 12316 -10770
rect 12360 -10804 12376 -10770
rect 12300 -10820 12376 -10804
rect 12322 -11134 12356 -10820
rect 12300 -11150 12376 -11134
rect 12300 -11184 12316 -11150
rect 12360 -11184 12376 -11150
rect 12300 -11190 12376 -11184
rect 12410 -11222 12444 -10732
rect 12525 -10772 12559 -10732
rect 12592 -10770 12668 -10764
rect 12592 -10772 12608 -10770
rect 12525 -10804 12608 -10772
rect 12652 -10772 12668 -10770
rect 12700 -10772 12734 -10732
rect 12652 -10804 12734 -10772
rect 12525 -10806 12734 -10804
rect 12592 -10820 12668 -10806
rect 12613 -11134 12647 -10820
rect 12592 -11150 12668 -11134
rect 12592 -11184 12608 -11150
rect 12652 -11184 12668 -11150
rect 12592 -11190 12668 -11184
rect 10766 -11234 10812 -11222
rect 10766 -11490 10772 -11234
rect 10806 -11490 10812 -11234
rect 9072 -11510 9148 -11494
rect 9250 -11510 9326 -11494
rect 10766 -11502 10812 -11490
rect 10944 -11234 10990 -11222
rect 10944 -11490 10950 -11234
rect 10984 -11490 10990 -11234
rect 10944 -11502 10990 -11490
rect 11058 -11234 11104 -11222
rect 11058 -11490 11064 -11234
rect 11098 -11490 11104 -11234
rect 11058 -11502 11104 -11490
rect 11236 -11234 11282 -11222
rect 11236 -11490 11242 -11234
rect 11276 -11490 11282 -11234
rect 11236 -11502 11282 -11490
rect 11350 -11234 11396 -11222
rect 11350 -11490 11356 -11234
rect 11390 -11490 11396 -11234
rect 11350 -11502 11396 -11490
rect 11528 -11234 11574 -11222
rect 11528 -11490 11534 -11234
rect 11568 -11490 11574 -11234
rect 11528 -11502 11574 -11490
rect 11642 -11234 11688 -11222
rect 11642 -11490 11648 -11234
rect 11682 -11490 11688 -11234
rect 11642 -11502 11688 -11490
rect 11820 -11234 11866 -11222
rect 11820 -11490 11826 -11234
rect 11860 -11490 11866 -11234
rect 11820 -11502 11866 -11490
rect 11934 -11234 11980 -11222
rect 11934 -11490 11940 -11234
rect 11974 -11490 11980 -11234
rect 11934 -11502 11980 -11490
rect 12112 -11234 12158 -11222
rect 12112 -11490 12118 -11234
rect 12152 -11490 12158 -11234
rect 12112 -11502 12158 -11490
rect 12226 -11234 12272 -11222
rect 12226 -11490 12232 -11234
rect 12266 -11490 12272 -11234
rect 12226 -11502 12272 -11490
rect 12404 -11234 12450 -11222
rect 12404 -11490 12410 -11234
rect 12444 -11490 12450 -11234
rect 12404 -11502 12450 -11490
rect 12518 -11234 12564 -11222
rect 12518 -11490 12524 -11234
rect 12558 -11490 12564 -11234
rect 12518 -11502 12564 -11490
rect 12696 -11234 12742 -11222
rect 12696 -11490 12702 -11234
rect 12736 -11490 12742 -11234
rect 12696 -11502 12742 -11490
rect 9072 -11544 9088 -11510
rect 9132 -11544 9148 -11510
rect 9072 -11550 9148 -11544
rect 9182 -11544 9266 -11510
rect 9310 -11544 9394 -11510
rect 9182 -11582 9216 -11544
rect 9250 -11550 9326 -11544
rect 9360 -11582 9394 -11544
rect 10840 -11540 10916 -11534
rect 10840 -11574 10856 -11540
rect 10900 -11574 10916 -11540
rect 6506 -11594 6552 -11582
rect 6506 -11850 6512 -11594
rect 6546 -11850 6552 -11594
rect 6506 -11862 6552 -11850
rect 6684 -11594 6730 -11582
rect 6684 -11850 6690 -11594
rect 6724 -11850 6730 -11594
rect 6684 -11862 6730 -11850
rect 6862 -11594 6908 -11582
rect 6862 -11850 6868 -11594
rect 6902 -11850 6908 -11594
rect 6862 -11862 6908 -11850
rect 7040 -11594 7086 -11582
rect 7040 -11850 7046 -11594
rect 7080 -11850 7086 -11594
rect 7040 -11862 7086 -11850
rect 7218 -11594 7264 -11582
rect 7218 -11850 7224 -11594
rect 7258 -11850 7264 -11594
rect 7218 -11862 7264 -11850
rect 7396 -11594 7442 -11582
rect 7396 -11850 7402 -11594
rect 7436 -11850 7442 -11594
rect 7396 -11862 7442 -11850
rect 7574 -11594 7620 -11582
rect 7574 -11850 7580 -11594
rect 7614 -11850 7620 -11594
rect 7574 -11862 7620 -11850
rect 7752 -11594 7798 -11582
rect 7752 -11850 7758 -11594
rect 7792 -11850 7798 -11594
rect 7752 -11862 7798 -11850
rect 7930 -11594 7976 -11582
rect 7930 -11850 7936 -11594
rect 7970 -11850 7976 -11594
rect 7930 -11862 7976 -11850
rect 8108 -11594 8154 -11582
rect 8108 -11850 8114 -11594
rect 8148 -11850 8154 -11594
rect 8108 -11862 8154 -11850
rect 8286 -11594 8332 -11582
rect 8286 -11850 8292 -11594
rect 8326 -11850 8332 -11594
rect 8286 -11862 8332 -11850
rect 8464 -11594 8510 -11582
rect 8464 -11850 8470 -11594
rect 8504 -11850 8510 -11594
rect 8464 -11862 8510 -11850
rect 8642 -11594 8688 -11582
rect 8642 -11850 8648 -11594
rect 8682 -11850 8688 -11594
rect 8642 -11862 8688 -11850
rect 8820 -11594 8866 -11582
rect 8820 -11850 8826 -11594
rect 8860 -11850 8866 -11594
rect 8820 -11862 8866 -11850
rect 8998 -11594 9044 -11582
rect 8998 -11850 9004 -11594
rect 9038 -11850 9044 -11594
rect 8998 -11862 9044 -11850
rect 9176 -11594 9222 -11582
rect 9176 -11850 9182 -11594
rect 9216 -11850 9222 -11594
rect 9176 -11862 9222 -11850
rect 9354 -11594 9400 -11582
rect 10840 -11590 10916 -11574
rect 9354 -11850 9360 -11594
rect 9394 -11850 9400 -11594
rect 11063 -11674 11097 -11502
rect 11132 -11540 11208 -11534
rect 11132 -11574 11148 -11540
rect 11192 -11574 11208 -11540
rect 11132 -11590 11208 -11574
rect 11043 -11727 11053 -11674
rect 11106 -11727 11116 -11674
rect 11356 -11675 11390 -11502
rect 11424 -11540 11500 -11534
rect 11424 -11574 11440 -11540
rect 11484 -11574 11500 -11540
rect 11424 -11590 11500 -11574
rect 11648 -11674 11682 -11502
rect 11716 -11540 11792 -11534
rect 11716 -11574 11732 -11540
rect 11776 -11574 11792 -11540
rect 11716 -11590 11792 -11574
rect 11940 -11674 11974 -11502
rect 12008 -11540 12084 -11534
rect 12008 -11574 12024 -11540
rect 12068 -11574 12084 -11540
rect 12008 -11590 12084 -11574
rect 12233 -11674 12267 -11502
rect 12300 -11540 12376 -11534
rect 12300 -11574 12316 -11540
rect 12360 -11574 12376 -11540
rect 12300 -11590 12376 -11574
rect 12525 -11541 12559 -11502
rect 12592 -11540 12668 -11534
rect 12592 -11541 12608 -11540
rect 12525 -11574 12608 -11541
rect 12652 -11541 12668 -11540
rect 12701 -11541 12735 -11502
rect 12652 -11574 12735 -11541
rect 12525 -11575 12735 -11574
rect 12592 -11590 12668 -11575
rect 11337 -11728 11347 -11675
rect 11400 -11728 11410 -11675
rect 11628 -11727 11638 -11674
rect 11691 -11727 11701 -11674
rect 11921 -11727 11931 -11674
rect 11984 -11727 11994 -11674
rect 12213 -11727 12223 -11674
rect 12276 -11727 12286 -11674
rect 13012 -11726 13022 -11673
rect 13075 -11726 13085 -11673
rect 9354 -11862 9400 -11850
rect 6511 -11900 6545 -11862
rect 6580 -11900 6656 -11894
rect 6688 -11900 6722 -11862
rect 6758 -11900 6834 -11894
rect 6868 -11900 6902 -11862
rect 6511 -11934 6596 -11900
rect 6640 -11934 6774 -11900
rect 6818 -11934 6902 -11900
rect 6580 -11950 6656 -11934
rect 6758 -11950 6834 -11934
rect 6868 -12040 6902 -11934
rect 6936 -11900 7012 -11894
rect 6936 -11934 6952 -11900
rect 6996 -11934 7012 -11900
rect 6936 -11950 7012 -11934
rect 7114 -11900 7190 -11894
rect 7114 -11934 7130 -11900
rect 7174 -11934 7190 -11900
rect 7114 -11950 7190 -11934
rect 7224 -12040 7258 -11862
rect 7292 -11900 7368 -11894
rect 7292 -11934 7308 -11900
rect 7352 -11934 7368 -11900
rect 7292 -11950 7368 -11934
rect 7470 -11900 7546 -11894
rect 7470 -11934 7486 -11900
rect 7530 -11934 7546 -11900
rect 7470 -11950 7546 -11934
rect 7580 -12040 7614 -11862
rect 7648 -11900 7724 -11894
rect 7648 -11934 7664 -11900
rect 7708 -11934 7724 -11900
rect 7648 -11950 7724 -11934
rect 7826 -11900 7902 -11894
rect 7826 -11934 7842 -11900
rect 7886 -11934 7902 -11900
rect 7826 -11950 7902 -11934
rect 7936 -12040 7970 -11862
rect 8004 -11900 8080 -11894
rect 8004 -11934 8020 -11900
rect 8064 -11934 8080 -11900
rect 8004 -11950 8080 -11934
rect 8182 -11900 8258 -11894
rect 8182 -11934 8198 -11900
rect 8242 -11934 8258 -11900
rect 8182 -11950 8258 -11934
rect 8292 -12040 8326 -11862
rect 8360 -11900 8436 -11894
rect 8360 -11934 8376 -11900
rect 8420 -11934 8436 -11900
rect 8360 -11950 8436 -11934
rect 8538 -11900 8614 -11894
rect 8538 -11934 8554 -11900
rect 8598 -11934 8614 -11900
rect 8538 -11950 8614 -11934
rect 8648 -12040 8682 -11862
rect 8716 -11900 8792 -11894
rect 8716 -11934 8732 -11900
rect 8776 -11934 8792 -11900
rect 8716 -11950 8792 -11934
rect 8894 -11900 8970 -11894
rect 8894 -11934 8910 -11900
rect 8954 -11934 8970 -11900
rect 8894 -11950 8970 -11934
rect 9072 -11900 9148 -11894
rect 9072 -11934 9088 -11900
rect 9132 -11934 9148 -11900
rect 9072 -11950 9148 -11934
rect 8912 -11985 8946 -11950
rect 9095 -11985 9129 -11950
rect 9182 -11985 9216 -11862
rect 9250 -11900 9326 -11894
rect 9250 -11934 9266 -11900
rect 9310 -11934 9326 -11900
rect 9250 -11950 9326 -11934
rect 8912 -12019 9216 -11985
rect 6868 -12074 8682 -12040
rect 5027 -13349 5037 -13296
rect 5090 -13349 5100 -13296
rect 5524 -13349 5534 -13296
rect 5587 -13349 5597 -13296
rect 5021 -13486 5031 -13433
rect 5084 -13486 5094 -13433
rect 4895 -14598 4905 -14545
rect 4958 -14598 4968 -14545
rect 4229 -14979 4239 -14926
rect 4292 -14979 4302 -14926
rect 3947 -15047 4023 -15032
rect 3879 -15048 4091 -15047
rect 3879 -15081 3963 -15048
rect 3879 -15120 3913 -15081
rect 3947 -15082 3963 -15081
rect 4007 -15081 4091 -15048
rect 4007 -15082 4023 -15081
rect 3947 -15088 4023 -15082
rect 4057 -15120 4091 -15081
rect -2179 -15132 -2133 -15120
rect -2179 -15388 -2173 -15132
rect -2139 -15388 -2133 -15132
rect -2179 -15400 -2133 -15388
rect -2001 -15132 -1955 -15120
rect -2001 -15388 -1995 -15132
rect -1961 -15388 -1955 -15132
rect -2001 -15400 -1955 -15388
rect -1823 -15132 -1777 -15120
rect -1823 -15388 -1817 -15132
rect -1783 -15388 -1777 -15132
rect -1823 -15400 -1777 -15388
rect -1645 -15132 -1599 -15120
rect -1645 -15388 -1639 -15132
rect -1605 -15388 -1599 -15132
rect -1645 -15400 -1599 -15388
rect -1467 -15132 -1421 -15120
rect -1467 -15388 -1461 -15132
rect -1427 -15388 -1421 -15132
rect -1467 -15400 -1421 -15388
rect -1289 -15132 -1243 -15120
rect -1289 -15388 -1283 -15132
rect -1249 -15388 -1243 -15132
rect -1289 -15400 -1243 -15388
rect -1111 -15132 -1065 -15120
rect -1111 -15388 -1105 -15132
rect -1071 -15388 -1065 -15132
rect -1111 -15400 -1065 -15388
rect -933 -15132 -887 -15120
rect -933 -15388 -927 -15132
rect -893 -15388 -887 -15132
rect -933 -15400 -887 -15388
rect -755 -15132 -709 -15120
rect -755 -15388 -749 -15132
rect -715 -15388 -709 -15132
rect -755 -15400 -709 -15388
rect -577 -15132 -531 -15120
rect -577 -15388 -571 -15132
rect -537 -15388 -531 -15132
rect -577 -15400 -531 -15388
rect -399 -15132 -353 -15120
rect -399 -15388 -393 -15132
rect -359 -15388 -353 -15132
rect -399 -15400 -353 -15388
rect -221 -15132 -175 -15120
rect -221 -15388 -215 -15132
rect -181 -15388 -175 -15132
rect -221 -15400 -175 -15388
rect -43 -15132 3 -15120
rect -43 -15388 -37 -15132
rect -3 -15388 3 -15132
rect -43 -15400 3 -15388
rect 135 -15132 181 -15120
rect 135 -15388 141 -15132
rect 175 -15388 181 -15132
rect 135 -15400 181 -15388
rect 313 -15132 359 -15120
rect 313 -15388 319 -15132
rect 353 -15388 359 -15132
rect 313 -15400 359 -15388
rect 491 -15132 537 -15120
rect 491 -15388 497 -15132
rect 531 -15388 537 -15132
rect 491 -15400 537 -15388
rect 669 -15132 715 -15120
rect 669 -15388 675 -15132
rect 709 -15388 715 -15132
rect 669 -15400 715 -15388
rect 847 -15132 893 -15120
rect 847 -15388 853 -15132
rect 887 -15388 893 -15132
rect 847 -15400 893 -15388
rect 1025 -15132 1071 -15120
rect 1025 -15388 1031 -15132
rect 1065 -15388 1071 -15132
rect 1025 -15400 1071 -15388
rect 1203 -15132 1249 -15120
rect 1203 -15388 1209 -15132
rect 1243 -15388 1249 -15132
rect 1203 -15400 1249 -15388
rect 1381 -15132 1427 -15120
rect 1381 -15388 1387 -15132
rect 1421 -15388 1427 -15132
rect 1381 -15400 1427 -15388
rect 1559 -15132 1605 -15120
rect 1559 -15388 1565 -15132
rect 1599 -15388 1605 -15132
rect 1559 -15400 1605 -15388
rect 1737 -15132 1783 -15120
rect 1737 -15388 1743 -15132
rect 1777 -15388 1783 -15132
rect 1737 -15400 1783 -15388
rect 1915 -15132 1961 -15120
rect 1915 -15388 1921 -15132
rect 1955 -15388 1961 -15132
rect 1915 -15400 1961 -15388
rect 2093 -15132 2139 -15120
rect 2093 -15388 2099 -15132
rect 2133 -15388 2139 -15132
rect 2093 -15400 2139 -15388
rect 2271 -15132 2317 -15120
rect 2271 -15388 2277 -15132
rect 2311 -15388 2317 -15132
rect 2271 -15400 2317 -15388
rect 2449 -15132 2495 -15120
rect 2449 -15388 2455 -15132
rect 2489 -15388 2495 -15132
rect 2449 -15400 2495 -15388
rect 2627 -15132 2673 -15120
rect 2627 -15388 2633 -15132
rect 2667 -15388 2673 -15132
rect 2627 -15400 2673 -15388
rect 2805 -15132 2851 -15120
rect 2805 -15388 2811 -15132
rect 2845 -15388 2851 -15132
rect 2805 -15400 2851 -15388
rect 2983 -15132 3029 -15120
rect 2983 -15388 2989 -15132
rect 3023 -15388 3029 -15132
rect 2983 -15400 3029 -15388
rect 3161 -15132 3207 -15120
rect 3161 -15388 3167 -15132
rect 3201 -15388 3207 -15132
rect 3161 -15400 3207 -15388
rect 3339 -15132 3385 -15120
rect 3339 -15388 3345 -15132
rect 3379 -15388 3385 -15132
rect 3339 -15400 3385 -15388
rect 3517 -15132 3563 -15120
rect 3517 -15388 3523 -15132
rect 3557 -15388 3563 -15132
rect 3517 -15400 3563 -15388
rect 3695 -15132 3741 -15120
rect 3695 -15388 3701 -15132
rect 3735 -15388 3741 -15132
rect 3695 -15400 3741 -15388
rect 3873 -15132 3919 -15120
rect 3873 -15388 3879 -15132
rect 3913 -15388 3919 -15132
rect 3873 -15400 3919 -15388
rect 4051 -15132 4097 -15120
rect 4051 -15388 4057 -15132
rect 4091 -15388 4097 -15132
rect 4051 -15400 4097 -15388
rect -2105 -15438 -2029 -15432
rect -2105 -15472 -2089 -15438
rect -2045 -15472 -2029 -15438
rect -2105 -15488 -2029 -15472
rect -2457 -15874 -2447 -15821
rect -2394 -15874 -2384 -15821
rect -1995 -15822 -1961 -15400
rect -1927 -15438 -1851 -15432
rect -1927 -15472 -1911 -15438
rect -1867 -15472 -1851 -15438
rect -1927 -15488 -1851 -15472
rect -2015 -15875 -2005 -15822
rect -1952 -15875 -1942 -15822
rect -2105 -16048 -2029 -16032
rect -2105 -16050 -2089 -16048
rect -2173 -16082 -2089 -16050
rect -2045 -16050 -2029 -16048
rect -1995 -16050 -1961 -15875
rect -1906 -15933 -1872 -15488
rect -1925 -15986 -1915 -15933
rect -1862 -15986 -1852 -15933
rect -2045 -16082 -1961 -16050
rect -2173 -16084 -1961 -16082
rect -2173 -16120 -2139 -16084
rect -2105 -16088 -2029 -16084
rect -1995 -16120 -1961 -16084
rect -1927 -16048 -1851 -16032
rect -1927 -16082 -1911 -16048
rect -1867 -16082 -1851 -16048
rect -1927 -16088 -1851 -16082
rect -1817 -16120 -1783 -15400
rect -1749 -15438 -1673 -15432
rect -1749 -15472 -1733 -15438
rect -1689 -15472 -1673 -15438
rect -1749 -15488 -1673 -15472
rect -1728 -15933 -1694 -15488
rect -1639 -15822 -1605 -15400
rect -1571 -15438 -1495 -15432
rect -1571 -15472 -1555 -15438
rect -1511 -15472 -1495 -15438
rect -1571 -15488 -1495 -15472
rect -1659 -15875 -1649 -15822
rect -1596 -15875 -1586 -15822
rect -1748 -15986 -1738 -15933
rect -1685 -15986 -1675 -15933
rect -1749 -16048 -1673 -16032
rect -1749 -16082 -1733 -16048
rect -1689 -16082 -1673 -16048
rect -1749 -16088 -1673 -16082
rect -1639 -16120 -1605 -15875
rect -1550 -15933 -1516 -15488
rect -1570 -15986 -1560 -15933
rect -1507 -15986 -1497 -15933
rect -1571 -16048 -1495 -16032
rect -1571 -16082 -1555 -16048
rect -1511 -16082 -1495 -16048
rect -1571 -16088 -1495 -16082
rect -1461 -16120 -1427 -15400
rect -1393 -15438 -1317 -15432
rect -1393 -15472 -1377 -15438
rect -1333 -15472 -1317 -15438
rect -1393 -15488 -1317 -15472
rect -1372 -15933 -1338 -15488
rect -1283 -15822 -1249 -15400
rect -1215 -15438 -1139 -15432
rect -1215 -15472 -1199 -15438
rect -1155 -15472 -1139 -15438
rect -1215 -15488 -1139 -15472
rect -1303 -15875 -1293 -15822
rect -1240 -15875 -1230 -15822
rect -1392 -15986 -1382 -15933
rect -1329 -15986 -1319 -15933
rect -1393 -16048 -1317 -16032
rect -1393 -16082 -1377 -16048
rect -1333 -16082 -1317 -16048
rect -1393 -16088 -1317 -16082
rect -1283 -16120 -1249 -15875
rect -1194 -15933 -1160 -15488
rect -1214 -15986 -1204 -15933
rect -1151 -15986 -1141 -15933
rect -1215 -16048 -1139 -16032
rect -1215 -16082 -1199 -16048
rect -1155 -16082 -1139 -16048
rect -1215 -16088 -1139 -16082
rect -1104 -16120 -1070 -15400
rect -1037 -15438 -961 -15432
rect -1037 -15472 -1021 -15438
rect -977 -15472 -961 -15438
rect -1037 -15488 -961 -15472
rect -1015 -15933 -981 -15488
rect -927 -15822 -893 -15400
rect -859 -15438 -783 -15432
rect -859 -15472 -843 -15438
rect -799 -15472 -783 -15438
rect -859 -15488 -783 -15472
rect -947 -15875 -937 -15822
rect -884 -15875 -874 -15822
rect -1035 -15986 -1025 -15933
rect -972 -15986 -962 -15933
rect -1037 -16048 -961 -16032
rect -1037 -16082 -1021 -16048
rect -977 -16082 -961 -16048
rect -1037 -16088 -961 -16082
rect -927 -16120 -893 -15875
rect -857 -15986 -847 -15933
rect -794 -15986 -784 -15933
rect -838 -16032 -804 -15986
rect -859 -16048 -783 -16032
rect -859 -16082 -843 -16048
rect -799 -16082 -783 -16048
rect -859 -16088 -783 -16082
rect -749 -16120 -715 -15400
rect -681 -15438 -605 -15432
rect -681 -15472 -665 -15438
rect -621 -15472 -605 -15438
rect -681 -15488 -605 -15472
rect -571 -15822 -537 -15400
rect -503 -15438 -427 -15432
rect -503 -15472 -487 -15438
rect -443 -15472 -427 -15438
rect -503 -15488 -427 -15472
rect -591 -15875 -581 -15822
rect -528 -15875 -518 -15822
rect -680 -15986 -670 -15933
rect -617 -15986 -607 -15933
rect -660 -16032 -626 -15986
rect -681 -16048 -605 -16032
rect -681 -16082 -665 -16048
rect -621 -16082 -605 -16048
rect -681 -16088 -605 -16082
rect -571 -16120 -537 -15875
rect -501 -15986 -491 -15933
rect -438 -15986 -428 -15933
rect -482 -16032 -448 -15986
rect -503 -16048 -427 -16032
rect -503 -16082 -487 -16048
rect -443 -16082 -427 -16048
rect -503 -16088 -427 -16082
rect -393 -16120 -359 -15400
rect -325 -15438 -249 -15432
rect -325 -15472 -309 -15438
rect -265 -15472 -249 -15438
rect -325 -15488 -249 -15472
rect -215 -15822 -181 -15400
rect -147 -15438 -71 -15432
rect -147 -15472 -131 -15438
rect -87 -15472 -71 -15438
rect -147 -15488 -71 -15472
rect -235 -15875 -225 -15822
rect -172 -15875 -162 -15822
rect -323 -15986 -313 -15933
rect -260 -15986 -250 -15933
rect -304 -16032 -270 -15986
rect -325 -16048 -249 -16032
rect -325 -16082 -309 -16048
rect -265 -16082 -249 -16048
rect -325 -16088 -249 -16082
rect -215 -16120 -181 -15875
rect -146 -15986 -136 -15933
rect -83 -15986 -73 -15933
rect -126 -16032 -92 -15986
rect -147 -16048 -71 -16032
rect -147 -16082 -131 -16048
rect -87 -16082 -71 -16048
rect -147 -16088 -71 -16082
rect -37 -16120 -3 -15400
rect 31 -15438 107 -15432
rect 31 -15472 47 -15438
rect 91 -15472 107 -15438
rect 31 -15488 107 -15472
rect 141 -15821 175 -15400
rect 209 -15438 285 -15432
rect 209 -15472 225 -15438
rect 269 -15472 285 -15438
rect 209 -15488 285 -15472
rect 122 -15874 132 -15821
rect 185 -15874 195 -15821
rect 33 -15986 43 -15933
rect 96 -15986 106 -15933
rect 52 -16032 86 -15986
rect 31 -16048 107 -16032
rect 31 -16082 47 -16048
rect 91 -16082 107 -16048
rect 31 -16088 107 -16082
rect 141 -16120 175 -15874
rect 230 -15933 264 -15488
rect 211 -15986 221 -15933
rect 274 -15986 284 -15933
rect 209 -16048 285 -16032
rect 209 -16082 225 -16048
rect 269 -16082 285 -16048
rect 209 -16088 285 -16082
rect 319 -16120 353 -15400
rect 387 -15438 463 -15432
rect 387 -15472 403 -15438
rect 447 -15472 463 -15438
rect 387 -15488 463 -15472
rect 408 -15933 442 -15488
rect 497 -15822 531 -15400
rect 565 -15438 641 -15432
rect 565 -15472 581 -15438
rect 625 -15472 641 -15438
rect 565 -15488 641 -15472
rect 477 -15875 487 -15822
rect 540 -15875 550 -15822
rect 388 -15986 398 -15933
rect 451 -15986 461 -15933
rect 387 -16048 463 -16032
rect 387 -16082 403 -16048
rect 447 -16082 463 -16048
rect 387 -16088 463 -16082
rect 497 -16120 531 -15875
rect 585 -15933 619 -15488
rect 565 -15986 575 -15933
rect 628 -15986 638 -15933
rect 565 -16048 641 -16032
rect 565 -16082 581 -16048
rect 625 -16082 641 -16048
rect 565 -16088 641 -16082
rect 675 -16120 709 -15400
rect 743 -15438 819 -15432
rect 743 -15472 759 -15438
rect 803 -15472 819 -15438
rect 743 -15488 819 -15472
rect 764 -15933 798 -15488
rect 853 -15822 887 -15400
rect 921 -15438 997 -15432
rect 921 -15472 937 -15438
rect 981 -15472 997 -15438
rect 921 -15488 997 -15472
rect 833 -15875 843 -15822
rect 896 -15875 906 -15822
rect 745 -15986 755 -15933
rect 808 -15986 818 -15933
rect 743 -16048 819 -16032
rect 743 -16082 759 -16048
rect 803 -16082 819 -16048
rect 743 -16088 819 -16082
rect 853 -16120 887 -15875
rect 941 -15933 975 -15488
rect 921 -15986 931 -15933
rect 984 -15986 994 -15933
rect 921 -16048 997 -16032
rect 921 -16082 937 -16048
rect 981 -16082 997 -16048
rect 921 -16088 997 -16082
rect 1031 -16120 1065 -15400
rect 1099 -15438 1175 -15432
rect 1099 -15472 1115 -15438
rect 1159 -15472 1175 -15438
rect 1099 -15488 1175 -15472
rect 1120 -15933 1154 -15488
rect 1209 -15822 1243 -15400
rect 1277 -15438 1353 -15432
rect 1277 -15472 1293 -15438
rect 1337 -15472 1353 -15438
rect 1277 -15488 1353 -15472
rect 1191 -15875 1201 -15822
rect 1254 -15875 1264 -15822
rect 1100 -15986 1110 -15933
rect 1163 -15986 1173 -15933
rect 1099 -16048 1175 -16032
rect 1099 -16082 1115 -16048
rect 1159 -16082 1175 -16048
rect 1099 -16088 1175 -16082
rect 1209 -16120 1243 -15875
rect 1279 -15986 1289 -15933
rect 1342 -15986 1352 -15933
rect 1298 -16032 1332 -15986
rect 1277 -16048 1353 -16032
rect 1277 -16082 1293 -16048
rect 1337 -16082 1353 -16048
rect 1277 -16088 1353 -16082
rect 1387 -16120 1421 -15400
rect 1455 -15438 1531 -15432
rect 1455 -15472 1471 -15438
rect 1515 -15472 1531 -15438
rect 1455 -15488 1531 -15472
rect 1565 -15822 1599 -15400
rect 1633 -15438 1709 -15432
rect 1633 -15472 1649 -15438
rect 1693 -15472 1709 -15438
rect 1633 -15488 1709 -15472
rect 1545 -15875 1555 -15822
rect 1608 -15875 1618 -15822
rect 1456 -15986 1466 -15933
rect 1519 -15986 1529 -15933
rect 1476 -16032 1510 -15986
rect 1455 -16048 1531 -16032
rect 1455 -16082 1471 -16048
rect 1515 -16082 1531 -16048
rect 1455 -16088 1531 -16082
rect 1565 -16120 1599 -15875
rect 1633 -15986 1643 -15933
rect 1696 -15986 1706 -15933
rect 1653 -16032 1687 -15986
rect 1633 -16048 1709 -16032
rect 1633 -16082 1649 -16048
rect 1693 -16082 1709 -16048
rect 1633 -16088 1709 -16082
rect 1744 -16120 1778 -15400
rect 1811 -15438 1887 -15432
rect 1811 -15472 1827 -15438
rect 1871 -15472 1887 -15438
rect 1811 -15488 1887 -15472
rect 1921 -15822 1955 -15400
rect 1989 -15438 2065 -15432
rect 1989 -15472 2005 -15438
rect 2049 -15472 2065 -15438
rect 1989 -15488 2065 -15472
rect 1900 -15875 1910 -15822
rect 1963 -15875 1973 -15822
rect 1812 -15986 1822 -15933
rect 1875 -15986 1885 -15933
rect 1832 -16032 1866 -15986
rect 1811 -16048 1887 -16032
rect 1811 -16082 1827 -16048
rect 1871 -16082 1887 -16048
rect 1811 -16088 1887 -16082
rect 1921 -16120 1955 -15875
rect 1990 -15986 2000 -15933
rect 2053 -15986 2063 -15933
rect 2010 -16032 2044 -15986
rect 1989 -16048 2065 -16032
rect 1989 -16082 2005 -16048
rect 2049 -16082 2065 -16048
rect 1989 -16088 2065 -16082
rect 2100 -16120 2134 -15400
rect 2167 -15438 2243 -15432
rect 2167 -15472 2183 -15438
rect 2227 -15472 2243 -15438
rect 2167 -15488 2243 -15472
rect 2277 -15822 2311 -15400
rect 2345 -15438 2421 -15432
rect 2345 -15472 2361 -15438
rect 2405 -15472 2421 -15438
rect 2345 -15488 2421 -15472
rect 2257 -15875 2267 -15822
rect 2320 -15875 2330 -15822
rect 2169 -15986 2179 -15933
rect 2232 -15986 2242 -15933
rect 2189 -16032 2223 -15986
rect 2167 -16048 2243 -16032
rect 2167 -16082 2183 -16048
rect 2227 -16082 2243 -16048
rect 2167 -16088 2243 -16082
rect 2277 -16120 2311 -15875
rect 2366 -15933 2400 -15488
rect 2346 -15986 2356 -15933
rect 2409 -15986 2419 -15933
rect 2345 -16048 2421 -16032
rect 2345 -16082 2361 -16048
rect 2405 -16082 2421 -16048
rect 2345 -16088 2421 -16082
rect 2455 -16120 2489 -15400
rect 2523 -15438 2599 -15432
rect 2523 -15472 2539 -15438
rect 2583 -15472 2599 -15438
rect 2523 -15488 2599 -15472
rect 2544 -15933 2578 -15488
rect 2633 -15822 2667 -15400
rect 2701 -15438 2777 -15432
rect 2701 -15472 2717 -15438
rect 2761 -15472 2777 -15438
rect 2701 -15488 2777 -15472
rect 2614 -15875 2624 -15822
rect 2677 -15875 2687 -15822
rect 2524 -15986 2534 -15933
rect 2587 -15986 2597 -15933
rect 2523 -16048 2599 -16032
rect 2523 -16082 2539 -16048
rect 2583 -16082 2599 -16048
rect 2523 -16088 2599 -16082
rect 2633 -16120 2667 -15875
rect 2722 -15933 2756 -15488
rect 2702 -15986 2712 -15933
rect 2765 -15986 2775 -15933
rect 2701 -16048 2777 -16032
rect 2701 -16082 2717 -16048
rect 2761 -16082 2777 -16048
rect 2701 -16088 2777 -16082
rect 2811 -16120 2845 -15400
rect 2879 -15438 2955 -15432
rect 2879 -15472 2895 -15438
rect 2939 -15472 2955 -15438
rect 2879 -15488 2955 -15472
rect 2900 -15933 2934 -15488
rect 2989 -15822 3023 -15400
rect 3057 -15438 3133 -15432
rect 3057 -15472 3073 -15438
rect 3117 -15472 3133 -15438
rect 3057 -15488 3133 -15472
rect 2969 -15875 2979 -15822
rect 3032 -15875 3042 -15822
rect 2881 -15986 2891 -15933
rect 2944 -15986 2954 -15933
rect 2879 -16048 2955 -16032
rect 2879 -16082 2895 -16048
rect 2939 -16082 2955 -16048
rect 2879 -16088 2955 -16082
rect 2989 -16120 3023 -15875
rect 3078 -15933 3112 -15488
rect 3058 -15986 3068 -15933
rect 3121 -15986 3131 -15933
rect 3057 -16048 3133 -16032
rect 3057 -16082 3073 -16048
rect 3117 -16082 3133 -16048
rect 3057 -16088 3133 -16082
rect 3167 -16120 3201 -15400
rect 3235 -15438 3311 -15432
rect 3235 -15472 3251 -15438
rect 3295 -15472 3311 -15438
rect 3235 -15488 3311 -15472
rect 3256 -15933 3290 -15488
rect 3345 -15822 3379 -15400
rect 3413 -15438 3489 -15432
rect 3413 -15472 3429 -15438
rect 3473 -15472 3489 -15438
rect 3413 -15488 3489 -15472
rect 3325 -15875 3335 -15822
rect 3388 -15875 3398 -15822
rect 3237 -15986 3247 -15933
rect 3300 -15986 3310 -15933
rect 3235 -16048 3311 -16032
rect 3235 -16082 3251 -16048
rect 3295 -16082 3311 -16048
rect 3235 -16088 3311 -16082
rect 3345 -16120 3379 -15875
rect 3414 -15986 3424 -15933
rect 3477 -15986 3487 -15933
rect 3434 -16032 3468 -15986
rect 3413 -16048 3489 -16032
rect 3413 -16082 3429 -16048
rect 3473 -16082 3489 -16048
rect 3413 -16088 3489 -16082
rect 3524 -16120 3558 -15400
rect 3591 -15438 3667 -15432
rect 3591 -15472 3607 -15438
rect 3651 -15472 3667 -15438
rect 3591 -15488 3667 -15472
rect 3701 -15822 3735 -15400
rect 3769 -15438 3845 -15432
rect 3769 -15472 3785 -15438
rect 3829 -15472 3845 -15438
rect 3769 -15488 3845 -15472
rect 3682 -15875 3692 -15822
rect 3745 -15875 3755 -15822
rect 3593 -15986 3603 -15933
rect 3656 -15986 3666 -15933
rect 3612 -16032 3646 -15986
rect 3591 -16048 3667 -16032
rect 3591 -16082 3607 -16048
rect 3651 -16082 3667 -16048
rect 3591 -16088 3667 -16082
rect 3701 -16120 3735 -15875
rect 3770 -15986 3780 -15933
rect 3833 -15986 3843 -15933
rect 3790 -16032 3824 -15986
rect 3769 -16048 3845 -16032
rect 3769 -16082 3785 -16048
rect 3829 -16082 3845 -16048
rect 3769 -16088 3845 -16082
rect 3879 -16047 3913 -15400
rect 3947 -15438 4023 -15432
rect 3947 -15472 3963 -15438
rect 4007 -15472 4023 -15438
rect 3947 -15488 4023 -15472
rect 4238 -15539 4291 -14979
rect 4228 -15592 4238 -15539
rect 4291 -15592 4301 -15539
rect 5031 -15540 5084 -13486
rect 5390 -13598 5400 -13545
rect 5453 -13598 5463 -13545
rect 5132 -13847 5142 -13794
rect 5195 -13847 5205 -13794
rect 5142 -14658 5195 -13847
rect 5133 -14711 5143 -14658
rect 5196 -14711 5206 -14658
rect 3947 -16047 4023 -16032
rect 3879 -16048 4090 -16047
rect 3879 -16081 3963 -16048
rect 3879 -16120 3913 -16081
rect 3947 -16082 3963 -16081
rect 4007 -16081 4090 -16048
rect 4007 -16082 4023 -16081
rect 3947 -16088 4023 -16082
rect 4056 -16120 4090 -16081
rect -2179 -16132 -2133 -16120
rect -3945 -16347 -3935 -16295
rect -3883 -16347 -3873 -16295
rect -4180 -16410 -4104 -16394
rect -4180 -16444 -4164 -16410
rect -4120 -16444 -4104 -16410
rect -4180 -16450 -4104 -16444
rect -6034 -16494 -5988 -16482
rect -6034 -16750 -6028 -16494
rect -5994 -16750 -5988 -16494
rect -6034 -16762 -5988 -16750
rect -5856 -16494 -5810 -16482
rect -5856 -16750 -5850 -16494
rect -5816 -16750 -5810 -16494
rect -5856 -16762 -5810 -16750
rect -5678 -16494 -5632 -16482
rect -5678 -16750 -5672 -16494
rect -5638 -16750 -5632 -16494
rect -5678 -16762 -5632 -16750
rect -5500 -16494 -5454 -16482
rect -5500 -16750 -5494 -16494
rect -5460 -16750 -5454 -16494
rect -5500 -16762 -5454 -16750
rect -5322 -16494 -5276 -16482
rect -5322 -16750 -5316 -16494
rect -5282 -16750 -5276 -16494
rect -5322 -16762 -5276 -16750
rect -5144 -16494 -5098 -16482
rect -5144 -16750 -5138 -16494
rect -5104 -16750 -5098 -16494
rect -5144 -16762 -5098 -16750
rect -4966 -16494 -4920 -16482
rect -4966 -16750 -4960 -16494
rect -4926 -16750 -4920 -16494
rect -4966 -16762 -4920 -16750
rect -4788 -16494 -4742 -16482
rect -4788 -16750 -4782 -16494
rect -4748 -16750 -4742 -16494
rect -4788 -16762 -4742 -16750
rect -4610 -16494 -4564 -16482
rect -4610 -16750 -4604 -16494
rect -4570 -16750 -4564 -16494
rect -4610 -16762 -4564 -16750
rect -4432 -16494 -4386 -16482
rect -4432 -16750 -4426 -16494
rect -4392 -16750 -4386 -16494
rect -4432 -16762 -4386 -16750
rect -4254 -16494 -4208 -16482
rect -4254 -16750 -4248 -16494
rect -4214 -16750 -4208 -16494
rect -4254 -16762 -4208 -16750
rect -4076 -16494 -4030 -16482
rect -4076 -16750 -4070 -16494
rect -4036 -16750 -4030 -16494
rect -4076 -16762 -4030 -16750
rect -6028 -16886 -5994 -16762
rect -5960 -16800 -5884 -16794
rect -5960 -16834 -5944 -16800
rect -5900 -16834 -5884 -16800
rect -5960 -16850 -5884 -16834
rect -5939 -16886 -5905 -16850
rect -5850 -16886 -5816 -16762
rect -5782 -16800 -5706 -16794
rect -5782 -16834 -5766 -16800
rect -5722 -16834 -5706 -16800
rect -5782 -16850 -5706 -16834
rect -5672 -16886 -5638 -16762
rect -5604 -16800 -5528 -16794
rect -5604 -16834 -5588 -16800
rect -5544 -16834 -5528 -16800
rect -5604 -16850 -5528 -16834
rect -6028 -16920 -5816 -16886
rect -5850 -17007 -5816 -16920
rect -5692 -16939 -5682 -16886
rect -5629 -16939 -5619 -16886
rect -6169 -17060 -6159 -17007
rect -6106 -17060 -6096 -17007
rect -5869 -17060 -5859 -17007
rect -5806 -17060 -5796 -17007
rect -5494 -17118 -5460 -16762
rect -5426 -16800 -5350 -16794
rect -5426 -16834 -5410 -16800
rect -5366 -16834 -5350 -16800
rect -5426 -16850 -5350 -16834
rect -5316 -16886 -5282 -16762
rect -5248 -16800 -5172 -16794
rect -5248 -16834 -5232 -16800
rect -5188 -16834 -5172 -16800
rect -5248 -16850 -5172 -16834
rect -5336 -16939 -5326 -16886
rect -5273 -16939 -5263 -16886
rect -5138 -17007 -5104 -16762
rect -5070 -16800 -4994 -16794
rect -5070 -16834 -5054 -16800
rect -5010 -16834 -4994 -16800
rect -5070 -16850 -4994 -16834
rect -4960 -16886 -4926 -16762
rect -4892 -16800 -4816 -16794
rect -4892 -16834 -4876 -16800
rect -4832 -16834 -4816 -16800
rect -4892 -16850 -4816 -16834
rect -4980 -16939 -4970 -16886
rect -4917 -16939 -4907 -16886
rect -5158 -17060 -5148 -17007
rect -5095 -17060 -5085 -17007
rect -5514 -17171 -5504 -17118
rect -5451 -17171 -5441 -17118
rect -7605 -17251 -7329 -17250
rect -4970 -17251 -4917 -16939
rect -4782 -17118 -4748 -16762
rect -4714 -16800 -4638 -16794
rect -4714 -16834 -4698 -16800
rect -4654 -16834 -4638 -16800
rect -4714 -16850 -4638 -16834
rect -4604 -16886 -4570 -16762
rect -4536 -16800 -4460 -16794
rect -4536 -16834 -4520 -16800
rect -4476 -16834 -4460 -16800
rect -4536 -16850 -4460 -16834
rect -4624 -16939 -4614 -16886
rect -4561 -16939 -4551 -16886
rect -4426 -17007 -4392 -16762
rect -4358 -16800 -4282 -16794
rect -4358 -16834 -4342 -16800
rect -4298 -16834 -4282 -16800
rect -4358 -16850 -4282 -16834
rect -4248 -16886 -4214 -16762
rect -4180 -16800 -4104 -16794
rect -4180 -16834 -4164 -16800
rect -4120 -16834 -4104 -16800
rect -4180 -16850 -4104 -16834
rect -4159 -16886 -4125 -16850
rect -4070 -16886 -4036 -16762
rect -4268 -16939 -4258 -16886
rect -4205 -16939 -4036 -16886
rect -4447 -17060 -4437 -17007
rect -4384 -17060 -4374 -17007
rect -3935 -17118 -3883 -16347
rect -2179 -16388 -2173 -16132
rect -2139 -16388 -2133 -16132
rect -2179 -16400 -2133 -16388
rect -2001 -16132 -1955 -16120
rect -2001 -16388 -1995 -16132
rect -1961 -16388 -1955 -16132
rect -2001 -16400 -1955 -16388
rect -1823 -16132 -1777 -16120
rect -1823 -16388 -1817 -16132
rect -1783 -16388 -1777 -16132
rect -1823 -16400 -1777 -16388
rect -1645 -16132 -1599 -16120
rect -1645 -16388 -1639 -16132
rect -1605 -16388 -1599 -16132
rect -1645 -16400 -1599 -16388
rect -1467 -16132 -1421 -16120
rect -1467 -16388 -1461 -16132
rect -1427 -16388 -1421 -16132
rect -1467 -16400 -1421 -16388
rect -1289 -16132 -1243 -16120
rect -1289 -16388 -1283 -16132
rect -1249 -16388 -1243 -16132
rect -1289 -16400 -1243 -16388
rect -1111 -16132 -1065 -16120
rect -1111 -16388 -1105 -16132
rect -1071 -16388 -1065 -16132
rect -1111 -16400 -1065 -16388
rect -933 -16132 -887 -16120
rect -933 -16388 -927 -16132
rect -893 -16388 -887 -16132
rect -933 -16400 -887 -16388
rect -755 -16132 -709 -16120
rect -755 -16388 -749 -16132
rect -715 -16388 -709 -16132
rect -755 -16400 -709 -16388
rect -577 -16132 -531 -16120
rect -577 -16388 -571 -16132
rect -537 -16388 -531 -16132
rect -577 -16400 -531 -16388
rect -399 -16132 -353 -16120
rect -399 -16388 -393 -16132
rect -359 -16388 -353 -16132
rect -399 -16400 -353 -16388
rect -221 -16132 -175 -16120
rect -221 -16388 -215 -16132
rect -181 -16388 -175 -16132
rect -221 -16400 -175 -16388
rect -43 -16132 3 -16120
rect -43 -16388 -37 -16132
rect -3 -16388 3 -16132
rect -43 -16400 3 -16388
rect 135 -16132 181 -16120
rect 135 -16388 141 -16132
rect 175 -16388 181 -16132
rect 135 -16400 181 -16388
rect 313 -16132 359 -16120
rect 313 -16388 319 -16132
rect 353 -16388 359 -16132
rect 313 -16400 359 -16388
rect 491 -16132 537 -16120
rect 491 -16388 497 -16132
rect 531 -16388 537 -16132
rect 491 -16400 537 -16388
rect 669 -16132 715 -16120
rect 669 -16388 675 -16132
rect 709 -16388 715 -16132
rect 669 -16400 715 -16388
rect 847 -16132 893 -16120
rect 847 -16388 853 -16132
rect 887 -16388 893 -16132
rect 847 -16400 893 -16388
rect 1025 -16132 1071 -16120
rect 1025 -16388 1031 -16132
rect 1065 -16388 1071 -16132
rect 1025 -16400 1071 -16388
rect 1203 -16132 1249 -16120
rect 1203 -16388 1209 -16132
rect 1243 -16388 1249 -16132
rect 1203 -16400 1249 -16388
rect 1381 -16132 1427 -16120
rect 1381 -16388 1387 -16132
rect 1421 -16388 1427 -16132
rect 1381 -16400 1427 -16388
rect 1559 -16132 1605 -16120
rect 1559 -16388 1565 -16132
rect 1599 -16388 1605 -16132
rect 1559 -16400 1605 -16388
rect 1737 -16132 1783 -16120
rect 1737 -16388 1743 -16132
rect 1777 -16388 1783 -16132
rect 1737 -16400 1783 -16388
rect 1915 -16132 1961 -16120
rect 1915 -16388 1921 -16132
rect 1955 -16388 1961 -16132
rect 1915 -16400 1961 -16388
rect 2093 -16132 2139 -16120
rect 2093 -16388 2099 -16132
rect 2133 -16388 2139 -16132
rect 2093 -16400 2139 -16388
rect 2271 -16132 2317 -16120
rect 2271 -16388 2277 -16132
rect 2311 -16388 2317 -16132
rect 2271 -16400 2317 -16388
rect 2449 -16132 2495 -16120
rect 2449 -16388 2455 -16132
rect 2489 -16388 2495 -16132
rect 2449 -16400 2495 -16388
rect 2627 -16132 2673 -16120
rect 2627 -16388 2633 -16132
rect 2667 -16388 2673 -16132
rect 2627 -16400 2673 -16388
rect 2805 -16132 2851 -16120
rect 2805 -16388 2811 -16132
rect 2845 -16388 2851 -16132
rect 2805 -16400 2851 -16388
rect 2983 -16132 3029 -16120
rect 2983 -16388 2989 -16132
rect 3023 -16388 3029 -16132
rect 2983 -16400 3029 -16388
rect 3161 -16132 3207 -16120
rect 3161 -16388 3167 -16132
rect 3201 -16388 3207 -16132
rect 3161 -16400 3207 -16388
rect 3339 -16132 3385 -16120
rect 3339 -16388 3345 -16132
rect 3379 -16388 3385 -16132
rect 3339 -16400 3385 -16388
rect 3517 -16132 3563 -16120
rect 3517 -16388 3523 -16132
rect 3557 -16388 3563 -16132
rect 3517 -16400 3563 -16388
rect 3695 -16132 3741 -16120
rect 3695 -16388 3701 -16132
rect 3735 -16388 3741 -16132
rect 3695 -16400 3741 -16388
rect 3873 -16132 3919 -16120
rect 3873 -16388 3879 -16132
rect 3913 -16388 3919 -16132
rect 3873 -16400 3919 -16388
rect 4051 -16132 4097 -16120
rect 4051 -16388 4057 -16132
rect 4091 -16388 4097 -16132
rect 4051 -16400 4097 -16388
rect -2105 -16438 -2029 -16432
rect -2105 -16472 -2089 -16438
rect -2045 -16472 -2029 -16438
rect -2105 -16488 -2029 -16472
rect -1927 -16438 -1851 -16432
rect -1927 -16472 -1911 -16438
rect -1867 -16472 -1851 -16438
rect -1927 -16488 -1851 -16472
rect -1906 -16542 -1872 -16488
rect -1927 -16595 -1917 -16542
rect -1864 -16595 -1854 -16542
rect -1817 -16665 -1783 -16400
rect -1749 -16438 -1673 -16432
rect -1749 -16472 -1733 -16438
rect -1689 -16472 -1673 -16438
rect -1749 -16488 -1673 -16472
rect -1571 -16438 -1495 -16432
rect -1571 -16472 -1555 -16438
rect -1511 -16472 -1495 -16438
rect -1571 -16488 -1495 -16472
rect -1728 -16542 -1694 -16488
rect -1550 -16541 -1516 -16488
rect -1748 -16595 -1738 -16542
rect -1685 -16595 -1675 -16542
rect -1571 -16594 -1561 -16541
rect -1508 -16594 -1498 -16541
rect -1837 -16718 -1827 -16665
rect -1774 -16718 -1764 -16665
rect -1461 -16666 -1427 -16400
rect -1393 -16438 -1317 -16432
rect -1393 -16472 -1377 -16438
rect -1333 -16472 -1317 -16438
rect -1393 -16488 -1317 -16472
rect -1215 -16438 -1139 -16432
rect -1215 -16472 -1199 -16438
rect -1155 -16472 -1139 -16438
rect -1215 -16488 -1139 -16472
rect -1372 -16543 -1338 -16488
rect -1194 -16542 -1160 -16488
rect -1391 -16596 -1381 -16543
rect -1328 -16596 -1318 -16543
rect -1214 -16595 -1204 -16542
rect -1151 -16595 -1141 -16542
rect -1104 -16665 -1070 -16400
rect -1037 -16438 -961 -16432
rect -1037 -16472 -1021 -16438
rect -977 -16472 -961 -16438
rect -1037 -16488 -961 -16472
rect -859 -16438 -783 -16432
rect -859 -16472 -843 -16438
rect -799 -16472 -783 -16438
rect -859 -16488 -783 -16472
rect -1016 -16542 -982 -16488
rect -1036 -16595 -1026 -16542
rect -973 -16595 -963 -16542
rect -749 -16664 -715 -16400
rect -681 -16438 -605 -16432
rect -681 -16472 -665 -16438
rect -621 -16472 -605 -16438
rect -681 -16488 -605 -16472
rect -503 -16438 -427 -16432
rect -503 -16472 -487 -16438
rect -443 -16472 -427 -16438
rect -503 -16488 -427 -16472
rect -1481 -16719 -1471 -16666
rect -1418 -16719 -1408 -16666
rect -1124 -16718 -1114 -16665
rect -1061 -16718 -1051 -16665
rect -769 -16717 -759 -16664
rect -706 -16717 -696 -16664
rect -393 -16665 -359 -16400
rect -325 -16438 -249 -16432
rect -325 -16472 -309 -16438
rect -265 -16472 -249 -16438
rect -325 -16488 -249 -16472
rect -147 -16438 -71 -16432
rect -147 -16472 -131 -16438
rect -87 -16472 -71 -16438
rect -147 -16488 -71 -16472
rect -37 -16665 -3 -16400
rect 31 -16438 107 -16432
rect 31 -16472 47 -16438
rect 91 -16472 107 -16438
rect 31 -16488 107 -16472
rect 209 -16438 285 -16432
rect 209 -16472 225 -16438
rect 269 -16472 285 -16438
rect 209 -16488 285 -16472
rect 230 -16542 264 -16488
rect 210 -16595 220 -16542
rect 273 -16595 283 -16542
rect -413 -16718 -403 -16665
rect -350 -16718 -340 -16665
rect -57 -16718 -47 -16665
rect 6 -16718 16 -16665
rect 319 -16666 353 -16400
rect 387 -16438 463 -16432
rect 387 -16472 403 -16438
rect 447 -16472 463 -16438
rect 387 -16488 463 -16472
rect 565 -16438 641 -16432
rect 565 -16472 581 -16438
rect 625 -16472 641 -16438
rect 565 -16488 641 -16472
rect 408 -16542 442 -16488
rect 586 -16542 620 -16488
rect 387 -16595 397 -16542
rect 450 -16595 460 -16542
rect 566 -16595 576 -16542
rect 629 -16595 639 -16542
rect 675 -16665 709 -16400
rect 743 -16438 819 -16432
rect 743 -16472 759 -16438
rect 803 -16472 819 -16438
rect 743 -16488 819 -16472
rect 921 -16438 997 -16432
rect 921 -16472 937 -16438
rect 981 -16472 997 -16438
rect 921 -16488 997 -16472
rect 765 -16542 799 -16488
rect 943 -16542 977 -16488
rect 745 -16595 755 -16542
rect 808 -16595 818 -16542
rect 923 -16595 933 -16542
rect 986 -16595 996 -16542
rect 1031 -16665 1065 -16400
rect 1099 -16438 1175 -16432
rect 1099 -16472 1115 -16438
rect 1159 -16472 1175 -16438
rect 1099 -16488 1175 -16472
rect 1277 -16438 1353 -16432
rect 1277 -16472 1293 -16438
rect 1337 -16472 1353 -16438
rect 1277 -16488 1353 -16472
rect 1120 -16542 1154 -16488
rect 1101 -16595 1111 -16542
rect 1164 -16595 1174 -16542
rect 1387 -16665 1421 -16400
rect 1455 -16438 1531 -16432
rect 1455 -16472 1471 -16438
rect 1515 -16472 1531 -16438
rect 1455 -16488 1531 -16472
rect 1633 -16438 1709 -16432
rect 1633 -16472 1649 -16438
rect 1693 -16472 1709 -16438
rect 1633 -16488 1709 -16472
rect 1744 -16665 1778 -16400
rect 1811 -16438 1887 -16432
rect 1811 -16472 1827 -16438
rect 1871 -16472 1887 -16438
rect 1811 -16488 1887 -16472
rect 1989 -16438 2065 -16432
rect 1989 -16472 2005 -16438
rect 2049 -16472 2065 -16438
rect 1989 -16488 2065 -16472
rect 2100 -16664 2134 -16400
rect 2167 -16438 2243 -16432
rect 2167 -16472 2183 -16438
rect 2227 -16472 2243 -16438
rect 2167 -16488 2243 -16472
rect 2345 -16438 2421 -16432
rect 2345 -16472 2361 -16438
rect 2405 -16472 2421 -16438
rect 2345 -16488 2421 -16472
rect 2366 -16542 2400 -16488
rect 2346 -16595 2356 -16542
rect 2409 -16595 2419 -16542
rect 299 -16719 309 -16666
rect 362 -16719 372 -16666
rect 655 -16718 665 -16665
rect 718 -16718 728 -16665
rect 835 -16718 845 -16665
rect 898 -16718 908 -16665
rect 1011 -16718 1021 -16665
rect 1074 -16718 1084 -16665
rect 1367 -16718 1377 -16665
rect 1430 -16718 1440 -16665
rect 1725 -16718 1735 -16665
rect 1788 -16718 1798 -16665
rect 2080 -16717 2090 -16664
rect 2143 -16717 2153 -16664
rect 2455 -16665 2489 -16400
rect 2523 -16438 2599 -16432
rect 2523 -16472 2539 -16438
rect 2583 -16472 2599 -16438
rect 2523 -16488 2599 -16472
rect 2701 -16438 2777 -16432
rect 2701 -16472 2717 -16438
rect 2761 -16472 2777 -16438
rect 2701 -16488 2777 -16472
rect 2544 -16542 2578 -16488
rect 2722 -16541 2756 -16488
rect 2524 -16595 2534 -16542
rect 2587 -16595 2597 -16542
rect 2703 -16594 2713 -16541
rect 2766 -16594 2776 -16541
rect 2811 -16665 2845 -16400
rect 2879 -16438 2955 -16432
rect 2879 -16472 2895 -16438
rect 2939 -16472 2955 -16438
rect 2879 -16488 2955 -16472
rect 3057 -16438 3133 -16432
rect 3057 -16472 3073 -16438
rect 3117 -16472 3133 -16438
rect 3057 -16488 3133 -16472
rect 2901 -16542 2935 -16488
rect 3079 -16542 3113 -16488
rect 2881 -16595 2891 -16542
rect 2944 -16595 2954 -16542
rect 3060 -16595 3070 -16542
rect 3123 -16595 3133 -16542
rect 3167 -16664 3201 -16400
rect 3235 -16438 3311 -16432
rect 3235 -16472 3251 -16438
rect 3295 -16472 3311 -16438
rect 3235 -16488 3311 -16472
rect 3413 -16438 3489 -16432
rect 3413 -16472 3429 -16438
rect 3473 -16472 3489 -16438
rect 3413 -16488 3489 -16472
rect 3257 -16542 3291 -16488
rect 3239 -16595 3249 -16542
rect 3302 -16595 3312 -16542
rect 2435 -16718 2445 -16665
rect 2498 -16718 2508 -16665
rect 2791 -16718 2801 -16665
rect 2854 -16718 2864 -16665
rect 3147 -16717 3157 -16664
rect 3210 -16717 3220 -16664
rect 3524 -16666 3558 -16400
rect 3591 -16438 3667 -16432
rect 3591 -16472 3607 -16438
rect 3651 -16472 3667 -16438
rect 3591 -16488 3667 -16472
rect 3769 -16438 3845 -16432
rect 3769 -16472 3785 -16438
rect 3829 -16472 3845 -16438
rect 3769 -16488 3845 -16472
rect 3879 -16665 3913 -16400
rect 3947 -16438 4023 -16432
rect 3947 -16472 3963 -16438
rect 4007 -16472 4023 -16438
rect 3947 -16488 4023 -16472
rect 4238 -16542 4291 -15592
rect 5021 -15593 5031 -15540
rect 5084 -15593 5094 -15540
rect 4228 -16595 4238 -16542
rect 4291 -16595 4301 -16542
rect -4802 -17171 -4792 -17118
rect -4739 -17171 -4729 -17118
rect -3945 -17170 -3935 -17118
rect -3883 -17170 -3873 -17118
rect 846 -17251 899 -16718
rect 3504 -16719 3514 -16666
rect 3567 -16719 3577 -16666
rect 3858 -16718 3868 -16665
rect 3921 -16718 3931 -16665
rect 5031 -16782 5084 -15593
rect 5400 -15653 5453 -13598
rect 5534 -13672 5587 -13349
rect 5524 -13725 5534 -13672
rect 5587 -13725 5597 -13672
rect 6912 -13922 6946 -12074
rect 8940 -13486 8950 -13433
rect 9003 -13486 9013 -13433
rect 9295 -13486 9305 -13433
rect 9358 -13486 9368 -13433
rect 8762 -13609 8772 -13556
rect 8825 -13609 8835 -13556
rect 7516 -13725 7526 -13672
rect 7579 -13725 7589 -13672
rect 7338 -13849 7348 -13796
rect 7401 -13849 7411 -13796
rect 5823 -13975 5833 -13922
rect 5886 -13975 5896 -13922
rect 6003 -13975 6013 -13922
rect 6066 -13975 6076 -13922
rect 5843 -14032 5877 -13975
rect 6022 -14032 6056 -13975
rect 6180 -13976 6190 -13923
rect 6243 -13976 6253 -13923
rect 6359 -13975 6369 -13922
rect 6422 -13975 6432 -13922
rect 6200 -14032 6234 -13976
rect 6378 -14032 6412 -13975
rect 6537 -13976 6547 -13923
rect 6600 -13976 6610 -13923
rect 6715 -13975 6725 -13922
rect 6778 -13975 6788 -13922
rect 6892 -13975 6902 -13922
rect 6955 -13975 6965 -13922
rect 6556 -14032 6590 -13976
rect 6734 -14032 6768 -13975
rect 6912 -14032 6946 -13975
rect 5645 -14048 5721 -14032
rect 5823 -14048 5899 -14032
rect 5577 -14082 5661 -14048
rect 5705 -14082 5790 -14048
rect 5577 -14120 5611 -14082
rect 5645 -14088 5721 -14082
rect 5756 -14120 5790 -14082
rect 5823 -14082 5839 -14048
rect 5883 -14082 5899 -14048
rect 5823 -14088 5899 -14082
rect 6001 -14048 6077 -14032
rect 6001 -14082 6017 -14048
rect 6061 -14082 6077 -14048
rect 6001 -14088 6077 -14082
rect 6179 -14048 6255 -14032
rect 6179 -14082 6195 -14048
rect 6239 -14082 6255 -14048
rect 6179 -14088 6255 -14082
rect 6357 -14048 6433 -14032
rect 6357 -14082 6373 -14048
rect 6417 -14082 6433 -14048
rect 6357 -14088 6433 -14082
rect 6535 -14048 6611 -14032
rect 6535 -14082 6551 -14048
rect 6595 -14082 6611 -14048
rect 6535 -14088 6611 -14082
rect 6713 -14048 6789 -14032
rect 6713 -14082 6729 -14048
rect 6773 -14082 6789 -14048
rect 6713 -14088 6789 -14082
rect 6891 -14048 6967 -14032
rect 6891 -14082 6907 -14048
rect 6951 -14082 6967 -14048
rect 6891 -14088 6967 -14082
rect 7069 -14048 7145 -14032
rect 7247 -14048 7323 -14032
rect 7069 -14082 7085 -14048
rect 7129 -14082 7263 -14048
rect 7307 -14082 7323 -14048
rect 7069 -14088 7145 -14082
rect 7179 -14120 7213 -14082
rect 7247 -14088 7323 -14082
rect 7357 -14120 7391 -13849
rect 7427 -13975 7437 -13922
rect 7490 -13975 7500 -13922
rect 7446 -14032 7480 -13975
rect 7425 -14048 7501 -14032
rect 7425 -14082 7441 -14048
rect 7485 -14082 7501 -14048
rect 7425 -14088 7501 -14082
rect 7535 -14120 7569 -13725
rect 7872 -13726 7882 -13673
rect 7935 -13726 7945 -13673
rect 8228 -13724 8238 -13671
rect 8291 -13724 8301 -13671
rect 7694 -13848 7704 -13795
rect 7757 -13848 7767 -13795
rect 7605 -13975 7615 -13922
rect 7668 -13975 7678 -13922
rect 7624 -14032 7658 -13975
rect 7603 -14048 7679 -14032
rect 7603 -14082 7619 -14048
rect 7663 -14082 7679 -14048
rect 7603 -14088 7679 -14082
rect 7713 -14120 7747 -13848
rect 7783 -13976 7793 -13923
rect 7846 -13976 7856 -13923
rect 7802 -14032 7836 -13976
rect 7781 -14048 7857 -14032
rect 7781 -14082 7797 -14048
rect 7841 -14082 7857 -14048
rect 7781 -14088 7857 -14082
rect 7892 -14120 7926 -13726
rect 8051 -13849 8061 -13796
rect 8114 -13849 8124 -13796
rect 7960 -13975 7970 -13922
rect 8023 -13975 8033 -13922
rect 7980 -14032 8014 -13975
rect 7959 -14048 8035 -14032
rect 7959 -14082 7975 -14048
rect 8019 -14082 8035 -14048
rect 7959 -14088 8035 -14082
rect 8069 -14120 8103 -13849
rect 8138 -13975 8148 -13922
rect 8201 -13975 8211 -13922
rect 8158 -14032 8192 -13975
rect 8137 -14048 8213 -14032
rect 8137 -14082 8153 -14048
rect 8197 -14082 8213 -14048
rect 8137 -14088 8213 -14082
rect 8248 -14120 8282 -13724
rect 8405 -13849 8415 -13796
rect 8468 -13849 8478 -13796
rect 8316 -13975 8326 -13922
rect 8379 -13975 8389 -13922
rect 8336 -14032 8370 -13975
rect 8315 -14048 8391 -14032
rect 8315 -14082 8331 -14048
rect 8375 -14082 8391 -14048
rect 8315 -14088 8391 -14082
rect 8425 -14120 8459 -13849
rect 8493 -14048 8569 -14032
rect 8671 -14048 8747 -14032
rect 8493 -14082 8509 -14048
rect 8553 -14082 8687 -14048
rect 8731 -14082 8747 -14048
rect 8493 -14088 8569 -14082
rect 8603 -14120 8637 -14082
rect 8671 -14088 8747 -14082
rect 8781 -14120 8815 -13609
rect 8851 -13975 8861 -13922
rect 8914 -13975 8924 -13922
rect 8871 -14032 8905 -13975
rect 8849 -14048 8925 -14032
rect 8849 -14082 8865 -14048
rect 8909 -14082 8925 -14048
rect 8849 -14088 8925 -14082
rect 8960 -14120 8994 -13486
rect 9117 -13609 9127 -13556
rect 9180 -13609 9190 -13556
rect 9028 -13975 9038 -13922
rect 9091 -13975 9101 -13922
rect 9048 -14032 9082 -13975
rect 9027 -14048 9103 -14032
rect 9027 -14082 9043 -14048
rect 9087 -14082 9103 -14048
rect 9027 -14088 9103 -14082
rect 9137 -14120 9171 -13609
rect 9207 -13975 9217 -13922
rect 9270 -13975 9280 -13922
rect 9227 -14032 9261 -13975
rect 9205 -14048 9281 -14032
rect 9205 -14082 9221 -14048
rect 9265 -14082 9281 -14048
rect 9205 -14088 9281 -14082
rect 9315 -14120 9349 -13486
rect 9473 -13609 9483 -13556
rect 9536 -13609 9546 -13556
rect 9384 -13975 9394 -13922
rect 9447 -13975 9457 -13922
rect 9404 -14032 9438 -13975
rect 9383 -14048 9459 -14032
rect 9383 -14082 9399 -14048
rect 9443 -14082 9459 -14048
rect 9383 -14088 9459 -14082
rect 9493 -14120 9527 -13609
rect 11432 -13725 11442 -13672
rect 11495 -13725 11505 -13672
rect 11788 -13725 11798 -13672
rect 11851 -13725 11861 -13672
rect 11254 -13849 11264 -13796
rect 11317 -13849 11327 -13796
rect 9919 -13976 9929 -13923
rect 9982 -13976 9992 -13923
rect 10098 -13975 10108 -13922
rect 10161 -13975 10171 -13922
rect 9938 -14032 9972 -13976
rect 10117 -14032 10151 -13975
rect 10274 -13976 10284 -13923
rect 10337 -13976 10347 -13923
rect 10452 -13976 10462 -13923
rect 10515 -13976 10525 -13923
rect 10630 -13975 10640 -13922
rect 10693 -13975 10703 -13922
rect 10294 -14032 10328 -13976
rect 10472 -14032 10506 -13976
rect 10650 -14032 10684 -13975
rect 10809 -13976 10819 -13923
rect 10872 -13976 10882 -13923
rect 10828 -14032 10862 -13976
rect 9561 -14048 9637 -14032
rect 9739 -14048 9815 -14032
rect 9561 -14082 9577 -14048
rect 9621 -14082 9755 -14048
rect 9799 -14082 9815 -14048
rect 9561 -14088 9637 -14082
rect 9671 -14120 9705 -14082
rect 9739 -14088 9815 -14082
rect 9917 -14048 9993 -14032
rect 9917 -14082 9933 -14048
rect 9977 -14082 9993 -14048
rect 9917 -14088 9993 -14082
rect 10095 -14048 10171 -14032
rect 10095 -14082 10111 -14048
rect 10155 -14082 10171 -14048
rect 10095 -14088 10171 -14082
rect 10273 -14048 10349 -14032
rect 10273 -14082 10289 -14048
rect 10333 -14082 10349 -14048
rect 10273 -14088 10349 -14082
rect 10451 -14048 10527 -14032
rect 10451 -14082 10467 -14048
rect 10511 -14082 10527 -14048
rect 10451 -14088 10527 -14082
rect 10629 -14048 10705 -14032
rect 10629 -14082 10645 -14048
rect 10689 -14082 10705 -14048
rect 10629 -14088 10705 -14082
rect 10807 -14048 10883 -14032
rect 10807 -14082 10823 -14048
rect 10867 -14082 10883 -14048
rect 10807 -14088 10883 -14082
rect 10985 -14048 11061 -14032
rect 11163 -14048 11239 -14032
rect 10985 -14082 11001 -14048
rect 11045 -14082 11179 -14048
rect 11223 -14082 11239 -14048
rect 10985 -14088 11061 -14082
rect 11095 -14120 11129 -14082
rect 11163 -14088 11239 -14082
rect 11273 -14120 11307 -13849
rect 11343 -13975 11353 -13922
rect 11406 -13975 11416 -13922
rect 11362 -14032 11396 -13975
rect 11341 -14048 11417 -14032
rect 11341 -14082 11357 -14048
rect 11401 -14082 11417 -14048
rect 11341 -14088 11417 -14082
rect 11452 -14120 11486 -13725
rect 11610 -13850 11620 -13797
rect 11673 -13850 11683 -13797
rect 11520 -13975 11530 -13922
rect 11583 -13975 11593 -13922
rect 11540 -14032 11574 -13975
rect 11519 -14048 11595 -14032
rect 11519 -14082 11535 -14048
rect 11579 -14082 11595 -14048
rect 11519 -14088 11595 -14082
rect 11630 -14120 11664 -13850
rect 11699 -13975 11709 -13922
rect 11762 -13975 11772 -13922
rect 11719 -14032 11753 -13975
rect 11697 -14048 11773 -14032
rect 11697 -14082 11713 -14048
rect 11757 -14082 11773 -14048
rect 11697 -14088 11773 -14082
rect 11807 -14120 11841 -13725
rect 12142 -13726 12152 -13673
rect 12205 -13726 12215 -13673
rect 12499 -13725 12509 -13672
rect 12562 -13725 12572 -13672
rect 11967 -13849 11977 -13796
rect 12030 -13849 12040 -13796
rect 11876 -13976 11886 -13923
rect 11939 -13976 11949 -13923
rect 11895 -14032 11929 -13976
rect 11875 -14048 11951 -14032
rect 11875 -14082 11891 -14048
rect 11935 -14082 11951 -14048
rect 11875 -14088 11951 -14082
rect 11986 -14120 12020 -13849
rect 12054 -13975 12064 -13922
rect 12117 -13975 12127 -13922
rect 12073 -14032 12107 -13975
rect 12053 -14048 12129 -14032
rect 12053 -14082 12069 -14048
rect 12113 -14082 12129 -14048
rect 12053 -14088 12129 -14082
rect 12162 -14120 12196 -13726
rect 12324 -13849 12334 -13796
rect 12387 -13849 12397 -13796
rect 12232 -13976 12242 -13923
rect 12295 -13976 12305 -13923
rect 12252 -14032 12286 -13976
rect 12231 -14048 12307 -14032
rect 12231 -14082 12247 -14048
rect 12291 -14082 12307 -14048
rect 12231 -14088 12307 -14082
rect 12342 -14120 12376 -13849
rect 12410 -13975 12420 -13922
rect 12473 -13975 12483 -13922
rect 12430 -14032 12464 -13975
rect 12409 -14048 12485 -14032
rect 12409 -14082 12425 -14048
rect 12469 -14082 12485 -14048
rect 12409 -14088 12485 -14082
rect 12519 -14048 12553 -13725
rect 12587 -14048 12663 -14032
rect 12519 -14082 12603 -14048
rect 12647 -14082 12731 -14048
rect 12519 -14120 12553 -14082
rect 12587 -14088 12663 -14082
rect 12697 -14120 12731 -14082
rect 5571 -14132 5617 -14120
rect 5571 -14388 5577 -14132
rect 5611 -14388 5617 -14132
rect 5571 -14400 5617 -14388
rect 5749 -14132 5795 -14120
rect 5749 -14388 5755 -14132
rect 5789 -14388 5795 -14132
rect 5749 -14400 5795 -14388
rect 5927 -14132 5973 -14120
rect 5927 -14388 5933 -14132
rect 5967 -14388 5973 -14132
rect 5927 -14400 5973 -14388
rect 6105 -14132 6151 -14120
rect 6105 -14388 6111 -14132
rect 6145 -14388 6151 -14132
rect 6105 -14400 6151 -14388
rect 6283 -14132 6329 -14120
rect 6283 -14388 6289 -14132
rect 6323 -14388 6329 -14132
rect 6283 -14400 6329 -14388
rect 6461 -14132 6507 -14120
rect 6461 -14388 6467 -14132
rect 6501 -14388 6507 -14132
rect 6461 -14400 6507 -14388
rect 6639 -14132 6685 -14120
rect 6639 -14388 6645 -14132
rect 6679 -14388 6685 -14132
rect 6639 -14400 6685 -14388
rect 6817 -14132 6863 -14120
rect 6817 -14388 6823 -14132
rect 6857 -14388 6863 -14132
rect 6817 -14400 6863 -14388
rect 6995 -14132 7041 -14120
rect 6995 -14388 7001 -14132
rect 7035 -14388 7041 -14132
rect 6995 -14400 7041 -14388
rect 7173 -14132 7219 -14120
rect 7173 -14388 7179 -14132
rect 7213 -14388 7219 -14132
rect 7173 -14400 7219 -14388
rect 7351 -14132 7397 -14120
rect 7351 -14388 7357 -14132
rect 7391 -14388 7397 -14132
rect 7351 -14400 7397 -14388
rect 7529 -14132 7575 -14120
rect 7529 -14388 7535 -14132
rect 7569 -14388 7575 -14132
rect 7529 -14400 7575 -14388
rect 7707 -14132 7753 -14120
rect 7707 -14388 7713 -14132
rect 7747 -14388 7753 -14132
rect 7707 -14400 7753 -14388
rect 7885 -14132 7931 -14120
rect 7885 -14388 7891 -14132
rect 7925 -14388 7931 -14132
rect 7885 -14400 7931 -14388
rect 8063 -14132 8109 -14120
rect 8063 -14388 8069 -14132
rect 8103 -14388 8109 -14132
rect 8063 -14400 8109 -14388
rect 8241 -14132 8287 -14120
rect 8241 -14388 8247 -14132
rect 8281 -14388 8287 -14132
rect 8241 -14400 8287 -14388
rect 8419 -14132 8465 -14120
rect 8419 -14388 8425 -14132
rect 8459 -14388 8465 -14132
rect 8419 -14400 8465 -14388
rect 8597 -14132 8643 -14120
rect 8597 -14388 8603 -14132
rect 8637 -14388 8643 -14132
rect 8597 -14400 8643 -14388
rect 8775 -14132 8821 -14120
rect 8775 -14388 8781 -14132
rect 8815 -14388 8821 -14132
rect 8775 -14400 8821 -14388
rect 8953 -14132 8999 -14120
rect 8953 -14388 8959 -14132
rect 8993 -14388 8999 -14132
rect 8953 -14400 8999 -14388
rect 9131 -14132 9177 -14120
rect 9131 -14388 9137 -14132
rect 9171 -14388 9177 -14132
rect 9131 -14400 9177 -14388
rect 9309 -14132 9355 -14120
rect 9309 -14388 9315 -14132
rect 9349 -14388 9355 -14132
rect 9309 -14400 9355 -14388
rect 9487 -14132 9533 -14120
rect 9487 -14388 9493 -14132
rect 9527 -14388 9533 -14132
rect 9487 -14400 9533 -14388
rect 9665 -14132 9711 -14120
rect 9665 -14388 9671 -14132
rect 9705 -14388 9711 -14132
rect 9665 -14400 9711 -14388
rect 9843 -14132 9889 -14120
rect 9843 -14388 9849 -14132
rect 9883 -14388 9889 -14132
rect 9843 -14400 9889 -14388
rect 10021 -14132 10067 -14120
rect 10021 -14388 10027 -14132
rect 10061 -14388 10067 -14132
rect 10021 -14400 10067 -14388
rect 10199 -14132 10245 -14120
rect 10199 -14388 10205 -14132
rect 10239 -14388 10245 -14132
rect 10199 -14400 10245 -14388
rect 10377 -14132 10423 -14120
rect 10377 -14388 10383 -14132
rect 10417 -14388 10423 -14132
rect 10377 -14400 10423 -14388
rect 10555 -14132 10601 -14120
rect 10555 -14388 10561 -14132
rect 10595 -14388 10601 -14132
rect 10555 -14400 10601 -14388
rect 10733 -14132 10779 -14120
rect 10733 -14388 10739 -14132
rect 10773 -14388 10779 -14132
rect 10733 -14400 10779 -14388
rect 10911 -14132 10957 -14120
rect 10911 -14388 10917 -14132
rect 10951 -14388 10957 -14132
rect 10911 -14400 10957 -14388
rect 11089 -14132 11135 -14120
rect 11089 -14388 11095 -14132
rect 11129 -14388 11135 -14132
rect 11089 -14400 11135 -14388
rect 11267 -14132 11313 -14120
rect 11267 -14388 11273 -14132
rect 11307 -14388 11313 -14132
rect 11267 -14400 11313 -14388
rect 11445 -14132 11491 -14120
rect 11445 -14388 11451 -14132
rect 11485 -14388 11491 -14132
rect 11445 -14400 11491 -14388
rect 11623 -14132 11669 -14120
rect 11623 -14388 11629 -14132
rect 11663 -14388 11669 -14132
rect 11623 -14400 11669 -14388
rect 11801 -14132 11847 -14120
rect 11801 -14388 11807 -14132
rect 11841 -14388 11847 -14132
rect 11801 -14400 11847 -14388
rect 11979 -14132 12025 -14120
rect 11979 -14388 11985 -14132
rect 12019 -14388 12025 -14132
rect 11979 -14400 12025 -14388
rect 12157 -14132 12203 -14120
rect 12157 -14388 12163 -14132
rect 12197 -14388 12203 -14132
rect 12157 -14400 12203 -14388
rect 12335 -14132 12381 -14120
rect 12335 -14388 12341 -14132
rect 12375 -14388 12381 -14132
rect 12335 -14400 12381 -14388
rect 12513 -14132 12559 -14120
rect 12513 -14388 12519 -14132
rect 12553 -14388 12559 -14132
rect 12513 -14400 12559 -14388
rect 12691 -14132 12737 -14120
rect 12691 -14388 12697 -14132
rect 12731 -14388 12737 -14132
rect 12691 -14400 12737 -14388
rect 5645 -14438 5721 -14432
rect 5645 -14472 5661 -14438
rect 5705 -14472 5721 -14438
rect 5645 -14488 5721 -14472
rect 5756 -14545 5790 -14400
rect 5823 -14438 5899 -14432
rect 5823 -14472 5839 -14438
rect 5883 -14472 5899 -14438
rect 5823 -14488 5899 -14472
rect 5736 -14598 5746 -14545
rect 5799 -14598 5809 -14545
rect 5843 -15032 5877 -14488
rect 5933 -14658 5967 -14400
rect 6001 -14438 6077 -14432
rect 6001 -14472 6017 -14438
rect 6061 -14472 6077 -14438
rect 6001 -14488 6077 -14472
rect 5914 -14711 5924 -14658
rect 5977 -14711 5987 -14658
rect 6022 -15032 6056 -14488
rect 6111 -14545 6145 -14400
rect 6179 -14438 6255 -14432
rect 6179 -14472 6195 -14438
rect 6239 -14472 6255 -14438
rect 6179 -14488 6255 -14472
rect 6091 -14598 6101 -14545
rect 6154 -14598 6164 -14545
rect 6200 -15032 6234 -14488
rect 6289 -14658 6323 -14400
rect 6357 -14438 6433 -14432
rect 6357 -14472 6373 -14438
rect 6417 -14472 6433 -14438
rect 6357 -14488 6433 -14472
rect 6269 -14711 6279 -14658
rect 6332 -14711 6342 -14658
rect 6378 -15032 6412 -14488
rect 6468 -14545 6502 -14400
rect 6535 -14438 6611 -14432
rect 6535 -14472 6551 -14438
rect 6595 -14472 6611 -14438
rect 6535 -14488 6611 -14472
rect 6449 -14598 6459 -14545
rect 6512 -14598 6522 -14545
rect 6557 -15032 6591 -14488
rect 6645 -14658 6679 -14400
rect 6713 -14438 6789 -14432
rect 6713 -14472 6729 -14438
rect 6773 -14472 6789 -14438
rect 6713 -14488 6789 -14472
rect 6823 -14545 6857 -14400
rect 6891 -14438 6967 -14432
rect 6891 -14472 6907 -14438
rect 6951 -14472 6967 -14438
rect 6891 -14488 6967 -14472
rect 6803 -14598 6813 -14545
rect 6866 -14598 6876 -14545
rect 7000 -14658 7034 -14400
rect 7069 -14438 7145 -14432
rect 7069 -14472 7085 -14438
rect 7129 -14472 7145 -14438
rect 7069 -14488 7145 -14472
rect 6626 -14711 6636 -14658
rect 6689 -14711 6699 -14658
rect 6981 -14711 6991 -14658
rect 7044 -14711 7054 -14658
rect 7179 -14749 7213 -14400
rect 7247 -14438 7323 -14432
rect 7247 -14472 7263 -14438
rect 7307 -14472 7323 -14438
rect 7247 -14488 7323 -14472
rect 6822 -14783 7213 -14749
rect 5645 -15047 5721 -15032
rect 5575 -15048 5789 -15047
rect 5575 -15081 5661 -15048
rect 5575 -15120 5609 -15081
rect 5645 -15082 5661 -15081
rect 5705 -15081 5789 -15048
rect 5705 -15082 5721 -15081
rect 5645 -15088 5721 -15082
rect 5755 -15120 5789 -15081
rect 5823 -15048 5899 -15032
rect 5823 -15082 5839 -15048
rect 5883 -15082 5899 -15048
rect 5823 -15088 5899 -15082
rect 6001 -15048 6077 -15032
rect 6001 -15082 6017 -15048
rect 6061 -15082 6077 -15048
rect 6001 -15088 6077 -15082
rect 6179 -15048 6255 -15032
rect 6179 -15082 6195 -15048
rect 6239 -15082 6255 -15048
rect 6179 -15088 6255 -15082
rect 6357 -15048 6433 -15032
rect 6357 -15082 6373 -15048
rect 6417 -15082 6433 -15048
rect 6357 -15088 6433 -15082
rect 6535 -15048 6611 -15032
rect 6535 -15082 6551 -15048
rect 6595 -15082 6611 -15048
rect 6535 -15088 6611 -15082
rect 6713 -15048 6789 -15032
rect 6713 -15082 6729 -15048
rect 6773 -15082 6789 -15048
rect 6713 -15088 6789 -15082
rect 6822 -15120 6856 -14783
rect 7357 -14824 7391 -14400
rect 7425 -14438 7501 -14432
rect 7425 -14472 7441 -14438
rect 7485 -14472 7501 -14438
rect 7425 -14488 7501 -14472
rect 6983 -14877 6993 -14824
rect 7046 -14877 7056 -14824
rect 7337 -14877 7347 -14824
rect 7400 -14877 7410 -14824
rect 6891 -15048 6967 -15032
rect 6891 -15082 6907 -15048
rect 6951 -15082 6967 -15048
rect 6891 -15088 6967 -15082
rect 7002 -15120 7036 -14877
rect 7070 -14976 7080 -14923
rect 7133 -14976 7143 -14923
rect 7090 -15032 7124 -14976
rect 7250 -14977 7260 -14924
rect 7313 -14977 7323 -14924
rect 7269 -15032 7303 -14977
rect 7069 -15048 7145 -15032
rect 7069 -15082 7085 -15048
rect 7129 -15082 7145 -15048
rect 7069 -15088 7145 -15082
rect 7247 -15048 7323 -15032
rect 7247 -15082 7263 -15048
rect 7307 -15082 7323 -15048
rect 7247 -15088 7323 -15082
rect 7357 -15120 7391 -14877
rect 7447 -14923 7481 -14488
rect 7429 -14976 7439 -14923
rect 7492 -14976 7502 -14923
rect 7447 -15032 7481 -14976
rect 7425 -15048 7501 -15032
rect 7425 -15082 7441 -15048
rect 7485 -15082 7501 -15048
rect 7425 -15088 7501 -15082
rect 7535 -15120 7569 -14400
rect 7603 -14438 7679 -14432
rect 7603 -14472 7619 -14438
rect 7663 -14472 7679 -14438
rect 7603 -14488 7679 -14472
rect 7781 -14438 7857 -14432
rect 7781 -14472 7797 -14438
rect 7841 -14472 7857 -14438
rect 7781 -14488 7857 -14472
rect 7959 -14438 8035 -14432
rect 7959 -14472 7975 -14438
rect 8019 -14472 8035 -14438
rect 7959 -14488 8035 -14472
rect 8137 -14438 8213 -14432
rect 8137 -14472 8153 -14438
rect 8197 -14472 8213 -14438
rect 8137 -14488 8213 -14472
rect 8315 -14438 8391 -14432
rect 8315 -14472 8331 -14438
rect 8375 -14472 8391 -14438
rect 8315 -14488 8391 -14472
rect 8493 -14438 8569 -14432
rect 8493 -14472 8509 -14438
rect 8553 -14472 8569 -14438
rect 8493 -14488 8569 -14472
rect 8671 -14438 8747 -14432
rect 8671 -14472 8687 -14438
rect 8731 -14472 8747 -14438
rect 8671 -14488 8747 -14472
rect 8849 -14438 8925 -14432
rect 8849 -14472 8865 -14438
rect 8909 -14472 8925 -14438
rect 8849 -14488 8925 -14472
rect 9027 -14438 9103 -14432
rect 9027 -14472 9043 -14438
rect 9087 -14472 9103 -14438
rect 9027 -14488 9103 -14472
rect 9205 -14438 9281 -14432
rect 9205 -14472 9221 -14438
rect 9265 -14472 9281 -14438
rect 9205 -14488 9281 -14472
rect 9383 -14438 9459 -14432
rect 9383 -14472 9399 -14438
rect 9443 -14472 9459 -14438
rect 9383 -14488 9459 -14472
rect 9561 -14438 9637 -14432
rect 9561 -14472 9577 -14438
rect 9621 -14472 9637 -14438
rect 9561 -14488 9637 -14472
rect 9739 -14438 9815 -14432
rect 9739 -14472 9755 -14438
rect 9799 -14472 9815 -14438
rect 9739 -14488 9815 -14472
rect 7625 -15032 7659 -14488
rect 7694 -14878 7704 -14825
rect 7757 -14878 7767 -14825
rect 7603 -15048 7679 -15032
rect 7603 -15082 7619 -15048
rect 7663 -15082 7679 -15048
rect 7603 -15088 7679 -15082
rect 7714 -15120 7748 -14878
rect 7802 -15032 7836 -14488
rect 8226 -14598 8236 -14545
rect 8289 -14598 8299 -14545
rect 8050 -14874 8060 -14821
rect 8113 -14874 8123 -14821
rect 7781 -15048 7857 -15032
rect 7781 -15082 7797 -15048
rect 7841 -15082 7857 -15048
rect 7781 -15088 7857 -15082
rect 7959 -15048 8035 -15032
rect 7959 -15082 7975 -15048
rect 8019 -15082 8035 -15048
rect 7959 -15088 8035 -15082
rect 8069 -15120 8103 -14874
rect 8137 -15048 8213 -15032
rect 8137 -15082 8153 -15048
rect 8197 -15082 8213 -15048
rect 8137 -15088 8213 -15082
rect 8247 -15120 8281 -14598
rect 8336 -14923 8370 -14488
rect 8407 -14710 8417 -14657
rect 8470 -14710 8480 -14657
rect 8317 -14976 8327 -14923
rect 8380 -14976 8390 -14923
rect 8336 -15032 8370 -14976
rect 8315 -15048 8391 -15032
rect 8315 -15082 8331 -15048
rect 8375 -15082 8391 -15048
rect 8315 -15088 8391 -15082
rect 8426 -15120 8460 -14710
rect 8514 -14806 8548 -14488
rect 8585 -14598 8595 -14545
rect 8648 -14598 8658 -14545
rect 8494 -14859 8504 -14806
rect 8557 -14859 8567 -14806
rect 8514 -14871 8548 -14859
rect 8495 -14977 8505 -14924
rect 8558 -14977 8568 -14924
rect 8514 -15032 8548 -14977
rect 8493 -15048 8569 -15032
rect 8493 -15082 8509 -15048
rect 8553 -15082 8569 -15048
rect 8493 -15088 8569 -15082
rect 8604 -15120 8638 -14598
rect 8762 -14711 8772 -14658
rect 8825 -14711 8835 -14658
rect 8692 -14924 8726 -14923
rect 8673 -14977 8683 -14924
rect 8736 -14977 8746 -14924
rect 8692 -15032 8726 -14977
rect 8671 -15048 8747 -15032
rect 8671 -15082 8687 -15048
rect 8731 -15082 8747 -15048
rect 8671 -15088 8747 -15082
rect 8781 -15120 8815 -14711
rect 8870 -15032 8904 -14488
rect 8940 -14599 8950 -14546
rect 9003 -14599 9013 -14546
rect 8849 -15048 8925 -15032
rect 8849 -15082 8865 -15048
rect 8909 -15082 8925 -15048
rect 8849 -15088 8925 -15082
rect 8960 -15120 8994 -14599
rect 9048 -15032 9082 -14488
rect 9117 -14712 9127 -14659
rect 9180 -14712 9190 -14659
rect 9027 -15048 9103 -15032
rect 9027 -15082 9043 -15048
rect 9087 -15082 9103 -15048
rect 9027 -15088 9103 -15082
rect 9137 -15120 9171 -14712
rect 9226 -15032 9260 -14488
rect 9294 -14598 9304 -14545
rect 9357 -14598 9367 -14545
rect 9205 -15048 9281 -15032
rect 9205 -15082 9221 -15048
rect 9265 -15082 9281 -15048
rect 9205 -15088 9281 -15082
rect 9314 -15120 9348 -14598
rect 9404 -15032 9438 -14488
rect 9651 -14598 9661 -14545
rect 9714 -14598 9724 -14545
rect 9473 -14711 9483 -14658
rect 9536 -14711 9546 -14658
rect 9383 -15048 9459 -15032
rect 9383 -15082 9399 -15048
rect 9443 -15082 9459 -15048
rect 9383 -15088 9459 -15082
rect 9493 -15120 9527 -14711
rect 9562 -14976 9572 -14923
rect 9625 -14976 9635 -14923
rect 9582 -15032 9616 -14976
rect 9561 -15048 9637 -15032
rect 9561 -15082 9577 -15048
rect 9621 -15082 9637 -15048
rect 9561 -15088 9637 -15082
rect 9671 -15120 9705 -14598
rect 9763 -14806 9797 -14488
rect 9848 -14659 9882 -14400
rect 9917 -14438 9993 -14432
rect 9917 -14472 9933 -14438
rect 9977 -14472 9993 -14438
rect 9917 -14488 9993 -14472
rect 9827 -14712 9837 -14659
rect 9890 -14712 9900 -14659
rect 9743 -14859 9753 -14806
rect 9806 -14859 9816 -14806
rect 9763 -14871 9797 -14859
rect 9740 -14976 9750 -14923
rect 9803 -14976 9813 -14923
rect 9760 -15032 9794 -14976
rect 9739 -15048 9815 -15032
rect 9739 -15082 9755 -15048
rect 9799 -15082 9815 -15048
rect 9739 -15088 9815 -15082
rect 9848 -15120 9882 -14712
rect 9939 -14923 9973 -14488
rect 10026 -14545 10060 -14400
rect 10095 -14438 10171 -14432
rect 10095 -14472 10111 -14438
rect 10155 -14472 10171 -14438
rect 10095 -14488 10171 -14472
rect 10006 -14598 10016 -14545
rect 10069 -14598 10079 -14545
rect 9919 -14976 9929 -14923
rect 9982 -14976 9992 -14923
rect 9939 -15032 9973 -14976
rect 9917 -15048 9993 -15032
rect 9917 -15082 9933 -15048
rect 9977 -15082 9993 -15048
rect 9917 -15088 9993 -15082
rect 10026 -15120 10060 -14598
rect 10205 -14658 10239 -14400
rect 10273 -14438 10349 -14432
rect 10273 -14472 10289 -14438
rect 10333 -14472 10349 -14438
rect 10273 -14488 10349 -14472
rect 10383 -14546 10417 -14400
rect 10451 -14438 10527 -14432
rect 10451 -14472 10467 -14438
rect 10511 -14472 10527 -14438
rect 10451 -14488 10527 -14472
rect 10363 -14599 10373 -14546
rect 10426 -14599 10436 -14546
rect 10186 -14711 10196 -14658
rect 10249 -14711 10259 -14658
rect 10185 -14875 10195 -14822
rect 10248 -14875 10258 -14822
rect 10095 -15048 10171 -15032
rect 10095 -15082 10111 -15048
rect 10155 -15082 10171 -15048
rect 10095 -15088 10171 -15082
rect 10205 -15120 10239 -14875
rect 10472 -15032 10506 -14488
rect 10560 -14658 10594 -14400
rect 10629 -14438 10705 -14432
rect 10629 -14472 10645 -14438
rect 10689 -14472 10705 -14438
rect 10629 -14488 10705 -14472
rect 10540 -14711 10550 -14658
rect 10603 -14711 10613 -14658
rect 10542 -14868 10552 -14815
rect 10605 -14868 10615 -14815
rect 10273 -15048 10349 -15032
rect 10273 -15082 10289 -15048
rect 10333 -15082 10349 -15048
rect 10273 -15088 10349 -15082
rect 10451 -15048 10527 -15032
rect 10451 -15082 10467 -15048
rect 10511 -15082 10527 -15048
rect 10451 -15088 10527 -15082
rect 10561 -15120 10595 -14868
rect 10650 -15032 10684 -14488
rect 10738 -14545 10772 -14400
rect 10807 -14438 10883 -14432
rect 10807 -14472 10823 -14438
rect 10867 -14472 10883 -14438
rect 10807 -14488 10883 -14472
rect 10719 -14598 10729 -14545
rect 10782 -14598 10792 -14545
rect 10828 -14923 10862 -14488
rect 10917 -14658 10951 -14400
rect 10985 -14438 11061 -14432
rect 10985 -14472 11001 -14438
rect 11045 -14472 11061 -14438
rect 10985 -14488 11061 -14472
rect 11096 -14658 11130 -14400
rect 11163 -14438 11239 -14432
rect 11163 -14472 11179 -14438
rect 11223 -14472 11239 -14438
rect 11163 -14488 11239 -14472
rect 10898 -14711 10908 -14658
rect 10961 -14711 10971 -14658
rect 11077 -14711 11087 -14658
rect 11140 -14711 11150 -14658
rect 10898 -14866 10908 -14813
rect 10961 -14866 10971 -14813
rect 11273 -14815 11307 -14400
rect 11341 -14438 11417 -14432
rect 11341 -14472 11357 -14438
rect 11401 -14472 11417 -14438
rect 11341 -14488 11417 -14472
rect 11519 -14438 11595 -14432
rect 11519 -14472 11535 -14438
rect 11579 -14472 11595 -14438
rect 11519 -14488 11595 -14472
rect 11697 -14438 11773 -14432
rect 11697 -14472 11713 -14438
rect 11757 -14472 11773 -14438
rect 11697 -14488 11773 -14472
rect 11875 -14438 11951 -14432
rect 11875 -14472 11891 -14438
rect 11935 -14472 11951 -14438
rect 11875 -14488 11951 -14472
rect 12053 -14438 12129 -14432
rect 12053 -14472 12069 -14438
rect 12113 -14472 12129 -14438
rect 12053 -14488 12129 -14472
rect 12231 -14438 12307 -14432
rect 12231 -14472 12247 -14438
rect 12291 -14472 12307 -14438
rect 12231 -14488 12307 -14472
rect 12409 -14438 12485 -14432
rect 12409 -14472 12425 -14438
rect 12469 -14472 12485 -14438
rect 12409 -14488 12485 -14472
rect 12587 -14438 12663 -14432
rect 12587 -14472 12603 -14438
rect 12647 -14472 12663 -14438
rect 12587 -14488 12663 -14472
rect 11430 -14709 11440 -14656
rect 11493 -14709 11503 -14656
rect 10809 -14976 10819 -14923
rect 10872 -14976 10882 -14923
rect 10828 -15032 10862 -14976
rect 10629 -15048 10705 -15032
rect 10629 -15082 10645 -15048
rect 10689 -15082 10705 -15048
rect 10629 -15088 10705 -15082
rect 10807 -15048 10883 -15032
rect 10807 -15082 10823 -15048
rect 10867 -15082 10883 -15048
rect 10807 -15088 10883 -15082
rect 10916 -15120 10950 -14866
rect 11254 -14868 11264 -14815
rect 11317 -14868 11327 -14815
rect 10986 -14976 10996 -14923
rect 11049 -14976 11059 -14923
rect 11165 -14976 11175 -14923
rect 11228 -14976 11238 -14923
rect 11006 -15032 11040 -14976
rect 11184 -15032 11218 -14976
rect 10985 -15048 11061 -15032
rect 10985 -15082 11001 -15048
rect 11045 -15082 11061 -15048
rect 10985 -15088 11061 -15082
rect 11163 -15048 11239 -15032
rect 11163 -15082 11179 -15048
rect 11223 -15082 11239 -15048
rect 11163 -15088 11239 -15082
rect 11273 -15120 11307 -14868
rect 11341 -15048 11417 -15032
rect 11341 -15082 11357 -15048
rect 11401 -15082 11417 -15048
rect 11341 -15088 11417 -15082
rect 11451 -15120 11485 -14709
rect 11717 -15032 11751 -14488
rect 11897 -15032 11931 -14488
rect 12075 -15032 12109 -14488
rect 12253 -15032 12287 -14488
rect 12430 -15032 12464 -14488
rect 11519 -15048 11595 -15032
rect 11519 -15082 11535 -15048
rect 11579 -15082 11595 -15048
rect 11519 -15088 11595 -15082
rect 11697 -15048 11773 -15032
rect 11697 -15082 11713 -15048
rect 11757 -15082 11773 -15048
rect 11697 -15088 11773 -15082
rect 11875 -15048 11951 -15032
rect 11875 -15082 11891 -15048
rect 11935 -15082 11951 -15048
rect 11875 -15088 11951 -15082
rect 12053 -15048 12129 -15032
rect 12053 -15082 12069 -15048
rect 12113 -15082 12129 -15048
rect 12053 -15088 12129 -15082
rect 12231 -15048 12307 -15032
rect 12231 -15082 12247 -15048
rect 12291 -15082 12307 -15048
rect 12231 -15088 12307 -15082
rect 12409 -15048 12485 -15032
rect 12409 -15082 12425 -15048
rect 12469 -15082 12485 -15048
rect 12587 -15048 12663 -15032
rect 12587 -15049 12603 -15048
rect 12409 -15088 12485 -15082
rect 12520 -15082 12603 -15049
rect 12647 -15049 12663 -15048
rect 12647 -15082 12730 -15049
rect 12520 -15083 12730 -15082
rect 12520 -15120 12554 -15083
rect 12587 -15088 12663 -15083
rect 12696 -15120 12730 -15083
rect 5571 -15132 5617 -15120
rect 5571 -15388 5577 -15132
rect 5611 -15388 5617 -15132
rect 5571 -15400 5617 -15388
rect 5749 -15132 5795 -15120
rect 5749 -15388 5755 -15132
rect 5789 -15388 5795 -15132
rect 5749 -15400 5795 -15388
rect 5927 -15132 5973 -15120
rect 5927 -15388 5933 -15132
rect 5967 -15388 5973 -15132
rect 5927 -15400 5973 -15388
rect 6105 -15132 6151 -15120
rect 6105 -15388 6111 -15132
rect 6145 -15388 6151 -15132
rect 6105 -15400 6151 -15388
rect 6283 -15132 6329 -15120
rect 6283 -15388 6289 -15132
rect 6323 -15388 6329 -15132
rect 6283 -15400 6329 -15388
rect 6461 -15132 6507 -15120
rect 6461 -15388 6467 -15132
rect 6501 -15388 6507 -15132
rect 6461 -15400 6507 -15388
rect 6639 -15132 6685 -15120
rect 6639 -15388 6645 -15132
rect 6679 -15388 6685 -15132
rect 6639 -15400 6685 -15388
rect 6817 -15132 6863 -15120
rect 6817 -15388 6823 -15132
rect 6857 -15388 6863 -15132
rect 6817 -15400 6863 -15388
rect 6995 -15132 7041 -15120
rect 6995 -15388 7001 -15132
rect 7035 -15388 7041 -15132
rect 6995 -15400 7041 -15388
rect 7173 -15132 7219 -15120
rect 7173 -15388 7179 -15132
rect 7213 -15388 7219 -15132
rect 7173 -15400 7219 -15388
rect 7351 -15132 7397 -15120
rect 7351 -15388 7357 -15132
rect 7391 -15388 7397 -15132
rect 7351 -15400 7397 -15388
rect 7529 -15132 7575 -15120
rect 7529 -15388 7535 -15132
rect 7569 -15388 7575 -15132
rect 7529 -15400 7575 -15388
rect 7707 -15132 7753 -15120
rect 7707 -15388 7713 -15132
rect 7747 -15388 7753 -15132
rect 7707 -15400 7753 -15388
rect 7885 -15132 7931 -15120
rect 7885 -15388 7891 -15132
rect 7925 -15388 7931 -15132
rect 7885 -15400 7931 -15388
rect 8063 -15132 8109 -15120
rect 8063 -15388 8069 -15132
rect 8103 -15388 8109 -15132
rect 8063 -15400 8109 -15388
rect 8241 -15132 8287 -15120
rect 8241 -15388 8247 -15132
rect 8281 -15388 8287 -15132
rect 8241 -15400 8287 -15388
rect 8419 -15132 8465 -15120
rect 8419 -15388 8425 -15132
rect 8459 -15388 8465 -15132
rect 8419 -15400 8465 -15388
rect 8597 -15132 8643 -15120
rect 8597 -15388 8603 -15132
rect 8637 -15388 8643 -15132
rect 8597 -15400 8643 -15388
rect 8775 -15132 8821 -15120
rect 8775 -15388 8781 -15132
rect 8815 -15388 8821 -15132
rect 8775 -15400 8821 -15388
rect 8953 -15132 8999 -15120
rect 8953 -15388 8959 -15132
rect 8993 -15388 8999 -15132
rect 8953 -15400 8999 -15388
rect 9131 -15132 9177 -15120
rect 9131 -15388 9137 -15132
rect 9171 -15388 9177 -15132
rect 9131 -15400 9177 -15388
rect 9309 -15132 9355 -15120
rect 9309 -15388 9315 -15132
rect 9349 -15388 9355 -15132
rect 9309 -15400 9355 -15388
rect 9487 -15132 9533 -15120
rect 9487 -15388 9493 -15132
rect 9527 -15388 9533 -15132
rect 9487 -15400 9533 -15388
rect 9665 -15132 9711 -15120
rect 9665 -15388 9671 -15132
rect 9705 -15388 9711 -15132
rect 9665 -15400 9711 -15388
rect 9843 -15132 9889 -15120
rect 9843 -15388 9849 -15132
rect 9883 -15388 9889 -15132
rect 9843 -15400 9889 -15388
rect 10021 -15132 10067 -15120
rect 10021 -15388 10027 -15132
rect 10061 -15388 10067 -15132
rect 10021 -15400 10067 -15388
rect 10199 -15132 10245 -15120
rect 10199 -15388 10205 -15132
rect 10239 -15388 10245 -15132
rect 10199 -15400 10245 -15388
rect 10377 -15132 10423 -15120
rect 10377 -15388 10383 -15132
rect 10417 -15388 10423 -15132
rect 10377 -15400 10423 -15388
rect 10555 -15132 10601 -15120
rect 10555 -15388 10561 -15132
rect 10595 -15388 10601 -15132
rect 10555 -15400 10601 -15388
rect 10733 -15132 10779 -15120
rect 10733 -15388 10739 -15132
rect 10773 -15388 10779 -15132
rect 10733 -15400 10779 -15388
rect 10911 -15132 10957 -15120
rect 10911 -15388 10917 -15132
rect 10951 -15388 10957 -15132
rect 10911 -15400 10957 -15388
rect 11089 -15132 11135 -15120
rect 11089 -15388 11095 -15132
rect 11129 -15388 11135 -15132
rect 11089 -15400 11135 -15388
rect 11267 -15132 11313 -15120
rect 11267 -15388 11273 -15132
rect 11307 -15388 11313 -15132
rect 11267 -15400 11313 -15388
rect 11445 -15132 11491 -15120
rect 11445 -15388 11451 -15132
rect 11485 -15388 11491 -15132
rect 11445 -15400 11491 -15388
rect 11623 -15132 11669 -15120
rect 11623 -15388 11629 -15132
rect 11663 -15388 11669 -15132
rect 11623 -15400 11669 -15388
rect 11801 -15132 11847 -15120
rect 11801 -15388 11807 -15132
rect 11841 -15388 11847 -15132
rect 11801 -15400 11847 -15388
rect 11979 -15132 12025 -15120
rect 11979 -15388 11985 -15132
rect 12019 -15388 12025 -15132
rect 11979 -15400 12025 -15388
rect 12157 -15132 12203 -15120
rect 12157 -15388 12163 -15132
rect 12197 -15388 12203 -15132
rect 12157 -15400 12203 -15388
rect 12335 -15132 12381 -15120
rect 12335 -15388 12341 -15132
rect 12375 -15388 12381 -15132
rect 12335 -15400 12381 -15388
rect 12513 -15132 12559 -15120
rect 12513 -15388 12519 -15132
rect 12553 -15388 12559 -15132
rect 12513 -15400 12559 -15388
rect 12691 -15132 12737 -15120
rect 12691 -15388 12697 -15132
rect 12731 -15388 12737 -15132
rect 12691 -15400 12737 -15388
rect 5645 -15438 5721 -15432
rect 5645 -15472 5661 -15438
rect 5705 -15472 5721 -15438
rect 5645 -15488 5721 -15472
rect 5755 -15539 5789 -15400
rect 5823 -15438 5899 -15432
rect 5823 -15472 5839 -15438
rect 5883 -15472 5899 -15438
rect 5823 -15488 5899 -15472
rect 5735 -15592 5745 -15539
rect 5798 -15592 5808 -15539
rect 5390 -15706 5400 -15653
rect 5453 -15706 5463 -15653
rect 5400 -16667 5453 -15706
rect 5737 -15803 5747 -15750
rect 5800 -15803 5810 -15750
rect 5645 -16048 5721 -16032
rect 5645 -16082 5661 -16048
rect 5705 -16082 5721 -16048
rect 5645 -16088 5721 -16082
rect 5756 -16120 5790 -15803
rect 5844 -16032 5878 -15488
rect 5933 -15652 5967 -15400
rect 6001 -15438 6077 -15432
rect 6001 -15472 6017 -15438
rect 6061 -15472 6077 -15438
rect 6001 -15488 6077 -15472
rect 5913 -15705 5923 -15652
rect 5976 -15705 5986 -15652
rect 5911 -16001 5921 -15948
rect 5974 -16001 5984 -15948
rect 5823 -16048 5899 -16032
rect 5823 -16082 5839 -16048
rect 5883 -16082 5899 -16048
rect 5823 -16088 5899 -16082
rect 5931 -16120 5965 -16001
rect 6022 -16032 6056 -15488
rect 6111 -15539 6145 -15400
rect 6179 -15438 6255 -15432
rect 6179 -15472 6195 -15438
rect 6239 -15472 6255 -15438
rect 6179 -15488 6255 -15472
rect 6091 -15592 6101 -15539
rect 6154 -15592 6164 -15539
rect 6091 -15802 6101 -15749
rect 6154 -15802 6164 -15749
rect 6001 -16048 6077 -16032
rect 6001 -16082 6017 -16048
rect 6061 -16082 6077 -16048
rect 6001 -16088 6077 -16082
rect 6112 -16120 6146 -15802
rect 6201 -16032 6235 -15488
rect 6289 -15652 6323 -15400
rect 6357 -15438 6433 -15432
rect 6357 -15472 6373 -15438
rect 6417 -15472 6433 -15438
rect 6357 -15488 6433 -15472
rect 6269 -15705 6279 -15652
rect 6332 -15705 6342 -15652
rect 6269 -16001 6279 -15948
rect 6332 -16001 6342 -15948
rect 6179 -16048 6255 -16032
rect 6179 -16082 6195 -16048
rect 6239 -16082 6255 -16048
rect 6179 -16088 6255 -16082
rect 6288 -16120 6322 -16001
rect 6379 -16032 6413 -15488
rect 6468 -15539 6502 -15400
rect 6535 -15438 6611 -15432
rect 6535 -15472 6551 -15438
rect 6595 -15472 6611 -15438
rect 6535 -15488 6611 -15472
rect 6448 -15592 6458 -15539
rect 6511 -15592 6521 -15539
rect 6446 -15803 6456 -15750
rect 6509 -15803 6519 -15750
rect 6357 -16048 6433 -16032
rect 6357 -16082 6373 -16048
rect 6417 -16082 6433 -16048
rect 6357 -16088 6433 -16082
rect 6467 -16120 6501 -15803
rect 6556 -16032 6590 -15488
rect 6645 -15652 6679 -15400
rect 6713 -15438 6789 -15432
rect 6822 -15438 6857 -15400
rect 6891 -15438 6967 -15432
rect 6713 -15472 6729 -15438
rect 6773 -15472 6907 -15438
rect 6951 -15472 6967 -15438
rect 6713 -15488 6789 -15472
rect 6625 -15705 6635 -15652
rect 6688 -15705 6698 -15652
rect 6703 -15804 6713 -15751
rect 6766 -15804 6776 -15751
rect 6624 -16001 6634 -15948
rect 6687 -16001 6697 -15948
rect 6734 -15956 6768 -15804
rect 6822 -15851 6856 -15472
rect 6891 -15488 6967 -15472
rect 6803 -15904 6813 -15851
rect 6866 -15904 6876 -15851
rect 7002 -15951 7036 -15400
rect 7069 -15438 7145 -15432
rect 7069 -15472 7085 -15438
rect 7129 -15472 7145 -15438
rect 7069 -15488 7145 -15472
rect 7179 -15750 7213 -15400
rect 7247 -15438 7323 -15432
rect 7247 -15472 7263 -15438
rect 7307 -15472 7323 -15438
rect 7247 -15488 7323 -15472
rect 7425 -15438 7501 -15432
rect 7425 -15472 7441 -15438
rect 7485 -15472 7501 -15438
rect 7425 -15488 7501 -15472
rect 7159 -15803 7169 -15750
rect 7222 -15803 7232 -15750
rect 7159 -15905 7169 -15852
rect 7222 -15905 7232 -15852
rect 6734 -15990 6858 -15956
rect 6535 -16048 6611 -16032
rect 6535 -16082 6551 -16048
rect 6595 -16082 6611 -16048
rect 6535 -16088 6611 -16082
rect 6644 -16120 6678 -16001
rect 6713 -16048 6789 -16032
rect 6713 -16082 6729 -16048
rect 6773 -16082 6789 -16048
rect 6713 -16088 6789 -16082
rect 6824 -16120 6858 -15990
rect 6984 -16004 6994 -15951
rect 7047 -16004 7057 -15951
rect 6891 -16048 6967 -16032
rect 6891 -16082 6907 -16048
rect 6951 -16082 6967 -16048
rect 6891 -16088 6967 -16082
rect 7002 -16120 7036 -16004
rect 7069 -16048 7145 -16032
rect 7069 -16082 7085 -16048
rect 7129 -16082 7145 -16048
rect 7069 -16088 7145 -16082
rect 7178 -16120 7212 -15905
rect 7447 -16032 7481 -15488
rect 7536 -15749 7570 -15400
rect 7603 -15438 7679 -15432
rect 7603 -15472 7619 -15438
rect 7663 -15472 7679 -15438
rect 7603 -15488 7679 -15472
rect 7781 -15438 7857 -15432
rect 7781 -15472 7797 -15438
rect 7841 -15472 7857 -15438
rect 7781 -15488 7857 -15472
rect 7516 -15802 7526 -15749
rect 7579 -15802 7589 -15749
rect 7516 -16006 7526 -15953
rect 7579 -16006 7589 -15953
rect 7247 -16048 7323 -16032
rect 7247 -16082 7263 -16048
rect 7307 -16082 7323 -16048
rect 7247 -16088 7323 -16082
rect 7425 -16048 7501 -16032
rect 7425 -16082 7441 -16048
rect 7485 -16082 7501 -16048
rect 7425 -16088 7501 -16082
rect 7535 -16120 7569 -16006
rect 7624 -16032 7658 -15488
rect 7803 -16032 7837 -15488
rect 7891 -15749 7925 -15400
rect 7959 -15438 8035 -15432
rect 8069 -15438 8103 -15400
rect 8137 -15438 8213 -15432
rect 7959 -15472 7975 -15438
rect 8019 -15472 8153 -15438
rect 8197 -15472 8213 -15438
rect 7959 -15488 8035 -15472
rect 7872 -15802 7882 -15749
rect 7935 -15802 7945 -15749
rect 8069 -15851 8103 -15472
rect 8137 -15488 8213 -15472
rect 8050 -15904 8060 -15851
rect 8113 -15904 8123 -15851
rect 8247 -15952 8281 -15400
rect 8315 -15438 8391 -15432
rect 8315 -15472 8331 -15438
rect 8375 -15472 8391 -15438
rect 8315 -15488 8391 -15472
rect 7871 -16005 7881 -15952
rect 7934 -16005 7944 -15952
rect 8227 -16005 8237 -15952
rect 8290 -16005 8300 -15952
rect 7603 -16048 7679 -16032
rect 7603 -16082 7619 -16048
rect 7663 -16082 7679 -16048
rect 7603 -16088 7679 -16082
rect 7781 -16048 7857 -16032
rect 7781 -16082 7797 -16048
rect 7841 -16082 7857 -16048
rect 7781 -16088 7857 -16082
rect 7891 -16120 7925 -16005
rect 7959 -16048 8035 -16032
rect 7959 -16082 7975 -16048
rect 8019 -16082 8035 -16048
rect 7959 -16088 8035 -16082
rect 8137 -16048 8213 -16032
rect 8137 -16082 8153 -16048
rect 8197 -16082 8213 -16048
rect 8137 -16088 8213 -16082
rect 8247 -16120 8281 -16005
rect 8336 -16032 8370 -15488
rect 8315 -16048 8391 -16032
rect 8315 -16082 8331 -16048
rect 8375 -16082 8391 -16048
rect 8315 -16088 8391 -16082
rect 8426 -16120 8460 -15400
rect 8493 -15438 8569 -15432
rect 8493 -15472 8509 -15438
rect 8553 -15472 8569 -15438
rect 8493 -15488 8569 -15472
rect 8671 -15438 8747 -15432
rect 8671 -15472 8687 -15438
rect 8731 -15472 8747 -15438
rect 8671 -15488 8747 -15472
rect 8849 -15438 8925 -15432
rect 8849 -15472 8865 -15438
rect 8909 -15472 8925 -15438
rect 8849 -15488 8925 -15472
rect 9027 -15438 9103 -15432
rect 9027 -15472 9043 -15438
rect 9087 -15472 9103 -15438
rect 9027 -15488 9103 -15472
rect 9205 -15438 9281 -15432
rect 9205 -15472 9221 -15438
rect 9265 -15472 9281 -15438
rect 9205 -15488 9281 -15472
rect 9383 -15438 9459 -15432
rect 9383 -15472 9399 -15438
rect 9443 -15472 9459 -15438
rect 9383 -15488 9459 -15472
rect 9561 -15438 9637 -15432
rect 9561 -15472 9577 -15438
rect 9621 -15472 9637 -15438
rect 9561 -15488 9637 -15472
rect 9739 -15438 9815 -15432
rect 9739 -15472 9755 -15438
rect 9799 -15472 9815 -15438
rect 9739 -15488 9815 -15472
rect 9917 -15438 9993 -15432
rect 9917 -15472 9933 -15438
rect 9977 -15472 9993 -15438
rect 9917 -15488 9993 -15472
rect 10095 -15438 10171 -15432
rect 10205 -15438 10239 -15400
rect 10273 -15438 10349 -15432
rect 10095 -15472 10111 -15438
rect 10155 -15472 10289 -15438
rect 10333 -15472 10349 -15438
rect 10095 -15488 10171 -15472
rect 8583 -15905 8593 -15852
rect 8646 -15905 8656 -15852
rect 8493 -16048 8569 -16032
rect 8493 -16082 8509 -16048
rect 8553 -16082 8569 -16048
rect 8493 -16088 8569 -16082
rect 8603 -16120 8637 -15905
rect 8870 -16032 8904 -15488
rect 9049 -16032 9083 -15488
rect 9226 -16032 9260 -15488
rect 9404 -16032 9438 -15488
rect 9653 -15905 9663 -15852
rect 9716 -15905 9726 -15852
rect 8671 -16048 8747 -16032
rect 8671 -16082 8687 -16048
rect 8731 -16082 8747 -16048
rect 8671 -16088 8747 -16082
rect 8849 -16048 8925 -16032
rect 8849 -16082 8865 -16048
rect 8909 -16082 8925 -16048
rect 8849 -16088 8925 -16082
rect 9027 -16048 9103 -16032
rect 9027 -16082 9043 -16048
rect 9087 -16082 9103 -16048
rect 9027 -16088 9103 -16082
rect 9205 -16048 9281 -16032
rect 9205 -16082 9221 -16048
rect 9265 -16082 9281 -16048
rect 9205 -16088 9281 -16082
rect 9383 -16048 9459 -16032
rect 9383 -16082 9399 -16048
rect 9443 -16082 9459 -16048
rect 9383 -16088 9459 -16082
rect 9561 -16048 9637 -16032
rect 9561 -16082 9577 -16048
rect 9621 -16082 9637 -16048
rect 9561 -16088 9637 -16082
rect 9672 -16120 9706 -15905
rect 9939 -16032 9973 -15488
rect 10205 -15852 10239 -15472
rect 10273 -15488 10349 -15472
rect 10383 -15751 10417 -15400
rect 10451 -15438 10527 -15432
rect 10451 -15472 10467 -15438
rect 10511 -15472 10527 -15438
rect 10451 -15488 10527 -15472
rect 10629 -15438 10705 -15432
rect 10629 -15472 10645 -15438
rect 10689 -15472 10705 -15438
rect 10629 -15488 10705 -15472
rect 10363 -15804 10373 -15751
rect 10426 -15804 10436 -15751
rect 10184 -15905 10194 -15852
rect 10247 -15905 10257 -15852
rect 10472 -16032 10506 -15488
rect 10650 -16032 10684 -15488
rect 10739 -15750 10773 -15400
rect 10807 -15438 10883 -15432
rect 10807 -15472 10823 -15438
rect 10867 -15472 10883 -15438
rect 10807 -15488 10883 -15472
rect 10720 -15803 10730 -15750
rect 10783 -15803 10793 -15750
rect 9739 -16048 9815 -16032
rect 9739 -16082 9755 -16048
rect 9799 -16082 9815 -16048
rect 9739 -16088 9815 -16082
rect 9917 -16048 9993 -16032
rect 9917 -16082 9933 -16048
rect 9977 -16082 9993 -16048
rect 9917 -16088 9993 -16082
rect 10095 -16048 10171 -16032
rect 10095 -16082 10111 -16048
rect 10155 -16082 10171 -16048
rect 10095 -16088 10171 -16082
rect 10273 -16048 10349 -16032
rect 10273 -16082 10289 -16048
rect 10333 -16082 10349 -16048
rect 10273 -16088 10349 -16082
rect 10451 -16048 10527 -16032
rect 10451 -16082 10467 -16048
rect 10511 -16082 10527 -16048
rect 10451 -16088 10527 -16082
rect 10629 -16048 10705 -16032
rect 10629 -16082 10645 -16048
rect 10689 -16082 10705 -16048
rect 10629 -16088 10705 -16082
rect 10739 -16120 10773 -15803
rect 10828 -16032 10862 -15488
rect 10807 -16048 10883 -16032
rect 10807 -16082 10823 -16048
rect 10867 -16082 10883 -16048
rect 10807 -16088 10883 -16082
rect 10916 -16120 10950 -15400
rect 10985 -15438 11061 -15432
rect 10985 -15472 11001 -15438
rect 11045 -15472 11061 -15438
rect 10985 -15488 11061 -15472
rect 11095 -15750 11129 -15400
rect 11163 -15438 11239 -15432
rect 11163 -15472 11179 -15438
rect 11223 -15472 11239 -15438
rect 11163 -15488 11239 -15472
rect 11341 -15438 11417 -15432
rect 11451 -15438 11485 -15400
rect 11519 -15438 11595 -15432
rect 11341 -15472 11357 -15438
rect 11401 -15472 11535 -15438
rect 11579 -15472 11595 -15438
rect 11341 -15488 11417 -15472
rect 11076 -15803 11086 -15750
rect 11139 -15803 11149 -15750
rect 11451 -15841 11485 -15472
rect 11519 -15488 11595 -15472
rect 11629 -15652 11663 -15400
rect 11697 -15438 11773 -15432
rect 11697 -15472 11713 -15438
rect 11757 -15472 11773 -15438
rect 11697 -15488 11773 -15472
rect 11609 -15705 11619 -15652
rect 11672 -15705 11682 -15652
rect 11629 -15706 11663 -15705
rect 11074 -15905 11084 -15852
rect 11137 -15905 11147 -15852
rect 11430 -15894 11440 -15841
rect 11493 -15894 11503 -15841
rect 11451 -15902 11485 -15894
rect 10985 -16048 11061 -16032
rect 10985 -16082 11001 -16048
rect 11045 -16082 11061 -16048
rect 10985 -16088 11061 -16082
rect 11094 -16120 11128 -15905
rect 11431 -16005 11441 -15952
rect 11494 -16005 11504 -15952
rect 11163 -16048 11239 -16032
rect 11163 -16082 11179 -16048
rect 11223 -16082 11239 -16048
rect 11163 -16088 11239 -16082
rect 11341 -16048 11417 -16032
rect 11341 -16082 11357 -16048
rect 11401 -16082 11417 -16048
rect 11341 -16088 11417 -16082
rect 11451 -16120 11485 -16005
rect 11718 -16032 11752 -15488
rect 11808 -15540 11842 -15400
rect 11875 -15438 11951 -15432
rect 11875 -15472 11891 -15438
rect 11935 -15472 11951 -15438
rect 11875 -15488 11951 -15472
rect 11788 -15593 11798 -15540
rect 11851 -15593 11861 -15540
rect 11787 -16005 11797 -15952
rect 11850 -16005 11860 -15952
rect 11519 -16048 11595 -16032
rect 11519 -16082 11535 -16048
rect 11579 -16082 11595 -16048
rect 11519 -16088 11595 -16082
rect 11697 -16048 11773 -16032
rect 11697 -16082 11713 -16048
rect 11757 -16082 11773 -16048
rect 11697 -16088 11773 -16082
rect 11806 -16120 11840 -16005
rect 11897 -16032 11931 -15488
rect 11985 -15652 12019 -15400
rect 12053 -15438 12129 -15432
rect 12053 -15472 12069 -15438
rect 12113 -15472 12129 -15438
rect 12053 -15488 12129 -15472
rect 11965 -15705 11975 -15652
rect 12028 -15705 12038 -15652
rect 12074 -16032 12108 -15488
rect 12165 -15539 12199 -15400
rect 12231 -15438 12307 -15432
rect 12231 -15472 12247 -15438
rect 12291 -15472 12307 -15438
rect 12231 -15488 12307 -15472
rect 12145 -15592 12155 -15539
rect 12208 -15592 12218 -15539
rect 12144 -16005 12154 -15952
rect 12207 -16005 12217 -15952
rect 11875 -16048 11951 -16032
rect 11875 -16082 11891 -16048
rect 11935 -16082 11951 -16048
rect 11875 -16088 11951 -16082
rect 12053 -16048 12129 -16032
rect 12053 -16082 12069 -16048
rect 12113 -16082 12129 -16048
rect 12053 -16088 12129 -16082
rect 12163 -16120 12197 -16005
rect 12252 -16032 12286 -15488
rect 12342 -15652 12376 -15400
rect 12409 -15438 12485 -15432
rect 12409 -15472 12425 -15438
rect 12469 -15472 12485 -15438
rect 12409 -15488 12485 -15472
rect 12322 -15705 12332 -15652
rect 12385 -15705 12395 -15652
rect 12431 -16032 12465 -15488
rect 12520 -15539 12554 -15400
rect 12587 -15438 12663 -15432
rect 12587 -15472 12603 -15438
rect 12647 -15472 12663 -15438
rect 12587 -15488 12663 -15472
rect 12501 -15592 12511 -15539
rect 12564 -15592 12574 -15539
rect 12501 -16005 12511 -15952
rect 12564 -16005 12574 -15952
rect 12231 -16048 12307 -16032
rect 12231 -16082 12247 -16048
rect 12291 -16082 12307 -16048
rect 12231 -16088 12307 -16082
rect 12409 -16048 12485 -16032
rect 12409 -16082 12425 -16048
rect 12469 -16082 12485 -16048
rect 12409 -16088 12485 -16082
rect 12520 -16120 12554 -16005
rect 12587 -16048 12663 -16032
rect 12587 -16082 12603 -16048
rect 12647 -16082 12663 -16048
rect 12587 -16088 12663 -16082
rect 5571 -16132 5617 -16120
rect 5571 -16388 5577 -16132
rect 5611 -16388 5617 -16132
rect 5571 -16400 5617 -16388
rect 5749 -16132 5795 -16120
rect 5749 -16388 5755 -16132
rect 5789 -16388 5795 -16132
rect 5749 -16400 5795 -16388
rect 5927 -16132 5973 -16120
rect 5927 -16388 5933 -16132
rect 5967 -16388 5973 -16132
rect 5927 -16400 5973 -16388
rect 6105 -16132 6151 -16120
rect 6105 -16388 6111 -16132
rect 6145 -16388 6151 -16132
rect 6105 -16400 6151 -16388
rect 6283 -16132 6329 -16120
rect 6283 -16388 6289 -16132
rect 6323 -16388 6329 -16132
rect 6283 -16400 6329 -16388
rect 6461 -16132 6507 -16120
rect 6461 -16388 6467 -16132
rect 6501 -16388 6507 -16132
rect 6461 -16400 6507 -16388
rect 6639 -16132 6685 -16120
rect 6639 -16388 6645 -16132
rect 6679 -16388 6685 -16132
rect 6639 -16400 6685 -16388
rect 6817 -16132 6863 -16120
rect 6817 -16388 6823 -16132
rect 6857 -16388 6863 -16132
rect 6817 -16400 6863 -16388
rect 6995 -16132 7041 -16120
rect 6995 -16388 7001 -16132
rect 7035 -16388 7041 -16132
rect 6995 -16400 7041 -16388
rect 7173 -16132 7219 -16120
rect 7173 -16388 7179 -16132
rect 7213 -16388 7219 -16132
rect 7173 -16400 7219 -16388
rect 7351 -16132 7397 -16120
rect 7351 -16388 7357 -16132
rect 7391 -16388 7397 -16132
rect 7351 -16400 7397 -16388
rect 7529 -16132 7575 -16120
rect 7529 -16388 7535 -16132
rect 7569 -16388 7575 -16132
rect 7529 -16400 7575 -16388
rect 7707 -16132 7753 -16120
rect 7707 -16388 7713 -16132
rect 7747 -16388 7753 -16132
rect 7707 -16400 7753 -16388
rect 7885 -16132 7931 -16120
rect 7885 -16388 7891 -16132
rect 7925 -16388 7931 -16132
rect 7885 -16400 7931 -16388
rect 8063 -16132 8109 -16120
rect 8063 -16388 8069 -16132
rect 8103 -16388 8109 -16132
rect 8063 -16400 8109 -16388
rect 8241 -16132 8287 -16120
rect 8241 -16388 8247 -16132
rect 8281 -16388 8287 -16132
rect 8241 -16400 8287 -16388
rect 8419 -16132 8465 -16120
rect 8419 -16388 8425 -16132
rect 8459 -16388 8465 -16132
rect 8419 -16400 8465 -16388
rect 8597 -16132 8643 -16120
rect 8597 -16388 8603 -16132
rect 8637 -16388 8643 -16132
rect 8597 -16400 8643 -16388
rect 8775 -16132 8821 -16120
rect 8775 -16388 8781 -16132
rect 8815 -16388 8821 -16132
rect 8775 -16400 8821 -16388
rect 8953 -16132 8999 -16120
rect 8953 -16388 8959 -16132
rect 8993 -16388 8999 -16132
rect 8953 -16400 8999 -16388
rect 9131 -16132 9177 -16120
rect 9131 -16388 9137 -16132
rect 9171 -16388 9177 -16132
rect 9131 -16400 9177 -16388
rect 9309 -16132 9355 -16120
rect 9309 -16388 9315 -16132
rect 9349 -16388 9355 -16132
rect 9309 -16400 9355 -16388
rect 9487 -16132 9533 -16120
rect 9487 -16388 9493 -16132
rect 9527 -16388 9533 -16132
rect 9487 -16400 9533 -16388
rect 9665 -16132 9711 -16120
rect 9665 -16388 9671 -16132
rect 9705 -16388 9711 -16132
rect 9665 -16400 9711 -16388
rect 9843 -16132 9889 -16120
rect 9843 -16388 9849 -16132
rect 9883 -16388 9889 -16132
rect 9843 -16400 9889 -16388
rect 10021 -16132 10067 -16120
rect 10021 -16388 10027 -16132
rect 10061 -16388 10067 -16132
rect 10021 -16400 10067 -16388
rect 10199 -16132 10245 -16120
rect 10199 -16388 10205 -16132
rect 10239 -16388 10245 -16132
rect 10199 -16400 10245 -16388
rect 10377 -16132 10423 -16120
rect 10377 -16388 10383 -16132
rect 10417 -16388 10423 -16132
rect 10377 -16400 10423 -16388
rect 10555 -16132 10601 -16120
rect 10555 -16388 10561 -16132
rect 10595 -16388 10601 -16132
rect 10555 -16400 10601 -16388
rect 10733 -16132 10779 -16120
rect 10733 -16388 10739 -16132
rect 10773 -16388 10779 -16132
rect 10733 -16400 10779 -16388
rect 10911 -16132 10957 -16120
rect 10911 -16388 10917 -16132
rect 10951 -16388 10957 -16132
rect 10911 -16400 10957 -16388
rect 11089 -16132 11135 -16120
rect 11089 -16388 11095 -16132
rect 11129 -16388 11135 -16132
rect 11089 -16400 11135 -16388
rect 11267 -16132 11313 -16120
rect 11267 -16388 11273 -16132
rect 11307 -16388 11313 -16132
rect 11267 -16400 11313 -16388
rect 11445 -16132 11491 -16120
rect 11445 -16388 11451 -16132
rect 11485 -16388 11491 -16132
rect 11445 -16400 11491 -16388
rect 11623 -16132 11669 -16120
rect 11623 -16388 11629 -16132
rect 11663 -16388 11669 -16132
rect 11623 -16400 11669 -16388
rect 11801 -16132 11847 -16120
rect 11801 -16388 11807 -16132
rect 11841 -16388 11847 -16132
rect 11801 -16400 11847 -16388
rect 11979 -16132 12025 -16120
rect 11979 -16388 11985 -16132
rect 12019 -16388 12025 -16132
rect 11979 -16400 12025 -16388
rect 12157 -16132 12203 -16120
rect 12157 -16388 12163 -16132
rect 12197 -16388 12203 -16132
rect 12157 -16400 12203 -16388
rect 12335 -16132 12381 -16120
rect 12335 -16388 12341 -16132
rect 12375 -16388 12381 -16132
rect 12335 -16400 12381 -16388
rect 12513 -16132 12559 -16120
rect 12513 -16388 12519 -16132
rect 12553 -16388 12559 -16132
rect 12513 -16400 12559 -16388
rect 12691 -16132 12737 -16120
rect 12691 -16388 12697 -16132
rect 12731 -16388 12737 -16132
rect 12691 -16400 12737 -16388
rect 5576 -16438 5610 -16400
rect 5645 -16438 5721 -16432
rect 5756 -16438 5790 -16400
rect 5576 -16472 5661 -16438
rect 5705 -16472 5790 -16438
rect 5823 -16438 5899 -16432
rect 5823 -16472 5839 -16438
rect 5883 -16472 5899 -16438
rect 5645 -16488 5721 -16472
rect 5823 -16488 5899 -16472
rect 6001 -16438 6077 -16432
rect 6001 -16472 6017 -16438
rect 6061 -16472 6077 -16438
rect 6001 -16488 6077 -16472
rect 6179 -16438 6255 -16432
rect 6179 -16472 6195 -16438
rect 6239 -16472 6255 -16438
rect 6179 -16488 6255 -16472
rect 6357 -16438 6433 -16432
rect 6357 -16472 6373 -16438
rect 6417 -16472 6433 -16438
rect 6357 -16488 6433 -16472
rect 6535 -16438 6611 -16432
rect 6535 -16472 6551 -16438
rect 6595 -16472 6611 -16438
rect 6535 -16488 6611 -16472
rect 6713 -16438 6789 -16432
rect 6713 -16472 6729 -16438
rect 6773 -16472 6789 -16438
rect 6713 -16488 6789 -16472
rect 6891 -16438 6967 -16432
rect 6891 -16472 6907 -16438
rect 6951 -16472 6967 -16438
rect 6891 -16488 6967 -16472
rect 7069 -16438 7145 -16432
rect 7178 -16438 7212 -16400
rect 7247 -16438 7323 -16432
rect 7069 -16472 7085 -16438
rect 7129 -16472 7263 -16438
rect 7307 -16472 7323 -16438
rect 7069 -16488 7145 -16472
rect 7247 -16488 7323 -16472
rect 6557 -16544 6591 -16488
rect 6735 -16544 6769 -16488
rect 6538 -16597 6548 -16544
rect 6601 -16597 6611 -16544
rect 6716 -16597 6726 -16544
rect 6779 -16597 6789 -16544
rect 6912 -16545 6946 -16488
rect 6893 -16598 6903 -16545
rect 6956 -16598 6966 -16545
rect 5389 -16720 5399 -16667
rect 5452 -16720 5462 -16667
rect 5021 -16835 5031 -16782
rect 5084 -16835 5094 -16782
rect 7357 -16890 7391 -16400
rect 7425 -16438 7501 -16432
rect 7425 -16472 7441 -16438
rect 7485 -16472 7501 -16438
rect 7425 -16488 7501 -16472
rect 7603 -16438 7679 -16432
rect 7603 -16472 7619 -16438
rect 7663 -16472 7679 -16438
rect 7603 -16488 7679 -16472
rect 7713 -16890 7747 -16400
rect 7781 -16438 7857 -16432
rect 7781 -16472 7797 -16438
rect 7841 -16472 7857 -16438
rect 7781 -16488 7857 -16472
rect 7959 -16438 8035 -16432
rect 7959 -16472 7975 -16438
rect 8019 -16472 8035 -16438
rect 7959 -16488 8035 -16472
rect 7980 -16545 8014 -16488
rect 7960 -16598 7970 -16545
rect 8023 -16598 8033 -16545
rect 8069 -16890 8103 -16400
rect 8137 -16438 8213 -16432
rect 8137 -16472 8153 -16438
rect 8197 -16472 8213 -16438
rect 8137 -16488 8213 -16472
rect 8315 -16438 8391 -16432
rect 8315 -16472 8331 -16438
rect 8375 -16472 8391 -16438
rect 8315 -16488 8391 -16472
rect 8158 -16544 8192 -16488
rect 8139 -16597 8149 -16544
rect 8202 -16597 8212 -16544
rect 8426 -16890 8460 -16400
rect 8493 -16438 8569 -16432
rect 8603 -16438 8637 -16400
rect 8671 -16438 8747 -16432
rect 8493 -16472 8509 -16438
rect 8553 -16472 8687 -16438
rect 8731 -16472 8747 -16438
rect 8493 -16488 8569 -16472
rect 8671 -16488 8747 -16472
rect 8781 -16666 8815 -16400
rect 8849 -16438 8925 -16432
rect 8849 -16472 8865 -16438
rect 8909 -16472 8925 -16438
rect 8849 -16488 8925 -16472
rect 8761 -16719 8771 -16666
rect 8824 -16719 8834 -16666
rect 8960 -16782 8994 -16400
rect 9027 -16438 9103 -16432
rect 9027 -16472 9043 -16438
rect 9087 -16472 9103 -16438
rect 9027 -16488 9103 -16472
rect 9138 -16666 9172 -16400
rect 9205 -16438 9281 -16432
rect 9205 -16472 9221 -16438
rect 9265 -16472 9281 -16438
rect 9205 -16488 9281 -16472
rect 9118 -16719 9128 -16666
rect 9181 -16719 9191 -16666
rect 9315 -16782 9349 -16400
rect 9383 -16438 9459 -16432
rect 9383 -16472 9399 -16438
rect 9443 -16472 9459 -16438
rect 9383 -16488 9459 -16472
rect 9493 -16666 9527 -16400
rect 9561 -16438 9637 -16432
rect 9672 -16438 9706 -16400
rect 9739 -16438 9815 -16432
rect 9561 -16472 9577 -16438
rect 9621 -16472 9755 -16438
rect 9799 -16472 9815 -16438
rect 9561 -16488 9637 -16472
rect 9474 -16719 9484 -16666
rect 9537 -16719 9547 -16666
rect 8940 -16835 8950 -16782
rect 9003 -16835 9013 -16782
rect 9295 -16835 9305 -16782
rect 9358 -16835 9368 -16782
rect 7337 -16943 7347 -16890
rect 7400 -16943 7410 -16890
rect 7694 -16943 7704 -16890
rect 7757 -16943 7767 -16890
rect 8050 -16943 8060 -16890
rect 8113 -16943 8123 -16890
rect 8406 -16943 8416 -16890
rect 8469 -16943 8479 -16890
rect 9672 -17251 9706 -16472
rect 9739 -16488 9815 -16472
rect 9848 -16666 9882 -16400
rect 9917 -16438 9993 -16432
rect 9917 -16472 9933 -16438
rect 9977 -16472 9993 -16438
rect 9917 -16488 9993 -16472
rect 9938 -16544 9972 -16488
rect 9919 -16597 9929 -16544
rect 9982 -16597 9992 -16544
rect 9828 -16719 9838 -16666
rect 9891 -16719 9901 -16666
rect 10028 -16781 10062 -16400
rect 10095 -16438 10171 -16432
rect 10095 -16472 10111 -16438
rect 10155 -16472 10171 -16438
rect 10095 -16488 10171 -16472
rect 10117 -16545 10151 -16488
rect 10097 -16598 10107 -16545
rect 10160 -16598 10170 -16545
rect 10205 -16665 10239 -16400
rect 10273 -16438 10349 -16432
rect 10273 -16472 10289 -16438
rect 10333 -16472 10349 -16438
rect 10273 -16488 10349 -16472
rect 10296 -16545 10330 -16488
rect 10277 -16598 10287 -16545
rect 10340 -16598 10350 -16545
rect 10185 -16718 10195 -16665
rect 10248 -16718 10258 -16665
rect 10383 -16781 10417 -16400
rect 10451 -16438 10527 -16432
rect 10451 -16472 10467 -16438
rect 10511 -16472 10527 -16438
rect 10451 -16488 10527 -16472
rect 10561 -16665 10595 -16400
rect 10629 -16438 10705 -16432
rect 10629 -16472 10645 -16438
rect 10689 -16472 10705 -16438
rect 10629 -16488 10705 -16472
rect 10540 -16718 10550 -16665
rect 10603 -16718 10613 -16665
rect 10739 -16779 10773 -16400
rect 10807 -16438 10883 -16432
rect 10807 -16472 10823 -16438
rect 10867 -16472 10883 -16438
rect 10807 -16488 10883 -16472
rect 10917 -16665 10951 -16400
rect 10985 -16437 11061 -16432
rect 11094 -16437 11128 -16400
rect 11163 -16437 11239 -16432
rect 10985 -16438 11239 -16437
rect 10985 -16472 11001 -16438
rect 11045 -16471 11179 -16438
rect 11045 -16472 11061 -16471
rect 10985 -16488 11061 -16472
rect 11163 -16472 11179 -16471
rect 11223 -16472 11239 -16438
rect 11163 -16488 11239 -16472
rect 10897 -16718 10907 -16665
rect 10960 -16718 10970 -16665
rect 10007 -16834 10017 -16781
rect 10070 -16834 10080 -16781
rect 10364 -16834 10374 -16781
rect 10427 -16834 10437 -16781
rect 10721 -16832 10731 -16779
rect 10784 -16832 10794 -16779
rect 11273 -16890 11307 -16400
rect 11341 -16438 11417 -16432
rect 11341 -16472 11357 -16438
rect 11401 -16472 11417 -16438
rect 11341 -16488 11417 -16472
rect 11519 -16438 11595 -16432
rect 11519 -16472 11535 -16438
rect 11579 -16472 11595 -16438
rect 11519 -16488 11595 -16472
rect 11362 -16545 11396 -16488
rect 11342 -16598 11352 -16545
rect 11405 -16598 11415 -16545
rect 11540 -16546 11574 -16488
rect 11520 -16599 11530 -16546
rect 11583 -16599 11593 -16546
rect 11630 -16890 11664 -16400
rect 11697 -16438 11773 -16432
rect 11697 -16472 11713 -16438
rect 11757 -16472 11773 -16438
rect 11697 -16488 11773 -16472
rect 11875 -16438 11951 -16432
rect 11875 -16472 11891 -16438
rect 11935 -16472 11951 -16438
rect 11875 -16488 11951 -16472
rect 11718 -16545 11752 -16488
rect 11699 -16598 11709 -16545
rect 11762 -16598 11772 -16545
rect 11985 -16889 12019 -16400
rect 12053 -16438 12129 -16432
rect 12053 -16472 12069 -16438
rect 12113 -16472 12129 -16438
rect 12053 -16488 12129 -16472
rect 12231 -16438 12307 -16432
rect 12231 -16472 12247 -16438
rect 12291 -16472 12307 -16438
rect 12231 -16488 12307 -16472
rect 12340 -16889 12374 -16400
rect 12409 -16438 12485 -16432
rect 12409 -16472 12425 -16438
rect 12469 -16472 12485 -16438
rect 12409 -16488 12485 -16472
rect 12520 -16440 12554 -16400
rect 12587 -16438 12663 -16432
rect 12587 -16440 12603 -16438
rect 12520 -16472 12603 -16440
rect 12647 -16440 12663 -16438
rect 12698 -16440 12732 -16400
rect 12647 -16472 12732 -16440
rect 12520 -16474 12732 -16472
rect 12587 -16488 12663 -16474
rect 11253 -16943 11263 -16890
rect 11316 -16943 11326 -16890
rect 11610 -16943 11620 -16890
rect 11673 -16943 11683 -16890
rect 11965 -16942 11975 -16889
rect 12028 -16942 12038 -16889
rect 12321 -16942 12331 -16889
rect 12384 -16942 12394 -16889
rect 13022 -17251 13075 -11726
rect -7605 -17459 13720 -17251
rect -7605 -17559 -7323 -17459
rect 13384 -17527 13720 -17459
rect 13384 -17559 13719 -17527
rect -7605 -17587 13719 -17559
<< via1 >>
rect -5867 -1963 -5814 -1910
rect -5689 -1963 -5636 -1910
rect -5510 -1963 -5457 -1910
rect -5333 -1963 -5280 -1910
rect -5155 -1963 -5102 -1910
rect -4976 -1963 -4923 -1910
rect -4799 -1963 -4746 -1910
rect -4621 -1963 -4568 -1910
rect -4443 -1963 -4390 -1910
rect -4265 -1963 -4212 -1910
rect -4086 -1963 -4033 -1910
rect -3909 -1963 -3856 -1910
rect -1109 -1963 -1056 -1910
rect -6498 -2582 -6445 -2529
rect -6625 -3454 -6572 -3401
rect -6044 -2833 -5991 -2780
rect -5777 -2583 -5724 -2530
rect -5866 -2833 -5813 -2780
rect -5421 -2721 -5368 -2668
rect -5066 -2583 -5013 -2530
rect -4710 -2721 -4657 -2668
rect -4354 -2583 -4301 -2530
rect -3998 -2721 -3945 -2668
rect -3908 -2833 -3855 -2780
rect -1109 -2478 -1056 -2425
rect -752 -2478 -699 -2425
rect -2624 -2611 -2571 -2558
rect -1285 -2611 -1232 -2558
rect -3298 -2721 -3245 -2668
rect -3731 -2833 -3678 -2780
rect -6134 -3454 -6081 -3401
rect -6498 -3693 -6445 -3640
rect -5777 -3569 -5724 -3516
rect -5422 -3693 -5369 -3640
rect -5066 -3454 -5013 -3401
rect -4710 -3454 -4657 -3401
rect -4353 -3693 -4300 -3640
rect -3998 -3569 -3945 -3516
rect -3642 -3454 -3589 -3401
rect -3131 -3454 -3078 -3401
rect -3298 -3569 -3245 -3516
rect -6498 -4324 -6445 -4271
rect -6134 -4443 -6081 -4390
rect -5778 -4324 -5725 -4271
rect -5422 -4559 -5369 -4506
rect -5066 -4443 -5013 -4390
rect -4709 -4443 -4656 -4390
rect -4353 -4559 -4300 -4506
rect -3998 -4324 -3945 -4271
rect -3642 -4443 -3589 -4390
rect -3298 -4559 -3245 -4506
rect -6498 -5194 -6445 -5141
rect -6625 -5375 -6572 -5322
rect -6134 -5285 -6081 -5232
rect -5777 -5468 -5724 -5415
rect -5422 -5194 -5369 -5141
rect -5066 -5286 -5013 -5233
rect -4710 -5375 -4657 -5322
rect -4353 -5194 -4300 -5141
rect -3997 -5468 -3944 -5415
rect -3642 -5372 -3589 -5319
rect -3130 -5286 -3077 -5233
rect -1197 -2718 -1144 -2665
rect -930 -2611 -877 -2558
rect -1019 -2718 -966 -2665
rect -841 -2718 -788 -2665
rect -129 -2718 -76 -2665
rect 50 -2718 103 -2665
rect 227 -2718 280 -2665
rect 1919 -2479 1972 -2426
rect 2275 -2479 2328 -2426
rect 940 -2718 993 -2665
rect 1117 -2718 1170 -2665
rect 1295 -2718 1348 -2665
rect 2097 -2607 2150 -2554
rect 2007 -2718 2060 -2665
rect 2186 -2718 2239 -2665
rect 3193 -2480 3246 -2427
rect 2453 -2607 2506 -2554
rect 2363 -2718 2416 -2665
rect -1645 -3510 -1584 -3449
rect -2004 -4465 -1951 -4412
rect -2624 -5377 -2571 -5324
rect -3298 -5469 -3245 -5416
rect -5956 -6069 -5903 -6016
rect -5601 -6069 -5548 -6016
rect -5778 -6184 -5725 -6131
rect -5244 -6069 -5191 -6016
rect -5065 -6184 -5012 -6131
rect -6498 -6301 -6445 -6248
rect -5421 -6301 -5368 -6248
rect -4888 -6069 -4835 -6016
rect -4710 -6301 -4657 -6248
rect -4532 -6069 -4479 -6016
rect -4175 -6069 -4122 -6016
rect -4354 -6184 -4301 -6131
rect -3820 -6069 -3767 -6016
rect -2624 -6060 -2571 -6007
rect -3298 -6184 -3245 -6131
rect -3998 -6300 -3945 -6247
rect -4786 -6431 -4733 -6378
rect -1876 -5285 -1823 -5232
rect -1286 -3624 -1233 -3571
rect -1108 -3509 -1055 -3456
rect -929 -3624 -876 -3571
rect -484 -3354 -431 -3301
rect -750 -3509 -697 -3456
rect -396 -3509 -343 -3456
rect -573 -3624 -520 -3571
rect -217 -3624 -164 -3571
rect 583 -3354 636 -3301
rect -39 -3509 14 -3456
rect 317 -3509 370 -3456
rect 850 -3509 903 -3456
rect 1206 -3509 1259 -3456
rect 1654 -3354 1707 -3301
rect 1562 -3509 1615 -3456
rect 1919 -3509 1972 -3456
rect 1384 -3617 1437 -3564
rect 1741 -3617 1794 -3564
rect 2097 -3617 2150 -3564
rect 2275 -3509 2328 -3456
rect 2451 -3617 2504 -3564
rect -841 -4245 -788 -4192
rect -662 -4245 -609 -4192
rect -483 -4245 -430 -4192
rect -306 -4245 -253 -4192
rect 407 -4245 460 -4192
rect 317 -4357 370 -4304
rect 583 -4245 636 -4192
rect 495 -4465 548 -4412
rect 761 -4245 814 -4192
rect 673 -4357 726 -4304
rect 850 -4465 903 -4412
rect 1474 -4245 1527 -4192
rect 1652 -4245 1705 -4192
rect 1830 -4245 1883 -4192
rect 2008 -4245 2061 -4192
rect 2538 -4327 2599 -4266
rect 2746 -4507 2807 -4446
rect -1287 -5150 -1234 -5097
rect -1646 -5339 -1585 -5278
rect -1105 -5266 -1052 -5213
rect -929 -5150 -876 -5097
rect -572 -5150 -519 -5097
rect -218 -5150 -165 -5097
rect -751 -5266 -698 -5213
rect -396 -5266 -343 -5213
rect -41 -5266 12 -5213
rect 316 -5266 369 -5213
rect -128 -5433 -75 -5380
rect 50 -5433 103 -5380
rect 228 -5433 281 -5380
rect 850 -5266 903 -5213
rect 1207 -5266 1260 -5213
rect 940 -5434 993 -5381
rect 1119 -5433 1172 -5380
rect 1385 -5146 1438 -5093
rect 1296 -5433 1349 -5380
rect 1740 -5146 1793 -5093
rect 1563 -5266 1616 -5213
rect 1917 -5266 1970 -5213
rect 2096 -5146 2149 -5093
rect 2274 -5266 2327 -5213
rect 2453 -5146 2506 -5093
rect -1876 -6417 -1823 -6364
rect -1282 -6417 -1229 -6364
rect -928 -6417 -876 -6365
rect -1110 -6532 -1057 -6479
rect -752 -6532 -699 -6479
rect 227 -6303 280 -6250
rect 942 -6303 995 -6250
rect 2096 -6060 2149 -6007
rect 2452 -6060 2505 -6007
rect 1918 -6177 1971 -6124
rect 2275 -6177 2328 -6124
rect 3194 -4857 3246 -4805
rect 4771 -4857 4823 -4805
rect 2879 -6417 2931 -6365
rect 5037 -5059 5090 -5006
rect 4905 -5265 4958 -5212
rect -753 -6651 -700 -6598
rect 4772 -6650 4825 -6597
rect -2003 -6767 -1950 -6714
rect 4770 -6944 4823 -6891
rect 4906 -6942 4959 -6889
rect 5038 -6940 5091 -6887
rect -3873 -7743 -3821 -7691
rect -3731 -7837 -3679 -7785
rect -3541 -7840 -3489 -7788
rect -5502 -12324 -5449 -12271
rect -6077 -12565 -6024 -12512
rect -5626 -12565 -5573 -12512
rect -6223 -13115 -6170 -13062
rect -6426 -13905 -6373 -13852
rect -5000 -12325 -4947 -12272
rect -4502 -12324 -4449 -12271
rect -5376 -12441 -5323 -12388
rect -5127 -12441 -5074 -12388
rect -4877 -12565 -4824 -12512
rect -4627 -12565 -4574 -12512
rect -4377 -12441 -4324 -12388
rect -3928 -12442 -3875 -12389
rect -5751 -13115 -5698 -13062
rect -5251 -13242 -5198 -13189
rect -4752 -13115 -4699 -13062
rect -4251 -13242 -4198 -13189
rect -6077 -13798 -6024 -13745
rect -5376 -13798 -5323 -13745
rect -5626 -13905 -5573 -13852
rect -5730 -14010 -5677 -13957
rect -5126 -13798 -5073 -13745
rect -4877 -13905 -4824 -13852
rect -4376 -13798 -4323 -13745
rect -4627 -13905 -4574 -13852
rect -4752 -14010 -4699 -13957
rect -3788 -13242 -3735 -13189
rect -3928 -13905 -3875 -13852
rect -3788 -14010 -3735 -13957
rect -6223 -14108 -6170 -14055
rect -5250 -14108 -5197 -14055
rect -4250 -14108 -4197 -14055
rect -6159 -14848 -6106 -14795
rect -5860 -14848 -5807 -14795
rect -5504 -14954 -5451 -14901
rect -5147 -14848 -5094 -14795
rect -4791 -14954 -4738 -14901
rect -4436 -14848 -4383 -14795
rect 4771 -7907 4824 -7854
rect 4906 -7905 4959 -7852
rect 5037 -7903 5090 -7850
rect -3382 -7986 -3329 -7933
rect -1382 -7975 -1329 -7922
rect -3542 -13242 -3489 -13189
rect -1203 -7976 -1150 -7923
rect -1025 -7975 -972 -7922
rect -848 -7975 -795 -7922
rect -670 -7975 -617 -7922
rect -490 -7975 -437 -7922
rect 755 -7975 808 -7922
rect 932 -7975 985 -7922
rect 1112 -7975 1165 -7922
rect 1289 -7976 1342 -7923
rect 1467 -7975 1520 -7922
rect 1644 -7975 1697 -7922
rect 2890 -7975 2943 -7922
rect 3069 -7975 3122 -7922
rect 3247 -7975 3300 -7922
rect 3424 -7975 3477 -7922
rect 3603 -7976 3656 -7923
rect 3778 -7975 3831 -7922
rect 4208 -7976 4261 -7923
rect -1916 -8587 -1863 -8534
rect -1739 -8587 -1686 -8534
rect -1826 -8706 -1773 -8653
rect -2447 -8820 -2394 -8767
rect -2005 -8820 -1952 -8767
rect -1558 -8587 -1505 -8534
rect -1382 -8587 -1329 -8534
rect -1470 -8706 -1417 -8653
rect -1648 -8820 -1595 -8767
rect -1203 -8587 -1150 -8534
rect -1293 -8820 -1240 -8767
rect -1026 -8587 -973 -8534
rect -1115 -8706 -1062 -8653
rect -848 -8587 -795 -8534
rect -936 -8820 -883 -8767
rect -670 -8587 -617 -8534
rect -758 -8706 -705 -8653
rect -491 -8587 -438 -8534
rect -580 -8819 -527 -8766
rect -314 -8587 -261 -8534
rect -402 -8706 -349 -8653
rect -136 -8587 -83 -8534
rect 42 -8587 95 -8534
rect -47 -8706 6 -8653
rect -225 -8820 -172 -8767
rect 221 -8587 274 -8534
rect 398 -8587 451 -8534
rect 310 -8706 363 -8653
rect 132 -8821 185 -8768
rect 577 -8587 630 -8534
rect 754 -8587 807 -8534
rect 666 -8706 719 -8653
rect 489 -8819 542 -8766
rect 932 -8587 985 -8534
rect 843 -8819 896 -8766
rect 1111 -8587 1164 -8534
rect 1022 -8706 1075 -8653
rect 1289 -8587 1342 -8534
rect 1201 -8820 1254 -8767
rect 1466 -8587 1519 -8534
rect 1377 -8706 1430 -8653
rect 1644 -8587 1697 -8534
rect 1556 -8820 1609 -8767
rect 1822 -8587 1875 -8534
rect 1733 -8706 1786 -8653
rect 2000 -8587 2053 -8534
rect 2178 -8587 2231 -8534
rect 2090 -8706 2143 -8653
rect 1911 -8820 1964 -8767
rect 2357 -8587 2410 -8534
rect 2534 -8587 2587 -8534
rect 2446 -8706 2499 -8653
rect 2267 -8820 2320 -8767
rect 2712 -8587 2765 -8534
rect 2890 -8587 2943 -8534
rect 2802 -8706 2855 -8653
rect 2624 -8820 2677 -8767
rect 3068 -8587 3121 -8534
rect 2980 -8820 3033 -8767
rect 3246 -8587 3299 -8534
rect 3158 -8706 3211 -8653
rect 3424 -8587 3477 -8534
rect 3336 -8820 3389 -8767
rect 3602 -8587 3655 -8534
rect 3513 -8706 3566 -8653
rect 3781 -8587 3834 -8534
rect 3692 -8820 3745 -8767
rect 3869 -8706 3922 -8653
rect -2315 -9978 -2262 -9925
rect -2447 -12325 -2394 -12272
rect -3382 -14108 -3329 -14055
rect -3936 -14954 -3883 -14901
rect -6159 -15535 -6106 -15482
rect -5860 -15641 -5807 -15588
rect -5504 -15534 -5451 -15481
rect -5148 -15642 -5095 -15589
rect -4792 -15534 -4739 -15481
rect -4435 -15641 -4383 -15589
rect -3935 -15641 -3883 -15589
rect -6159 -16246 -6106 -16193
rect -5860 -16347 -5807 -16294
rect -5504 -16246 -5451 -16193
rect -5148 -16347 -5095 -16294
rect -4792 -16246 -4739 -16193
rect -4436 -16347 -4383 -16294
rect -1916 -9599 -1863 -9546
rect -1916 -9978 -1863 -9925
rect -1738 -9599 -1685 -9546
rect -1738 -9979 -1685 -9926
rect -1558 -9599 -1505 -9546
rect -1560 -9978 -1507 -9925
rect -1382 -9977 -1329 -9924
rect -312 -9599 -259 -9546
rect -314 -9978 -261 -9925
rect -136 -9598 -83 -9545
rect -136 -9979 -83 -9926
rect 42 -9599 95 -9546
rect 43 -9978 96 -9925
rect 222 -9598 275 -9545
rect 220 -9978 273 -9925
rect 399 -9599 452 -9546
rect 398 -9978 451 -9925
rect 577 -9599 630 -9546
rect 576 -9978 629 -9925
rect 2178 -9600 2231 -9547
rect 2357 -9599 2410 -9546
rect 2356 -9978 2409 -9925
rect 2534 -9599 2587 -9546
rect 2534 -9978 2587 -9925
rect 2713 -9599 2766 -9546
rect 2712 -9979 2765 -9926
rect 2891 -9978 2944 -9925
rect 3069 -9978 3122 -9925
rect 3246 -9978 3299 -9925
rect 4771 -9367 4824 -9314
rect 4208 -9599 4261 -9546
rect -1827 -10961 -1774 -10908
rect -1470 -10961 -1417 -10908
rect -1114 -10961 -1061 -10908
rect -758 -10961 -705 -10908
rect -402 -10961 -349 -10908
rect -46 -10961 7 -10908
rect 309 -10961 362 -10908
rect 665 -10961 718 -10908
rect 931 -10961 984 -10908
rect 1199 -10961 1252 -10908
rect 1556 -10961 1609 -10908
rect 1913 -10961 1966 -10908
rect 2268 -10961 2321 -10908
rect 2623 -10961 2676 -10908
rect 2980 -10961 3033 -10908
rect 3335 -10961 3388 -10908
rect 3692 -10961 3745 -10908
rect -2004 -11690 -1951 -11637
rect -1915 -11972 -1862 -11919
rect -1649 -11581 -1596 -11528
rect -1738 -11972 -1685 -11919
rect -1559 -11972 -1506 -11919
rect -1293 -11581 -1240 -11528
rect -1381 -11972 -1328 -11919
rect -1203 -11972 -1150 -11919
rect -937 -11581 -884 -11528
rect -1025 -11972 -972 -11919
rect -848 -11972 -795 -11919
rect -580 -11690 -527 -11637
rect -670 -11972 -617 -11919
rect -492 -11972 -439 -11919
rect -224 -11810 -171 -11757
rect -314 -11972 -261 -11919
rect -136 -11972 -83 -11919
rect 131 -11810 184 -11757
rect 42 -11972 95 -11919
rect 220 -11972 273 -11919
rect 487 -11810 540 -11757
rect 399 -11972 452 -11919
rect 577 -11972 630 -11919
rect 1377 -11581 1430 -11528
rect 1288 -11972 1341 -11919
rect 1468 -11972 1521 -11919
rect 1733 -11581 1786 -11528
rect 1644 -11973 1697 -11920
rect 1823 -11972 1876 -11919
rect 2089 -11581 2142 -11528
rect 2000 -11972 2053 -11919
rect 2178 -11972 2231 -11919
rect 2446 -11690 2499 -11637
rect 2357 -11972 2410 -11919
rect 2534 -11972 2587 -11919
rect 2800 -11810 2853 -11757
rect 2713 -11972 2766 -11919
rect 2890 -11972 2943 -11919
rect 3157 -11810 3210 -11757
rect 3068 -11972 3121 -11919
rect 3247 -11972 3300 -11919
rect 3513 -11810 3566 -11757
rect 3425 -11972 3478 -11919
rect 3603 -11972 3656 -11919
rect 3871 -11691 3924 -11638
rect 3781 -11972 3834 -11919
rect -2005 -12595 -1952 -12542
rect -1649 -12595 -1596 -12542
rect -1294 -12707 -1241 -12654
rect -937 -12836 -884 -12783
rect -582 -12706 -529 -12653
rect -224 -12836 -171 -12783
rect 130 -12706 183 -12653
rect 486 -12837 539 -12784
rect 1378 -12836 1431 -12783
rect 1735 -12707 1788 -12654
rect 2088 -12835 2141 -12782
rect 2445 -12706 2498 -12653
rect 2801 -12835 2854 -12782
rect 3158 -12705 3211 -12652
rect 3514 -12595 3567 -12542
rect 3871 -12595 3924 -12542
rect -2004 -13598 -1951 -13545
rect -1648 -13725 -1595 -13672
rect -581 -13598 -528 -13545
rect -1291 -13725 -1238 -13672
rect -937 -13725 -884 -13672
rect -225 -13847 -172 -13794
rect 133 -13847 186 -13794
rect 487 -13848 540 -13795
rect 1379 -13725 1432 -13672
rect 1732 -13725 1785 -13672
rect 2091 -13725 2144 -13672
rect 2446 -13598 2499 -13545
rect 2802 -13847 2855 -13794
rect 3157 -13848 3210 -13795
rect 3870 -13598 3923 -13545
rect 3512 -13847 3565 -13794
rect -2315 -14596 -2262 -14543
rect -1381 -14596 -1328 -14543
rect -1204 -14596 -1151 -14543
rect -1026 -14596 -973 -14543
rect -848 -14596 -795 -14543
rect -847 -14979 -794 -14926
rect -669 -14596 -616 -14543
rect -669 -14979 -616 -14926
rect -491 -14596 -438 -14543
rect -491 -14979 -438 -14926
rect -314 -14980 -261 -14927
rect -137 -14979 -84 -14926
rect 43 -14979 96 -14926
rect 1288 -14596 1341 -14543
rect 1289 -14980 1342 -14927
rect 1466 -14596 1519 -14543
rect 1467 -14979 1520 -14926
rect 1644 -14596 1697 -14543
rect 1644 -14979 1697 -14926
rect 1823 -14595 1876 -14542
rect 1822 -14979 1875 -14926
rect 2000 -14596 2053 -14543
rect 1999 -14979 2052 -14926
rect 2178 -14596 2231 -14543
rect 2180 -14979 2233 -14926
rect 3246 -14597 3299 -14544
rect 3424 -14596 3477 -14543
rect 3425 -14979 3478 -14926
rect 3602 -14596 3655 -14543
rect 3603 -14979 3656 -14926
rect 3781 -14596 3834 -14543
rect 3780 -14979 3833 -14926
rect 5184 -7908 5237 -7855
rect 5337 -7903 5390 -7850
rect 5185 -8687 5237 -8635
rect 11054 -8769 11107 -8716
rect 11345 -8769 11398 -8716
rect 11638 -8769 11691 -8716
rect 11932 -8769 11985 -8716
rect 12222 -8769 12275 -8716
rect 6769 -9367 6822 -9314
rect 6679 -9598 6732 -9545
rect 6947 -9368 7000 -9315
rect 7126 -9368 7179 -9315
rect 7303 -9366 7356 -9313
rect 7482 -9366 7535 -9313
rect 7659 -9368 7712 -9315
rect 7837 -9367 7890 -9314
rect 8015 -9368 8068 -9315
rect 8194 -9367 8247 -9314
rect 8371 -9367 8424 -9314
rect 8549 -9367 8602 -9314
rect 8727 -9368 8780 -9315
rect 8906 -9367 8959 -9314
rect 11144 -9427 11197 -9374
rect 11436 -9428 11489 -9375
rect 11728 -9428 11781 -9375
rect 12020 -9429 12073 -9376
rect 12312 -9428 12365 -9375
rect 5337 -9978 5390 -9925
rect 6680 -10366 6733 -10313
rect 6858 -10520 6911 -10467
rect 7214 -10519 7267 -10466
rect 7571 -10519 7624 -10466
rect 7927 -10519 7980 -10466
rect 8283 -10520 8336 -10467
rect 8638 -10519 8691 -10466
rect 9171 -10367 9224 -10314
rect 8995 -10520 9048 -10467
rect 7037 -11419 7090 -11366
rect 7393 -11419 7446 -11366
rect 7748 -11420 7801 -11367
rect 8103 -11419 8156 -11366
rect 8461 -11419 8514 -11366
rect 8817 -11419 8870 -11366
rect 11053 -11727 11106 -11674
rect 11347 -11728 11400 -11675
rect 11638 -11727 11691 -11674
rect 11931 -11727 11984 -11674
rect 12223 -11727 12276 -11674
rect 13022 -11726 13075 -11673
rect 5037 -13349 5090 -13296
rect 5534 -13349 5587 -13296
rect 5031 -13486 5084 -13433
rect 4905 -14598 4958 -14545
rect 4239 -14979 4292 -14926
rect -2447 -15874 -2394 -15821
rect -2005 -15875 -1952 -15822
rect -1915 -15986 -1862 -15933
rect -1649 -15875 -1596 -15822
rect -1738 -15986 -1685 -15933
rect -1560 -15986 -1507 -15933
rect -1293 -15875 -1240 -15822
rect -1382 -15986 -1329 -15933
rect -1204 -15986 -1151 -15933
rect -937 -15875 -884 -15822
rect -1025 -15986 -972 -15933
rect -847 -15986 -794 -15933
rect -581 -15875 -528 -15822
rect -670 -15986 -617 -15933
rect -491 -15986 -438 -15933
rect -225 -15875 -172 -15822
rect -313 -15986 -260 -15933
rect -136 -15986 -83 -15933
rect 132 -15874 185 -15821
rect 43 -15986 96 -15933
rect 221 -15986 274 -15933
rect 487 -15875 540 -15822
rect 398 -15986 451 -15933
rect 575 -15986 628 -15933
rect 843 -15875 896 -15822
rect 755 -15986 808 -15933
rect 931 -15986 984 -15933
rect 1201 -15875 1254 -15822
rect 1110 -15986 1163 -15933
rect 1289 -15986 1342 -15933
rect 1555 -15875 1608 -15822
rect 1466 -15986 1519 -15933
rect 1643 -15986 1696 -15933
rect 1910 -15875 1963 -15822
rect 1822 -15986 1875 -15933
rect 2000 -15986 2053 -15933
rect 2267 -15875 2320 -15822
rect 2179 -15986 2232 -15933
rect 2356 -15986 2409 -15933
rect 2624 -15875 2677 -15822
rect 2534 -15986 2587 -15933
rect 2712 -15986 2765 -15933
rect 2979 -15875 3032 -15822
rect 2891 -15986 2944 -15933
rect 3068 -15986 3121 -15933
rect 3335 -15875 3388 -15822
rect 3247 -15986 3300 -15933
rect 3424 -15986 3477 -15933
rect 3692 -15875 3745 -15822
rect 3603 -15986 3656 -15933
rect 3780 -15986 3833 -15933
rect 4238 -15592 4291 -15539
rect 5400 -13598 5453 -13545
rect 5142 -13847 5195 -13794
rect 5143 -14711 5196 -14658
rect -3935 -16347 -3883 -16295
rect -5682 -16939 -5629 -16886
rect -6159 -17060 -6106 -17007
rect -5859 -17060 -5806 -17007
rect -5326 -16939 -5273 -16886
rect -4970 -16939 -4917 -16886
rect -5148 -17060 -5095 -17007
rect -5504 -17171 -5451 -17118
rect -4614 -16939 -4561 -16886
rect -4258 -16939 -4205 -16886
rect -4437 -17060 -4384 -17007
rect -1917 -16595 -1864 -16542
rect -1738 -16595 -1685 -16542
rect -1561 -16594 -1508 -16541
rect -1827 -16718 -1774 -16665
rect -1381 -16596 -1328 -16543
rect -1204 -16595 -1151 -16542
rect -1026 -16595 -973 -16542
rect -1471 -16719 -1418 -16666
rect -1114 -16718 -1061 -16665
rect -759 -16717 -706 -16664
rect 220 -16595 273 -16542
rect -403 -16718 -350 -16665
rect -47 -16718 6 -16665
rect 397 -16595 450 -16542
rect 576 -16595 629 -16542
rect 755 -16595 808 -16542
rect 933 -16595 986 -16542
rect 1111 -16595 1164 -16542
rect 2356 -16595 2409 -16542
rect 309 -16719 362 -16666
rect 665 -16718 718 -16665
rect 845 -16718 898 -16665
rect 1021 -16718 1074 -16665
rect 1377 -16718 1430 -16665
rect 1735 -16718 1788 -16665
rect 2090 -16717 2143 -16664
rect 2534 -16595 2587 -16542
rect 2713 -16594 2766 -16541
rect 2891 -16595 2944 -16542
rect 3070 -16595 3123 -16542
rect 3249 -16595 3302 -16542
rect 2445 -16718 2498 -16665
rect 2801 -16718 2854 -16665
rect 3157 -16717 3210 -16664
rect 5031 -15593 5084 -15540
rect 4238 -16595 4291 -16542
rect -4792 -17171 -4739 -17118
rect -3935 -17170 -3883 -17118
rect 3514 -16719 3567 -16666
rect 3868 -16718 3921 -16665
rect 5534 -13725 5587 -13672
rect 8950 -13486 9003 -13433
rect 9305 -13486 9358 -13433
rect 8772 -13609 8825 -13556
rect 7526 -13725 7579 -13672
rect 7348 -13849 7401 -13796
rect 5833 -13975 5886 -13922
rect 6013 -13975 6066 -13922
rect 6190 -13976 6243 -13923
rect 6369 -13975 6422 -13922
rect 6547 -13976 6600 -13923
rect 6725 -13975 6778 -13922
rect 6902 -13975 6955 -13922
rect 7437 -13975 7490 -13922
rect 7882 -13726 7935 -13673
rect 8238 -13724 8291 -13671
rect 7704 -13848 7757 -13795
rect 7615 -13975 7668 -13922
rect 7793 -13976 7846 -13923
rect 8061 -13849 8114 -13796
rect 7970 -13975 8023 -13922
rect 8148 -13975 8201 -13922
rect 8415 -13849 8468 -13796
rect 8326 -13975 8379 -13922
rect 8861 -13975 8914 -13922
rect 9127 -13609 9180 -13556
rect 9038 -13975 9091 -13922
rect 9217 -13975 9270 -13922
rect 9483 -13609 9536 -13556
rect 9394 -13975 9447 -13922
rect 11442 -13725 11495 -13672
rect 11798 -13725 11851 -13672
rect 11264 -13849 11317 -13796
rect 9929 -13976 9982 -13923
rect 10108 -13975 10161 -13922
rect 10284 -13976 10337 -13923
rect 10462 -13976 10515 -13923
rect 10640 -13975 10693 -13922
rect 10819 -13976 10872 -13923
rect 11353 -13975 11406 -13922
rect 11620 -13850 11673 -13797
rect 11530 -13975 11583 -13922
rect 11709 -13975 11762 -13922
rect 12152 -13726 12205 -13673
rect 12509 -13725 12562 -13672
rect 11977 -13849 12030 -13796
rect 11886 -13976 11939 -13923
rect 12064 -13975 12117 -13922
rect 12334 -13849 12387 -13796
rect 12242 -13976 12295 -13923
rect 12420 -13975 12473 -13922
rect 5746 -14598 5799 -14545
rect 5924 -14711 5977 -14658
rect 6101 -14598 6154 -14545
rect 6279 -14711 6332 -14658
rect 6459 -14598 6512 -14545
rect 6813 -14598 6866 -14545
rect 6636 -14711 6689 -14658
rect 6991 -14711 7044 -14658
rect 6993 -14877 7046 -14824
rect 7347 -14877 7400 -14824
rect 7080 -14976 7133 -14923
rect 7260 -14977 7313 -14924
rect 7439 -14976 7492 -14923
rect 7704 -14878 7757 -14825
rect 8236 -14598 8289 -14545
rect 8060 -14874 8113 -14821
rect 8417 -14710 8470 -14657
rect 8327 -14976 8380 -14923
rect 8595 -14598 8648 -14545
rect 8504 -14859 8557 -14806
rect 8505 -14977 8558 -14924
rect 8772 -14711 8825 -14658
rect 8683 -14977 8736 -14924
rect 8950 -14599 9003 -14546
rect 9127 -14712 9180 -14659
rect 9304 -14598 9357 -14545
rect 9661 -14598 9714 -14545
rect 9483 -14711 9536 -14658
rect 9572 -14976 9625 -14923
rect 9837 -14712 9890 -14659
rect 9753 -14859 9806 -14806
rect 9750 -14976 9803 -14923
rect 10016 -14598 10069 -14545
rect 9929 -14976 9982 -14923
rect 10373 -14599 10426 -14546
rect 10196 -14711 10249 -14658
rect 10195 -14875 10248 -14822
rect 10550 -14711 10603 -14658
rect 10552 -14868 10605 -14815
rect 10729 -14598 10782 -14545
rect 10908 -14711 10961 -14658
rect 11087 -14711 11140 -14658
rect 10908 -14866 10961 -14813
rect 11440 -14709 11493 -14656
rect 10819 -14976 10872 -14923
rect 11264 -14868 11317 -14815
rect 10996 -14976 11049 -14923
rect 11175 -14976 11228 -14923
rect 5745 -15592 5798 -15539
rect 5400 -15706 5453 -15653
rect 5747 -15803 5800 -15750
rect 5923 -15705 5976 -15652
rect 5921 -16001 5974 -15948
rect 6101 -15592 6154 -15539
rect 6101 -15802 6154 -15749
rect 6279 -15705 6332 -15652
rect 6279 -16001 6332 -15948
rect 6458 -15592 6511 -15539
rect 6456 -15803 6509 -15750
rect 6635 -15705 6688 -15652
rect 6713 -15804 6766 -15751
rect 6634 -16001 6687 -15948
rect 6813 -15904 6866 -15851
rect 7169 -15803 7222 -15750
rect 7169 -15905 7222 -15852
rect 6994 -16004 7047 -15951
rect 7526 -15802 7579 -15749
rect 7526 -16006 7579 -15953
rect 7882 -15802 7935 -15749
rect 8060 -15904 8113 -15851
rect 7881 -16005 7934 -15952
rect 8237 -16005 8290 -15952
rect 8593 -15905 8646 -15852
rect 9663 -15905 9716 -15852
rect 10373 -15804 10426 -15751
rect 10194 -15905 10247 -15852
rect 10730 -15803 10783 -15750
rect 11086 -15803 11139 -15750
rect 11619 -15705 11672 -15652
rect 11084 -15905 11137 -15852
rect 11440 -15894 11493 -15841
rect 11441 -16005 11494 -15952
rect 11798 -15593 11851 -15540
rect 11797 -16005 11850 -15952
rect 11975 -15705 12028 -15652
rect 12155 -15592 12208 -15539
rect 12154 -16005 12207 -15952
rect 12332 -15705 12385 -15652
rect 12511 -15592 12564 -15539
rect 12511 -16005 12564 -15952
rect 6548 -16597 6601 -16544
rect 6726 -16597 6779 -16544
rect 6903 -16598 6956 -16545
rect 5399 -16720 5452 -16667
rect 5031 -16835 5084 -16782
rect 7970 -16598 8023 -16545
rect 8149 -16597 8202 -16544
rect 8771 -16719 8824 -16666
rect 9128 -16719 9181 -16666
rect 9484 -16719 9537 -16666
rect 8950 -16835 9003 -16782
rect 9305 -16835 9358 -16782
rect 7347 -16943 7400 -16890
rect 7704 -16943 7757 -16890
rect 8060 -16943 8113 -16890
rect 8416 -16943 8469 -16890
rect 9929 -16597 9982 -16544
rect 9838 -16719 9891 -16666
rect 10107 -16598 10160 -16545
rect 10287 -16598 10340 -16545
rect 10195 -16718 10248 -16665
rect 10550 -16718 10603 -16665
rect 10907 -16718 10960 -16665
rect 10017 -16834 10070 -16781
rect 10374 -16834 10427 -16781
rect 10731 -16832 10784 -16779
rect 11352 -16598 11405 -16545
rect 11530 -16599 11583 -16546
rect 11709 -16598 11762 -16545
rect 11263 -16943 11316 -16890
rect 11620 -16943 11673 -16890
rect 11975 -16942 12028 -16889
rect 12331 -16942 12384 -16889
<< metal2 >>
rect -5867 -1910 -5814 -1900
rect -5689 -1910 -5636 -1900
rect -5510 -1910 -5457 -1900
rect -5333 -1910 -5280 -1900
rect -5155 -1910 -5102 -1900
rect -4976 -1910 -4923 -1900
rect -4799 -1910 -4746 -1900
rect -4621 -1910 -4568 -1900
rect -4443 -1910 -4390 -1900
rect -4265 -1910 -4212 -1900
rect -4086 -1910 -4033 -1900
rect -3909 -1910 -3856 -1900
rect -1109 -1910 -1056 -1900
rect -5814 -1963 -5689 -1910
rect -5636 -1963 -5510 -1910
rect -5457 -1963 -5333 -1910
rect -5280 -1963 -5155 -1910
rect -5102 -1963 -4976 -1910
rect -4923 -1963 -4799 -1910
rect -4746 -1963 -4621 -1910
rect -4568 -1963 -4443 -1910
rect -4390 -1963 -4265 -1910
rect -4212 -1963 -4086 -1910
rect -4033 -1963 -3909 -1910
rect -3856 -1963 -1109 -1910
rect -5867 -1973 -5814 -1963
rect -5689 -1973 -5636 -1963
rect -5510 -1973 -5457 -1963
rect -5333 -1973 -5280 -1963
rect -5155 -1973 -5102 -1963
rect -4976 -1973 -4923 -1963
rect -4799 -1973 -4746 -1963
rect -4621 -1973 -4568 -1963
rect -4443 -1973 -4390 -1963
rect -4265 -1973 -4212 -1963
rect -4086 -1973 -4033 -1963
rect -3909 -1973 -3856 -1963
rect -1109 -1973 -1056 -1963
rect -1109 -2425 -1056 -2415
rect -752 -2425 -699 -2415
rect -1056 -2478 -752 -2425
rect -1109 -2488 -1056 -2478
rect -752 -2488 -699 -2478
rect 1919 -2426 1972 -2416
rect 2275 -2426 2328 -2416
rect 3193 -2426 3246 -2417
rect 1972 -2479 2275 -2426
rect 2328 -2427 3246 -2426
rect 2328 -2479 3193 -2427
rect 1919 -2489 1972 -2479
rect 2275 -2489 2328 -2479
rect 3193 -2490 3246 -2480
rect -6498 -2529 -6445 -2519
rect -5777 -2529 -5724 -2520
rect -6445 -2530 -5724 -2529
rect -5066 -2530 -5013 -2520
rect -4354 -2530 -4301 -2520
rect -6445 -2582 -5777 -2530
rect -6498 -2592 -6445 -2582
rect -5724 -2583 -5066 -2530
rect -5013 -2583 -4354 -2530
rect -5777 -2593 -5724 -2583
rect -5066 -2593 -5013 -2583
rect -4354 -2593 -4301 -2583
rect -2624 -2558 -2571 -2548
rect -1285 -2558 -1232 -2548
rect -930 -2558 -877 -2548
rect -2571 -2611 -1285 -2558
rect -1232 -2611 -930 -2558
rect -2624 -2621 -2571 -2611
rect -1285 -2621 -1232 -2611
rect -930 -2621 -877 -2611
rect 2097 -2554 2150 -2544
rect 2453 -2554 2506 -2544
rect 2150 -2607 2453 -2554
rect 2097 -2617 2150 -2607
rect 2453 -2617 2506 -2607
rect -5421 -2668 -5368 -2658
rect -4710 -2668 -4657 -2658
rect -3998 -2668 -3945 -2658
rect -3298 -2668 -3245 -2658
rect -5368 -2721 -4710 -2668
rect -4657 -2721 -3998 -2668
rect -3945 -2721 -3298 -2668
rect -5421 -2731 -5368 -2721
rect -4710 -2731 -4657 -2721
rect -3998 -2731 -3945 -2721
rect -3298 -2731 -3245 -2721
rect -1197 -2665 -1144 -2655
rect -1019 -2665 -966 -2655
rect -841 -2665 -788 -2655
rect -129 -2665 -76 -2655
rect 50 -2665 103 -2655
rect 227 -2665 280 -2655
rect 940 -2665 993 -2655
rect 1117 -2665 1170 -2655
rect 1295 -2665 1348 -2655
rect 2007 -2665 2060 -2655
rect 2186 -2665 2239 -2655
rect 2363 -2665 2416 -2655
rect -1144 -2718 -1019 -2665
rect -966 -2718 -841 -2665
rect -788 -2718 -129 -2665
rect -76 -2718 50 -2665
rect 103 -2718 227 -2665
rect 280 -2718 940 -2665
rect 993 -2718 1117 -2665
rect 1170 -2718 1295 -2665
rect 1348 -2718 2007 -2665
rect 2060 -2718 2186 -2665
rect 2239 -2718 2363 -2665
rect -1197 -2728 -1144 -2718
rect -1019 -2728 -966 -2718
rect -841 -2728 -788 -2718
rect -129 -2728 -76 -2718
rect 50 -2728 103 -2718
rect 227 -2728 280 -2718
rect 940 -2728 993 -2718
rect 1117 -2728 1170 -2718
rect 1295 -2728 1348 -2718
rect 2007 -2728 2060 -2718
rect 2186 -2728 2239 -2718
rect 2363 -2728 2416 -2718
rect -6044 -2780 -5991 -2770
rect -5866 -2780 -5813 -2770
rect -5991 -2833 -5866 -2780
rect -6044 -2843 -5991 -2833
rect -5866 -2843 -5813 -2833
rect -3908 -2780 -3855 -2770
rect -3731 -2780 -3678 -2770
rect -3855 -2833 -3731 -2780
rect -3908 -2843 -3855 -2833
rect -3731 -2843 -3678 -2833
rect -484 -3301 -431 -3291
rect 583 -3301 636 -3291
rect 1654 -3301 1707 -3291
rect -431 -3354 583 -3301
rect 636 -3354 1654 -3301
rect -484 -3364 -431 -3354
rect 583 -3364 636 -3354
rect 1654 -3364 1707 -3354
rect -6625 -3401 -6572 -3391
rect -6134 -3401 -6081 -3391
rect -5066 -3401 -5013 -3391
rect -6572 -3454 -6134 -3401
rect -6081 -3454 -5066 -3401
rect -6625 -3464 -6572 -3454
rect -6134 -3464 -6081 -3454
rect -5066 -3464 -5013 -3454
rect -4710 -3401 -4657 -3391
rect -3642 -3401 -3589 -3391
rect -3131 -3401 -3078 -3391
rect -4657 -3454 -3642 -3401
rect -3589 -3454 -3131 -3401
rect -4710 -3464 -4657 -3454
rect -3642 -3464 -3589 -3454
rect -3131 -3464 -3078 -3454
rect -1645 -3449 -1584 -3439
rect -5777 -3516 -5724 -3506
rect -3998 -3516 -3945 -3506
rect -3298 -3516 -3245 -3506
rect -5724 -3569 -3998 -3516
rect -3945 -3569 -3298 -3516
rect -1108 -3456 -1055 -3446
rect -750 -3456 -697 -3446
rect -396 -3456 -343 -3446
rect -39 -3456 14 -3446
rect 317 -3456 370 -3446
rect -1584 -3509 -1108 -3456
rect -1055 -3509 -750 -3456
rect -697 -3509 -396 -3456
rect -343 -3509 -39 -3456
rect 14 -3509 317 -3456
rect -1645 -3520 -1584 -3510
rect -1108 -3519 -1055 -3509
rect -750 -3519 -697 -3509
rect -396 -3519 -343 -3509
rect -39 -3519 14 -3509
rect 317 -3519 370 -3509
rect 850 -3456 903 -3446
rect 1206 -3456 1259 -3446
rect 1562 -3456 1615 -3446
rect 1919 -3456 1972 -3446
rect 2275 -3456 2328 -3446
rect 3019 -3452 3080 -3442
rect 903 -3509 1206 -3456
rect 1259 -3509 1562 -3456
rect 1615 -3509 1919 -3456
rect 1972 -3509 2275 -3456
rect 2328 -3509 3019 -3456
rect 850 -3519 903 -3509
rect 1206 -3519 1259 -3509
rect 1562 -3519 1615 -3509
rect 1919 -3519 1972 -3509
rect 2275 -3519 2328 -3509
rect 3080 -3509 3891 -3456
rect 3019 -3523 3080 -3513
rect -5777 -3579 -5724 -3569
rect -3998 -3579 -3945 -3569
rect -3298 -3579 -3245 -3569
rect -1286 -3571 -1233 -3561
rect -929 -3571 -876 -3561
rect -573 -3571 -520 -3561
rect -217 -3571 -164 -3561
rect -1702 -3624 -1286 -3571
rect -1233 -3624 -929 -3571
rect -876 -3624 -573 -3571
rect -520 -3624 -217 -3571
rect -6498 -3640 -6445 -3630
rect -5422 -3640 -5369 -3630
rect -4353 -3640 -4300 -3630
rect -1702 -3640 -1649 -3624
rect -1286 -3634 -1233 -3624
rect -929 -3634 -876 -3624
rect -573 -3634 -520 -3624
rect -217 -3634 -164 -3624
rect 1384 -3564 1437 -3554
rect 1741 -3564 1794 -3554
rect 2097 -3564 2150 -3554
rect 2451 -3564 2504 -3554
rect 1437 -3617 1741 -3564
rect 1794 -3617 2097 -3564
rect 2150 -3617 2451 -3564
rect 1384 -3627 1437 -3617
rect 1741 -3627 1794 -3617
rect 2097 -3627 2150 -3617
rect 2451 -3627 2504 -3617
rect -6445 -3693 -5422 -3640
rect -5369 -3693 -4353 -3640
rect -4300 -3693 -1649 -3640
rect -6498 -3703 -6445 -3693
rect -5422 -3703 -5369 -3693
rect -4353 -3703 -4300 -3693
rect -2546 -3928 -2485 -3693
rect -2546 -3999 -2485 -3989
rect -841 -4192 -788 -4182
rect -662 -4192 -609 -4182
rect -483 -4192 -430 -4182
rect -306 -4192 -253 -4182
rect 407 -4192 460 -4182
rect 583 -4192 636 -4182
rect 761 -4192 814 -4182
rect 1474 -4192 1527 -4182
rect 1652 -4192 1705 -4182
rect 1830 -4192 1883 -4182
rect 2008 -4192 2061 -4182
rect -788 -4245 -662 -4192
rect -609 -4245 -483 -4192
rect -430 -4245 -306 -4192
rect -253 -4245 407 -4192
rect 460 -4245 583 -4192
rect 636 -4245 761 -4192
rect 814 -4245 1474 -4192
rect 1527 -4245 1652 -4192
rect 1705 -4245 1830 -4192
rect 1883 -4245 2008 -4192
rect -841 -4255 -788 -4245
rect -662 -4255 -609 -4245
rect -483 -4255 -430 -4245
rect -306 -4255 -253 -4245
rect 407 -4255 460 -4245
rect 583 -4255 636 -4245
rect 761 -4255 814 -4245
rect 1474 -4255 1527 -4245
rect 1652 -4255 1705 -4245
rect 1830 -4255 1883 -4245
rect 2008 -4255 2061 -4245
rect -6498 -4271 -6445 -4261
rect -5778 -4271 -5725 -4261
rect -3998 -4271 -3945 -4261
rect -6445 -4324 -5778 -4271
rect -5725 -4324 -3998 -4271
rect 2538 -4266 2599 -4256
rect 317 -4304 370 -4294
rect 673 -4304 726 -4294
rect -6498 -4334 -6445 -4324
rect -5778 -4334 -5725 -4324
rect -3998 -4334 -3945 -4324
rect -2357 -4357 317 -4304
rect 370 -4357 673 -4304
rect 2538 -4337 2599 -4327
rect -6134 -4390 -6081 -4380
rect -5066 -4390 -5013 -4380
rect -4709 -4390 -4656 -4380
rect -3642 -4390 -3589 -4380
rect -2357 -4390 -2304 -4357
rect 317 -4367 370 -4357
rect 673 -4367 726 -4357
rect -6081 -4443 -5066 -4390
rect -5013 -4443 -4709 -4390
rect -4656 -4443 -3642 -4390
rect -3589 -4443 -2304 -4390
rect -2004 -4412 -1951 -4402
rect 495 -4412 548 -4402
rect 850 -4412 903 -4402
rect -6134 -4453 -6081 -4443
rect -5066 -4453 -5013 -4443
rect -4709 -4453 -4656 -4443
rect -3642 -4453 -3589 -4443
rect -1951 -4465 495 -4412
rect 548 -4465 850 -4412
rect -2004 -4475 -1951 -4465
rect 495 -4475 548 -4465
rect 850 -4475 903 -4465
rect 2746 -4446 2807 -4436
rect -5422 -4506 -5369 -4496
rect -4353 -4506 -4300 -4496
rect -3298 -4506 -3245 -4496
rect -2385 -4505 -2324 -4495
rect -5369 -4559 -4353 -4506
rect -4300 -4559 -3298 -4506
rect -3245 -4559 -2385 -4506
rect -5422 -4569 -5369 -4559
rect -4353 -4569 -4300 -4559
rect -3298 -4569 -3245 -4559
rect 2746 -4517 2807 -4507
rect -2385 -4576 -2324 -4566
rect 3194 -4805 3246 -4795
rect 4771 -4805 4823 -4795
rect 3246 -4857 4771 -4805
rect 3194 -4867 3246 -4857
rect 4771 -4867 4823 -4857
rect 3021 -5002 3082 -4992
rect 5037 -5006 5090 -4996
rect 4985 -5007 5037 -5006
rect 3082 -5059 5037 -5007
rect 3021 -5073 3082 -5063
rect 5037 -5069 5090 -5059
rect -2385 -5093 -2324 -5083
rect -6498 -5141 -6445 -5131
rect -5422 -5141 -5369 -5131
rect -6445 -5187 -5422 -5147
rect -6498 -5204 -6445 -5194
rect -4353 -5141 -4300 -5131
rect -5369 -5188 -4353 -5148
rect -5422 -5204 -5369 -5194
rect -1287 -5097 -1234 -5087
rect -929 -5097 -876 -5087
rect -572 -5097 -519 -5087
rect -218 -5097 -165 -5087
rect -2324 -5150 -1287 -5097
rect -1234 -5150 -929 -5097
rect -876 -5150 -572 -5097
rect -519 -5150 -218 -5097
rect 1385 -5093 1438 -5083
rect 1740 -5093 1793 -5083
rect 2096 -5093 2149 -5083
rect 2453 -5093 2506 -5083
rect -2385 -5164 -2324 -5154
rect -1287 -5160 -1234 -5150
rect -929 -5160 -876 -5150
rect -572 -5160 -519 -5150
rect -218 -5160 -165 -5150
rect 311 -5148 372 -5138
rect -4353 -5204 -4300 -5194
rect -1105 -5213 -1052 -5203
rect -751 -5213 -698 -5203
rect -396 -5213 -343 -5203
rect -41 -5213 12 -5203
rect 1438 -5146 1740 -5093
rect 1793 -5146 2096 -5093
rect 2149 -5146 2453 -5093
rect 1385 -5156 1438 -5146
rect 1740 -5156 1793 -5146
rect 2096 -5156 2149 -5146
rect 2453 -5156 2506 -5146
rect 311 -5213 372 -5209
rect -6134 -5232 -6081 -5222
rect -5066 -5233 -5013 -5223
rect -6081 -5279 -5066 -5239
rect -6134 -5295 -6081 -5285
rect -3130 -5233 -3077 -5223
rect -5013 -5279 -3130 -5239
rect -5066 -5296 -5013 -5286
rect -1876 -5232 -1823 -5222
rect -3077 -5279 -1876 -5239
rect -3130 -5296 -3077 -5286
rect -1052 -5266 -751 -5213
rect -698 -5266 -396 -5213
rect -343 -5266 -41 -5213
rect 12 -5266 316 -5213
rect 369 -5219 372 -5213
rect 846 -5213 903 -5203
rect 1207 -5213 1260 -5203
rect 1563 -5213 1616 -5203
rect 1917 -5213 1970 -5203
rect 2274 -5213 2327 -5203
rect 4905 -5212 4958 -5202
rect -1876 -5295 -1823 -5285
rect -1646 -5278 -1585 -5268
rect -1105 -5276 -1052 -5266
rect -751 -5276 -698 -5266
rect -396 -5276 -343 -5266
rect -41 -5276 12 -5266
rect 316 -5276 369 -5266
rect 846 -5266 850 -5213
rect 903 -5266 1207 -5213
rect 1260 -5266 1563 -5213
rect 1616 -5266 1917 -5213
rect 1970 -5266 2274 -5213
rect 2327 -5265 4905 -5213
rect 2327 -5266 4958 -5265
rect -6625 -5322 -6572 -5312
rect -4710 -5322 -4657 -5312
rect -6572 -5369 -4710 -5329
rect -6625 -5385 -6572 -5375
rect -3642 -5319 -3589 -5309
rect -4657 -5369 -3642 -5329
rect -4710 -5385 -4657 -5375
rect -2624 -5324 -2571 -5314
rect -3589 -5369 -2624 -5329
rect -3642 -5382 -3589 -5372
rect -1646 -5349 -1585 -5339
rect 846 -5278 907 -5266
rect 1207 -5276 1260 -5266
rect 1563 -5276 1616 -5266
rect 1917 -5276 1970 -5266
rect 2274 -5276 2327 -5266
rect 4905 -5275 4958 -5266
rect 846 -5349 907 -5339
rect -2624 -5387 -2571 -5377
rect -128 -5380 -75 -5370
rect 50 -5380 103 -5370
rect 228 -5380 281 -5370
rect 940 -5380 993 -5371
rect 1119 -5380 1172 -5370
rect 1296 -5380 1349 -5370
rect -5777 -5415 -5724 -5405
rect -3997 -5415 -3944 -5405
rect -5724 -5462 -3997 -5422
rect -5777 -5478 -5724 -5468
rect -3298 -5416 -3245 -5406
rect -3944 -5462 -3298 -5422
rect -3997 -5478 -3944 -5468
rect -75 -5433 50 -5380
rect 103 -5433 228 -5380
rect 281 -5381 1119 -5380
rect 281 -5433 940 -5381
rect -128 -5443 -75 -5433
rect 50 -5443 103 -5433
rect 228 -5443 281 -5433
rect 993 -5433 1119 -5381
rect 1172 -5433 1296 -5380
rect 940 -5444 993 -5434
rect 1119 -5443 1172 -5433
rect 1296 -5443 1349 -5433
rect -3298 -5479 -3245 -5469
rect -5956 -6016 -5903 -6006
rect -5601 -6016 -5548 -6006
rect -5244 -6016 -5191 -6006
rect -4888 -6016 -4835 -6006
rect -4532 -6016 -4479 -6006
rect -4175 -6016 -4122 -6006
rect -3820 -6016 -3767 -6006
rect -5903 -6069 -5601 -6016
rect -5548 -6069 -5244 -6016
rect -5191 -6069 -4888 -6016
rect -4835 -6069 -4532 -6016
rect -4479 -6069 -4175 -6016
rect -4122 -6069 -3820 -6016
rect -5956 -6079 -5903 -6069
rect -5601 -6079 -5548 -6069
rect -5244 -6079 -5191 -6069
rect -4888 -6079 -4835 -6069
rect -4532 -6079 -4479 -6069
rect -4175 -6079 -4122 -6069
rect -3820 -6079 -3767 -6069
rect -2624 -6007 -2571 -5997
rect 2096 -6007 2149 -5997
rect 2452 -6007 2505 -5997
rect -2571 -6060 2096 -6007
rect 2149 -6060 2452 -6007
rect -2624 -6070 -2571 -6060
rect 2096 -6070 2149 -6060
rect 2452 -6070 2505 -6060
rect -5778 -6131 -5725 -6121
rect -5065 -6131 -5012 -6121
rect -4354 -6131 -4301 -6121
rect -3298 -6131 -3245 -6121
rect 1918 -6124 1971 -6114
rect 2275 -6124 2328 -6114
rect -2821 -6125 1918 -6124
rect -5725 -6184 -5065 -6131
rect -5012 -6184 -4354 -6131
rect -4301 -6184 -3298 -6131
rect -5778 -6194 -5725 -6184
rect -5065 -6194 -5012 -6184
rect -4354 -6194 -4301 -6184
rect -3298 -6194 -3245 -6184
rect -2856 -6177 1918 -6125
rect 1971 -6177 2275 -6124
rect -6498 -6248 -6445 -6238
rect -5421 -6248 -5368 -6238
rect -4710 -6248 -4657 -6238
rect -3998 -6247 -3945 -6237
rect -6445 -6301 -5421 -6248
rect -5368 -6301 -4710 -6248
rect -4657 -6300 -3998 -6248
rect -4657 -6301 -3945 -6300
rect -6498 -6311 -6445 -6301
rect -5421 -6311 -5368 -6301
rect -4710 -6311 -4657 -6301
rect -3998 -6310 -3945 -6301
rect -4786 -6378 -4733 -6368
rect -2856 -6401 -2803 -6177
rect 1918 -6187 1971 -6177
rect 2275 -6187 2328 -6177
rect -3874 -6408 -2803 -6401
rect -4733 -6431 -2803 -6408
rect -4786 -6454 -2803 -6431
rect -2702 -6250 -2649 -6249
rect 227 -6250 280 -6240
rect 942 -6250 995 -6240
rect -2702 -6303 227 -6250
rect 280 -6303 942 -6250
rect -4786 -6461 -3820 -6454
rect -3874 -7691 -3821 -6461
rect -2702 -6542 -2649 -6303
rect 227 -6313 280 -6303
rect 942 -6313 995 -6303
rect -1876 -6364 -1823 -6354
rect -1282 -6364 -1229 -6354
rect -1823 -6417 -1282 -6364
rect -1229 -6365 -1177 -6364
rect -928 -6365 -876 -6355
rect 2879 -6365 2931 -6355
rect -1229 -6417 -928 -6365
rect -876 -6417 2879 -6365
rect -1876 -6427 -1823 -6417
rect -1282 -6427 -1229 -6417
rect -928 -6427 -876 -6417
rect 2879 -6427 2931 -6417
rect -1110 -6479 -1057 -6469
rect -752 -6479 -699 -6469
rect -1057 -6532 -752 -6479
rect -1110 -6542 -1057 -6532
rect -752 -6542 -699 -6532
rect -3874 -7743 -3873 -7691
rect -3873 -7753 -3821 -7743
rect -3731 -6595 -2649 -6542
rect -3731 -7785 -3678 -6595
rect -753 -6598 -700 -6588
rect 4772 -6597 4825 -6587
rect -700 -6650 4772 -6598
rect -700 -6651 4825 -6650
rect -753 -6661 -700 -6651
rect 4772 -6660 4825 -6651
rect -2003 -6714 -1950 -6704
rect -1950 -6767 5237 -6714
rect -2003 -6777 -1950 -6767
rect -3545 -6806 -3484 -6796
rect -3545 -6877 -3484 -6867
rect -3679 -7837 -3678 -7785
rect -3541 -7788 -3489 -6877
rect 4770 -6891 4823 -6881
rect -3386 -6979 -3325 -6969
rect 4770 -6996 4823 -6944
rect 4906 -6889 4959 -6879
rect 4906 -6994 4959 -6942
rect -3386 -7050 -3325 -7040
rect -3731 -7847 -3679 -7837
rect -3541 -7850 -3489 -7840
rect -3382 -7933 -3329 -7050
rect 4771 -7844 4823 -6996
rect 4907 -7842 4959 -6994
rect 5038 -6887 5091 -6877
rect 5038 -7840 5091 -6940
rect 4771 -7854 4824 -7844
rect -1382 -7922 -1329 -7912
rect -1203 -7922 -1150 -7913
rect -1025 -7922 -972 -7912
rect -848 -7922 -795 -7912
rect -670 -7922 -617 -7912
rect -490 -7922 -437 -7912
rect 755 -7922 808 -7912
rect 932 -7922 985 -7912
rect 1112 -7922 1165 -7912
rect 1289 -7922 1342 -7913
rect 1467 -7922 1520 -7912
rect 1644 -7922 1697 -7912
rect 2890 -7922 2943 -7912
rect 3069 -7922 3122 -7912
rect 3247 -7922 3300 -7912
rect 3424 -7922 3477 -7912
rect 3603 -7922 3656 -7913
rect 3778 -7922 3831 -7912
rect -1329 -7923 -1025 -7922
rect -1329 -7975 -1203 -7923
rect -1382 -7985 -1329 -7975
rect -1150 -7975 -1025 -7923
rect -972 -7975 -848 -7922
rect -795 -7975 -670 -7922
rect -617 -7975 -490 -7922
rect -437 -7975 755 -7922
rect 808 -7975 932 -7922
rect 985 -7975 1112 -7922
rect 1165 -7923 1467 -7922
rect 1165 -7975 1289 -7923
rect -1203 -7986 -1150 -7976
rect -1025 -7985 -972 -7975
rect -848 -7985 -795 -7975
rect -670 -7985 -617 -7975
rect -490 -7985 -437 -7975
rect 755 -7985 808 -7975
rect 932 -7985 985 -7975
rect 1112 -7985 1165 -7975
rect 1342 -7975 1467 -7923
rect 1520 -7975 1644 -7922
rect 1697 -7975 2890 -7922
rect 2943 -7975 3069 -7922
rect 3122 -7975 3247 -7922
rect 3300 -7975 3424 -7922
rect 3477 -7923 3778 -7922
rect 3477 -7975 3603 -7923
rect 1289 -7986 1342 -7976
rect 1467 -7985 1520 -7975
rect 1644 -7985 1697 -7975
rect 2890 -7985 2943 -7975
rect 3069 -7985 3122 -7975
rect 3247 -7985 3300 -7975
rect 3424 -7985 3477 -7975
rect 3656 -7975 3778 -7923
rect 4208 -7923 4261 -7913
rect 4771 -7917 4824 -7907
rect 4906 -7852 4959 -7842
rect 4906 -7915 4959 -7905
rect 5037 -7850 5091 -7840
rect 5090 -7898 5091 -7850
rect 5184 -7855 5237 -6767
rect 5037 -7913 5090 -7903
rect 5184 -7918 5237 -7908
rect 5337 -7850 5390 -6425
rect 5337 -7913 5390 -7903
rect 3831 -7975 4208 -7923
rect 3603 -7986 3656 -7976
rect 3778 -7976 4208 -7975
rect 3778 -7985 3831 -7976
rect 4208 -7986 4261 -7976
rect -3382 -7996 -3329 -7986
rect -1916 -8534 -1863 -8524
rect -1739 -8534 -1686 -8524
rect -1558 -8534 -1505 -8524
rect -1382 -8534 -1329 -8524
rect -1203 -8534 -1150 -8524
rect -1026 -8534 -973 -8524
rect -848 -8534 -795 -8524
rect -670 -8534 -617 -8524
rect -491 -8534 -438 -8524
rect -314 -8534 -261 -8524
rect -136 -8534 -83 -8524
rect 42 -8534 95 -8524
rect 221 -8534 274 -8524
rect 398 -8534 451 -8524
rect 577 -8534 630 -8524
rect 754 -8534 807 -8524
rect 932 -8534 985 -8524
rect 1111 -8534 1164 -8524
rect 1289 -8534 1342 -8524
rect 1466 -8534 1519 -8524
rect 1644 -8534 1697 -8524
rect 1822 -8534 1875 -8524
rect 2000 -8534 2053 -8524
rect 2178 -8534 2231 -8524
rect 2357 -8534 2410 -8524
rect 2534 -8534 2587 -8524
rect 2712 -8534 2765 -8524
rect 2890 -8534 2943 -8524
rect 3068 -8534 3121 -8524
rect 3246 -8534 3299 -8524
rect 3424 -8534 3477 -8524
rect 3602 -8534 3655 -8524
rect 3781 -8534 3834 -8524
rect -1863 -8587 -1739 -8534
rect -1686 -8587 -1558 -8534
rect -1505 -8587 -1382 -8534
rect -1329 -8587 -1203 -8534
rect -1150 -8587 -1026 -8534
rect -973 -8587 -848 -8534
rect -795 -8587 -670 -8534
rect -617 -8587 -491 -8534
rect -438 -8587 -314 -8534
rect -261 -8587 -136 -8534
rect -83 -8587 42 -8534
rect 95 -8587 221 -8534
rect 274 -8587 398 -8534
rect 451 -8587 577 -8534
rect 630 -8587 754 -8534
rect 807 -8587 932 -8534
rect 985 -8587 1111 -8534
rect 1164 -8587 1289 -8534
rect 1342 -8587 1466 -8534
rect 1519 -8587 1644 -8534
rect 1697 -8587 1822 -8534
rect 1875 -8587 2000 -8534
rect 2053 -8587 2178 -8534
rect 2231 -8587 2357 -8534
rect 2410 -8587 2534 -8534
rect 2587 -8587 2712 -8534
rect 2765 -8587 2890 -8534
rect 2943 -8587 3068 -8534
rect 3121 -8587 3246 -8534
rect 3299 -8587 3424 -8534
rect 3477 -8587 3602 -8534
rect 3655 -8587 3781 -8534
rect -1916 -8597 -1863 -8587
rect -1739 -8597 -1686 -8587
rect -1558 -8597 -1505 -8587
rect -1382 -8597 -1329 -8587
rect -1203 -8597 -1150 -8587
rect -1026 -8597 -973 -8587
rect -848 -8597 -795 -8587
rect -670 -8597 -617 -8587
rect -491 -8597 -438 -8587
rect -314 -8597 -261 -8587
rect -136 -8597 -83 -8587
rect 42 -8597 95 -8587
rect 221 -8597 274 -8587
rect 398 -8597 451 -8587
rect 577 -8597 630 -8587
rect 754 -8597 807 -8587
rect 932 -8597 985 -8587
rect 1111 -8597 1164 -8587
rect 1289 -8597 1342 -8587
rect 1466 -8597 1519 -8587
rect 1644 -8597 1697 -8587
rect 1822 -8597 1875 -8587
rect 2000 -8597 2053 -8587
rect 2178 -8597 2231 -8587
rect 2357 -8597 2410 -8587
rect 2534 -8597 2587 -8587
rect 2712 -8597 2765 -8587
rect 2890 -8597 2943 -8587
rect 3068 -8597 3121 -8587
rect 3246 -8597 3299 -8587
rect 3424 -8597 3477 -8587
rect 3602 -8597 3655 -8587
rect 3781 -8597 3834 -8587
rect 5185 -8633 5237 -8625
rect 5185 -8635 10564 -8633
rect -1826 -8653 -1773 -8643
rect -1470 -8653 -1417 -8643
rect -1115 -8653 -1062 -8643
rect -758 -8653 -705 -8643
rect -402 -8653 -349 -8643
rect -47 -8653 6 -8643
rect 310 -8653 363 -8643
rect 666 -8653 719 -8643
rect 1022 -8653 1075 -8643
rect 1377 -8653 1430 -8643
rect 1733 -8653 1786 -8643
rect 2090 -8653 2143 -8643
rect 2446 -8653 2499 -8643
rect 2802 -8653 2855 -8643
rect 3158 -8653 3211 -8643
rect 3513 -8653 3566 -8643
rect 3869 -8653 3922 -8643
rect -1773 -8706 -1470 -8653
rect -1417 -8706 -1115 -8653
rect -1062 -8706 -758 -8653
rect -705 -8706 -402 -8653
rect -349 -8706 -47 -8653
rect 6 -8706 310 -8653
rect 363 -8706 666 -8653
rect 719 -8706 1022 -8653
rect 1075 -8706 1377 -8653
rect 1430 -8706 1733 -8653
rect 1786 -8706 2090 -8653
rect 2143 -8706 2446 -8653
rect 2499 -8706 2802 -8653
rect 2855 -8706 3158 -8653
rect 3211 -8706 3513 -8653
rect 3566 -8706 3869 -8653
rect 5237 -8685 10564 -8635
rect 5185 -8697 5237 -8687
rect -1826 -8716 -1773 -8706
rect -1470 -8716 -1417 -8706
rect -1115 -8716 -1062 -8706
rect -758 -8716 -705 -8706
rect -402 -8716 -349 -8706
rect -47 -8716 6 -8706
rect 310 -8716 363 -8706
rect 666 -8716 719 -8706
rect 1022 -8716 1075 -8706
rect 1377 -8716 1430 -8706
rect 1733 -8716 1786 -8706
rect 2090 -8716 2143 -8706
rect 2446 -8716 2499 -8706
rect 2802 -8716 2855 -8706
rect 3158 -8716 3211 -8706
rect 3513 -8716 3566 -8706
rect 3869 -8716 3922 -8706
rect 10512 -8716 10564 -8685
rect 11054 -8716 11107 -8706
rect 11345 -8716 11398 -8706
rect 11638 -8716 11691 -8706
rect 11932 -8716 11985 -8706
rect 12222 -8716 12275 -8706
rect -2447 -8767 -2394 -8757
rect -2005 -8767 -1952 -8757
rect -1648 -8767 -1595 -8757
rect -1293 -8767 -1240 -8757
rect -936 -8767 -883 -8757
rect -580 -8766 -527 -8756
rect -2394 -8820 -2005 -8767
rect -1952 -8820 -1648 -8767
rect -1595 -8820 -1293 -8767
rect -1240 -8820 -936 -8767
rect -883 -8819 -580 -8767
rect -225 -8767 -172 -8757
rect 132 -8767 185 -8758
rect 489 -8766 542 -8756
rect -527 -8819 -225 -8767
rect -883 -8820 -225 -8819
rect -172 -8768 489 -8767
rect -172 -8820 132 -8768
rect -2447 -8830 -2394 -8820
rect -2005 -8830 -1952 -8820
rect -1648 -8830 -1595 -8820
rect -1293 -8830 -1240 -8820
rect -936 -8830 -883 -8820
rect -580 -8829 -527 -8820
rect -225 -8830 -172 -8820
rect 185 -8819 489 -8768
rect 843 -8766 896 -8756
rect 542 -8819 843 -8767
rect 1201 -8767 1254 -8757
rect 1556 -8767 1609 -8757
rect 1911 -8767 1964 -8757
rect 2267 -8767 2320 -8757
rect 2624 -8767 2677 -8757
rect 2980 -8767 3033 -8757
rect 3336 -8767 3389 -8757
rect 3692 -8767 3745 -8757
rect 896 -8819 1201 -8767
rect 185 -8820 1201 -8819
rect 1254 -8820 1556 -8767
rect 1609 -8820 1911 -8767
rect 1964 -8820 2267 -8767
rect 2320 -8820 2624 -8767
rect 2677 -8820 2980 -8767
rect 3033 -8820 3336 -8767
rect 3389 -8820 3692 -8767
rect 10512 -8768 11054 -8716
rect 10584 -8769 11054 -8768
rect 11107 -8769 11345 -8716
rect 11398 -8769 11638 -8716
rect 11691 -8769 11932 -8716
rect 11985 -8769 12222 -8716
rect 11054 -8779 11107 -8769
rect 11345 -8779 11398 -8769
rect 11638 -8779 11691 -8769
rect 11932 -8779 11985 -8769
rect 12222 -8779 12275 -8769
rect 132 -8831 185 -8821
rect 489 -8829 542 -8820
rect 843 -8829 896 -8820
rect 1201 -8830 1254 -8820
rect 1556 -8830 1609 -8820
rect 1911 -8830 1964 -8820
rect 2267 -8830 2320 -8820
rect 2624 -8830 2677 -8820
rect 2980 -8830 3033 -8820
rect 3336 -8830 3389 -8820
rect 3692 -8830 3745 -8820
rect 4771 -9314 4824 -9304
rect 6769 -9314 6822 -9304
rect 6947 -9314 7000 -9305
rect 7126 -9314 7179 -9305
rect 7303 -9313 7356 -9303
rect 4824 -9367 6769 -9314
rect 6822 -9315 7303 -9314
rect 6822 -9367 6947 -9315
rect 4771 -9377 4824 -9367
rect 6769 -9377 6822 -9367
rect 7000 -9367 7126 -9315
rect 6947 -9378 7000 -9368
rect 7179 -9366 7303 -9315
rect 7482 -9313 7535 -9303
rect 7356 -9366 7482 -9314
rect 7659 -9314 7712 -9305
rect 7837 -9314 7890 -9304
rect 8015 -9314 8068 -9305
rect 8194 -9314 8247 -9304
rect 8371 -9314 8424 -9304
rect 8549 -9314 8602 -9304
rect 8727 -9314 8780 -9305
rect 8906 -9314 8959 -9304
rect 7535 -9315 7837 -9314
rect 7535 -9366 7659 -9315
rect 7179 -9367 7659 -9366
rect 7126 -9378 7179 -9368
rect 7303 -9376 7356 -9367
rect 7482 -9376 7535 -9367
rect 7712 -9367 7837 -9315
rect 7890 -9315 8194 -9314
rect 7890 -9367 8015 -9315
rect 7659 -9378 7712 -9368
rect 7837 -9377 7890 -9367
rect 8068 -9367 8194 -9315
rect 8247 -9367 8371 -9314
rect 8424 -9367 8549 -9314
rect 8602 -9315 8906 -9314
rect 8602 -9367 8727 -9315
rect 8015 -9378 8068 -9368
rect 8194 -9377 8247 -9367
rect 8371 -9377 8424 -9367
rect 8549 -9377 8602 -9367
rect 8780 -9367 8906 -9315
rect 8727 -9378 8780 -9368
rect 8906 -9377 8959 -9367
rect 11144 -9374 11197 -9364
rect 11436 -9375 11489 -9365
rect 11728 -9375 11781 -9365
rect 12020 -9375 12073 -9366
rect 12312 -9375 12365 -9365
rect 11197 -9427 11436 -9375
rect 11144 -9428 11436 -9427
rect 11489 -9428 11728 -9375
rect 11781 -9376 12312 -9375
rect 11781 -9428 12020 -9376
rect 11144 -9437 11197 -9428
rect 11436 -9438 11489 -9428
rect 11728 -9438 11781 -9428
rect 12073 -9428 12312 -9376
rect 12020 -9439 12073 -9429
rect 12312 -9438 12365 -9428
rect -1916 -9546 -1863 -9536
rect -1738 -9546 -1685 -9536
rect -1558 -9546 -1505 -9536
rect -312 -9546 -259 -9536
rect -136 -9545 -83 -9535
rect -1863 -9599 -1738 -9546
rect -1685 -9599 -1558 -9546
rect -1505 -9599 -312 -9546
rect -259 -9598 -136 -9546
rect 42 -9546 95 -9536
rect 222 -9545 275 -9535
rect -83 -9598 42 -9546
rect -259 -9599 42 -9598
rect 95 -9598 222 -9546
rect 399 -9546 452 -9536
rect 577 -9546 630 -9536
rect 2178 -9546 2231 -9537
rect 2357 -9546 2410 -9536
rect 2534 -9546 2587 -9536
rect 2713 -9546 2766 -9536
rect 4208 -9546 4261 -9536
rect 6679 -9545 6732 -9535
rect 275 -9598 399 -9546
rect 95 -9599 399 -9598
rect 452 -9599 577 -9546
rect 630 -9547 2357 -9546
rect 630 -9599 2178 -9547
rect -1916 -9609 -1863 -9599
rect -1738 -9609 -1685 -9599
rect -1558 -9609 -1505 -9599
rect -312 -9609 -259 -9599
rect -136 -9608 -83 -9599
rect 42 -9609 95 -9599
rect 222 -9608 275 -9599
rect 399 -9609 452 -9599
rect 577 -9609 630 -9599
rect 2231 -9599 2357 -9547
rect 2410 -9599 2534 -9546
rect 2587 -9599 2713 -9546
rect 2766 -9599 4208 -9546
rect 4261 -9598 6679 -9546
rect 4261 -9599 6732 -9598
rect 2178 -9610 2231 -9600
rect 2357 -9609 2410 -9599
rect 2534 -9609 2587 -9599
rect 2713 -9609 2766 -9599
rect 4208 -9609 4261 -9599
rect 6679 -9608 6732 -9599
rect -2315 -9925 -2262 -9915
rect -1916 -9925 -1863 -9915
rect -1738 -9925 -1685 -9916
rect -1560 -9925 -1507 -9915
rect -1382 -9924 -1329 -9914
rect -2262 -9978 -1916 -9925
rect -1863 -9926 -1560 -9925
rect -1863 -9978 -1738 -9926
rect -2315 -9988 -2262 -9978
rect -1916 -9988 -1863 -9978
rect -1685 -9978 -1560 -9926
rect -1507 -9977 -1382 -9925
rect -314 -9925 -261 -9915
rect -136 -9925 -83 -9916
rect 43 -9925 96 -9915
rect 220 -9925 273 -9915
rect 398 -9925 451 -9915
rect 576 -9925 629 -9915
rect 2356 -9925 2409 -9915
rect 2534 -9925 2587 -9915
rect 2712 -9925 2765 -9916
rect 2891 -9925 2944 -9915
rect 3069 -9925 3122 -9915
rect 3246 -9925 3299 -9915
rect 5337 -9925 5390 -9915
rect -1329 -9977 -314 -9925
rect -1507 -9978 -314 -9977
rect -261 -9926 43 -9925
rect -261 -9978 -136 -9926
rect -1738 -9989 -1685 -9979
rect -1560 -9988 -1507 -9978
rect -1382 -9987 -1329 -9978
rect -314 -9988 -261 -9978
rect -83 -9978 43 -9926
rect 96 -9978 220 -9925
rect 273 -9978 398 -9925
rect 451 -9978 576 -9925
rect 629 -9978 2356 -9925
rect 2409 -9978 2534 -9925
rect 2587 -9926 2891 -9925
rect 2587 -9978 2712 -9926
rect -136 -9989 -83 -9979
rect 43 -9988 96 -9978
rect 220 -9988 273 -9978
rect 398 -9988 451 -9978
rect 576 -9988 629 -9978
rect 2356 -9988 2409 -9978
rect 2534 -9988 2587 -9978
rect 2765 -9978 2891 -9926
rect 2944 -9978 3069 -9925
rect 3122 -9978 3246 -9925
rect 3299 -9978 5337 -9925
rect 2712 -9989 2765 -9979
rect 2891 -9988 2944 -9978
rect 3069 -9988 3122 -9978
rect 3246 -9988 3299 -9978
rect 5337 -9988 5390 -9978
rect 6680 -10313 6733 -10303
rect 9171 -10313 9224 -10304
rect 6733 -10314 9224 -10313
rect 6733 -10366 9171 -10314
rect 6680 -10376 6733 -10366
rect 9171 -10377 9224 -10367
rect 6858 -10466 6911 -10457
rect 7214 -10466 7267 -10456
rect 7571 -10466 7624 -10456
rect 7927 -10466 7980 -10456
rect 8283 -10466 8336 -10457
rect 8638 -10466 8691 -10456
rect 8995 -10466 9048 -10457
rect 6858 -10467 7214 -10466
rect 6911 -10519 7214 -10467
rect 7267 -10519 7571 -10466
rect 7624 -10519 7927 -10466
rect 7980 -10467 8638 -10466
rect 7980 -10519 8283 -10467
rect 6858 -10530 6911 -10520
rect 7214 -10529 7267 -10519
rect 7571 -10529 7624 -10519
rect 7927 -10529 7980 -10519
rect 8336 -10519 8638 -10467
rect 8691 -10467 9048 -10466
rect 8691 -10519 8995 -10467
rect 8283 -10530 8336 -10520
rect 8638 -10529 8691 -10519
rect 8995 -10530 9048 -10520
rect -1827 -10908 -1774 -10898
rect -1470 -10908 -1417 -10898
rect -1114 -10908 -1061 -10898
rect -758 -10908 -705 -10898
rect -402 -10908 -349 -10898
rect -46 -10908 7 -10898
rect 309 -10908 362 -10898
rect 665 -10908 718 -10898
rect 931 -10908 984 -10898
rect 1199 -10908 1252 -10898
rect 1556 -10908 1609 -10898
rect 1913 -10908 1966 -10898
rect 2268 -10908 2321 -10898
rect 2623 -10908 2676 -10898
rect 2980 -10908 3033 -10898
rect 3335 -10908 3388 -10898
rect 3692 -10908 3745 -10898
rect -1774 -10961 -1470 -10908
rect -1417 -10961 -1114 -10908
rect -1061 -10961 -758 -10908
rect -705 -10961 -402 -10908
rect -349 -10961 -46 -10908
rect 7 -10961 309 -10908
rect 362 -10961 665 -10908
rect 718 -10961 931 -10908
rect 984 -10961 1199 -10908
rect 1252 -10961 1556 -10908
rect 1609 -10961 1913 -10908
rect 1966 -10961 2268 -10908
rect 2321 -10961 2623 -10908
rect 2676 -10961 2980 -10908
rect 3033 -10961 3335 -10908
rect 3388 -10961 3692 -10908
rect -1827 -10971 -1774 -10961
rect -1470 -10971 -1417 -10961
rect -1114 -10971 -1061 -10961
rect -758 -10971 -705 -10961
rect -402 -10971 -349 -10961
rect -46 -10971 7 -10961
rect 309 -10971 362 -10961
rect 665 -10971 718 -10961
rect 931 -10971 984 -10961
rect 1199 -10971 1252 -10961
rect 1556 -10971 1609 -10961
rect 1913 -10971 1966 -10961
rect 2268 -10971 2321 -10961
rect 2623 -10971 2676 -10961
rect 2980 -10971 3033 -10961
rect 3335 -10971 3388 -10961
rect 3692 -10971 3745 -10961
rect 7037 -11366 7090 -11356
rect 7393 -11366 7446 -11356
rect 7748 -11366 7801 -11357
rect 8103 -11366 8156 -11356
rect 8461 -11366 8514 -11356
rect 8817 -11366 8870 -11356
rect 7090 -11419 7393 -11366
rect 7446 -11367 8103 -11366
rect 7446 -11419 7748 -11367
rect 7037 -11429 7090 -11419
rect 7393 -11429 7446 -11419
rect 7801 -11419 8103 -11367
rect 8156 -11419 8461 -11366
rect 8514 -11419 8817 -11366
rect 7748 -11430 7801 -11420
rect 8103 -11429 8156 -11419
rect 8461 -11429 8514 -11419
rect 8817 -11429 8870 -11419
rect -1649 -11528 -1596 -11518
rect -1293 -11528 -1240 -11518
rect -937 -11528 -884 -11518
rect 1377 -11528 1430 -11518
rect 1733 -11528 1786 -11518
rect 2089 -11528 2142 -11518
rect -1596 -11581 -1293 -11528
rect -1240 -11581 -937 -11528
rect -884 -11581 1377 -11528
rect 1430 -11581 1733 -11528
rect 1786 -11581 2089 -11528
rect -1649 -11591 -1596 -11581
rect -1293 -11591 -1240 -11581
rect -937 -11591 -884 -11581
rect 1377 -11591 1430 -11581
rect 1733 -11591 1786 -11581
rect 2089 -11591 2142 -11581
rect -2004 -11637 -1951 -11627
rect -580 -11637 -527 -11627
rect 2446 -11637 2499 -11627
rect 3871 -11637 3924 -11628
rect -1951 -11690 -580 -11637
rect -527 -11690 2446 -11637
rect 2499 -11638 3924 -11637
rect 2499 -11690 3871 -11638
rect -2004 -11700 -1951 -11690
rect -580 -11700 -527 -11690
rect 2446 -11700 2499 -11690
rect 3871 -11701 3924 -11691
rect 11053 -11674 11106 -11664
rect 11347 -11674 11400 -11665
rect 11638 -11674 11691 -11664
rect 11931 -11674 11984 -11664
rect 12223 -11674 12276 -11664
rect 13022 -11673 13075 -11663
rect 11106 -11675 11638 -11674
rect 11106 -11727 11347 -11675
rect 11053 -11737 11106 -11727
rect 11400 -11727 11638 -11675
rect 11691 -11727 11931 -11674
rect 11984 -11727 12223 -11674
rect 12276 -11726 13022 -11674
rect 12276 -11727 13075 -11726
rect 11347 -11738 11400 -11728
rect 11638 -11737 11691 -11727
rect 11931 -11737 11984 -11727
rect 12223 -11737 12276 -11727
rect 13022 -11736 13075 -11727
rect -224 -11757 -171 -11747
rect 131 -11757 184 -11747
rect 487 -11757 540 -11747
rect 2800 -11757 2853 -11747
rect 3157 -11757 3210 -11747
rect 3513 -11757 3566 -11747
rect -171 -11810 131 -11757
rect 184 -11810 487 -11757
rect 540 -11810 2800 -11757
rect 2853 -11810 3157 -11757
rect 3210 -11810 3513 -11757
rect -224 -11820 -171 -11810
rect 131 -11820 184 -11810
rect 487 -11820 540 -11810
rect 2800 -11820 2853 -11810
rect 3157 -11820 3210 -11810
rect 3513 -11820 3566 -11810
rect -1915 -11919 -1862 -11909
rect -1738 -11919 -1685 -11909
rect -1559 -11919 -1506 -11909
rect -1381 -11919 -1328 -11909
rect -1203 -11919 -1150 -11909
rect -1025 -11919 -972 -11909
rect -848 -11919 -795 -11909
rect -670 -11919 -617 -11909
rect -492 -11919 -439 -11909
rect -314 -11919 -261 -11909
rect -136 -11919 -83 -11909
rect 42 -11919 95 -11909
rect 220 -11919 273 -11909
rect 399 -11919 452 -11909
rect 577 -11919 630 -11909
rect 1288 -11919 1341 -11909
rect 1468 -11919 1521 -11909
rect 1644 -11919 1697 -11910
rect 1823 -11919 1876 -11909
rect 2000 -11919 2053 -11909
rect 2178 -11919 2231 -11909
rect 2357 -11919 2410 -11909
rect 2534 -11919 2587 -11909
rect 2713 -11919 2766 -11909
rect 2890 -11919 2943 -11909
rect 3068 -11919 3121 -11909
rect 3247 -11919 3300 -11909
rect 3425 -11919 3478 -11909
rect 3603 -11919 3656 -11909
rect 3781 -11919 3834 -11909
rect -1862 -11972 -1738 -11919
rect -1685 -11972 -1559 -11919
rect -1506 -11972 -1381 -11919
rect -1328 -11972 -1203 -11919
rect -1150 -11972 -1025 -11919
rect -972 -11972 -848 -11919
rect -795 -11972 -670 -11919
rect -617 -11972 -492 -11919
rect -439 -11972 -314 -11919
rect -261 -11972 -136 -11919
rect -83 -11972 42 -11919
rect 95 -11972 220 -11919
rect 273 -11972 399 -11919
rect 452 -11972 577 -11919
rect 630 -11972 1288 -11919
rect 1341 -11972 1468 -11919
rect 1521 -11920 1823 -11919
rect 1521 -11972 1644 -11920
rect -1915 -11982 -1862 -11972
rect -1738 -11982 -1685 -11972
rect -1559 -11982 -1506 -11972
rect -1381 -11982 -1328 -11972
rect -1203 -11982 -1150 -11972
rect -1025 -11982 -972 -11972
rect -848 -11982 -795 -11972
rect -670 -11982 -617 -11972
rect -492 -11982 -439 -11972
rect -314 -11982 -261 -11972
rect -136 -11982 -83 -11972
rect 42 -11982 95 -11972
rect 220 -11982 273 -11972
rect 399 -11982 452 -11972
rect 577 -11982 630 -11972
rect 1288 -11982 1341 -11972
rect 1468 -11982 1521 -11972
rect 1697 -11972 1823 -11920
rect 1876 -11972 2000 -11919
rect 2053 -11972 2178 -11919
rect 2231 -11972 2357 -11919
rect 2410 -11972 2534 -11919
rect 2587 -11972 2713 -11919
rect 2766 -11972 2890 -11919
rect 2943 -11972 3068 -11919
rect 3121 -11972 3247 -11919
rect 3300 -11972 3425 -11919
rect 3478 -11972 3603 -11919
rect 3656 -11972 3781 -11919
rect 1644 -11983 1697 -11973
rect 1823 -11982 1876 -11972
rect 2000 -11982 2053 -11972
rect 2178 -11982 2231 -11972
rect 2357 -11982 2410 -11972
rect 2534 -11982 2587 -11972
rect 2713 -11982 2766 -11972
rect 2890 -11982 2943 -11972
rect 3068 -11982 3121 -11972
rect 3247 -11982 3300 -11972
rect 3425 -11982 3478 -11972
rect 3603 -11982 3656 -11972
rect 3781 -11982 3834 -11972
rect -5502 -12271 -5449 -12261
rect -5000 -12271 -4947 -12262
rect -4502 -12271 -4449 -12261
rect -5449 -12272 -4502 -12271
rect -5449 -12324 -5000 -12272
rect -5502 -12334 -5449 -12324
rect -4947 -12324 -4502 -12272
rect -2447 -12272 -2394 -12262
rect -4449 -12324 -2447 -12272
rect -5000 -12335 -4947 -12325
rect -4502 -12325 -2447 -12324
rect -4502 -12334 -4449 -12325
rect -2447 -12335 -2394 -12325
rect -5376 -12388 -5323 -12378
rect -5127 -12388 -5074 -12378
rect -4377 -12388 -4324 -12378
rect -3928 -12388 -3875 -12379
rect -5323 -12441 -5127 -12388
rect -5074 -12441 -4377 -12388
rect -4324 -12389 -3875 -12388
rect -4324 -12441 -3928 -12389
rect -5376 -12451 -5323 -12441
rect -5127 -12451 -5074 -12441
rect -4377 -12451 -4324 -12441
rect -3928 -12452 -3875 -12442
rect -6077 -12512 -6024 -12502
rect -5626 -12512 -5573 -12502
rect -4877 -12512 -4824 -12502
rect -4627 -12512 -4574 -12502
rect -6024 -12565 -5626 -12512
rect -5573 -12565 -4877 -12512
rect -4824 -12565 -4627 -12512
rect -6077 -12575 -6024 -12565
rect -5626 -12575 -5573 -12565
rect -4877 -12575 -4824 -12565
rect -4627 -12575 -4574 -12565
rect -2005 -12542 -1952 -12532
rect -1649 -12542 -1596 -12532
rect 3514 -12542 3567 -12532
rect 3871 -12542 3924 -12532
rect -1952 -12595 -1649 -12542
rect -1596 -12544 -1284 -12542
rect -1250 -12544 3514 -12542
rect -1596 -12595 3514 -12544
rect 3567 -12595 3871 -12542
rect -2005 -12605 -1952 -12595
rect -1649 -12605 -1596 -12595
rect 3514 -12605 3567 -12595
rect 3871 -12605 3924 -12595
rect -1294 -12653 -1241 -12644
rect -582 -12653 -529 -12643
rect 130 -12653 183 -12643
rect 1735 -12653 1788 -12644
rect 2445 -12653 2498 -12643
rect 3158 -12652 3211 -12642
rect -1294 -12654 -582 -12653
rect -1241 -12706 -582 -12654
rect -529 -12706 130 -12653
rect 183 -12654 2445 -12653
rect 183 -12706 1735 -12654
rect -1294 -12717 -1241 -12707
rect -582 -12716 -529 -12706
rect 130 -12716 183 -12706
rect 1788 -12706 2445 -12654
rect 2498 -12705 3158 -12653
rect 2498 -12706 3211 -12705
rect 1735 -12717 1788 -12707
rect 2445 -12716 2498 -12706
rect 3158 -12715 3211 -12706
rect -937 -12783 -884 -12773
rect -224 -12783 -171 -12773
rect 486 -12783 539 -12774
rect 1378 -12783 1431 -12773
rect 2088 -12782 2141 -12772
rect -884 -12836 -224 -12783
rect -171 -12784 1378 -12783
rect -171 -12836 486 -12784
rect -937 -12846 -884 -12836
rect -224 -12846 -171 -12836
rect 539 -12836 1378 -12784
rect 1431 -12835 2088 -12783
rect 2801 -12782 2854 -12772
rect 2141 -12835 2801 -12783
rect 1431 -12836 2854 -12835
rect 486 -12847 539 -12837
rect 1378 -12846 1431 -12836
rect 2088 -12845 2141 -12836
rect 2801 -12845 2854 -12836
rect -6223 -13062 -6170 -13052
rect -5751 -13062 -5698 -13052
rect -4752 -13062 -4699 -13052
rect -6170 -13115 -5751 -13062
rect -5698 -13115 -4752 -13062
rect -6223 -13125 -6170 -13115
rect -5751 -13125 -5698 -13115
rect -4752 -13125 -4699 -13115
rect -5251 -13189 -5198 -13179
rect -4251 -13189 -4198 -13179
rect -3788 -13189 -3735 -13179
rect -3542 -13189 -3489 -13179
rect -5198 -13242 -4251 -13189
rect -4198 -13242 -3788 -13189
rect -3735 -13242 -3542 -13189
rect -5251 -13252 -5198 -13242
rect -4251 -13252 -4198 -13242
rect -3788 -13252 -3735 -13242
rect -3542 -13252 -3489 -13242
rect 5037 -13296 5090 -13286
rect 5534 -13296 5587 -13286
rect 5090 -13349 5534 -13296
rect 5037 -13359 5090 -13349
rect 5534 -13359 5587 -13349
rect 5031 -13433 5084 -13423
rect 8950 -13433 9003 -13423
rect 9305 -13433 9358 -13423
rect 5084 -13486 8950 -13433
rect 9003 -13486 9305 -13433
rect 5031 -13496 5084 -13486
rect 8950 -13496 9003 -13486
rect 9305 -13496 9358 -13486
rect -2004 -13545 -1951 -13535
rect -581 -13545 -528 -13535
rect 2446 -13545 2499 -13535
rect 3870 -13545 3923 -13535
rect 5400 -13545 5453 -13535
rect -1951 -13598 -581 -13545
rect -528 -13598 2446 -13545
rect 2499 -13598 3870 -13545
rect 3923 -13598 5400 -13545
rect 5453 -13556 8828 -13545
rect 9127 -13556 9180 -13546
rect 9483 -13556 9536 -13546
rect 5453 -13598 8772 -13556
rect -2004 -13608 -1951 -13598
rect -581 -13608 -528 -13598
rect 2446 -13608 2499 -13598
rect 3870 -13608 3923 -13598
rect 5400 -13608 5453 -13598
rect 8825 -13609 9127 -13556
rect 9180 -13609 9483 -13556
rect 8772 -13619 8825 -13609
rect 9127 -13619 9180 -13609
rect 9483 -13619 9536 -13609
rect -1648 -13672 -1595 -13662
rect -1291 -13672 -1238 -13662
rect -937 -13672 -884 -13662
rect 1379 -13672 1432 -13662
rect 1732 -13672 1785 -13662
rect 2091 -13672 2144 -13662
rect 5534 -13672 5587 -13662
rect 7526 -13672 7579 -13662
rect 7882 -13672 7935 -13663
rect 8238 -13671 8291 -13661
rect -1595 -13725 -1291 -13672
rect -1238 -13725 -937 -13672
rect -884 -13725 1379 -13672
rect 1432 -13725 1732 -13672
rect 1785 -13725 2091 -13672
rect 2144 -13725 5323 -13672
rect -1648 -13735 -1595 -13725
rect -1291 -13735 -1238 -13725
rect -937 -13735 -884 -13725
rect 1379 -13735 1432 -13725
rect 1732 -13735 1785 -13725
rect 2091 -13735 2144 -13725
rect -6077 -13745 -6024 -13735
rect -5376 -13745 -5323 -13735
rect -5126 -13745 -5073 -13735
rect -4376 -13745 -4323 -13735
rect -6024 -13798 -5376 -13745
rect -5323 -13798 -5126 -13745
rect -5073 -13798 -4376 -13745
rect -6077 -13808 -6024 -13798
rect -5376 -13808 -5323 -13798
rect -5126 -13808 -5073 -13798
rect -4376 -13808 -4323 -13798
rect -225 -13794 -172 -13784
rect 133 -13794 186 -13784
rect 487 -13794 540 -13785
rect 2802 -13794 2855 -13784
rect 3157 -13794 3210 -13785
rect 3512 -13794 3565 -13784
rect 5142 -13794 5195 -13784
rect -6426 -13852 -6373 -13842
rect -5626 -13852 -5573 -13842
rect -4877 -13852 -4824 -13842
rect -4627 -13852 -4574 -13842
rect -3928 -13852 -3875 -13842
rect -6373 -13905 -5626 -13852
rect -5573 -13905 -4877 -13852
rect -4824 -13905 -4627 -13852
rect -4574 -13905 -3928 -13852
rect -172 -13847 133 -13794
rect 186 -13795 2802 -13794
rect 186 -13847 487 -13795
rect -225 -13857 -172 -13847
rect 133 -13857 186 -13847
rect 540 -13847 2802 -13795
rect 2855 -13795 3512 -13794
rect 2855 -13847 3157 -13795
rect 487 -13858 540 -13848
rect 2802 -13857 2855 -13847
rect 3210 -13847 3512 -13795
rect 3565 -13847 5142 -13794
rect 3157 -13858 3210 -13848
rect 3512 -13857 3565 -13847
rect 5142 -13857 5195 -13847
rect 5270 -13796 5323 -13725
rect 5587 -13725 7526 -13672
rect 7579 -13673 8238 -13672
rect 7579 -13725 7882 -13673
rect 5534 -13735 5587 -13725
rect 7526 -13735 7579 -13725
rect 7935 -13724 8238 -13673
rect 11442 -13672 11495 -13662
rect 11798 -13672 11851 -13662
rect 12152 -13672 12205 -13663
rect 12509 -13672 12562 -13662
rect 8291 -13724 11442 -13672
rect 7935 -13725 11442 -13724
rect 11495 -13725 11798 -13672
rect 11851 -13673 12509 -13672
rect 11851 -13725 12152 -13673
rect 7882 -13736 7935 -13726
rect 8238 -13734 8291 -13725
rect 11442 -13735 11495 -13725
rect 11798 -13735 11851 -13725
rect 12205 -13725 12509 -13673
rect 12152 -13736 12205 -13726
rect 12509 -13735 12562 -13725
rect 7348 -13796 7401 -13786
rect 7704 -13795 7757 -13785
rect 5270 -13849 7348 -13796
rect 7401 -13848 7704 -13796
rect 8061 -13796 8114 -13786
rect 8415 -13796 8468 -13786
rect 11264 -13796 11317 -13786
rect 11620 -13796 11673 -13787
rect 11977 -13796 12030 -13786
rect 12334 -13796 12387 -13786
rect 7757 -13848 8061 -13796
rect 7401 -13849 8061 -13848
rect 8114 -13849 8415 -13796
rect 8468 -13849 11264 -13796
rect 11317 -13797 11977 -13796
rect 11317 -13849 11620 -13797
rect 7348 -13859 7401 -13849
rect 7704 -13858 7757 -13849
rect 8061 -13859 8114 -13849
rect 8415 -13859 8468 -13849
rect 11264 -13859 11317 -13849
rect 11673 -13849 11977 -13797
rect 12030 -13849 12334 -13796
rect 11620 -13860 11673 -13850
rect 11977 -13859 12030 -13849
rect 12334 -13859 12387 -13849
rect -6426 -13915 -6373 -13905
rect -5626 -13915 -5573 -13905
rect -4877 -13915 -4824 -13905
rect -4627 -13915 -4574 -13905
rect -3928 -13915 -3875 -13905
rect 5833 -13922 5886 -13912
rect 6013 -13922 6066 -13912
rect 6190 -13922 6243 -13913
rect 6369 -13922 6422 -13912
rect 6547 -13922 6600 -13913
rect 6725 -13922 6778 -13912
rect 6902 -13922 6955 -13912
rect 7437 -13922 7490 -13912
rect 7615 -13922 7668 -13912
rect 7793 -13922 7846 -13913
rect 7970 -13922 8023 -13912
rect 8148 -13922 8201 -13912
rect 8326 -13922 8379 -13912
rect 8861 -13922 8914 -13912
rect 9038 -13922 9091 -13912
rect 9217 -13922 9270 -13912
rect 9394 -13922 9447 -13912
rect 9929 -13922 9982 -13913
rect 10108 -13922 10161 -13912
rect 10284 -13922 10337 -13913
rect 10462 -13922 10515 -13913
rect 10640 -13922 10693 -13912
rect 10819 -13922 10872 -13913
rect 11353 -13922 11406 -13912
rect 11530 -13922 11583 -13912
rect 11709 -13922 11762 -13912
rect 11886 -13922 11939 -13913
rect 12064 -13922 12117 -13912
rect 12242 -13922 12295 -13913
rect 12420 -13922 12473 -13912
rect -5730 -13957 -5677 -13947
rect -4752 -13957 -4699 -13947
rect -3788 -13957 -3735 -13947
rect -5677 -14010 -4752 -13957
rect -4699 -14010 -3788 -13957
rect 5886 -13975 6013 -13922
rect 6066 -13923 6369 -13922
rect 6066 -13975 6190 -13923
rect 5833 -13985 5886 -13975
rect 6013 -13985 6066 -13975
rect 6243 -13975 6369 -13923
rect 6422 -13923 6725 -13922
rect 6422 -13975 6547 -13923
rect 6190 -13986 6243 -13976
rect 6369 -13985 6422 -13975
rect 6600 -13975 6725 -13923
rect 6778 -13975 6902 -13922
rect 6955 -13975 7437 -13922
rect 7490 -13975 7615 -13922
rect 7668 -13923 7970 -13922
rect 7668 -13975 7793 -13923
rect 6547 -13986 6600 -13976
rect 6725 -13985 6778 -13975
rect 6902 -13985 6955 -13975
rect 7437 -13985 7490 -13975
rect 7615 -13985 7668 -13975
rect 7846 -13975 7970 -13923
rect 8023 -13975 8148 -13922
rect 8201 -13975 8326 -13922
rect 8379 -13975 8861 -13922
rect 8914 -13975 9038 -13922
rect 9091 -13975 9217 -13922
rect 9270 -13975 9394 -13922
rect 9447 -13923 10108 -13922
rect 9447 -13975 9929 -13923
rect 7793 -13986 7846 -13976
rect 7970 -13985 8023 -13975
rect 8148 -13985 8201 -13975
rect 8326 -13985 8379 -13975
rect 8861 -13985 8914 -13975
rect 9038 -13985 9091 -13975
rect 9217 -13985 9270 -13975
rect 9394 -13985 9447 -13975
rect 9982 -13975 10108 -13923
rect 10161 -13923 10640 -13922
rect 10161 -13975 10284 -13923
rect 9929 -13986 9982 -13976
rect 10108 -13985 10161 -13975
rect 10337 -13975 10462 -13923
rect 10284 -13986 10337 -13976
rect 10515 -13975 10640 -13923
rect 10693 -13923 11353 -13922
rect 10693 -13975 10819 -13923
rect 10462 -13986 10515 -13976
rect 10640 -13985 10693 -13975
rect 10872 -13975 11353 -13923
rect 11406 -13975 11530 -13922
rect 11583 -13975 11709 -13922
rect 11762 -13923 12064 -13922
rect 11762 -13975 11886 -13923
rect 10819 -13986 10872 -13976
rect 11353 -13985 11406 -13975
rect 11530 -13985 11583 -13975
rect 11709 -13985 11762 -13975
rect 11939 -13975 12064 -13923
rect 12117 -13923 12420 -13922
rect 12117 -13975 12242 -13923
rect 11886 -13986 11939 -13976
rect 12064 -13985 12117 -13975
rect 12295 -13975 12420 -13923
rect 12242 -13986 12295 -13976
rect 12420 -13985 12473 -13975
rect -5730 -14020 -5677 -14010
rect -4752 -14020 -4699 -14010
rect -3788 -14020 -3735 -14010
rect -6223 -14055 -6170 -14045
rect -5250 -14055 -5197 -14045
rect -4250 -14055 -4197 -14045
rect -3382 -14055 -3329 -14045
rect -6170 -14108 -5250 -14055
rect -5197 -14108 -4250 -14055
rect -4197 -14108 -3382 -14055
rect -6223 -14118 -6170 -14108
rect -5250 -14118 -5197 -14108
rect -4250 -14118 -4197 -14108
rect -3382 -14118 -3329 -14108
rect -2315 -14543 -2262 -14533
rect -1381 -14543 -1328 -14533
rect -1204 -14543 -1151 -14533
rect -1026 -14543 -973 -14533
rect -848 -14543 -795 -14533
rect -669 -14543 -616 -14533
rect -491 -14543 -438 -14533
rect 1288 -14543 1341 -14533
rect 1466 -14543 1519 -14533
rect 1644 -14543 1697 -14533
rect 1823 -14542 1876 -14532
rect -2262 -14596 -1381 -14543
rect -1328 -14596 -1204 -14543
rect -1151 -14596 -1026 -14543
rect -973 -14596 -848 -14543
rect -795 -14596 -669 -14543
rect -616 -14596 -491 -14543
rect -438 -14596 1288 -14543
rect 1341 -14596 1466 -14543
rect 1519 -14596 1644 -14543
rect 1697 -14595 1823 -14543
rect 2000 -14543 2053 -14533
rect 2178 -14543 2231 -14533
rect 3246 -14543 3299 -14534
rect 3424 -14543 3477 -14533
rect 3602 -14543 3655 -14533
rect 3781 -14543 3834 -14533
rect 1876 -14595 2000 -14543
rect 1697 -14596 2000 -14595
rect 2053 -14596 2178 -14543
rect 2231 -14544 3424 -14543
rect 2231 -14596 3246 -14544
rect -2315 -14606 -2262 -14596
rect -1381 -14606 -1328 -14596
rect -1204 -14606 -1151 -14596
rect -1026 -14606 -973 -14596
rect -848 -14606 -795 -14596
rect -669 -14606 -616 -14596
rect -491 -14606 -438 -14596
rect 1288 -14606 1341 -14596
rect 1466 -14606 1519 -14596
rect 1644 -14606 1697 -14596
rect 1823 -14605 1876 -14596
rect 2000 -14606 2053 -14596
rect 2178 -14606 2231 -14596
rect 3299 -14596 3424 -14544
rect 3477 -14596 3602 -14543
rect 3655 -14596 3781 -14543
rect 3246 -14607 3299 -14597
rect 3424 -14606 3477 -14596
rect 3602 -14606 3655 -14596
rect 3781 -14606 3834 -14596
rect 4905 -14545 4958 -14535
rect 5746 -14545 5799 -14535
rect 6101 -14545 6154 -14535
rect 6459 -14545 6512 -14535
rect 6813 -14545 6866 -14535
rect 8236 -14545 8289 -14535
rect 8595 -14545 8648 -14535
rect 8950 -14545 9003 -14536
rect 9304 -14545 9357 -14535
rect 9661 -14545 9714 -14535
rect 10016 -14545 10069 -14535
rect 10373 -14545 10426 -14536
rect 10729 -14545 10782 -14535
rect 4958 -14598 5746 -14545
rect 5799 -14598 6101 -14545
rect 6154 -14598 6459 -14545
rect 6512 -14598 6813 -14545
rect 6866 -14598 8236 -14545
rect 8289 -14598 8595 -14545
rect 8648 -14546 9304 -14545
rect 8648 -14598 8950 -14546
rect 4905 -14608 4958 -14598
rect 5746 -14608 5799 -14598
rect 6101 -14608 6154 -14598
rect 6459 -14608 6512 -14598
rect 6813 -14608 6866 -14598
rect 8236 -14608 8289 -14598
rect 8595 -14608 8648 -14598
rect 9003 -14598 9304 -14546
rect 9357 -14598 9661 -14545
rect 9714 -14598 10016 -14545
rect 10069 -14546 10729 -14545
rect 10069 -14598 10373 -14546
rect 8950 -14609 9003 -14599
rect 9304 -14608 9357 -14598
rect 9661 -14608 9714 -14598
rect 10016 -14608 10069 -14598
rect 10426 -14598 10729 -14546
rect 10373 -14609 10426 -14599
rect 10729 -14608 10782 -14598
rect 5143 -14658 5196 -14648
rect 5924 -14658 5977 -14648
rect 6279 -14658 6332 -14648
rect 6636 -14658 6689 -14648
rect 6991 -14658 7044 -14648
rect 8417 -14657 8470 -14647
rect 5196 -14711 5924 -14658
rect 5977 -14711 6279 -14658
rect 6332 -14711 6636 -14658
rect 6689 -14711 6991 -14658
rect 7044 -14710 8417 -14658
rect 8772 -14658 8825 -14648
rect 9127 -14658 9180 -14649
rect 9483 -14658 9536 -14648
rect 9837 -14658 9890 -14649
rect 10196 -14658 10249 -14648
rect 10550 -14658 10603 -14648
rect 10908 -14658 10961 -14648
rect 8470 -14710 8772 -14658
rect 7044 -14711 8772 -14710
rect 8825 -14659 9483 -14658
rect 8825 -14711 9127 -14659
rect 5143 -14721 5196 -14711
rect 5924 -14721 5977 -14711
rect 6279 -14721 6332 -14711
rect 6636 -14721 6689 -14711
rect 6991 -14721 7044 -14711
rect 8417 -14720 8470 -14711
rect 8772 -14721 8825 -14711
rect 9180 -14711 9483 -14659
rect 9536 -14659 10196 -14658
rect 9536 -14711 9837 -14659
rect 9127 -14722 9180 -14712
rect 9483 -14721 9536 -14711
rect 9890 -14711 10196 -14659
rect 10249 -14711 10550 -14658
rect 10603 -14711 10908 -14658
rect 9837 -14722 9890 -14712
rect 10196 -14721 10249 -14711
rect 10550 -14721 10603 -14711
rect 10908 -14721 10961 -14711
rect 11087 -14656 11140 -14648
rect 11440 -14656 11493 -14646
rect 11087 -14658 11440 -14656
rect 11140 -14708 11440 -14658
rect 11140 -14709 11192 -14708
rect 11087 -14721 11140 -14711
rect 11440 -14719 11493 -14709
rect -6159 -14795 -6106 -14785
rect -5860 -14795 -5807 -14785
rect -5147 -14795 -5094 -14785
rect -4436 -14795 -4383 -14785
rect -6106 -14848 -5860 -14795
rect -5807 -14848 -5147 -14795
rect -5094 -14848 -4436 -14795
rect 8504 -14806 8557 -14796
rect -6159 -14858 -6106 -14848
rect -5860 -14858 -5807 -14848
rect -5147 -14858 -5094 -14848
rect -4436 -14858 -4383 -14848
rect 6993 -14824 7046 -14814
rect 7347 -14824 7400 -14814
rect 7704 -14824 7757 -14815
rect 7046 -14877 7347 -14824
rect 7400 -14825 7757 -14824
rect 7400 -14877 7704 -14825
rect 6993 -14887 7046 -14877
rect 7347 -14887 7400 -14877
rect 7704 -14888 7757 -14878
rect 8060 -14821 8113 -14811
rect 8113 -14859 8504 -14821
rect 9753 -14806 9806 -14796
rect 8557 -14859 9753 -14821
rect 10195 -14821 10248 -14812
rect 9806 -14822 10248 -14821
rect 9806 -14859 10195 -14822
rect 8113 -14874 10195 -14859
rect 8060 -14884 8113 -14874
rect 10195 -14885 10248 -14875
rect 10552 -14814 10605 -14805
rect 10908 -14813 10961 -14803
rect 10552 -14815 10908 -14814
rect 10605 -14866 10908 -14815
rect 10961 -14814 11013 -14813
rect 11264 -14814 11317 -14805
rect 10961 -14815 11317 -14814
rect 10961 -14866 11264 -14815
rect 10552 -14878 10605 -14868
rect 10908 -14876 10961 -14866
rect 11264 -14878 11317 -14868
rect -5504 -14901 -5451 -14891
rect -4791 -14901 -4738 -14891
rect -3936 -14901 -3883 -14891
rect -5451 -14954 -4791 -14901
rect -4738 -14954 -3936 -14901
rect -5504 -14964 -5451 -14954
rect -4791 -14964 -4738 -14954
rect -3936 -14964 -3883 -14954
rect -847 -14926 -794 -14916
rect -669 -14926 -616 -14916
rect -491 -14926 -438 -14916
rect -314 -14926 -261 -14917
rect -137 -14926 -84 -14916
rect 43 -14926 96 -14916
rect 1289 -14926 1342 -14917
rect 1467 -14926 1520 -14916
rect 1644 -14926 1697 -14916
rect 1822 -14926 1875 -14916
rect 1999 -14926 2052 -14916
rect 2180 -14926 2233 -14916
rect 3425 -14926 3478 -14916
rect 3603 -14926 3656 -14916
rect 3780 -14926 3833 -14916
rect 4239 -14926 4292 -14916
rect -794 -14979 -669 -14926
rect -616 -14979 -491 -14926
rect -438 -14927 -137 -14926
rect -438 -14979 -314 -14927
rect -847 -14989 -794 -14979
rect -669 -14989 -616 -14979
rect -491 -14989 -438 -14979
rect -261 -14979 -137 -14927
rect -84 -14979 43 -14926
rect 96 -14927 1467 -14926
rect 96 -14979 1289 -14927
rect -314 -14990 -261 -14980
rect -137 -14989 -84 -14979
rect 43 -14989 96 -14979
rect 1342 -14979 1467 -14927
rect 1520 -14979 1644 -14926
rect 1697 -14979 1822 -14926
rect 1875 -14979 1999 -14926
rect 2052 -14979 2180 -14926
rect 2233 -14979 3425 -14926
rect 3478 -14979 3603 -14926
rect 3656 -14979 3780 -14926
rect 3833 -14979 4239 -14926
rect 1289 -14990 1342 -14980
rect 1467 -14989 1520 -14979
rect 1644 -14989 1697 -14979
rect 1822 -14989 1875 -14979
rect 1999 -14989 2052 -14979
rect 2180 -14989 2233 -14979
rect 3425 -14989 3478 -14979
rect 3603 -14989 3656 -14979
rect 3780 -14989 3833 -14979
rect 4239 -14989 4292 -14979
rect 7080 -14923 7133 -14913
rect 7260 -14923 7313 -14914
rect 7439 -14923 7492 -14913
rect 8327 -14923 8380 -14913
rect 8505 -14923 8558 -14914
rect 8683 -14923 8736 -14914
rect 9572 -14923 9625 -14913
rect 9750 -14923 9803 -14913
rect 9929 -14923 9982 -14913
rect 10819 -14923 10872 -14913
rect 10996 -14923 11049 -14913
rect 11175 -14923 11228 -14913
rect 7133 -14924 7439 -14923
rect 7133 -14976 7260 -14924
rect 7080 -14986 7133 -14976
rect 7313 -14976 7439 -14924
rect 7492 -14976 8327 -14923
rect 8380 -14924 9572 -14923
rect 8380 -14976 8505 -14924
rect 7260 -14987 7313 -14977
rect 7439 -14986 7492 -14976
rect 8327 -14986 8380 -14976
rect 8558 -14976 8683 -14924
rect 8505 -14987 8558 -14977
rect 8736 -14976 9572 -14924
rect 9625 -14976 9750 -14923
rect 9803 -14976 9929 -14923
rect 9982 -14976 10819 -14923
rect 10872 -14976 10996 -14923
rect 11049 -14976 11175 -14923
rect 8683 -14987 8736 -14977
rect 9572 -14986 9625 -14976
rect 9750 -14986 9803 -14976
rect 9929 -14986 9982 -14976
rect 10819 -14986 10872 -14976
rect 10996 -14986 11049 -14976
rect 11175 -14986 11228 -14976
rect -6159 -15481 -6106 -15472
rect -5504 -15481 -5451 -15471
rect -4792 -15481 -4739 -15471
rect -6159 -15482 -5504 -15481
rect -6106 -15534 -5504 -15482
rect -5451 -15534 -4792 -15481
rect -6159 -15545 -6106 -15535
rect -5504 -15544 -5451 -15534
rect -4792 -15544 -4739 -15534
rect 4238 -15539 4291 -15529
rect 5031 -15539 5084 -15530
rect 5745 -15539 5798 -15529
rect 6101 -15539 6154 -15529
rect 6458 -15539 6511 -15529
rect 11798 -15539 11851 -15530
rect 12155 -15539 12208 -15529
rect 12511 -15539 12564 -15529
rect -5860 -15588 -5807 -15578
rect -5148 -15589 -5095 -15579
rect -4435 -15589 -4383 -15579
rect -3935 -15589 -3883 -15579
rect -5807 -15641 -5148 -15589
rect -5860 -15651 -5807 -15641
rect -5095 -15641 -4435 -15589
rect -4383 -15641 -3935 -15589
rect 4291 -15540 5745 -15539
rect 4291 -15592 5031 -15540
rect 4238 -15602 4291 -15592
rect 5084 -15592 5745 -15540
rect 5798 -15592 6101 -15539
rect 6154 -15592 6458 -15539
rect 6511 -15540 12155 -15539
rect 6511 -15592 11798 -15540
rect 5031 -15603 5084 -15593
rect 5745 -15602 5798 -15592
rect 6101 -15602 6154 -15592
rect 6458 -15602 6511 -15592
rect 11851 -15592 12155 -15540
rect 12208 -15592 12511 -15539
rect 11798 -15603 11851 -15593
rect 12155 -15602 12208 -15592
rect 12511 -15602 12564 -15592
rect -5148 -15652 -5095 -15642
rect -4435 -15651 -4383 -15641
rect -3935 -15651 -3883 -15641
rect 5400 -15652 5453 -15643
rect 5923 -15652 5976 -15642
rect 6279 -15652 6332 -15642
rect 6635 -15652 6688 -15642
rect 11619 -15652 11672 -15642
rect 11975 -15652 12028 -15642
rect 12332 -15652 12385 -15642
rect 5400 -15653 5923 -15652
rect 5453 -15705 5923 -15653
rect 5976 -15705 6279 -15652
rect 6332 -15705 6635 -15652
rect 6688 -15705 11619 -15652
rect 11672 -15705 11975 -15652
rect 12028 -15705 12332 -15652
rect 5400 -15716 5453 -15706
rect 5923 -15715 5976 -15705
rect 6279 -15715 6332 -15705
rect 6635 -15715 6688 -15705
rect 11619 -15715 11672 -15705
rect 11975 -15715 12028 -15705
rect 12332 -15715 12385 -15705
rect 5747 -15750 5800 -15740
rect 6101 -15749 6154 -15739
rect 5800 -15802 6101 -15750
rect 6456 -15750 6509 -15740
rect 6713 -15750 6766 -15741
rect 7169 -15750 7222 -15740
rect 7526 -15749 7579 -15739
rect 6154 -15802 6456 -15750
rect 5800 -15803 6456 -15802
rect 6509 -15751 7169 -15750
rect 6509 -15803 6713 -15751
rect -2447 -15821 -2394 -15811
rect -2005 -15821 -1952 -15812
rect -2394 -15822 -1952 -15821
rect -1649 -15822 -1596 -15812
rect -1293 -15822 -1240 -15812
rect -937 -15822 -884 -15812
rect -581 -15822 -528 -15812
rect -225 -15822 -172 -15812
rect 132 -15821 185 -15811
rect -2394 -15874 -2005 -15822
rect -2447 -15884 -2394 -15874
rect -1952 -15875 -1649 -15822
rect -1596 -15875 -1293 -15822
rect -1240 -15875 -937 -15822
rect -884 -15875 -581 -15822
rect -528 -15875 -225 -15822
rect -172 -15874 132 -15822
rect 487 -15822 540 -15812
rect 843 -15822 896 -15812
rect 1201 -15822 1254 -15812
rect 1555 -15822 1608 -15812
rect 1910 -15822 1963 -15812
rect 2267 -15822 2320 -15812
rect 2624 -15822 2677 -15812
rect 2979 -15822 3032 -15812
rect 3335 -15822 3388 -15812
rect 3692 -15822 3745 -15812
rect 5747 -15813 5800 -15803
rect 6101 -15812 6154 -15803
rect 6456 -15813 6509 -15803
rect 6766 -15803 7169 -15751
rect 7222 -15802 7526 -15750
rect 7882 -15749 7935 -15739
rect 7579 -15802 7882 -15750
rect 10373 -15750 10426 -15741
rect 10730 -15750 10783 -15740
rect 11086 -15750 11139 -15740
rect 7935 -15751 10730 -15750
rect 7935 -15802 10373 -15751
rect 7222 -15803 10373 -15802
rect 6713 -15814 6766 -15804
rect 7169 -15813 7222 -15803
rect 7526 -15812 7579 -15803
rect 7882 -15812 7935 -15803
rect 10426 -15803 10730 -15751
rect 10783 -15803 11086 -15750
rect 10373 -15814 10426 -15804
rect 10730 -15813 10783 -15803
rect 11086 -15813 11139 -15803
rect 185 -15874 487 -15822
rect -172 -15875 487 -15874
rect 540 -15875 843 -15822
rect 896 -15875 1201 -15822
rect 1254 -15875 1555 -15822
rect 1608 -15875 1910 -15822
rect 1963 -15875 2267 -15822
rect 2320 -15875 2624 -15822
rect 2677 -15875 2979 -15822
rect 3032 -15875 3335 -15822
rect 3388 -15875 3692 -15822
rect 11440 -15841 11493 -15831
rect -2005 -15885 -1952 -15875
rect -1649 -15885 -1596 -15875
rect -1293 -15885 -1240 -15875
rect -937 -15885 -884 -15875
rect -581 -15885 -528 -15875
rect -225 -15885 -172 -15875
rect 132 -15884 185 -15875
rect 487 -15885 540 -15875
rect 843 -15885 896 -15875
rect 1201 -15885 1254 -15875
rect 1555 -15885 1608 -15875
rect 1910 -15885 1963 -15875
rect 2267 -15885 2320 -15875
rect 2624 -15885 2677 -15875
rect 2979 -15885 3032 -15875
rect 3335 -15885 3388 -15875
rect 3692 -15885 3745 -15875
rect 6813 -15851 6866 -15841
rect 7169 -15851 7222 -15842
rect 8060 -15851 8113 -15841
rect 8593 -15851 8646 -15842
rect 9663 -15851 9716 -15842
rect 10194 -15851 10247 -15842
rect 11084 -15851 11137 -15842
rect 6866 -15852 8060 -15851
rect 6866 -15904 7169 -15852
rect 6813 -15914 6866 -15904
rect 7222 -15904 8060 -15852
rect 8113 -15852 11440 -15851
rect 8113 -15904 8593 -15852
rect 7169 -15915 7222 -15905
rect 8060 -15914 8113 -15904
rect 8646 -15904 9663 -15852
rect 8593 -15915 8646 -15905
rect 9716 -15904 10194 -15852
rect 9663 -15915 9716 -15905
rect 10247 -15904 11084 -15852
rect 10194 -15915 10247 -15905
rect 11137 -15894 11440 -15852
rect 11137 -15904 11493 -15894
rect 11084 -15915 11137 -15905
rect -1915 -15933 -1862 -15923
rect -1738 -15933 -1685 -15923
rect -1560 -15933 -1507 -15923
rect -1382 -15933 -1329 -15923
rect -1204 -15933 -1151 -15923
rect -1025 -15933 -972 -15923
rect -847 -15933 -794 -15923
rect -670 -15933 -617 -15923
rect -491 -15933 -438 -15923
rect -313 -15933 -260 -15923
rect -136 -15933 -83 -15923
rect 43 -15933 96 -15923
rect 221 -15933 274 -15923
rect 398 -15933 451 -15923
rect 575 -15933 628 -15923
rect 755 -15933 808 -15923
rect 931 -15933 984 -15923
rect 1110 -15933 1163 -15923
rect 1289 -15933 1342 -15923
rect 1466 -15933 1519 -15923
rect 1643 -15933 1696 -15923
rect 1822 -15933 1875 -15923
rect 2000 -15933 2053 -15923
rect 2179 -15933 2232 -15923
rect 2356 -15933 2409 -15923
rect 2534 -15933 2587 -15923
rect 2712 -15933 2765 -15923
rect 2891 -15933 2944 -15923
rect 3068 -15933 3121 -15923
rect 3247 -15933 3300 -15923
rect 3424 -15933 3477 -15923
rect 3603 -15933 3656 -15923
rect 3780 -15933 3833 -15923
rect -1862 -15986 -1738 -15933
rect -1685 -15986 -1560 -15933
rect -1507 -15986 -1382 -15933
rect -1329 -15986 -1204 -15933
rect -1151 -15986 -1025 -15933
rect -972 -15986 -847 -15933
rect -794 -15986 -670 -15933
rect -617 -15986 -491 -15933
rect -438 -15986 -313 -15933
rect -260 -15986 -136 -15933
rect -83 -15986 43 -15933
rect 96 -15986 221 -15933
rect 274 -15986 398 -15933
rect 451 -15986 575 -15933
rect 628 -15986 755 -15933
rect 808 -15986 931 -15933
rect 984 -15986 1110 -15933
rect 1163 -15986 1289 -15933
rect 1342 -15986 1466 -15933
rect 1519 -15986 1643 -15933
rect 1696 -15986 1822 -15933
rect 1875 -15986 2000 -15933
rect 2053 -15986 2179 -15933
rect 2232 -15986 2356 -15933
rect 2409 -15986 2534 -15933
rect 2587 -15986 2712 -15933
rect 2765 -15986 2891 -15933
rect 2944 -15986 3068 -15933
rect 3121 -15986 3247 -15933
rect 3300 -15986 3424 -15933
rect 3477 -15986 3603 -15933
rect 3656 -15986 3780 -15933
rect -1915 -15996 -1862 -15986
rect -1738 -15996 -1685 -15986
rect -1560 -15996 -1507 -15986
rect -1382 -15996 -1329 -15986
rect -1204 -15996 -1151 -15986
rect -1025 -15996 -972 -15986
rect -847 -15996 -794 -15986
rect -670 -15996 -617 -15986
rect -491 -15996 -438 -15986
rect -313 -15996 -260 -15986
rect -136 -15996 -83 -15986
rect 43 -15996 96 -15986
rect 221 -15996 274 -15986
rect 398 -15996 451 -15986
rect 575 -15996 628 -15986
rect 755 -15996 808 -15986
rect 931 -15996 984 -15986
rect 1110 -15996 1163 -15986
rect 1289 -15996 1342 -15986
rect 1466 -15996 1519 -15986
rect 1643 -15996 1696 -15986
rect 1822 -15996 1875 -15986
rect 2000 -15996 2053 -15986
rect 2179 -15996 2232 -15986
rect 2356 -15996 2409 -15986
rect 2534 -15996 2587 -15986
rect 2712 -15996 2765 -15986
rect 2891 -15996 2944 -15986
rect 3068 -15996 3121 -15986
rect 3247 -15996 3300 -15986
rect 3424 -15996 3477 -15986
rect 3603 -15996 3656 -15986
rect 3780 -15996 3833 -15986
rect 5921 -15947 5974 -15938
rect 6279 -15947 6332 -15938
rect 6634 -15947 6687 -15938
rect 6994 -15947 7047 -15941
rect 5921 -15948 7047 -15947
rect 5974 -16000 6279 -15948
rect 5921 -16011 5974 -16001
rect 6332 -16000 6634 -15948
rect 6279 -16011 6332 -16001
rect 6687 -15951 7047 -15948
rect 6687 -16000 6994 -15951
rect 6634 -16011 6687 -16001
rect 6994 -16014 7047 -16004
rect 7526 -15952 7579 -15943
rect 7881 -15952 7934 -15942
rect 8237 -15952 8290 -15942
rect 11441 -15952 11494 -15942
rect 11797 -15952 11850 -15942
rect 12154 -15952 12207 -15942
rect 12511 -15952 12564 -15942
rect 7526 -15953 7881 -15952
rect 7579 -16005 7881 -15953
rect 7934 -16005 8237 -15952
rect 8290 -16005 11441 -15952
rect 11494 -16005 11797 -15952
rect 11850 -16005 12154 -15952
rect 12207 -16005 12511 -15952
rect 7526 -16016 7579 -16006
rect 7881 -16015 7934 -16005
rect 8237 -16015 8290 -16005
rect 11441 -16015 11494 -16005
rect 11797 -16015 11850 -16005
rect 12154 -16015 12207 -16005
rect 12511 -16015 12564 -16005
rect -6159 -16193 -6106 -16183
rect -5504 -16193 -5451 -16183
rect -4792 -16193 -4739 -16183
rect -6106 -16246 -5504 -16193
rect -5451 -16246 -4792 -16193
rect -6159 -16256 -6106 -16246
rect -5504 -16256 -5451 -16246
rect -4792 -16256 -4739 -16246
rect -5860 -16294 -5807 -16284
rect -5148 -16294 -5095 -16284
rect -4436 -16294 -4383 -16284
rect -3935 -16294 -3883 -16285
rect -5807 -16347 -5148 -16294
rect -5095 -16346 -4436 -16294
rect -5860 -16357 -5807 -16347
rect -5148 -16357 -5095 -16347
rect -4383 -16295 -3883 -16294
rect -4383 -16346 -3935 -16295
rect -4436 -16357 -4383 -16347
rect -3935 -16357 -3883 -16347
rect -1917 -16542 -1864 -16532
rect -1738 -16542 -1685 -16532
rect -1561 -16541 -1508 -16531
rect -1864 -16595 -1738 -16542
rect -1685 -16594 -1561 -16542
rect -1381 -16542 -1328 -16533
rect -1204 -16542 -1151 -16532
rect -1026 -16542 -973 -16532
rect 220 -16542 273 -16532
rect 397 -16542 450 -16532
rect 576 -16542 629 -16532
rect 755 -16542 808 -16532
rect 933 -16542 986 -16532
rect 1111 -16542 1164 -16532
rect 2356 -16542 2409 -16532
rect 2534 -16542 2587 -16532
rect 2713 -16541 2766 -16531
rect -1508 -16543 -1204 -16542
rect -1508 -16594 -1381 -16543
rect -1685 -16595 -1381 -16594
rect -1917 -16605 -1864 -16595
rect -1738 -16605 -1685 -16595
rect -1561 -16604 -1508 -16595
rect -1328 -16595 -1204 -16543
rect -1151 -16595 -1026 -16542
rect -973 -16595 220 -16542
rect 273 -16595 397 -16542
rect 450 -16595 576 -16542
rect 629 -16595 755 -16542
rect 808 -16595 933 -16542
rect 986 -16595 1111 -16542
rect 1164 -16595 2356 -16542
rect 2409 -16595 2534 -16542
rect 2587 -16594 2713 -16542
rect 2891 -16542 2944 -16532
rect 3070 -16542 3123 -16532
rect 3249 -16542 3302 -16532
rect 4238 -16542 4291 -16532
rect 2766 -16594 2891 -16542
rect 2587 -16595 2891 -16594
rect 2944 -16595 3070 -16542
rect 3123 -16595 3249 -16542
rect 3302 -16595 4238 -16542
rect -1381 -16606 -1328 -16596
rect -1204 -16605 -1151 -16595
rect -1026 -16605 -973 -16595
rect 220 -16605 273 -16595
rect 397 -16605 450 -16595
rect 576 -16605 629 -16595
rect 755 -16605 808 -16595
rect 933 -16605 986 -16595
rect 1111 -16605 1164 -16595
rect 2356 -16605 2409 -16595
rect 2534 -16605 2587 -16595
rect 2713 -16604 2766 -16595
rect 2891 -16605 2944 -16595
rect 3070 -16605 3123 -16595
rect 3249 -16605 3302 -16595
rect 4238 -16605 4291 -16595
rect 6548 -16544 6601 -16534
rect 6726 -16544 6779 -16534
rect 6601 -16597 6726 -16545
rect 6903 -16545 6956 -16535
rect 7970 -16545 8023 -16535
rect 8149 -16544 8202 -16534
rect 6779 -16597 6903 -16545
rect 6548 -16598 6903 -16597
rect 6956 -16598 7970 -16545
rect 8023 -16597 8149 -16545
rect 9929 -16544 9982 -16534
rect 8202 -16597 9929 -16545
rect 10107 -16545 10160 -16535
rect 10287 -16545 10340 -16535
rect 11352 -16545 11405 -16535
rect 11530 -16545 11583 -16536
rect 11709 -16545 11762 -16535
rect 9982 -16597 10107 -16545
rect 8023 -16598 10107 -16597
rect 10160 -16598 10287 -16545
rect 10340 -16598 11352 -16545
rect 11405 -16546 11709 -16545
rect 11405 -16598 11530 -16546
rect 6548 -16607 6601 -16598
rect 6726 -16607 6779 -16598
rect 6903 -16608 6956 -16598
rect 7970 -16608 8023 -16598
rect 8149 -16607 8202 -16598
rect 9929 -16607 9982 -16598
rect 10107 -16608 10160 -16598
rect 10287 -16608 10340 -16598
rect 11352 -16608 11405 -16598
rect 11583 -16598 11709 -16546
rect 11530 -16609 11583 -16599
rect 11709 -16608 11762 -16598
rect -1827 -16665 -1774 -16655
rect -1471 -16665 -1418 -16656
rect -1114 -16665 -1061 -16655
rect -759 -16664 -706 -16654
rect -1774 -16666 -1114 -16665
rect -1774 -16718 -1471 -16666
rect -1827 -16728 -1774 -16718
rect -1418 -16718 -1114 -16666
rect -1061 -16717 -759 -16665
rect -403 -16665 -350 -16655
rect -47 -16665 6 -16655
rect 309 -16665 362 -16656
rect 665 -16665 718 -16655
rect 845 -16665 898 -16655
rect 1021 -16665 1074 -16655
rect 1377 -16665 1430 -16655
rect 1735 -16665 1788 -16655
rect 2090 -16664 2143 -16654
rect -706 -16717 -403 -16665
rect -1061 -16718 -403 -16717
rect -350 -16718 -47 -16665
rect 6 -16666 665 -16665
rect 6 -16718 309 -16666
rect -1471 -16729 -1418 -16719
rect -1114 -16728 -1061 -16718
rect -759 -16727 -706 -16718
rect -403 -16728 -350 -16718
rect -47 -16728 6 -16718
rect 362 -16718 665 -16666
rect 718 -16718 845 -16665
rect 898 -16718 1021 -16665
rect 1074 -16718 1377 -16665
rect 1430 -16718 1735 -16665
rect 1788 -16717 2090 -16665
rect 2445 -16665 2498 -16655
rect 2801 -16665 2854 -16655
rect 3157 -16664 3210 -16654
rect 2143 -16717 2445 -16665
rect 1788 -16718 2445 -16717
rect 2498 -16718 2801 -16665
rect 2854 -16717 3157 -16665
rect 3514 -16665 3567 -16656
rect 3868 -16665 3921 -16655
rect 3210 -16666 3868 -16665
rect 3210 -16717 3514 -16666
rect 2854 -16718 3514 -16717
rect 309 -16729 362 -16719
rect 665 -16728 718 -16718
rect 845 -16728 898 -16718
rect 1021 -16728 1074 -16718
rect 1377 -16728 1430 -16718
rect 1735 -16728 1788 -16718
rect 2090 -16727 2143 -16718
rect 2445 -16728 2498 -16718
rect 2801 -16728 2854 -16718
rect 3157 -16727 3210 -16718
rect 3567 -16718 3868 -16666
rect 3514 -16729 3567 -16719
rect 3868 -16728 3921 -16718
rect 5399 -16666 5452 -16657
rect 8771 -16666 8824 -16656
rect 9128 -16666 9181 -16656
rect 9484 -16666 9537 -16656
rect 5399 -16667 8771 -16666
rect 5452 -16719 8771 -16667
rect 8824 -16719 9128 -16666
rect 9181 -16719 9484 -16666
rect 5399 -16730 5452 -16720
rect 8771 -16729 8824 -16719
rect 9128 -16729 9181 -16719
rect 9484 -16729 9537 -16719
rect 9838 -16665 9891 -16656
rect 10195 -16665 10248 -16655
rect 10550 -16665 10603 -16655
rect 10907 -16665 10960 -16655
rect 9838 -16666 10195 -16665
rect 9891 -16718 10195 -16666
rect 10248 -16718 10550 -16665
rect 10603 -16718 10907 -16665
rect 9838 -16729 9891 -16719
rect 10195 -16728 10248 -16718
rect 10550 -16728 10603 -16718
rect 10907 -16728 10960 -16718
rect 5031 -16782 5084 -16772
rect 8950 -16782 9003 -16772
rect 9305 -16782 9358 -16772
rect 5084 -16835 8950 -16782
rect 9003 -16835 9305 -16782
rect 5031 -16845 5084 -16835
rect 8950 -16845 9003 -16835
rect 9305 -16845 9358 -16835
rect 10017 -16780 10070 -16771
rect 10374 -16780 10427 -16771
rect 10731 -16779 10784 -16769
rect 10017 -16781 10731 -16780
rect 10070 -16833 10374 -16781
rect 10017 -16844 10070 -16834
rect 10427 -16832 10731 -16781
rect 10427 -16833 10784 -16832
rect 10374 -16844 10427 -16834
rect 10731 -16842 10784 -16833
rect -5682 -16886 -5629 -16876
rect -5326 -16886 -5273 -16876
rect -4970 -16886 -4917 -16876
rect -4614 -16886 -4561 -16876
rect -4258 -16886 -4205 -16876
rect -5629 -16939 -5326 -16886
rect -5273 -16939 -4970 -16886
rect -4917 -16939 -4614 -16886
rect -4561 -16939 -4258 -16886
rect -5682 -16949 -5629 -16939
rect -5326 -16949 -5273 -16939
rect -4970 -16949 -4917 -16939
rect -4614 -16949 -4561 -16939
rect -4258 -16949 -4205 -16939
rect 7347 -16890 7400 -16880
rect 7704 -16890 7757 -16880
rect 8060 -16890 8113 -16880
rect 8416 -16890 8469 -16880
rect 11263 -16890 11316 -16880
rect 11620 -16890 11673 -16880
rect 11975 -16889 12028 -16879
rect 7400 -16943 7704 -16890
rect 7757 -16943 8060 -16890
rect 8113 -16943 8416 -16890
rect 8469 -16943 11263 -16890
rect 11316 -16943 11620 -16890
rect 11673 -16942 11975 -16890
rect 12331 -16889 12384 -16879
rect 12028 -16942 12331 -16890
rect 11673 -16943 12384 -16942
rect 7347 -16953 7400 -16943
rect 7704 -16953 7757 -16943
rect 8060 -16953 8113 -16943
rect 8416 -16953 8469 -16943
rect 11263 -16953 11316 -16943
rect 11620 -16953 11673 -16943
rect 11975 -16952 12028 -16943
rect 12331 -16952 12384 -16943
rect -6159 -17007 -6106 -16997
rect -5859 -17007 -5806 -16997
rect -5148 -17007 -5095 -16997
rect -4437 -17007 -4384 -16997
rect -6106 -17060 -5859 -17007
rect -5806 -17060 -5148 -17007
rect -5095 -17060 -4437 -17007
rect -6159 -17070 -6106 -17060
rect -5859 -17070 -5806 -17060
rect -5148 -17070 -5095 -17060
rect -4437 -17070 -4384 -17060
rect -5504 -17118 -5451 -17108
rect -4792 -17118 -4739 -17108
rect -3935 -17118 -3883 -17108
rect -5451 -17170 -4792 -17118
rect -5504 -17181 -5451 -17171
rect -4739 -17170 -3935 -17118
rect -4792 -17181 -4739 -17171
rect -3935 -17180 -3883 -17170
<< via2 >>
rect 3019 -3513 3080 -3452
rect -2546 -3989 -2485 -3928
rect 2538 -4327 2599 -4266
rect -2385 -4566 -2324 -4505
rect 2746 -4507 2807 -4446
rect 3021 -5063 3082 -5002
rect -2385 -5154 -2324 -5093
rect 311 -5209 372 -5148
rect -1646 -5339 -1585 -5278
rect 846 -5339 907 -5278
rect -3545 -6867 -3484 -6806
rect -3386 -7040 -3325 -6979
<< metal3 >>
rect 3009 -3452 3090 -3447
rect 3009 -3513 3019 -3452
rect 3080 -3513 3090 -3452
rect 3009 -3518 3090 -3513
rect -2556 -3928 -2475 -3923
rect -2556 -3989 -2546 -3928
rect -2485 -3989 -2475 -3928
rect -2556 -3994 -2475 -3989
rect -2546 -4266 -2485 -3994
rect 2528 -4266 2609 -4261
rect -2546 -4327 2538 -4266
rect 2599 -4327 2609 -4266
rect -2546 -6637 -2485 -4327
rect 2528 -4332 2609 -4327
rect 2736 -4446 2817 -4441
rect -2385 -4500 2746 -4446
rect -2395 -4505 2746 -4500
rect -2395 -4566 -2385 -4505
rect -2324 -4507 2746 -4505
rect 2807 -4507 2817 -4446
rect -2324 -4566 -2314 -4507
rect 2736 -4512 2817 -4507
rect -2395 -4571 -2314 -4566
rect -2385 -5088 -2324 -4571
rect 3021 -4997 3082 -3518
rect 3011 -5002 3092 -4997
rect 3011 -5063 3021 -5002
rect 3082 -5063 3092 -5002
rect 3011 -5068 3092 -5063
rect -2395 -5093 -2314 -5088
rect -2395 -5154 -2385 -5093
rect -2324 -5154 -2314 -5093
rect -2395 -5159 -2314 -5154
rect 301 -5147 382 -5143
rect 3021 -5147 3082 -5068
rect 301 -5148 3082 -5147
rect -3545 -6698 -2485 -6637
rect -3545 -6801 -3484 -6698
rect -2385 -6786 -2324 -5159
rect 301 -5209 311 -5148
rect 372 -5208 3082 -5148
rect 372 -5209 382 -5208
rect 301 -5214 382 -5209
rect -1656 -5278 -1575 -5273
rect 836 -5278 917 -5273
rect -1656 -5339 -1646 -5278
rect -1585 -5339 846 -5278
rect 907 -5339 917 -5278
rect -1656 -5344 -1575 -5339
rect 836 -5344 917 -5339
rect -3555 -6806 -3474 -6801
rect -3555 -6867 -3545 -6806
rect -3484 -6867 -3474 -6806
rect -3555 -6872 -3474 -6867
rect -3386 -6847 -2324 -6786
rect -3386 -6974 -3325 -6847
rect -3396 -6979 -3315 -6974
rect -3396 -7040 -3386 -6979
rect -3325 -7040 -3315 -6979
rect -3396 -7045 -3315 -7040
<< labels >>
flabel metal2 3147 -3484 3147 -3484 1 FreeSans 1200 0 0 0 on
port 4 n
flabel metal2 3431 -5243 3431 -5243 1 FreeSans 1200 0 0 0 op
port 3 n
flabel metal2 5049 -9956 5049 -9956 1 FreeSans 1200 0 0 0 cmc
port 11 n
flabel metal1 4262 -15741 4262 -15741 1 FreeSans 1200 0 0 0 bias_a
port 7 n
flabel metal1 6929 -13167 6929 -13167 1 FreeSans 1200 0 0 0 bias_d
port 10 n
flabel metal2 10414 -8662 10414 -8662 1 FreeSans 1200 0 0 0 bias_e
port 6 n
flabel metal1 -7420 -1403 -7420 -1403 1 FreeSans 1200 0 0 0 VDD
port 12 n power bidirectional
flabel metal1 -7407 -17402 -7407 -17402 1 FreeSans 1200 0 0 0 VSS
port 13 n ground bidirectional
flabel metal1 -6957 -14245 -6957 -14245 1 FreeSans 1200 0 0 0 i_bias
port 5 n
flabel metal1 -3636 -12323 -3636 -12323 1 FreeSans 1200 0 0 0 bias_c
port 9 n
flabel metal1 -6950 -12541 -6950 -12541 1 FreeSans 1200 0 0 0 ip
port 1 n
flabel metal1 -6952 -13880 -6952 -13880 1 FreeSans 1200 0 0 0 in
port 2 n
flabel metal1 -4277 -7715 -4277 -7715 1 FreeSans 1200 0 0 0 bias_b
port 8 n
<< end >>
