* NGSPICE file created from analog_top.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_BRTJC6 a_n345_n500# a_1135_n588# a_n603_n588#
+ a_n1393_n588# a_n1609_n500# a_661_n588# a_n1135_n500# a_n977_n500# a_1293_n588#
+ a_n761_n588# a_n503_n500# a_n1551_n588# a_129_n500# a_n1293_n500# a_287_n500# a_n661_n500#
+ a_1451_n588# a_n1451_n500# a_919_n500# a_445_n500# a_1077_n500# a_29_n588# a_n129_n588#
+ a_603_n500# a_187_n588# a_1235_n500# a_n287_n588# a_761_n500# a_819_n588# a_345_n588#
+ a_n1077_n588# a_n29_n500# a_1393_n500# a_n919_n588# a_n1743_n722# a_n187_n500# a_977_n588#
+ a_n445_n588# a_503_n588# a_n1235_n588# a_1551_n500# a_n819_n500#
X0 a_n819_n500# a_n919_n588# a_n977_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n588# a_n819_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n588# a_761_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n588# a_n345_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n588# a_603_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n588# a_129_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n588# a_n1451_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n588# a_1235_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n588# a_n503_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n588# a_n29_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n588# a_287_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n588# a_n1609_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n588# a_1393_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n588# a_n1135_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_n503_n500# a_n603_n588# a_n661_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_1077_n500# a_977_n588# a_919_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n588# a_n187_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n588# a_445_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n588# a_n1293_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n588# a_1077_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CADZ46 a_n345_n500# a_n1609_n500# a_n1135_n500#
+ a_29_n597# a_n977_n500# a_n129_n597# a_187_n597# a_n503_n500# a_129_n500# a_n1293_n500#
+ a_n287_n597# a_819_n597# a_n1077_n597# a_287_n500# a_n661_n500# a_345_n597# a_n919_n597#
+ a_n1451_n500# a_977_n597# a_n445_n597# a_919_n500# a_n1235_n597# a_445_n500# a_503_n597#
+ w_n1809_n797# a_n603_n597# a_1077_n500# a_1135_n597# a_661_n597# a_n1393_n597# a_603_n500#
+ a_1293_n597# a_n761_n597# a_1235_n500# a_n1551_n597# a_761_n500# a_n29_n500# a_1451_n597#
+ a_1393_n500# a_n187_n500# a_1551_n500# a_n819_n500#
X0 a_n819_n500# a_n919_n597# a_n977_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n597# a_n819_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n597# a_761_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n597# a_n345_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n597# a_603_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n597# a_129_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n597# a_n1451_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n597# a_1235_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n597# a_n503_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n597# a_n29_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n597# a_287_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n597# a_n1609_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n597# a_1393_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n597# a_n1135_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_1077_n500# a_977_n597# a_919_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X15 a_n503_n500# a_n603_n597# a_n661_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n597# a_n187_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n597# a_445_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n597# a_n1293_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n597# a_1077_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
.ends

.subckt esd_cell esd VSS VDD
Xsky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0 VSS VSS VSS VSS VSS VSS esd VSS VSS VSS esd
+ VSS esd VSS VSS VSS VSS esd VSS esd esd VSS VSS VSS VSS VSS VSS esd VSS VSS VSS
+ VSS esd VSS VSS esd VSS VSS VSS VSS VSS esd sky130_fd_pr__nfet_g5v0d10v5_BRTJC6
Xsky130_fd_pr__pfet_g5v0d10v5_CADZ46_0 VDD VDD esd VDD VDD VDD VDD esd esd VDD VDD
+ VDD VDD VDD VDD VDD VDD esd VDD VDD VDD VDD esd VDD VDD VDD esd VDD VDD VDD VDD
+ VDD VDD VDD VDD esd VDD VDD esd esd VDD esd sky130_fd_pr__pfet_g5v0d10v5_CADZ46
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CEWQ64 c1_n260_n210# m3_n360_n310#
X0 c1_n260_n210# m3_n360_n310# sky130_fd_pr__cap_mim_m3_1 l=2.1e+06u w=2.1e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CGPBWM m3_n1031_n980# c1_n931_n880#
X0 c1_n931_n880# m3_n1031_n980# sky130_fd_pr__cap_mim_m3_1 l=8.8e+06u w=8.8e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136#
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
X0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt transmission_gate out en_b en VSS VDD in
Xsky130_fd_pr__pfet_01v8_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ sky130_fd_pr__pfet_01v8_UNG2NQ
Xsky130_fd_pr__nfet_01v8_6J4AMR_0 out in in out in in VSS out en in out out out sky130_fd_pr__nfet_01v8_6J4AMR
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_II a_n207_n140# a_n1039_n205# a_1275_n205# a_29_n205#
+ a_327_n140# a_n1275_n140# a_n683_n205# a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140#
+ a_1097_n205# a_1395_n140# a_n505_n205# a_n741_n140# a_563_n205# a_861_n140# a_919_n205#
+ a_n327_n205# a_n563_n140# a_385_n205# a_1217_n140# a_n1395_n205# a_683_n140# a_n919_n140#
+ a_n149_n205# w_n1489_n241# a_1039_n140# a_n385_n140# a_207_n205# a_n1217_n205# a_505_n140#
+ a_n1453_n140# a_n861_n205#
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1395_n140# a_1275_n205# a_1217_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_327_n140# a_207_n205# a_149_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_149_n140# a_29_n205# a_n29_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_861_n140# a_741_n205# a_683_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n207_n140# a_n327_n205# a_n385_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_1217_n140# a_1097_n205# a_1039_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n1275_n140# a_n1395_n205# a_n1453_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n205# a_n919_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1217_n205# a_n1275_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n205# a_505_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n205# a_861_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n29_n140# a_n149_n205# a_n207_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_n563_n140# a_n683_n205# a_n741_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FF a_20_n120# a_n78_n120# a_n33_n208# VSUBS
X0 a_20_n120# a_n33_n208# a_n78_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
.ends

.subckt sky130_fd_pr__nfet_01v8_DD a_1751_n140# a_n149_n194# a_1987_n194# a_n2819_n194#
+ a_n207_n140# a_n1809_n140# a_n2877_n140# a_207_n194# a_n2285_n194# a_1453_n194#
+ a_n1217_n194# a_n3353_n194# a_327_n140# a_n1275_n140# a_n2343_n140# a_2521_n194#
+ a_n861_n194# a_1573_n140# a_n3411_n140# a_2641_n140# a_n2699_n140# a_2877_n194#
+ a_1809_n194# a_2997_n140# a_n29_n140# a_n1039_n194# a_n3175_n194# a_1929_n140# a_149_n140#
+ a_n1097_n140# a_2343_n194# a_1275_n194# a_29_n194# a_n2107_n194# a_n2165_n140# a_n3233_n140#
+ a_3411_n194# a_n683_n194# a_1395_n140# a_3531_n140# a_2463_n140# a_n741_n140# a_2699_n194#
+ a_741_n194# a_n3589_n140# a_n1751_n194# a_861_n140# a_1097_n194# a_2819_n140# a_3233_n194#
+ a_2165_n194# a_n3055_n140# a_n505_n194# a_2285_n140# a_n563_n140# a_563_n194# a_3353_n140#
+ a_1217_n140# a_n1573_n194# a_n2641_n194# a_683_n140# a_n919_n140# a_n1631_n140#
+ a_919_n194# a_3055_n194# a_n2997_n194# a_n1987_n140# a_n327_n194# a_n1929_n194#
+ a_3175_n140# a_1039_n140# a_n385_n140# a_385_n194# a_2107_n140# a_n1395_n194# a_n2463_n194#
+ a_n3531_n194# a_505_n140# a_n1453_n140# a_1631_n194# a_n2521_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2165_n140# a_n2285_n194# a_n2343_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_3175_n140# a_3055_n194# a_2997_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n3233_n140# a_n3353_n194# a_n3411_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_2997_n140# a_2877_n194# a_2819_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1987_n140# a_n2107_n194# a_n2165_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1809_n140# a_n1929_n194# a_n1987_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n1453_n140# a_n1573_n194# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2463_n140# a_2343_n194# a_2285_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n2521_n140# a_n2641_n194# a_n2699_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_3531_n140# a_3411_n194# a_3353_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1751_n140# a_1631_n194# a_1573_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n3055_n140# a_n3175_n194# a_n3233_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_2819_n140# a_2699_n194# a_2641_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n2877_n140# a_n2997_n194# a_n3055_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_2285_n140# a_2165_n194# a_2107_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_n2699_n140# a_n2819_n194# a_n2877_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n2343_n140# a_n2463_n194# a_n2521_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_2107_n140# a_1987_n194# a_1929_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X31 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_3353_n140# a_3233_n194# a_3175_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_n3411_n140# a_n3531_n194# a_n3589_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X36 a_1573_n140# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_1929_n140# a_1809_n194# a_1751_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_n1631_n140# a_n1751_n194# a_n1809_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_2641_n140# a_2521_n194# a_2463_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_CC a_n1008_n140# a_2374_n140# a_1306_n140# a_n652_n140#
+ a_652_n194# a_n1662_n194# a_772_n140# a_n2730_n194# a_n1720_n140# a_n60_n194# a_2076_n194#
+ a_1008_n194# a_2196_n140# a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194#
+ a_n2552_n194# a_594_n140# a_n1542_n140# a_n2610_n140# a_1720_n194# a_1840_n140#
+ a_n238_n194# a_n2908_n194# a_3086_n140# a_n296_n140# a_n1898_n140# a_n2966_n140#
+ a_296_n194# a_2018_n140# a_60_n140# a_n1306_n194# a_n2374_n194# a_n1364_n140# a_1542_n194#
+ a_416_n140# a_n2432_n140# a_2610_n194# a_n950_n194# a_1662_n140# a_2730_n140# a_2966_n194#
+ a_1898_n194# a_n2788_n140# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194#
+ a_238_n140# a_n1186_n140# a_n2254_n140# a_2432_n194# a_1364_n194# a_n772_n194# a_2552_n140#
+ a_1484_n140# a_n830_n140# a_2788_n194# a_830_n194# a_n1840_n194# a_950_n140# a_n3086_n194#
+ a_2908_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_n3144_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2374_n140# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2788_n140# a_n2908_n194# a_n2966_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n2432_n140# a_n2552_n194# a_n2610_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2966_n140# a_n3086_n194# a_n3144_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_2730_n140# a_2610_n194# a_2552_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n2610_n140# a_n2730_n194# a_n2788_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n2254_n140# a_n2374_n194# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_3086_n140# a_2966_n194# a_2908_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_2552_n140# a_2432_n194# a_2374_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_2908_n140# a_2788_n194# a_2730_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_BB a_n1008_n140# a_n652_n140# a_652_n194# a_772_n140#
+ a_n60_n194# a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140#
+ a_296_n194# a_60_n140# a_416_n140# a_n950_n194# a_n118_n140# a_118_n194# a_238_n140#
+ a_n772_n194# a_n830_n140# a_830_n194# a_950_n140# a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__pfet_01v8_HH a_n1008_n140# a_n416_n205# a_1306_n140# a_n652_n140#
+ a_474_n205# a_n1484_n205# a_772_n140# a_n1720_n140# a_1720_n205# a_n238_n205# a_n474_n140#
+ a_296_n205# a_1128_n140# a_594_n140# a_1542_n205# a_n1306_n205# w_n2112_n240# a_n1542_n140#
+ a_n950_n205# a_1840_n140# a_1898_n205# a_n296_n140# a_n1898_n140# a_2018_n140# a_60_n140#
+ a_118_n205# a_n1128_n205# a_n1364_n140# a_1364_n205# a_416_n140# a_n772_n205# a_1662_n140#
+ a_830_n205# a_n1840_n205# a_n118_n140# a_1186_n205# a_n2018_n205# a_238_n140# a_n1186_n140#
+ a_n594_n205# a_1484_n140# a_n830_n140# a_652_n205# a_n1662_n205# a_950_n140# a_n60_n205#
+ a_n2076_n140# a_1008_n205#
X0 a_1662_n140# a_1542_n205# a_1484_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n205# a_n296_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n205# a_n830_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_2018_n140# a_1898_n205# a_1840_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1008_n140# a_n1128_n205# a_n1186_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_594_n140# a_474_n205# a_416_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_60_n140# a_n60_n205# a_n118_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1484_n140# a_1364_n205# a_1306_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1542_n140# a_n1662_n205# a_n1720_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_950_n140# a_830_n205# a_772_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n830_n140# a_n950_n205# a_n1008_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n474_n140# a_n594_n205# a_n652_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_1840_n140# a_1720_n205# a_1662_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_416_n140# a_296_n205# a_238_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1898_n140# a_n2018_n205# a_n2076_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n296_n140# a_n416_n205# a_n474_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n1720_n140# a_n1840_n205# a_n1898_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1306_n140# a_1186_n205# a_1128_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1364_n140# a_n1484_n205# a_n1542_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_238_n140# a_118_n205# a_60_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_1128_n140# a_1008_n205# a_950_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_n1186_n140# a_n1306_n205# a_n1364_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_772_n140# a_652_n205# a_594_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_GG a_n652_n140# a_652_n194# a_772_n140# a_n60_n194#
+ a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140# a_296_n194#
+ a_60_n140# a_416_n140# a_n118_n140# a_118_n194# a_238_n140# a_n772_n194# a_n830_n140#
+ a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_AA a_n149_n194# a_n207_n140# a_207_n194# a_n1217_n194#
+ a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140# a_n1097_n140#
+ a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194# a_861_n140#
+ a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140# a_n919_n140#
+ a_919_n194# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194# a_n1395_n194# a_505_n140#
+ a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_EE a_n352_n194# a_n60_n194# a_n644_n194# a_n936_n194#
+ a_n410_n140# a_n994_n140# a_n702_n140# a_n232_n140# a_n524_n140# a_524_n194# a_232_n194#
+ a_n816_n140# a_816_n194# a_644_n140# a_352_n140# a_936_n140# a_60_n140# a_174_n140#
+ a_466_n140# a_758_n140# a_n118_n140# VSUBS
X0 a_n232_n140# a_n352_n194# a_n410_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n524_n140# a_n644_n194# a_n702_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n816_n140# a_n936_n194# a_n994_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_352_n140# a_232_n194# a_174_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_644_n140# a_524_n194# a_466_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_936_n140# a_816_n194# a_758_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580#
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
.ends

.subckt sc_cmfb cmc on bias_a p2_b p1 cm VSS p2 VDD op p1_b
Xtransmission_gate_10 on p1_b p1 VSS VDD transmission_gate_3/out transmission_gate
Xtransmission_gate_11 op p1_b p1 VSS VDD transmission_gate_4/out transmission_gate
Xtransmission_gate_0 transmission_gate_7/in p1_b p1 VSS VDD cm transmission_gate
Xtransmission_gate_1 transmission_gate_6/in p1_b p1 VSS VDD cm transmission_gate
Xtransmission_gate_2 transmission_gate_8/in p1_b p1 VSS VDD bias_a transmission_gate
Xtransmission_gate_3 transmission_gate_3/out p2_b p2 VSS VDD cm transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in unit_cap_mim_m3m4
Xtransmission_gate_4 transmission_gate_4/out p2_b p2 VSS VDD cm transmission_gate
Xunit_cap_mim_m3m4_1 on cmc unit_cap_mim_m3m4
Xtransmission_gate_5 transmission_gate_9/in p2_b p2 VSS VDD bias_a transmission_gate
Xunit_cap_mim_m3m4_2 op cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ unit_cap_mim_m3m4
Xtransmission_gate_6 op p2_b p2 VSS VDD transmission_gate_6/in transmission_gate
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ unit_cap_mim_m3m4
Xtransmission_gate_7 on p2_b p2 VSS VDD transmission_gate_7/in transmission_gate
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_4 on cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc unit_cap_mim_m3m4
Xtransmission_gate_8 cmc p2_b p2 VSS VDD transmission_gate_8/in transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc unit_cap_mim_m3m4
Xtransmission_gate_9 cmc p1_b p1 VSS VDD transmission_gate_9/in transmission_gate
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ unit_cap_mim_m3m4
.ends

.subckt ota_w_test ip in p1 op i_bias cm bias_a bias_b bias_c bias_d cmc VDD VSS on
+ p2_b p1_b p2
Xsky130_fd_pr__pfet_01v8_lvt_II_2 m1_n6302_n3889# bias_b m1_n6302_n3889# bias_b VDD
+ m1_n6302_n3889# bias_b bias_b VDD m1_n6302_n3889# VDD bias_b m1_n6302_n3889# bias_b
+ VDD bias_b m1_n208_n2883# bias_b bias_b m1_1038_n2886# bias_b m1_n6302_n3889# m1_n6302_n3889#
+ VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b bias_b m1_1038_n2886# m1_n6302_n3889#
+ bias_b sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_lvt_FF_9 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_DD_2 m1_n947_n12836# bias_d VSS bias_d bias_a m1_n1659_n11581#
+ m1_n947_n12836# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# op on bias_d
+ bias_d on on op on bias_d VSS op m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n1659_n11581#
+ bias_d bias_d bias_d VSS m1_n947_n12836# m1_n947_n12836# op VSS m1_n947_n12836#
+ op m1_n1659_n11581# m1_n1659_n11581# bias_d bias_d on bias_d on bias_d m1_n1659_n11581#
+ bias_d bias_d on VSS op VSS VSS op on bias_d bias_d m1_n947_n12836# op op bias_d
+ bias_d bias_d VSS bias_d VSS m1_n1659_n11581# m1_n947_n12836# m1_n2176_n12171# VSS
+ m1_n1659_n11581# bias_d bias_d on VSS m1_n1659_n11581# bias_d m1_n947_n12836# VSS
+ sky130_fd_pr__nfet_01v8_DD
Xsky130_fd_pr__pfet_01v8_lvt_II_3 m1_2462_n3318# bias_b m1_2463_n5585# bias_b VDD
+ m1_2462_n3318# bias_b bias_b VDD m1_2463_n5585# VDD bias_b m1_2463_n5585# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2463_n5585# m1_2462_n3318#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2462_n3318#
+ bias_b sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__pfet_01v8_lvt_II_4 m1_1038_n2886# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_n208_n2883# VDD VDD VDD bias_b VDD bias_b m1_n208_n2883# bias_b bias_b
+ m1_n208_n2883# bias_b VDD VDD VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b VDD m1_1038_n2886#
+ VDD bias_b sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_CC_4 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a
+ VSS cmc VSS cmc cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc VSS cmc cmc VSS VSS m1_n5574_n13620# m1_n5574_n13620#
+ bias_a m1_n5574_n13620# VSS bias_a cmc VSS cmc VSS VSS bias_a bias_a m1_n5574_n13620#
+ m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620# m1_n5574_n13620#
+ m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a bias_a bias_a m1_n5574_n13620#
+ m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620# cmc cmc VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_5 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS
+ bias_a VSS VSS bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS VSS bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS VSS VSS cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS m1_n5574_n13620# bias_a
+ bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_6 VSS VSS VSS VSS bias_a bias_a m1_n947_n12836# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n1659_n11581# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n947_n12836# bias_a m1_n1659_n11581# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n1659_n11581# m1_n947_n12836# bias_a bias_a bias_a
+ m1_n1659_n11581# m1_n2176_n12171# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_10 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS
+ bias_a VSS cmc cmc bias_a VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS cmc bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_7 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n947_n12836# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n1659_n11581# m1_n2176_n12171# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n2176_n12171# m1_n1659_n11581# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_0 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias i_bias
+ i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__nfet_01v8_CC_11 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a
+ VSS cmc VSS bias_a bias_a cmc VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc VSS bias_a cmc VSS VSS m1_n5574_n13620# m1_n5574_n13620#
+ bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620# bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ cmc bias_a m1_n5574_n13620# m1_n5574_n13620# VSS cmc bias_a VSS m1_n5574_n13620#
+ bias_a cmc VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_8 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n947_n12836# m1_n947_n12836# bias_a m1_n1659_n11581# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n1659_n11581# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n1659_n11581# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n1659_n11581# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n947_n12836# m1_n2176_n12171# m1_n947_n12836# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_1 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__nfet_01v8_CC_9 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a
+ VSS cmc VSS VSS cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc VSS VSS cmc VSS VSS m1_n5574_n13620# m1_n5574_n13620#
+ bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# VSS cmc VSS VSS VSS bias_a cmc m1_n5574_n13620# m1_n5574_n13620#
+ m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a bias_a bias_a m1_n5574_n13620#
+ m1_n5574_n13620# VSS bias_a bias_a VSS m1_n5574_n13620# cmc cmc VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_2 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__nfet_01v8_CC_12 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS
+ bias_a VSS bias_a bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS bias_a bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS cmc bias_a VSS bias_a VSS VSS cmc cmc
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620# bias_a bias_a
+ cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS
+ m1_n5574_n13620# cmc cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc bias_a VSS
+ m1_n5574_n13620# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_3 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias i_bias
+ i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__pfet_01v8_HH_0 VDD bias_c m1_6690_n8907# op bias_c bias_c m1_1038_n2886#
+ bias_b bias_c VDD m1_n208_n2883# bias_c VDD on bias_c VDD VDD m1_2463_n5585# VDD
+ m1_2462_n3318# m1_2462_n3318# op m1_2463_n5585# m1_2462_n3318# VDD VDD VDD bias_b
+ bias_c m1_1038_n2886# bias_c m1_6690_n8907# VDD bias_c VDD VDD m1_2463_n5585# on
+ VDD bias_c m1_2462_n3318# m1_n208_n2883# bias_c bias_c VDD VDD m1_2463_n5585# VDD
+ sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__nfet_01v8_lvt_GG_0 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_10 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__pfet_01v8_HH_1 op VDD on op VDD bias_c m1_1038_n2886# op bias_c bias_c
+ VDD VDD m1_1038_n2886# on bias_c bias_c VDD m1_n208_n2883# bias_c m1_1038_n2886#
+ m1_1038_n2886# m1_n6302_n3889# m1_n208_n2883# m1_1038_n2886# m1_n6302_n3889# bias_c
+ bias_c op bias_c VDD bias_c on bias_c bias_c cm bias_c m1_n208_n2883# cm m1_n208_n2883#
+ VDD m1_1038_n2886# m1_n208_n2883# bias_c bias_c on bias_c m1_n208_n2883# bias_c
+ sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__nfet_01v8_AA_0 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_lvt_GG_1 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_11 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__pfet_01v8_HH_3 VDD bias_c bias_b on bias_c bias_c m1_n208_n2883# m1_6690_n8907#
+ bias_c VDD m1_1038_n2886# bias_c VDD op bias_c VDD VDD m1_2462_n3318# VDD m1_2463_n5585#
+ m1_2463_n5585# on m1_2462_n3318# m1_2463_n5585# VDD VDD VDD m1_6690_n8907# bias_c
+ m1_n208_n2883# bias_c bias_b VDD bias_c VDD VDD m1_2462_n3318# op VDD bias_c m1_2463_n5585#
+ m1_1038_n2886# bias_c bias_c VDD VDD m1_2462_n3318# VDD sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__pfet_01v8_HH_2 on VDD op on VDD bias_c m1_n208_n2883# on bias_c bias_c
+ VDD VDD m1_n208_n2883# op bias_c bias_c VDD m1_1038_n2886# bias_c m1_n208_n2883#
+ m1_n208_n2883# m1_n6302_n3889# m1_1038_n2886# m1_n208_n2883# m1_n6302_n3889# bias_c
+ bias_c on bias_c VDD bias_c op bias_c bias_c cm bias_c m1_1038_n2886# cm m1_1038_n2886#
+ VDD m1_n208_n2883# m1_1038_n2886# bias_c bias_c op bias_c m1_1038_n2886# bias_c
+ sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__nfet_01v8_lvt_GG_2 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_AA_1 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d bias_a m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_a m1_6690_n8907# bias_a VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_AA_2 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_a
+ m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_lvt_FF_12 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_GG_3 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_AA_3 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d
+ m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_lvt_FF_13 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_GG_4 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_14 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_15 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_GG_5 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_EE_0 cm cm cm cm cm cm cm m1_11534_n9706# m1_11242_n9716#
+ cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# cm cm cm cm VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_GG_6 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_EE_1 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490# m1_11534_n9706#
+ m1_11242_n9716# cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# m1_11940_n10482#
+ m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_GG_7 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_0 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_EE_2 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490# m1_11534_n11258#
+ m1_11244_n11260# cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260#
+ m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_FF_1 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_EE_3 cm cm cm cm VSS cm VSS m1_11534_n11258# m1_11244_n11260#
+ cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260# VSS VSS cm VSS
+ VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_FF_2 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsc_cmfb_0 cmc on bias_a p2_b p1 cm VSS p2 VDD op p1_b sc_cmfb
Xsky130_fd_pr__nfet_01v8_lvt_FF_3 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_4 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_5 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_6 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__pfet_01v8_lvt_II_0 m1_n208_n2883# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_1038_n2886# VDD VDD VDD bias_b VDD bias_b m1_1038_n2886# bias_b bias_b
+ m1_1038_n2886# bias_b VDD VDD VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b VDD m1_n208_n2883#
+ VDD bias_b sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_lvt_FF_7 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_DD_0 m1_n1659_n11581# bias_d VSS bias_d bias_a m1_n947_n12836#
+ m1_n1659_n11581# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# on op bias_d
+ bias_d op op on op bias_d VSS on m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n947_n12836#
+ bias_d bias_d bias_d VSS m1_n1659_n11581# m1_n1659_n11581# on VSS m1_n1659_n11581#
+ on m1_n947_n12836# m1_n947_n12836# bias_d bias_d op bias_d op bias_d m1_n947_n12836#
+ bias_d bias_d op VSS on VSS VSS on op bias_d bias_d m1_n1659_n11581# on on bias_d
+ bias_d bias_d VSS bias_d VSS m1_n947_n12836# m1_n1659_n11581# m1_n2176_n12171# VSS
+ m1_n947_n12836# bias_d bias_d op VSS m1_n947_n12836# bias_d m1_n1659_n11581# VSS
+ sky130_fd_pr__nfet_01v8_DD
Xsky130_fd_pr__pfet_01v8_lvt_II_1 m1_2463_n5585# bias_b m1_2462_n3318# bias_b VDD
+ m1_2463_n5585# bias_b bias_b VDD m1_2462_n3318# VDD bias_b m1_2462_n3318# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2462_n3318# m1_2463_n5585#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2463_n5585#
+ bias_b sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_lvt_FF_8 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_DD_1 m1_n947_n12836# bias_d bias_d bias_d op m1_n947_n12836#
+ m1_n2176_n12171# bias_d VSS bias_d VSS bias_d m1_n1659_n11581# on VSS bias_d bias_d
+ on bias_a bias_a bias_a bias_d bias_d bias_a m1_n1659_n11581# VSS bias_d on op VSS
+ VSS bias_d bias_d bias_d m1_n947_n12836# m1_n2176_n12171# bias_a bias_d m1_n947_n12836#
+ bias_a m1_n2176_n12171# m1_n1659_n11581# bias_d bias_d bias_a bias_d op VSS m1_n2176_n12171#
+ bias_d VSS bias_a bias_d VSS op bias_d bias_a on bias_d bias_d m1_n1659_n11581#
+ op on VSS bias_d bias_d on bias_d bias_d m1_n2176_n12171# VSS m1_n1659_n11581# bias_d
+ m1_n947_n12836# bias_d VSS bias_a op m1_n947_n12836# bias_d m1_n2176_n12171# VSS
+ sky130_fd_pr__nfet_01v8_DD
.ends

.subckt sky130_fd_sc_hd__clkinv_16 A VGND VPWR Y VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.0605e+12p pd=1.261e+07u as=1.0059e+12p ps=1.151e+07u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.515e+12p pd=3.103e+07u as=3.655e+12p ps=3.331e+07u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt onebit_dac v_b out v_lo v_hi v VSS VDD
Xtransmission_gate_0 out v_b v VSS VDD v_hi transmission_gate
Xtransmission_gate_1 out v v_b VSS VDD v_lo transmission_gate
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_VU7MNH a_n652_n140# a_652_n194# a_772_n140# a_n60_n194#
+ a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140# a_296_n194#
+ a_60_n140# a_416_n140# a_n118_n140# a_118_n194# a_238_n140# a_n772_n194# a_n830_n140#
+ a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_TRAZV8 a_20_n120# a_n78_n120# a_n33_n208# VSUBS
X0 a_20_n120# a_n33_n208# a_n78_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
.ends

.subckt sky130_fd_pr__nfet_01v8_BASQVB a_n1008_n140# a_n652_n140# a_652_n194# a_772_n140#
+ a_n60_n194# a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140#
+ a_296_n194# a_60_n140# a_416_n140# a_n950_n194# a_n118_n140# a_118_n194# a_238_n140#
+ a_n772_n194# a_n830_n140# a_830_n194# a_950_n140# a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_UFQYRB a_1751_n140# a_n149_n194# a_1987_n194# a_n2819_n194#
+ a_n207_n140# a_n1809_n140# a_n2877_n140# a_207_n194# a_n2285_n194# a_1453_n194#
+ a_n1217_n194# a_n3353_n194# a_327_n140# a_n1275_n140# a_n2343_n140# a_2521_n194#
+ a_n861_n194# a_1573_n140# a_n3411_n140# a_2641_n140# a_n2699_n140# a_2877_n194#
+ a_1809_n194# a_2997_n140# a_n29_n140# a_n1039_n194# a_n3175_n194# a_1929_n140# a_149_n140#
+ a_n1097_n140# a_2343_n194# a_1275_n194# a_29_n194# a_n2107_n194# a_n2165_n140# a_n3233_n140#
+ a_3411_n194# a_n683_n194# a_1395_n140# a_3531_n140# a_2463_n140# a_n741_n140# a_2699_n194#
+ a_741_n194# a_n3589_n140# a_n1751_n194# a_861_n140# a_1097_n194# a_2819_n140# a_3233_n194#
+ a_2165_n194# a_n3055_n140# a_n505_n194# a_2285_n140# a_n563_n140# a_563_n194# a_3353_n140#
+ a_1217_n140# a_n1573_n194# a_n2641_n194# a_683_n140# a_n919_n140# a_n1631_n140#
+ a_919_n194# a_3055_n194# a_n2997_n194# a_n1987_n140# a_n327_n194# a_n1929_n194#
+ a_3175_n140# a_1039_n140# a_n385_n140# a_385_n194# a_2107_n140# a_n1395_n194# a_n2463_n194#
+ a_n3531_n194# a_505_n140# a_n1453_n140# a_1631_n194# a_n2521_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2165_n140# a_n2285_n194# a_n2343_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_3175_n140# a_3055_n194# a_2997_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n3233_n140# a_n3353_n194# a_n3411_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_2997_n140# a_2877_n194# a_2819_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1987_n140# a_n2107_n194# a_n2165_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1809_n140# a_n1929_n194# a_n1987_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n1453_n140# a_n1573_n194# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2463_n140# a_2343_n194# a_2285_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n2521_n140# a_n2641_n194# a_n2699_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_3531_n140# a_3411_n194# a_3353_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1751_n140# a_1631_n194# a_1573_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n3055_n140# a_n3175_n194# a_n3233_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_2819_n140# a_2699_n194# a_2641_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n2877_n140# a_n2997_n194# a_n3055_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_2285_n140# a_2165_n194# a_2107_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_n2699_n140# a_n2819_n194# a_n2877_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n2343_n140# a_n2463_n194# a_n2521_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_2107_n140# a_1987_n194# a_1929_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X31 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_3353_n140# a_3233_n194# a_3175_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_n3411_n140# a_n3531_n194# a_n3589_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X36 a_1573_n140# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_1929_n140# a_1809_n194# a_1751_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_n1631_n140# a_n1751_n194# a_n1809_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_2641_n140# a_2521_n194# a_2463_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_7P4E2J a_n149_n194# a_n207_n140# a_207_n194# a_n1217_n194#
+ a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140# a_n1097_n140#
+ a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194# a_861_n140#
+ a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140# a_n919_n140#
+ a_919_n194# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194# a_n1395_n194# a_505_n140#
+ a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_KEEN2X a_n1008_n140# a_2374_n140# a_1306_n140# a_n652_n140#
+ a_652_n194# a_n1662_n194# a_772_n140# a_n2730_n194# a_n1720_n140# a_n60_n194# a_2076_n194#
+ a_1008_n194# a_2196_n140# a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194#
+ a_n2552_n194# a_594_n140# a_n1542_n140# a_n2610_n140# a_1720_n194# a_1840_n140#
+ a_n238_n194# a_n2908_n194# a_3086_n140# a_n296_n140# a_n1898_n140# a_n2966_n140#
+ a_296_n194# a_2018_n140# a_60_n140# a_n1306_n194# a_n2374_n194# a_n1364_n140# a_1542_n194#
+ a_416_n140# a_n2432_n140# a_2610_n194# a_n950_n194# a_1662_n140# a_2730_n140# a_2966_n194#
+ a_1898_n194# a_n2788_n140# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194#
+ a_238_n140# a_n1186_n140# a_n2254_n140# a_2432_n194# a_1364_n194# a_n772_n194# a_2552_n140#
+ a_1484_n140# a_n830_n140# a_2788_n194# a_830_n194# a_n1840_n194# a_950_n140# a_n3086_n194#
+ a_2908_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_n3144_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2374_n140# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2788_n140# a_n2908_n194# a_n2966_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n2432_n140# a_n2552_n194# a_n2610_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2966_n140# a_n3086_n194# a_n3144_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_2730_n140# a_2610_n194# a_2552_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n2610_n140# a_n2730_n194# a_n2788_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n2254_n140# a_n2374_n194# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_3086_n140# a_2966_n194# a_2908_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_2552_n140# a_2432_n194# a_2374_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_2908_n140# a_2788_n194# a_2730_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__nfet_01v8_VJ4JGY a_n352_n194# a_n60_n194# a_n644_n194# a_n936_n194#
+ a_n410_n140# a_n994_n140# a_n702_n140# a_n232_n140# a_n524_n140# a_524_n194# a_232_n194#
+ a_n816_n140# a_816_n194# a_644_n140# a_352_n140# a_936_n140# a_60_n140# a_174_n140#
+ a_466_n140# a_758_n140# a_n118_n140# VSUBS
X0 a_n232_n140# a_n352_n194# a_n410_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n524_n140# a_n644_n194# a_n702_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n816_n140# a_n936_n194# a_n994_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_352_n140# a_232_n194# a_174_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_644_n140# a_524_n194# a_466_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_936_n140# a_816_n194# a_758_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__pfet_01v8_E4DCBA a_n1008_n140# a_n416_n205# a_1306_n140# a_n652_n140#
+ a_474_n205# a_n1484_n205# a_772_n140# a_n1720_n140# a_1720_n205# a_n238_n205# a_n474_n140#
+ a_296_n205# a_1128_n140# a_594_n140# a_1542_n205# a_n1306_n205# a_n1542_n140# a_n950_n205#
+ w_n2112_n241# a_1840_n140# a_1898_n205# a_n296_n140# a_n1898_n140# a_2018_n140#
+ a_60_n140# a_118_n205# a_n1128_n205# a_n1364_n140# a_1364_n205# a_416_n140# a_n772_n205#
+ a_1662_n140# a_830_n205# a_n1840_n205# a_n118_n140# a_1186_n205# a_n2018_n205# a_238_n140#
+ a_n1186_n140# a_n594_n205# a_1484_n140# a_n830_n140# a_652_n205# a_n1662_n205# a_950_n140#
+ a_n60_n205# a_n2076_n140# a_1008_n205#
X0 a_1662_n140# a_1542_n205# a_1484_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n205# a_n296_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n205# a_n830_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_2018_n140# a_1898_n205# a_1840_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1008_n140# a_n1128_n205# a_n1186_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_594_n140# a_474_n205# a_416_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_60_n140# a_n60_n205# a_n118_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1484_n140# a_1364_n205# a_1306_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1542_n140# a_n1662_n205# a_n1720_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_950_n140# a_830_n205# a_772_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n830_n140# a_n950_n205# a_n1008_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n474_n140# a_n594_n205# a_n652_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_1840_n140# a_1720_n205# a_1662_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_416_n140# a_296_n205# a_238_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1898_n140# a_n2018_n205# a_n2076_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n296_n140# a_n416_n205# a_n474_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n1720_n140# a_n1840_n205# a_n1898_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1306_n140# a_1186_n205# a_1128_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1364_n140# a_n1484_n205# a_n1542_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_238_n140# a_118_n205# a_60_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_1128_n140# a_1008_n205# a_950_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_n1186_n140# a_n1306_n205# a_n1364_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_772_n140# a_652_n205# a_594_n140# w_n2112_n241# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6QKDBA a_n207_n140# a_n1039_n205# a_1275_n205#
+ a_29_n205# a_327_n140# a_n1275_n140# a_n683_n205# a_741_n205# a_n29_n140# a_149_n140#
+ a_n1097_n140# a_1097_n205# a_1395_n140# a_n505_n205# a_n741_n140# a_563_n205# a_861_n140#
+ a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_1217_n140# a_n1395_n205# a_683_n140#
+ a_n919_n140# a_n149_n205# w_n1489_n241# a_1039_n140# a_n385_n140# a_207_n205# a_n1217_n205#
+ a_505_n140# a_n1453_n140# a_n861_n205#
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1395_n140# a_1275_n205# a_1217_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_327_n140# a_207_n205# a_149_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_149_n140# a_29_n205# a_n29_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_861_n140# a_741_n205# a_683_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n207_n140# a_n327_n205# a_n385_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_1217_n140# a_1097_n205# a_1039_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n1275_n140# a_n1395_n205# a_n1453_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n205# a_n919_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1217_n205# a_n1275_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n205# a_505_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n205# a_861_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n29_n140# a_n149_n205# a_n207_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_n563_n140# a_n683_n205# a_n741_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
.ends

.subckt ota ip in op i_bias cm VSS on p2_b VDD p1_b p2 p1
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_0 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_1 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_2 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_3 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_4 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_0 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_1 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_5 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_2 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_BASQVB_0 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias
+ i_bias i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_6 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_3 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_0 m1_n1659_n11581# bias_d VSS bias_d bias_a m1_n947_n12836#
+ m1_n1659_n11581# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# on op bias_d
+ bias_d op op on op bias_d VSS on m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n947_n12836#
+ bias_d bias_d bias_d VSS m1_n1659_n11581# m1_n1659_n11581# on VSS m1_n1659_n11581#
+ on m1_n947_n12836# m1_n947_n12836# bias_d bias_d op bias_d op bias_d m1_n947_n12836#
+ bias_d bias_d op VSS on VSS VSS on op bias_d bias_d m1_n1659_n11581# on on bias_d
+ bias_d bias_d VSS bias_d VSS m1_n947_n12836# m1_n1659_n11581# m1_n2176_n12171# VSS
+ m1_n947_n12836# bias_d bias_d op VSS m1_n947_n12836# bias_d m1_n1659_n11581# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_1 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias
+ bias_c i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_7 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_4 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_1 m1_n947_n12836# bias_d bias_d bias_d op m1_n947_n12836#
+ m1_n2176_n12171# bias_d VSS bias_d VSS bias_d m1_n1659_n11581# on VSS bias_d bias_d
+ on bias_a bias_a bias_a bias_d bias_d bias_a m1_n1659_n11581# VSS bias_d on op VSS
+ VSS bias_d bias_d bias_d m1_n947_n12836# m1_n2176_n12171# bias_a bias_d m1_n947_n12836#
+ bias_a m1_n2176_n12171# m1_n1659_n11581# bias_d bias_d bias_a bias_d op VSS m1_n2176_n12171#
+ bias_d VSS bias_a bias_d VSS op bias_d bias_a on bias_d bias_d m1_n1659_n11581#
+ op on VSS bias_d bias_d on bias_d bias_d m1_n2176_n12171# VSS m1_n1659_n11581# bias_d
+ m1_n947_n12836# bias_d VSS bias_a op m1_n947_n12836# bias_d m1_n2176_n12171# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_2 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias
+ bias_c i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_5 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_2 m1_n947_n12836# bias_d VSS bias_d bias_a m1_n1659_n11581#
+ m1_n947_n12836# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# op on bias_d
+ bias_d on on op on bias_d VSS op m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n1659_n11581#
+ bias_d bias_d bias_d VSS m1_n947_n12836# m1_n947_n12836# op VSS m1_n947_n12836#
+ op m1_n1659_n11581# m1_n1659_n11581# bias_d bias_d on bias_d on bias_d m1_n1659_n11581#
+ bias_d bias_d on VSS op VSS VSS op on bias_d bias_d m1_n947_n12836# op op bias_d
+ bias_d bias_d VSS bias_d VSS m1_n1659_n11581# m1_n947_n12836# m1_n2176_n12171# VSS
+ m1_n1659_n11581# bias_d bias_d on VSS m1_n1659_n11581# bias_d m1_n947_n12836# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_3 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias
+ i_bias i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_10 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_11 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_6 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_12 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_7 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_7P4E2J_0 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_KEEN2X_10 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS cmc cmc bias_a VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS cmc bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_13 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_8 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_KEEN2X_11 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS bias_a bias_a cmc VSS m1_n5574_n13620# cmc VSS bias_a bias_a
+ cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS bias_a cmc VSS VSS
+ m1_n5574_n13620# m1_n5574_n13620# bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc
+ VSS VSS bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620#
+ bias_a bias_a cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# bias_a cmc
+ cmc VSS VSS m1_n5574_n13620# bias_a cmc bias_a m1_n5574_n13620# m1_n5574_n13620#
+ VSS cmc bias_a VSS m1_n5574_n13620# bias_a cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_7P4E2J_1 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d bias_a m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_a m1_6690_n8907# bias_a VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_9 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_14 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_7P4E2J_2 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_a
+ m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_7P4E2J_3 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d
+ m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_15 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_KEEN2X_12 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS bias_a bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# bias_a VSS bias_a bias_a VSS
+ VSS m1_n5574_n13620# m1_n5574_n13620# cmc m1_n5574_n13620# VSS cmc bias_a VSS bias_a
+ VSS VSS cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620#
+ bias_a bias_a cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc bias_a
+ bias_a VSS VSS m1_n5574_n13620# cmc cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS
+ cmc bias_a VSS m1_n5574_n13620# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_VJ4JGY_0 cm cm cm cm cm cm cm m1_11534_n9706# m1_11242_n9716#
+ cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# cm cm cm cm VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_1 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490#
+ m1_11534_n9706# m1_11242_n9716# cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711#
+ m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_2 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490#
+ m1_11534_n11258# m1_11244_n11260# cm cm cm cm m1_12410_n11263# m1_12118_n11263#
+ cm m1_11826_n11260# m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_3 cm cm cm cm VSS cm VSS m1_11534_n11258# m1_11244_n11260#
+ cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260# VSS VSS cm VSS
+ VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__pfet_01v8_E4DCBA_0 VDD bias_c m1_6690_n8907# op bias_c bias_c m1_1038_n2886#
+ bias_b bias_c VDD m1_n208_n2883# bias_c VDD on bias_c VDD m1_2463_n5585# VDD VDD
+ m1_2462_n3318# m1_2462_n3318# op m1_2463_n5585# m1_2462_n3318# VDD VDD VDD bias_b
+ bias_c m1_1038_n2886# bias_c m1_6690_n8907# VDD bias_c VDD VDD m1_2463_n5585# on
+ VDD bias_c m1_2462_n3318# m1_n208_n2883# bias_c bias_c VDD VDD m1_2463_n5585# VDD
+ sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_2 on VDD op on VDD bias_c m1_n208_n2883# on bias_c
+ bias_c VDD VDD m1_n208_n2883# op bias_c bias_c m1_1038_n2886# bias_c VDD m1_n208_n2883#
+ m1_n208_n2883# m1_n6302_n3889# m1_1038_n2886# m1_n208_n2883# m1_n6302_n3889# bias_c
+ bias_c on bias_c VDD bias_c op bias_c bias_c cm bias_c m1_1038_n2886# cm m1_1038_n2886#
+ VDD m1_n208_n2883# m1_1038_n2886# bias_c bias_c op bias_c m1_1038_n2886# bias_c
+ sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_1 op VDD on op VDD bias_c m1_1038_n2886# op bias_c
+ bias_c VDD VDD m1_1038_n2886# on bias_c bias_c m1_n208_n2883# bias_c VDD m1_1038_n2886#
+ m1_1038_n2886# m1_n6302_n3889# m1_n208_n2883# m1_1038_n2886# m1_n6302_n3889# bias_c
+ bias_c op bias_c VDD bias_c on bias_c bias_c cm bias_c m1_n208_n2883# cm m1_n208_n2883#
+ VDD m1_1038_n2886# m1_n208_n2883# bias_c bias_c on bias_c m1_n208_n2883# bias_c
+ sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_3 VDD bias_c bias_b on bias_c bias_c m1_n208_n2883#
+ m1_6690_n8907# bias_c VDD m1_1038_n2886# bias_c VDD op bias_c VDD m1_2462_n3318#
+ VDD VDD m1_2463_n5585# m1_2463_n5585# on m1_2462_n3318# m1_2463_n5585# VDD VDD VDD
+ m1_6690_n8907# bias_c m1_n208_n2883# bias_c bias_b VDD bias_c VDD VDD m1_2462_n3318#
+ op VDD bias_c m1_2463_n5585# m1_1038_n2886# bias_c bias_c VDD VDD m1_2462_n3318#
+ VDD sky130_fd_pr__pfet_01v8_E4DCBA
Xsc_cmfb_0 cmc on bias_a p2_b p1 cm VSS p2 VDD op p1_b sc_cmfb
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_0 m1_n208_n2883# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_1038_n2886# VDD VDD VDD bias_b VDD bias_b m1_1038_n2886# bias_b bias_b
+ m1_1038_n2886# bias_b VDD VDD VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b VDD m1_n208_n2883#
+ VDD bias_b sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_4 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS cmc cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS cmc cmc VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# bias_a m1_n5574_n13620# VSS bias_a cmc VSS cmc VSS VSS bias_a bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ bias_a bias_a m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_1 m1_2463_n5585# bias_b m1_2462_n3318# bias_b
+ VDD m1_2463_n5585# bias_b bias_b VDD m1_2462_n3318# VDD bias_b m1_2462_n3318# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2462_n3318# m1_2463_n5585#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2463_n5585#
+ bias_b sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_5 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS VSS bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS VSS bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS VSS VSS cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS m1_n5574_n13620# bias_a
+ bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_3 m1_2462_n3318# bias_b m1_2463_n5585# bias_b
+ VDD m1_2462_n3318# bias_b bias_b VDD m1_2463_n5585# VDD bias_b m1_2463_n5585# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2463_n5585# m1_2462_n3318#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2462_n3318#
+ bias_b sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_2 m1_n6302_n3889# bias_b m1_n6302_n3889# bias_b
+ VDD m1_n6302_n3889# bias_b bias_b VDD m1_n6302_n3889# VDD bias_b m1_n6302_n3889#
+ bias_b VDD bias_b m1_n208_n2883# bias_b bias_b m1_1038_n2886# bias_b m1_n6302_n3889#
+ m1_n6302_n3889# VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b bias_b m1_1038_n2886#
+ m1_n6302_n3889# bias_b sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_6 VSS VSS VSS VSS bias_a bias_a m1_n947_n12836# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n1659_n11581# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n947_n12836# bias_a m1_n1659_n11581# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n1659_n11581# m1_n947_n12836# bias_a bias_a bias_a
+ m1_n1659_n11581# m1_n2176_n12171# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_4 m1_1038_n2886# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_n208_n2883# VDD VDD VDD bias_b VDD bias_b m1_n208_n2883# bias_b bias_b
+ m1_n208_n2883# bias_b VDD VDD VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b VDD m1_1038_n2886#
+ VDD bias_b sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_7 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n947_n12836# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n1659_n11581# m1_n2176_n12171# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n2176_n12171# m1_n1659_n11581# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_KEEN2X_9 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS VSS cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS VSS cmc VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ bias_a bias_a m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a VSS m1_n5574_n13620#
+ cmc cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_KEEN2X_8 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n947_n12836# m1_n947_n12836# bias_a m1_n1659_n11581# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n1659_n11581# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n1659_n11581# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n1659_n11581# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n947_n12836# m1_n2176_n12171# m1_n947_n12836# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
.ends

.subckt sky130_fd_pr__nfet_01v8_E56BNL a_n33_32# a_15_n90# a_n73_n90# VSUBS
X0 a_15_n90# a_n33_32# a_n73_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt switch_5t out en_b en VDD in VSS
Xtransmission_gate_0 transmission_gate_1/in en_b en VSS VDD in transmission_gate
Xtransmission_gate_1 out en_b en VSS VDD transmission_gate_1/in transmission_gate
Xsky130_fd_pr__nfet_01v8_E56BNL_0 en_b transmission_gate_1/in VSS VSS sky130_fd_pr__nfet_01v8_E56BNL
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
.ends

.subckt a_mux2_en en s0 in0 VDD out VSS in1
Xswitch_5t_0 out switch_5t_1/en s0 VDD switch_5t_0/in VSS switch_5t
Xswitch_5t_1 out s0 switch_5t_1/en VDD switch_5t_1/in VSS switch_5t
Xtransmission_gate_0 switch_5t_1/in transmission_gate_1/en_b en VSS VDD in0 transmission_gate
Xtransmission_gate_1 switch_5t_0/in transmission_gate_1/en_b en VSS VDD in1 transmission_gate
Xsky130_fd_sc_hd__inv_1_0 transmission_gate_1/en_b en VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_1 switch_5t_1/en s0 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VPWR X VNB VPB
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=6.142e+11p pd=7.3e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=7.039e+11p ps=8e+06u w=420000u l=150000u
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=2.7965e+11p ps=3.21e+06u w=420000u l=150000u
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.8025e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=150000u
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_XAYTAL a_n129_n203# a_n173_n100# w_n311_n319#
X0 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=1.28e+12p pd=1.056e+07u as=0p ps=0u w=1e+06u l=150000u
X1 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VPWR X VNB VPB
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=6.517e+11p ps=5.37e+06u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=4.027e+11p pd=3.97e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__dfxbp_1 CLK D VGND VPWR Q Q_N VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=9.432e+11p ps=1.006e+07u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.32905e+12p pd=1.228e+07u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X6 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1059_315# a_1490_369# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X17 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23 Q_N a_1490_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q_N a_1490_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 VPWR a_1059_315# a_1490_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
.ends

.subckt clock_v2 clk p2d_b p2d p2_b p2 p1d_b p1d p1_b p1 Ad_b Ad A_b A Bd_b Bd B_b
+ B VDD VSS
Xsky130_fd_sc_hd__clkbuf_16_11 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD p1d_b VSS VDD
+ sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_248 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_237 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_226 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_215 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_204 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_12 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD p2d_b VSS VDD
+ sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_249 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_238 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_227 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_216 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_205 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_13 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD p2d VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_239 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_228 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_217 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_0 sky130_fd_sc_hd__clkinv_1_0/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_14 sky130_fd_sc_hd__clkinv_4_10/Y VSS VDD p2_b VSS VDD
+ sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_10 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_4_10/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_229 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_218 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_207 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_1 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_140 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_162 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_15 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD p2 VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_11 sky130_fd_sc_hd__nand2_4_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_219 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_208 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_2 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_209 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_3 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS VDD sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/A
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_165 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_2 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__nand2_4_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_190 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_5 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_111 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_166 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_180 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_4_3 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_6 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_168 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_157 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_193 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_160 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_171 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_182 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_8 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_4_4/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_158 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_150 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_161 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_172 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_183 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_194 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_5/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_159 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_195 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_140 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_162 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_6 sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/A
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_190 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_196 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_141 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_130 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_152 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_185 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_90 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_7 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_191 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_180 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_142 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_186 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_80 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_8 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__clkinv_4_8/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_121 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_110 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_143 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_132 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_154 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_165 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_198 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_187 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_92 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_9 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__clkinv_4_9/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_193 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_182 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_81 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_100 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_122 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_111 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_133 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_166 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_199 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_188 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_71 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_82 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_93 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_0 p2 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__mux2_1_0/S
+ sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS VDD sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_93 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_172 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_82 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_150 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_112 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_145 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_134 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_167 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_178 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_189 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_50 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_61 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_1 clk sky130_fd_sc_hd__dfxbp_1_1/D VSS VDD sky130_fd_sc_hd__nand2_1_1/A
+ sky130_fd_sc_hd__dfxbp_1_1/D VSS VDD sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_94 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_61 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_50 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_195 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_184 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_173 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_140 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_83 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_162 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_102 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_146 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_157 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_168 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_179 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_73 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_84 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_95 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_95 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_73 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_62 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_141 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_196 sky130_fd_sc_hd__clkinv_1_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_174 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_152 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_163 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_103 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_125 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_114 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_158 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_169 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_52 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_63 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_96 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_41 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_197 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_186 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_164 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_131 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_142 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD B VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_115 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_137 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_126 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_148 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_159 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_42 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_20 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_31 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_75 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_86 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_97 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_1/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_64 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_53 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_198 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_187 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_121 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_86 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_132 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_154 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD Bd VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_105 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_138 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_127 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_149 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_10 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_54 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_32 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_65 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_87 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_10 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_21 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_76 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_43 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_199 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_3/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_177 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_100 sky130_fd_sc_hd__clkinv_1_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_122 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD
+ sky130_fd_sc_hd__nand2_1_4/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_32 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD B_b VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_139 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_22 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_44 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_11 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_77 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_99 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_11 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_66 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_55 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_44 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_178 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_167 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_112 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_101 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_22 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_88 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_123 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_134 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD Bd_b VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_118 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_129 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_56 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_34 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_67 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_78 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_89 sky130_fd_sc_hd__clkinv_1_1/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A
+ VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_56 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_78 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_34 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_157 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_102 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_89 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_113 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_146 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_168 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_4 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD Ad_b VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_24 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_13 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_68 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_0/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_46 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_35 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_169 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_2/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_103 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_2/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_125 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_136 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_147 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_158 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_5 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD Ad VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_109 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_25 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_47 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_58 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_36 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_69 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_69 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_58 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_104 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_159 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_6 sky130_fd_sc_hd__clkinv_4_4/Y VSS VDD A_b VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_15 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_48 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_59 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_59 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_48 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_26 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_116 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_127 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_138 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_37 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_149 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_7 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD A VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_49 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_1/B VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_27 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_38 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_250 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_49 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_117 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_27 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_8 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD p1 VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_17 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_39 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_251 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_240 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_107 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_118 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_129 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_9 sky130_fd_sc_hd__clkinv_4_7/Y VSS VDD p1_b VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_1_0/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_18 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_29 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_252 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_241 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_230 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_18 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_108 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_1_1/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_253 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_242 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_231 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_220 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_109 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_1_3/A clk VSS VDD sky130_fd_sc_hd__nand2_4_3/A
+ VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_1_2/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_254 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_243 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_232 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_221 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_210 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/B
+ VSS VDD sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_255 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_244 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_233 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_222 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_211 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_200 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux2_1_0 Ad_b Bd_b sky130_fd_sc_hd__mux2_1_0/S VSS VDD sky130_fd_sc_hd__mux2_1_0/X
+ VSS VDD sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1_3/A
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_245 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_234 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_223 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_212 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_201 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_246 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_235 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_224 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_213 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_202 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_30 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_10 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD p1d VSS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_6 clk VSS VDD sky130_fd_sc_hd__nand2_1_2/A VSS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_247 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_236 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_225 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_214 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_203 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
.ends

.subckt sky130_fd_pr__nfet_01v8_E56BNL_AA a_n72_n90# a_16_n90# a_n32_32# VSUBS
X0 a_16_n90# a_n32_32# a_n72_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
.ends

.subckt switch_5t_AA out en_b en VDD in VSS
Xtransmission_gate_0 transmission_gate_1/in en_b en VSS VDD in transmission_gate
Xtransmission_gate_1 out en_b en VSS VDD transmission_gate_1/in transmission_gate
Xsky130_fd_pr__nfet_01v8_E56BNL_0 VSS transmission_gate_1/in en_b VSS sky130_fd_pr__nfet_01v8_E56BNL_AA
.ends

.subckt a_mux4_en s1 s0 in0 in2 in3 out en VSS in1 VDD
Xsky130_fd_sc_hd__inv_1_4 switch_5t_0/en switch_5t_0/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_5 switch_5t_2/en switch_5t_2/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_0 out switch_5t_0/en_b switch_5t_0/en VDD switch_5t_0/in VSS switch_5t_AA
Xsky130_fd_sc_hd__inv_1_6 switch_5t_3/en switch_5t_3/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_1 out switch_5t_1/en_b switch_5t_1/en VDD switch_5t_1/in VSS switch_5t_AA
Xsky130_fd_sc_hd__inv_1_8 transmission_gate_3/en_b en VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_2 out switch_5t_2/en_b switch_5t_2/en VDD switch_5t_2/in VSS switch_5t_AA
Xswitch_5t_3 out switch_5t_3/en_b switch_5t_3/en VDD switch_5t_3/in VSS switch_5t_AA
Xtransmission_gate_0 switch_5t_0/in transmission_gate_3/en_b en VSS VDD in0 transmission_gate
Xtransmission_gate_1 switch_5t_1/in transmission_gate_3/en_b en VSS VDD in1 transmission_gate
Xtransmission_gate_2 switch_5t_2/in transmission_gate_3/en_b en VSS VDD in2 transmission_gate
Xtransmission_gate_3 switch_5t_3/in transmission_gate_3/en_b en VSS VDD in3 transmission_gate
Xsky130_fd_sc_hd__nand2_1_0 s0 s1 VSS VDD switch_5t_3/en_b VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_1 s0 sky130_fd_sc_hd__inv_1_0/Y VSS VDD switch_5t_2/en_b
+ VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_2 s1 sky130_fd_sc_hd__inv_1_1/Y VSS VDD switch_5t_1/en_b
+ VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/Y
+ VSS VDD switch_5t_0/en_b VSS VDD sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/Y s0 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y s1 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 switch_5t_1/en switch_5t_1/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TABSMU c1_n1210_n1160# m3_n1310_n1260#
X0 c1_n1210_n1160# m3_n1310_n1260# sky130_fd_pr__cap_mim_m3_1 l=1.16e+07u w=1.16e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_VCQUSW a_n810_n632# a_1802_n632# a_n4080_n100# a_2640_n100#
+ a_2010_n100# a_3852_131# a_n3750_n632# a_n3120_n632# a_3600_n632# a_2594_n401# a_n88_n632#
+ a_n2866_n401# a_n2912_n100# a_n718_n632# a_n556_n729# a_2548_n100# a_n182_n100#
+ a_n3658_n632# a_n3028_n632# a_n3496_n729# a_2012_n632# a_2642_n632# a_n1140_n100#
+ a_n1770_n100# a_n1398_n197# a_2172_131# a_n812_n100# a_n4128_131# a_3224_n729# a_n766_n401#
+ a_3480_n100# a_n3122_n100# a_n3752_n100# a_240_n632# a_870_n632# a_n2448_131# a_3388_n100#
+ a_3434_n401# a_n3706_n401# a_3482_n632# a_492_131# a_1500_n632# a_4064_n729# a_n1650_n632#
+ a_n1020_n632# a_n768_131# a_n2238_n197# a_n1558_n632# a_n2610_n100# a_n1396_n729#
+ w_n4520_n851# a_750_n100# a_120_n100# a_1124_n729# a_n2490_n632# a_2340_n632# a_2970_n632#
+ a_1380_n100# a_658_n100# a_n510_n100# a_n1022_n100# a_n1652_n100# a_n138_n197# a_1288_n100#
+ a_n3450_n100# a_n3078_n197# a_n2398_n632# a_122_n632# a_752_n632# a_1334_n401# a_74_n401#
+ a_702_n197# a_1382_n632# a_n1606_n401# a_1962_n197# a_3012_131# a_n390_n632# a_1918_n100#
+ a_28_n100# a_3180_n632# a_n2492_n100# a_1332_131# a_n2236_n729# a_n298_n632# a_3810_n632#
+ a_2850_n100# a_2220_n100# a_n3960_n632# a_n3330_n632# a_2174_n401# a_n1608_131#
+ a_n928_n632# a_n2446_n401# a_n136_n729# a_n3868_n632# a_n3238_n632# a_2758_n100#
+ a_2128_n100# a_n392_n100# a_n3076_n729# a_2802_n197# a_2222_n632# a_2852_n632# a_n1350_n100#
+ a_n1980_n100# a_n4170_n632# a_4020_n632# a_n346_n401# a_3690_n100# a_3060_n100#
+ a_n3332_n100# a_n3962_n100# a_2592_131# a_450_n632# a_n3286_n401# a_3598_n100# a_n4078_n632#
+ a_1080_n632# a_3014_n401# a_n2868_131# a_3062_n632# a_3692_n632# a_n2190_n100# a_3642_n197#
+ a_n1860_n632# a_n1230_n632# a_1710_n632# a_n4172_n100# a_n2820_n100# a_n1768_n632#
+ a_n1138_n632# a_n1188_131# a_704_n729# a_n4126_n401# a_960_n100# a_330_n100# a_1964_n729#
+ a_1590_n100# a_282_n197# a_n2070_n632# a_2550_n632# a_n90_n100# a_n978_n197# a_n1186_n401#
+ a_868_n100# a_238_n100# a_n720_n100# a_n1232_n100# a_n1862_n100# a_914_n401# a_1498_n100#
+ a_n3030_n100# a_n3660_n100# a_n2700_n632# a_332_n632# a_962_n632# a_1542_n197# a_1592_n632#
+ a_n3918_n197# a_n2608_n632# a_3390_n632# a_n2072_n100# a_3432_131# a_n600_n632#
+ a_1752_131# a_2804_n729# a_n3540_n632# a_2430_n100# a_n2702_n100# a_n3708_131# a_n508_n632#
+ a_n2026_n401# a_2382_n197# a_2968_n100# a_2338_n100# a_n976_n729# a_n3448_n632#
+ a_n1560_n100# a_2432_n632# a_3644_n729# a_3270_n100# a_n602_n100# a_n2028_131# a_n3916_n729#
+ a_n3542_n100# a_660_n632# a_n1818_n197# a_3178_n100# a_1290_n632# a_3900_n100# a_3854_n401#
+ a_3222_n197# a_3272_n632# a_n348_131# a_30_n632# a_3808_n100# a_n1440_n632# a_1920_n632#
+ a_284_n729# a_n2658_n197# a_3902_n632# a_n2400_n100# a_n1978_n632# a_n1348_n632#
+ a_n3288_131# a_4110_n100# a_494_n401# a_540_n100# a_4062_n197# a_4018_n100# a_1544_n729#
+ a_n2280_n632# a_2130_n632# a_2760_n632# a_1170_n100# a_72_131# a_n300_n100# a_n930_n100#
+ a_n1442_n100# a_n558_n197# a_n1816_n729# a_448_n100# a_n3240_n100# a_n3870_n100#
+ a_n3498_n197# a_n2188_n632# a_4112_n632# a_1078_n100# a_1754_n401# a_1800_n100#
+ a_n2910_n632# a_542_n632# a_1122_n197# a_n180_n632# a_1172_n632# a_2384_n729# a_n2818_n632#
+ a_1708_n100# a_912_131# a_n2656_n729# a_n2282_n100#
X0 a_n90_n100# a_n138_n197# a_n182_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_330_n100# a_282_n197# a_238_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2 a_n3868_n632# a_n3916_n729# a_n3960_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X3 a_n1348_n632# a_n1396_n729# a_n1440_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X4 a_n3450_n100# a_n3498_n197# a_n3542_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X5 a_3480_n100# a_3432_131# a_3388_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X6 a_3062_n632# a_3014_n401# a_2970_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X7 a_542_n632# a_494_n401# a_450_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X8 a_2432_n632# a_2384_n729# a_2340_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X9 a_n1770_n100# a_n1818_n197# a_n1862_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X10 a_1800_n100# a_1752_131# a_1708_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X11 a_n508_n632# a_n556_n729# a_n600_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X12 a_1592_n632# a_1544_n729# a_1500_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X13 a_2222_n632# a_2174_n401# a_2130_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X14 a_540_n100# a_492_131# a_448_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X15 a_2220_n100# a_2172_131# a_2128_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X16 a_n3660_n100# a_n3708_131# a_n3752_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X17 a_n300_n100# a_n348_131# a_n392_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X18 a_3690_n100# a_3642_n197# a_3598_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X19 a_n3028_n632# a_n3076_n729# a_n3120_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X20 a_n2398_n632# a_n2446_n401# a_n2490_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X21 a_4110_n100# a_4062_n197# a_4018_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X22 a_n1558_n632# a_n1606_n401# a_n1650_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X23 a_n1980_n100# a_n2028_131# a_n2072_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X24 a_2010_n100# a_1962_n197# a_1918_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X25 a_3272_n632# a_3224_n729# a_3180_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X26 a_n510_n100# a_n558_n197# a_n602_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X27 a_750_n100# a_702_n197# a_658_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X28 a_752_n632# a_704_n729# a_660_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X29 a_2642_n632# a_2594_n401# a_2550_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X30 a_n3870_n100# a_n3918_n197# a_n3962_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X31 a_3900_n100# a_3852_131# a_3808_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X32 a_n4078_n632# a_n4126_n401# a_n4170_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X33 a_n718_n632# a_n766_n401# a_n810_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X34 a_1802_n632# a_1754_n401# a_1710_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X35 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=2.48e+12p pd=2.096e+07u as=0p ps=0u w=1e+06u l=150000u
X36 a_n3238_n632# a_n3286_n401# a_n3330_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X37 a_n2608_n632# a_n2656_n729# a_n2700_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X38 a_n2190_n100# a_n2238_n197# a_n2282_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X39 a_n720_n100# a_n768_131# a_n812_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X40 a_960_n100# a_912_131# a_868_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X41 a_n1768_n632# a_n1816_n729# a_n1860_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X42 a_4112_n632# a_4064_n729# a_4020_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X43 a_n4080_n100# a_n4128_131# a_n4172_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X44 a_2852_n632# a_2804_n729# a_2760_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X45 a_3482_n632# a_3434_n401# a_3390_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X46 a_962_n632# a_914_n401# a_870_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X47 a_n2400_n100# a_n2448_131# a_n2492_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X48 a_2430_n100# a_2382_n197# a_2338_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X49 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n928_n632# a_n976_n729# a_n1020_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X51 a_122_n632# a_74_n401# a_30_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X52 a_2012_n632# a_1964_n729# a_1920_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X53 a_n3448_n632# a_n3496_n729# a_n3540_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X54 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_n930_n100# a_n978_n197# a_n1022_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X56 a_n2818_n632# a_n2866_n401# a_n2910_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X57 a_n1140_n100# a_n1188_131# a_n1232_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X58 a_1170_n100# a_1122_n197# a_1078_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X59 a_n88_n632# a_n136_n729# a_n180_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X60 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n2610_n100# a_n2658_n197# a_n2702_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X62 a_2640_n100# a_2592_131# a_2548_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X63 a_1172_n632# a_1124_n729# a_1080_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X64 a_3692_n632# a_3644_n729# a_3600_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X65 a_n3030_n100# a_n3078_n197# a_n3122_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X66 a_3060_n100# a_3012_131# a_2968_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X67 a_n1978_n632# a_n2026_n401# a_n2070_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X68 a_n3658_n632# a_n3706_n401# a_n3750_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X69 a_n1138_n632# a_n1186_n401# a_n1230_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X70 a_n1350_n100# a_n1398_n197# a_n1442_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X71 a_1380_n100# a_1332_131# a_1288_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X72 a_n2820_n100# a_n2868_131# a_n2912_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X73 a_2850_n100# a_2802_n197# a_2758_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X74 a_332_n632# a_284_n729# a_240_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X75 a_n3240_n100# a_n3288_131# a_n3332_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X76 a_3270_n100# a_3222_n197# a_3178_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X77 a_n298_n632# a_n346_n401# a_n390_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X78 a_1382_n632# a_1334_n401# a_1290_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X79 a_3902_n632# a_3854_n401# a_3810_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X80 a_n1560_n100# a_n1608_131# a_n1652_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X81 a_120_n100# a_72_131# a_28_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X82 a_1590_n100# a_1542_n197# a_1498_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X83 a_n2188_n632# a_n2236_n729# a_n2280_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt latch_pmos_pair sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
Xsky130_fd_pr__pfet_01v8_VCQUSW_0 sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100# sky130_fd_pr__pfet_01v8_VCQUSW
.ends

.subckt sky130_fd_pr__pfet_01v8_VCG74W a_543_n100# a_159_n100# a_n609_n100# a_495_n197#
+ a_n705_n100# a_255_n100# a_n657_n197# a_n369_131# a_351_n100# a_n417_n100# a_n801_n100#
+ a_303_n197# a_n129_n100# a_n513_n100# a_n465_n197# a_n561_131# a_63_n100# a_n225_n100#
+ a_399_131# a_111_n197# a_n321_n100# a_n273_n197# a_15_131# a_n753_131# a_639_n100#
+ w_n1031_n319# a_591_131# a_207_131# a_735_n100# a_n33_n100# a_687_n197# a_447_n100#
+ a_n81_n197# a_n177_131#
X0 a_63_n100# a_15_131# a_n33_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n129_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_255_n100# a_207_131# a_159_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_351_n100# a_303_n197# a_255_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_543_n100# a_495_n197# a_447_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 w_n1031_n319# w_n1031_n319# a_735_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=5.24e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_159_n100# a_111_n197# a_63_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_447_n100# a_399_131# a_351_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_639_n100# a_591_131# a_543_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_735_n100# a_687_n197# a_639_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n801_n100# w_n1031_n319# w_n1031_n319# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_n513_n100# a_n561_131# a_n609_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_n321_n100# a_n369_131# a_n417_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_n225_n100# a_n273_n197# a_n321_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_n705_n100# a_n753_131# a_n801_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_n609_n100# a_n657_n197# a_n705_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n417_n100# a_n465_n197# a_n513_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n129_n100# a_n177_131# a_n225_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
.ends

.subckt precharge_pmos sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131#
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ sky130_fd_pr__pfet_01v8_VCG74W
.ends

.subckt current_tail a_543_n100# a_159_n100# a_n609_n100# a_n1569_n100# a_n705_n100#
+ a_255_n100# a_1407_n100# a_351_n100# a_n417_n100# a_n801_n100# a_1503_n100# a_1119_n100#
+ a_n1377_n100# a_n129_n100# a_n513_n100# a_1215_n100# a_63_n100# a_n1089_n100# a_n1473_n100#
+ a_n225_n100# a_1311_n100# a_927_n100# a_n1185_n100# a_n321_n100# a_1023_n100# a_639_n100#
+ a_n1281_n100# a_735_n100# a_n33_n100# a_n897_n100# a_831_n100# a_447_n100# a_n1521_122#
+ a_n993_n100# a_n1763_n274#
X0 a_n801_n100# a_n1521_122# a_n897_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n513_n100# a_n1521_122# a_n609_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n321_n100# a_n1521_122# a_n417_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n225_n100# a_n1521_122# a_n321_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_n897_n100# a_n1521_122# a_n993_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 a_n705_n100# a_n1521_122# a_n801_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n609_n100# a_n1521_122# a_n705_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n417_n100# a_n1521_122# a_n513_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n129_n100# a_n1521_122# a_n225_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_63_n100# a_n1521_122# a_n33_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_927_n100# a_n1521_122# a_831_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11 a_1023_n100# a_n1521_122# a_927_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1569_n100# a_n1763_n274# a_n1763_n274# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=6.2e+11p ps=5.24e+06u w=1e+06u l=150000u
X13 a_1119_n100# a_n1521_122# a_1023_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_1215_n100# a_n1521_122# a_1119_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_1311_n100# a_n1521_122# a_1215_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_1407_n100# a_n1521_122# a_1311_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_1503_n100# a_n1521_122# a_1407_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1763_n274# a_n1763_n274# a_1503_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n33_n100# a_n1521_122# a_n129_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_351_n100# a_n1521_122# a_255_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X21 a_159_n100# a_n1521_122# a_63_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22 a_255_n100# a_n1521_122# a_159_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_447_n100# a_n1521_122# a_351_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X24 a_543_n100# a_n1521_122# a_447_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X25 a_639_n100# a_n1521_122# a_543_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_735_n100# a_n1521_122# a_639_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_831_n100# a_n1521_122# a_735_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n1473_n100# a_n1521_122# a_n1569_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X29 a_n1377_n100# a_n1521_122# a_n1473_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X30 a_n1281_n100# a_n1521_122# a_n1377_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X31 a_n1185_n100# a_n1521_122# a_n1281_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X32 a_n1089_n100# a_n1521_122# a_n1185_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X33 a_n993_n100# a_n1521_122# a_n1089_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_J3WY8C a_n4080_n100# a_n1188_122# a_282_n188# a_n978_n188#
+ a_1542_n188# a_n3918_n188# a_3432_122# a_1752_122# a_n3708_122# a_2382_n188# a_4228_n100#
+ a_n2028_122# a_n1818_n188# a_3222_n188# a_n348_122# a_n2658_n188# a_n3288_122# a_4062_n188#
+ a_72_122# a_n558_n188# a_n3498_n188# a_1122_n188# a_912_122# a_n4172_n100# a_3852_122#
+ a_n1398_n188# a_2172_122# a_n4128_122# a_n2448_122# a_492_122# a_n768_122# a_n2238_n188#
+ a_n138_n188# a_n3078_n188# a_1962_n188# a_702_n188# a_3012_122# a_1332_122# a_n1608_122#
+ a_n4382_n100# a_2802_n188# a_2592_122# a_3642_n188# a_n2868_122# VSUBS
X0 a_n4080_n100# a_n1398_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=1.24e+13p pd=1.048e+08u as=1.24e+13p ps=1.048e+08u w=1e+06u l=150000u
X1 a_n4080_n100# a_1332_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n4080_n100# a_n2868_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n4080_n100# a_2802_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n4080_n100# a_n3288_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n4080_n100# a_3222_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n4080_n100# a_72_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n4080_n100# a_n1608_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n4080_n100# a_1542_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n4080_n100# a_n138_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n4080_n100# a_282_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n4080_n100# a_n3498_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n4080_n100# a_3432_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n4080_n100# a_n1818_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n4080_n100# a_1752_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n4080_n100# a_492_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n4080_n100# a_2172_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n4080_n100# a_n3708_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n4080_n100# a_n348_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n4080_n100# a_3642_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n4080_n100# a_4062_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n4080_n100# a_n2028_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n4080_n100# a_1962_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n4080_n100# a_702_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n4080_n100# a_n3918_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n4080_n100# a_n558_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n4080_n100# a_3852_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_4228_n100# a_4228_n100# a_4228_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X28 a_n4080_n100# a_n2238_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_n4080_n100# a_n768_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n4080_n100# a_912_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n4080_n100# a_n4128_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_n4080_n100# a_n2448_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_n4080_n100# a_2382_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_n4080_n100# a_n978_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n4382_n100# a_n4382_n100# a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X36 a_n4080_n100# a_n1188_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_n4080_n100# a_1122_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n4080_n100# a_n2658_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_n4080_n100# a_2592_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_n4080_n100# a_n3078_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_n4080_n100# a_3012_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt latch_nmos_pair sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
.ends

.subckt input_diff_pair sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_4 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_5 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_6 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_7 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
.ends

.subckt comparator_v2 outp outn ip VDD VSS in clk
Xlatch_pmos_pair_0 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD VDD VDD
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD latch_pmos_pair
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__buf_2_1/X outp VSS VDD outn VSS VDD sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__buf_2_0/X outn VSS VDD outp VSS VDD sky130_fd_sc_hd__nand2_4
Xsky130_fd_pr__pfet_01v8_VCG74W_1 li_940_3458# li_940_3458# li_940_3458# clk VDD VDD
+ clk clk li_940_3458# li_940_3458# li_940_3458# clk VDD VDD clk clk VDD li_940_3458#
+ clk clk VDD clk clk clk VDD VDD clk clk li_940_3458# li_940_3458# clk VDD clk clk
+ sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk VDD sky130_fd_sc_hd__buf_2_1/A clk
+ clk VDD clk clk clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ clk VDD clk clk sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_sc_hd__buf_2_0 sky130_fd_sc_hd__buf_2_0/A VSS VDD sky130_fd_sc_hd__buf_2_0/X
+ VSS VDD sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_1 sky130_fd_sc_hd__buf_2_1/A VSS VDD sky130_fd_sc_hd__buf_2_1/X
+ VSS VDD sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_0 clk sky130_fd_sc_hd__buf_2_0/A clk VDD VDD clk sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A clk sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A clk clk VDD VDD clk clk clk sky130_fd_sc_hd__buf_2_0/A
+ clk clk clk clk precharge_pmos
Xcurrent_tail_0 li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# VSS VSS VSS
+ li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS VSS VSS li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS li_n2324_818# li_n2324_818# VSS VSS VSS clk li_n2324_818# VSS current_tail
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_1 clk li_940_818# clk VDD VDD clk li_940_818# li_940_818# li_940_818#
+ clk li_940_818# VDD VDD clk VDD VDD clk clk li_940_818# VDD li_940_818# li_940_818#
+ clk clk VDD VDD clk clk clk li_940_818# clk clk clk clk precharge_pmos
Xlatch_nmos_pair_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A latch_nmos_pair
Xinput_diff_pair_0 ip ip ip in in VSS ip in in in in VSS li_940_3458# ip ip ip in
+ ip li_n2324_818# ip ip in ip ip ip in in in ip ip ip in ip in ip in ip in in ip
+ ip VSS ip ip in ip li_n2324_818# ip ip in in in ip ip ip in in in li_940_3458# in
+ in ip ip in ip in ip ip ip VSS ip in ip ip ip in in in ip ip in in ip in VSS ip
+ in in in in in ip in li_940_818# ip ip in ip ip li_n2324_818# in in ip ip ip in
+ ip ip ip ip in in in in in in VSS ip in in ip ip ip ip ip in in ip ip in in ip li_940_818#
+ ip ip in li_n2324_818# in in in VSS ip in in ip ip ip in ip ip ip in in ip in ip
+ in ip ip ip in in in in in VSS in ip li_n2324_818# ip ip in ip ip in ip ip in ip
+ ip li_940_3458# in in ip ip ip in in in ip ip in ip ip in in in VSS ip in VSS VSS
+ in in ip ip in in ip ip ip in in ip ip li_940_3458# in ip in ip ip in li_n2324_818#
+ ip in in in in in in ip ip in in ip ip ip ip VSS ip ip ip in in in in ip ip in ip
+ ip ip in in ip ip in in ip in in li_n2324_818# in in in in ip in in ip in ip li_940_818#
+ VSS ip ip ip ip in in ip ip VSS in in in ip in in ip ip ip in in ip in in VSS in
+ in li_n2324_818# ip in in in ip ip ip ip in in ip ip li_940_818# in ip ip in in
+ in ip in ip in ip ip ip in in in ip ip ip ip in in in ip ip in in in in ip VSS VSS
+ in in ip ip in in in input_diff_pair
.ends

.subckt sky130_fd_pr__nfet_01v8_CFEPS5 a_n275_n238# a_n129_n152# a_n173_n64#
X0 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=8.32e+11p pd=7.76e+06u as=0p ps=0u w=650000u l=150000u
X1 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt analog_top ip in rst_n i_bias_1 i_bias_2 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1
+ debug op a_probe_0 a_probe_1 a_probe_2 a_probe_3 clk d_probe_0 d_probe_1 d_probe_2
+ d_probe_3 d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1
+ VDD VSS
Xesd_cell_5 a_probe_0 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_2 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_18 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_29 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_20 ota_1/cm ota_1/p1_b ota_1/p1 VSS VDD transmission_gate_21/in
+ transmission_gate
Xtransmission_gate_31 transmission_gate_31/out clock_v2_0/p1d_b clock_v2_0/p1d VSS
+ VDD ip transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_70 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_19 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_21 ota_1/in ota_1/p2_b ota_1/p2 VSS VDD transmission_gate_21/in
+ transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_3 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_10 transmission_gate_5/in rst_n transmission_gate_26/en VSS VDD
+ ota_w_test_0/cm transmission_gate
Xesd_cell_6 a_probe_3 VSS VDD esd_cell
Xtransmission_gate_32 transmission_gate_32/out clock_v2_0/p1d_b clock_v2_0/p1d VSS
+ VDD in transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_71 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_60 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_4 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_22 ota_1/ip ota_1/p2_b ota_1/p2 VSS VDD transmission_gate_23/in
+ transmission_gate
Xtransmission_gate_11 transmission_gate_6/in rst_n transmission_gate_26/en VSS VDD
+ ota_w_test_0/cm transmission_gate
Xota_w_test_0 ota_w_test_0/ip ota_w_test_0/in ota_1/p1 ota_w_test_0/op i_bias_1 ota_w_test_0/cm
+ a_mux4_en_0/in0 a_mux4_en_1/in1 a_mux4_en_0/in1 a_mux4_en_0/in2 a_mux4_en_1/in2
+ VDD VSS ota_w_test_0/on ota_1/p2_b ota_1/p1_b ota_1/p2 ota_w_test
Xesd_cell_7 a_probe_2 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_50 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_61 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_23 ota_1/cm ota_1/p1_b ota_1/p1 VSS VDD transmission_gate_23/in
+ transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_5 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_12 a_mux2_en_0/in0 clock_v2_0/Ad_b clock_v2_0/Ad VSS VDD ota_w_test_0/op
+ transmission_gate
Xsky130_fd_sc_hd__clkinv_16_0 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD d_probe_3 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_51 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_62 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_40 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_6 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_24 ota_1/ip rst_n transmission_gate_26/en VSS VDD ota_1/cm transmission_gate
Xtransmission_gate_13 a_mux2_en_0/in1 clock_v2_0/Bd_b clock_v2_0/Bd VSS VDD ota_w_test_0/op
+ transmission_gate
Xsky130_fd_sc_hd__clkinv_16_1 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD d_probe_2 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_52 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_63 transmission_gate_21/in transmission_gate_19/out
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_30 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_41 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_25 ota_1/in rst_n transmission_gate_26/en VSS VDD ota_1/cm transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_7 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_14 a_mux2_en_0/in0 clock_v2_0/Bd_b clock_v2_0/Bd VSS VDD ota_w_test_0/on
+ transmission_gate
Xsky130_fd_sc_hd__clkinv_16_2 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD d_probe_1 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_20 transmission_gate_23/in transmission_gate_32/out
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_64 transmission_gate_21/in transmission_gate_31/out
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_31 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_42 sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_53 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_0 rst_n VSS VDD transmission_gate_26/en VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_26 ota_1/op rst_n transmission_gate_26/en VSS VDD ota_1/on transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_8 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_15 a_mux2_en_0/in1 clock_v2_0/Ad_b clock_v2_0/Ad VSS VDD ota_w_test_0/on
+ transmission_gate
Xsky130_fd_sc_hd__clkinv_16_3 sky130_fd_sc_hd__clkinv_4_4/Y VSS VDD d_probe_0 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_65 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_21 transmission_gate_23/in transmission_gate_19/in
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_43 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_10 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_32 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_54 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__mux4_1_0/X VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_9 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_27 transmission_gate_31/out clock_v2_0/p2d_b clock_v2_0/p2d VSS
+ VDD onebit_dac_1/out transmission_gate
Xtransmission_gate_16 a_mux2_en_0/in0 rst_n transmission_gate_26/en VSS VDD a_mux2_en_0/in1
+ transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_22 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_11 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_66 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_44 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_55 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_33 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__mux4_1_1/X VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_28 transmission_gate_0/out clock_v2_0/p2d_b clock_v2_0/p2d VSS
+ VDD onebit_dac_1/out transmission_gate
Xtransmission_gate_17 transmission_gate_19/out clock_v2_0/p1d_b clock_v2_0/p1d VSS
+ VDD a_mux2_en_0/in0 transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_67 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_12 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_45 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_34 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_23 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_56 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xonebit_dac_0 onebit_dac_1/v_b onebit_dac_0/out VDD VSS op VSS VDD onebit_dac
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__mux4_1_2/X VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_29 transmission_gate_32/out clock_v2_0/p2d_b clock_v2_0/p2d VSS
+ VDD onebit_dac_0/out transmission_gate
Xtransmission_gate_18 transmission_gate_19/in clock_v2_0/p1d_b clock_v2_0/p1d VSS
+ VDD a_mux2_en_0/in1 transmission_gate
Xota_1 ota_1/ip ota_1/in ota_1/op i_bias_2 ota_1/cm VSS ota_1/on ota_1/p2_b VDD ota_1/p1_b
+ ota_1/p2 ota_1/p1 ota
Xa_mux2_en_0 debug a_mod_grp_ctrl_0 a_mux2_en_0/in0 VDD a_probe_0 VSS a_mux2_en_0/in1
+ a_mux2_en
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_13 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_68 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_46 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_57 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_24 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xonebit_dac_1 onebit_dac_1/v_b onebit_dac_1/out VSS VDD op VSS VDD onebit_dac
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_35 sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__mux4_1_3/X VSS VDD sky130_fd_sc_hd__clkinv_4_4/Y
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_19 transmission_gate_19/out clock_v2_0/p2d_b clock_v2_0/p2d VSS
+ VDD transmission_gate_19/in transmission_gate
Xa_mux2_en_1 debug a_mod_grp_ctrl_0 ota_1/op VDD a_probe_1 VSS ota_1/on a_mux2_en
Xsky130_fd_sc_hd__mux4_1_0 clock_v2_0/p2d clock_v2_0/Bd clock_v2_0/p2d_b clock_v2_0/Bd_b
+ d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_0/X VSS VDD
+ sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_69 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_47 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_58 transmission_gate_21/in transmission_gate_19/out
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_14 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_25 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__pfet_01v8_hvt_XAYTAL_0 onebit_dac_1/v_b VDD VDD sky130_fd_pr__pfet_01v8_hvt_XAYTAL
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_36 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_2 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__mux4_1_1 clock_v2_0/p1d clock_v2_0/Ad clock_v2_0/p1d_b clock_v2_0/Ad_b
+ d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_1/X VSS VDD
+ sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_26 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_48 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_15 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_59 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_3 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_37 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__mux4_1_2 ota_1/p2 clock_v2_0/B ota_1/p2_b clock_v2_0/B_b d_clk_grp_1_ctrl_0
+ d_clk_grp_1_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_2/X VSS VDD sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_27 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_49 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_16 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_38 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_4 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_0 transmission_gate_0/out clock_v2_0/p1d_b clock_v2_0/p1d VSS VDD
+ ip transmission_gate
Xsky130_fd_sc_hd__mux4_1_3 ota_1/p1 clock_v2_0/A ota_1/p1_b clock_v2_0/A_b d_clk_grp_1_ctrl_0
+ d_clk_grp_1_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_3/X VSS VDD sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_17 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_28 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_39 ota_1/op ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_5 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_18 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_29 ota_1/on ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_1 transmission_gate_5/in ota_1/p2_b ota_1/p2 VSS VDD transmission_gate_8/in
+ transmission_gate
Xclock_v2_0 clk clock_v2_0/p2d_b clock_v2_0/p2d ota_1/p2_b ota_1/p2 clock_v2_0/p1d_b
+ clock_v2_0/p1d ota_1/p1_b ota_1/p1 clock_v2_0/Ad_b clock_v2_0/Ad clock_v2_0/A_b
+ clock_v2_0/A clock_v2_0/Bd_b clock_v2_0/Bd clock_v2_0/B_b clock_v2_0/B VDD VSS clock_v2
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_6 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_2 transmission_gate_2/out clock_v2_0/p1d_b clock_v2_0/p1d VSS VDD
+ in transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_19 transmission_gate_23/in transmission_gate_19/in
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_7 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_3 ota_w_test_0/in clock_v2_0/A_b clock_v2_0/A VSS VDD transmission_gate_5/in
+ transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_8 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_4 ota_w_test_0/in clock_v2_0/B_b clock_v2_0/B VSS VDD transmission_gate_6/in
+ transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_9 sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_5 ota_w_test_0/ip clock_v2_0/B_b clock_v2_0/B VSS VDD transmission_gate_5/in
+ transmission_gate
Xtransmission_gate_6 ota_w_test_0/ip clock_v2_0/A_b clock_v2_0/A VSS VDD transmission_gate_6/in
+ transmission_gate
Xtransmission_gate_7 transmission_gate_6/in ota_1/p2_b ota_1/p2 VSS VDD transmission_gate_9/in
+ transmission_gate
Xtransmission_gate_8 ota_w_test_0/cm ota_1/p1_b ota_1/p1 VSS VDD transmission_gate_8/in
+ transmission_gate
Xtransmission_gate_9 ota_w_test_0/cm ota_1/p1_b ota_1/p1 VSS VDD transmission_gate_9/in
+ transmission_gate
Xa_mux4_en_0 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1 a_mux4_en_0/in0 a_mux4_en_0/in2 a_mux4_en_0/in3
+ a_probe_3 debug VSS a_mux4_en_0/in1 VDD a_mux4_en
Xa_mux4_en_1 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1 ota_w_test_0/cm a_mux4_en_1/in2 a_mux4_en_1/in3
+ a_probe_2 debug VSS a_mux4_en_1/in1 VDD a_mux4_en
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_40 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_30 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_41 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_42 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_20 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_31 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_32 transmission_gate_9/in transmission_gate_2/out
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_10 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_21 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_43 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_44 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_33 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_11 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_22 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_45 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_34 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_12 transmission_gate_8/in transmission_gate_0/out
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_23 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_TABSMU_0 ota_1/on VSS sky130_fd_pr__cap_mim_m3_1_TABSMU
Xcomparator_v2_0 op onebit_dac_1/v_b ota_1/op VDD VSS ota_1/on ota_1/p1_b comparator_v2
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_46 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_35 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_13 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_24 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_0 in VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_TABSMU_1 ota_1/op VSS sky130_fd_pr__cap_mim_m3_1_TABSMU
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_47 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_36 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_25 sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_1 ip VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_14 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_37 transmission_gate_9/in transmission_gate_2/out
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_15 transmission_gate_6/in a_mux2_en_0/in1 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_26 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__nfet_01v8_CFEPS5_0 VSS onebit_dac_1/v_b VSS sky130_fd_pr__nfet_01v8_CFEPS5
Xesd_cell_2 i_bias_2 VSS VDD esd_cell
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_0 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_38 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_16 transmission_gate_5/in a_mux2_en_0/in0 sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_27 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_3 i_bias_1 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_17 transmission_gate_8/in transmission_gate_0/out
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_28 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_39 sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1031_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n931_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_4 a_probe_1 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_30 transmission_gate_2/out clock_v2_0/p2d_b clock_v2_0/p2d VSS
+ VDD onebit_dac_0/out transmission_gate
.ends

