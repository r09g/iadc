magic
tech sky130A
magscale 1 2
timestamp 1654572275
<< nmos >>
rect -3531 -140 -3411 140
rect -3353 -140 -3233 140
rect -3175 -140 -3055 140
rect -2997 -140 -2877 140
rect -2819 -140 -2699 140
rect -2641 -140 -2521 140
rect -2463 -140 -2343 140
rect -2285 -140 -2165 140
rect -2107 -140 -1987 140
rect -1929 -140 -1809 140
rect -1751 -140 -1631 140
rect -1573 -140 -1453 140
rect -1395 -140 -1275 140
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
rect 1275 -140 1395 140
rect 1453 -140 1573 140
rect 1631 -140 1751 140
rect 1809 -140 1929 140
rect 1987 -140 2107 140
rect 2165 -140 2285 140
rect 2343 -140 2463 140
rect 2521 -140 2641 140
rect 2699 -140 2819 140
rect 2877 -140 2997 140
rect 3055 -140 3175 140
rect 3233 -140 3353 140
rect 3411 -140 3531 140
<< ndiff >>
rect -3589 128 -3531 140
rect -3589 -128 -3577 128
rect -3543 -128 -3531 128
rect -3589 -140 -3531 -128
rect -3411 128 -3353 140
rect -3411 -128 -3399 128
rect -3365 -128 -3353 128
rect -3411 -140 -3353 -128
rect -3233 128 -3175 140
rect -3233 -128 -3221 128
rect -3187 -128 -3175 128
rect -3233 -140 -3175 -128
rect -3055 128 -2997 140
rect -3055 -128 -3043 128
rect -3009 -128 -2997 128
rect -3055 -140 -2997 -128
rect -2877 128 -2819 140
rect -2877 -128 -2865 128
rect -2831 -128 -2819 128
rect -2877 -140 -2819 -128
rect -2699 128 -2641 140
rect -2699 -128 -2687 128
rect -2653 -128 -2641 128
rect -2699 -140 -2641 -128
rect -2521 128 -2463 140
rect -2521 -128 -2509 128
rect -2475 -128 -2463 128
rect -2521 -140 -2463 -128
rect -2343 128 -2285 140
rect -2343 -128 -2331 128
rect -2297 -128 -2285 128
rect -2343 -140 -2285 -128
rect -2165 128 -2107 140
rect -2165 -128 -2153 128
rect -2119 -128 -2107 128
rect -2165 -140 -2107 -128
rect -1987 128 -1929 140
rect -1987 -128 -1975 128
rect -1941 -128 -1929 128
rect -1987 -140 -1929 -128
rect -1809 128 -1751 140
rect -1809 -128 -1797 128
rect -1763 -128 -1751 128
rect -1809 -140 -1751 -128
rect -1631 128 -1573 140
rect -1631 -128 -1619 128
rect -1585 -128 -1573 128
rect -1631 -140 -1573 -128
rect -1453 128 -1395 140
rect -1453 -128 -1441 128
rect -1407 -128 -1395 128
rect -1453 -140 -1395 -128
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
rect 1395 128 1453 140
rect 1395 -128 1407 128
rect 1441 -128 1453 128
rect 1395 -140 1453 -128
rect 1573 128 1631 140
rect 1573 -128 1585 128
rect 1619 -128 1631 128
rect 1573 -140 1631 -128
rect 1751 128 1809 140
rect 1751 -128 1763 128
rect 1797 -128 1809 128
rect 1751 -140 1809 -128
rect 1929 128 1987 140
rect 1929 -128 1941 128
rect 1975 -128 1987 128
rect 1929 -140 1987 -128
rect 2107 128 2165 140
rect 2107 -128 2119 128
rect 2153 -128 2165 128
rect 2107 -140 2165 -128
rect 2285 128 2343 140
rect 2285 -128 2297 128
rect 2331 -128 2343 128
rect 2285 -140 2343 -128
rect 2463 128 2521 140
rect 2463 -128 2475 128
rect 2509 -128 2521 128
rect 2463 -140 2521 -128
rect 2641 128 2699 140
rect 2641 -128 2653 128
rect 2687 -128 2699 128
rect 2641 -140 2699 -128
rect 2819 128 2877 140
rect 2819 -128 2831 128
rect 2865 -128 2877 128
rect 2819 -140 2877 -128
rect 2997 128 3055 140
rect 2997 -128 3009 128
rect 3043 -128 3055 128
rect 2997 -140 3055 -128
rect 3175 128 3233 140
rect 3175 -128 3187 128
rect 3221 -128 3233 128
rect 3175 -140 3233 -128
rect 3353 128 3411 140
rect 3353 -128 3365 128
rect 3399 -128 3411 128
rect 3353 -140 3411 -128
rect 3531 128 3589 140
rect 3531 -128 3543 128
rect 3577 -128 3589 128
rect 3531 -140 3589 -128
<< ndiffc >>
rect -3577 -128 -3543 128
rect -3399 -128 -3365 128
rect -3221 -128 -3187 128
rect -3043 -128 -3009 128
rect -2865 -128 -2831 128
rect -2687 -128 -2653 128
rect -2509 -128 -2475 128
rect -2331 -128 -2297 128
rect -2153 -128 -2119 128
rect -1975 -128 -1941 128
rect -1797 -128 -1763 128
rect -1619 -128 -1585 128
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
rect 1585 -128 1619 128
rect 1763 -128 1797 128
rect 1941 -128 1975 128
rect 2119 -128 2153 128
rect 2297 -128 2331 128
rect 2475 -128 2509 128
rect 2653 -128 2687 128
rect 2831 -128 2865 128
rect 3009 -128 3043 128
rect 3187 -128 3221 128
rect 3365 -128 3399 128
rect 3543 -128 3577 128
<< poly >>
rect -3509 212 -3433 228
rect -3509 194 -3493 212
rect -3531 178 -3493 194
rect -3449 194 -3433 212
rect -3331 212 -3255 228
rect -3331 194 -3315 212
rect -3449 178 -3411 194
rect -3531 140 -3411 178
rect -3353 178 -3315 194
rect -3271 194 -3255 212
rect -3153 212 -3077 228
rect -3153 194 -3137 212
rect -3271 178 -3233 194
rect -3353 140 -3233 178
rect -3175 178 -3137 194
rect -3093 194 -3077 212
rect -2975 212 -2899 228
rect -2975 194 -2959 212
rect -3093 178 -3055 194
rect -3175 140 -3055 178
rect -2997 178 -2959 194
rect -2915 194 -2899 212
rect -2797 212 -2721 228
rect -2797 194 -2781 212
rect -2915 178 -2877 194
rect -2997 140 -2877 178
rect -2819 178 -2781 194
rect -2737 194 -2721 212
rect -2619 212 -2543 228
rect -2619 194 -2603 212
rect -2737 178 -2699 194
rect -2819 140 -2699 178
rect -2641 178 -2603 194
rect -2559 194 -2543 212
rect -2441 212 -2365 228
rect -2441 194 -2425 212
rect -2559 178 -2521 194
rect -2641 140 -2521 178
rect -2463 178 -2425 194
rect -2381 194 -2365 212
rect -2263 212 -2187 228
rect -2263 194 -2247 212
rect -2381 178 -2343 194
rect -2463 140 -2343 178
rect -2285 178 -2247 194
rect -2203 194 -2187 212
rect -2085 212 -2009 228
rect -2085 194 -2069 212
rect -2203 178 -2165 194
rect -2285 140 -2165 178
rect -2107 178 -2069 194
rect -2025 194 -2009 212
rect -1907 212 -1831 228
rect -1907 194 -1891 212
rect -2025 178 -1987 194
rect -2107 140 -1987 178
rect -1929 178 -1891 194
rect -1847 194 -1831 212
rect -1729 212 -1653 228
rect -1729 194 -1713 212
rect -1847 178 -1809 194
rect -1929 140 -1809 178
rect -1751 178 -1713 194
rect -1669 194 -1653 212
rect -1551 212 -1475 228
rect -1551 194 -1535 212
rect -1669 178 -1631 194
rect -1751 140 -1631 178
rect -1573 178 -1535 194
rect -1491 194 -1475 212
rect -1373 212 -1297 228
rect -1373 194 -1357 212
rect -1491 178 -1453 194
rect -1573 140 -1453 178
rect -1395 178 -1357 194
rect -1313 194 -1297 212
rect -1195 212 -1119 228
rect -1195 194 -1179 212
rect -1313 178 -1275 194
rect -1395 140 -1275 178
rect -1217 178 -1179 194
rect -1135 194 -1119 212
rect -1017 212 -941 228
rect -1017 194 -1001 212
rect -1135 178 -1097 194
rect -1217 140 -1097 178
rect -1039 178 -1001 194
rect -957 194 -941 212
rect -839 212 -763 228
rect -839 194 -823 212
rect -957 178 -919 194
rect -1039 140 -919 178
rect -861 178 -823 194
rect -779 194 -763 212
rect -661 212 -585 228
rect -661 194 -645 212
rect -779 178 -741 194
rect -861 140 -741 178
rect -683 178 -645 194
rect -601 194 -585 212
rect -483 212 -407 228
rect -483 194 -467 212
rect -601 178 -563 194
rect -683 140 -563 178
rect -505 178 -467 194
rect -423 194 -407 212
rect -305 212 -229 228
rect -305 194 -289 212
rect -423 178 -385 194
rect -505 140 -385 178
rect -327 178 -289 194
rect -245 194 -229 212
rect -127 212 -51 228
rect -127 194 -111 212
rect -245 178 -207 194
rect -327 140 -207 178
rect -149 178 -111 194
rect -67 194 -51 212
rect 51 212 127 228
rect 51 194 67 212
rect -67 178 -29 194
rect -149 140 -29 178
rect 29 178 67 194
rect 111 194 127 212
rect 229 212 305 228
rect 229 194 245 212
rect 111 178 149 194
rect 29 140 149 178
rect 207 178 245 194
rect 289 194 305 212
rect 407 212 483 228
rect 407 194 423 212
rect 289 178 327 194
rect 207 140 327 178
rect 385 178 423 194
rect 467 194 483 212
rect 585 212 661 228
rect 585 194 601 212
rect 467 178 505 194
rect 385 140 505 178
rect 563 178 601 194
rect 645 194 661 212
rect 763 212 839 228
rect 763 194 779 212
rect 645 178 683 194
rect 563 140 683 178
rect 741 178 779 194
rect 823 194 839 212
rect 941 212 1017 228
rect 941 194 957 212
rect 823 178 861 194
rect 741 140 861 178
rect 919 178 957 194
rect 1001 194 1017 212
rect 1119 212 1195 228
rect 1119 194 1135 212
rect 1001 178 1039 194
rect 919 140 1039 178
rect 1097 178 1135 194
rect 1179 194 1195 212
rect 1297 212 1373 228
rect 1297 194 1313 212
rect 1179 178 1217 194
rect 1097 140 1217 178
rect 1275 178 1313 194
rect 1357 194 1373 212
rect 1475 212 1551 228
rect 1475 194 1491 212
rect 1357 178 1395 194
rect 1275 140 1395 178
rect 1453 178 1491 194
rect 1535 194 1551 212
rect 1653 212 1729 228
rect 1653 194 1669 212
rect 1535 178 1573 194
rect 1453 140 1573 178
rect 1631 178 1669 194
rect 1713 194 1729 212
rect 1831 212 1907 228
rect 1831 194 1847 212
rect 1713 178 1751 194
rect 1631 140 1751 178
rect 1809 178 1847 194
rect 1891 194 1907 212
rect 2009 212 2085 228
rect 2009 194 2025 212
rect 1891 178 1929 194
rect 1809 140 1929 178
rect 1987 178 2025 194
rect 2069 194 2085 212
rect 2187 212 2263 228
rect 2187 194 2203 212
rect 2069 178 2107 194
rect 1987 140 2107 178
rect 2165 178 2203 194
rect 2247 194 2263 212
rect 2365 212 2441 228
rect 2365 194 2381 212
rect 2247 178 2285 194
rect 2165 140 2285 178
rect 2343 178 2381 194
rect 2425 194 2441 212
rect 2543 212 2619 228
rect 2543 194 2559 212
rect 2425 178 2463 194
rect 2343 140 2463 178
rect 2521 178 2559 194
rect 2603 194 2619 212
rect 2721 212 2797 228
rect 2721 194 2737 212
rect 2603 178 2641 194
rect 2521 140 2641 178
rect 2699 178 2737 194
rect 2781 194 2797 212
rect 2899 212 2975 228
rect 2899 194 2915 212
rect 2781 178 2819 194
rect 2699 140 2819 178
rect 2877 178 2915 194
rect 2959 194 2975 212
rect 3077 212 3153 228
rect 3077 194 3093 212
rect 2959 178 2997 194
rect 2877 140 2997 178
rect 3055 178 3093 194
rect 3137 194 3153 212
rect 3255 212 3331 228
rect 3255 194 3271 212
rect 3137 178 3175 194
rect 3055 140 3175 178
rect 3233 178 3271 194
rect 3315 194 3331 212
rect 3433 212 3509 228
rect 3433 194 3449 212
rect 3315 178 3353 194
rect 3233 140 3353 178
rect 3411 178 3449 194
rect 3493 194 3509 212
rect 3493 178 3531 194
rect 3411 140 3531 178
rect -3531 -178 -3411 -140
rect -3531 -194 -3493 -178
rect -3509 -212 -3493 -194
rect -3449 -194 -3411 -178
rect -3353 -178 -3233 -140
rect -3353 -194 -3315 -178
rect -3449 -212 -3433 -194
rect -3509 -228 -3433 -212
rect -3331 -212 -3315 -194
rect -3271 -194 -3233 -178
rect -3175 -178 -3055 -140
rect -3175 -194 -3137 -178
rect -3271 -212 -3255 -194
rect -3331 -228 -3255 -212
rect -3153 -212 -3137 -194
rect -3093 -194 -3055 -178
rect -2997 -178 -2877 -140
rect -2997 -194 -2959 -178
rect -3093 -212 -3077 -194
rect -3153 -228 -3077 -212
rect -2975 -212 -2959 -194
rect -2915 -194 -2877 -178
rect -2819 -178 -2699 -140
rect -2819 -194 -2781 -178
rect -2915 -212 -2899 -194
rect -2975 -228 -2899 -212
rect -2797 -212 -2781 -194
rect -2737 -194 -2699 -178
rect -2641 -178 -2521 -140
rect -2641 -194 -2603 -178
rect -2737 -212 -2721 -194
rect -2797 -228 -2721 -212
rect -2619 -212 -2603 -194
rect -2559 -194 -2521 -178
rect -2463 -178 -2343 -140
rect -2463 -194 -2425 -178
rect -2559 -212 -2543 -194
rect -2619 -228 -2543 -212
rect -2441 -212 -2425 -194
rect -2381 -194 -2343 -178
rect -2285 -178 -2165 -140
rect -2285 -194 -2247 -178
rect -2381 -212 -2365 -194
rect -2441 -228 -2365 -212
rect -2263 -212 -2247 -194
rect -2203 -194 -2165 -178
rect -2107 -178 -1987 -140
rect -2107 -194 -2069 -178
rect -2203 -212 -2187 -194
rect -2263 -228 -2187 -212
rect -2085 -212 -2069 -194
rect -2025 -194 -1987 -178
rect -1929 -178 -1809 -140
rect -1929 -194 -1891 -178
rect -2025 -212 -2009 -194
rect -2085 -228 -2009 -212
rect -1907 -212 -1891 -194
rect -1847 -194 -1809 -178
rect -1751 -178 -1631 -140
rect -1751 -194 -1713 -178
rect -1847 -212 -1831 -194
rect -1907 -228 -1831 -212
rect -1729 -212 -1713 -194
rect -1669 -194 -1631 -178
rect -1573 -178 -1453 -140
rect -1573 -194 -1535 -178
rect -1669 -212 -1653 -194
rect -1729 -228 -1653 -212
rect -1551 -212 -1535 -194
rect -1491 -194 -1453 -178
rect -1395 -178 -1275 -140
rect -1395 -194 -1357 -178
rect -1491 -212 -1475 -194
rect -1551 -228 -1475 -212
rect -1373 -212 -1357 -194
rect -1313 -194 -1275 -178
rect -1217 -178 -1097 -140
rect -1217 -194 -1179 -178
rect -1313 -212 -1297 -194
rect -1373 -228 -1297 -212
rect -1195 -212 -1179 -194
rect -1135 -194 -1097 -178
rect -1039 -178 -919 -140
rect -1039 -194 -1001 -178
rect -1135 -212 -1119 -194
rect -1195 -228 -1119 -212
rect -1017 -212 -1001 -194
rect -957 -194 -919 -178
rect -861 -178 -741 -140
rect -861 -194 -823 -178
rect -957 -212 -941 -194
rect -1017 -228 -941 -212
rect -839 -212 -823 -194
rect -779 -194 -741 -178
rect -683 -178 -563 -140
rect -683 -194 -645 -178
rect -779 -212 -763 -194
rect -839 -228 -763 -212
rect -661 -212 -645 -194
rect -601 -194 -563 -178
rect -505 -178 -385 -140
rect -505 -194 -467 -178
rect -601 -212 -585 -194
rect -661 -228 -585 -212
rect -483 -212 -467 -194
rect -423 -194 -385 -178
rect -327 -178 -207 -140
rect -327 -194 -289 -178
rect -423 -212 -407 -194
rect -483 -228 -407 -212
rect -305 -212 -289 -194
rect -245 -194 -207 -178
rect -149 -178 -29 -140
rect -149 -194 -111 -178
rect -245 -212 -229 -194
rect -305 -228 -229 -212
rect -127 -212 -111 -194
rect -67 -194 -29 -178
rect 29 -178 149 -140
rect 29 -194 67 -178
rect -67 -212 -51 -194
rect -127 -228 -51 -212
rect 51 -212 67 -194
rect 111 -194 149 -178
rect 207 -178 327 -140
rect 207 -194 245 -178
rect 111 -212 127 -194
rect 51 -228 127 -212
rect 229 -212 245 -194
rect 289 -194 327 -178
rect 385 -178 505 -140
rect 385 -194 423 -178
rect 289 -212 305 -194
rect 229 -228 305 -212
rect 407 -212 423 -194
rect 467 -194 505 -178
rect 563 -178 683 -140
rect 563 -194 601 -178
rect 467 -212 483 -194
rect 407 -228 483 -212
rect 585 -212 601 -194
rect 645 -194 683 -178
rect 741 -178 861 -140
rect 741 -194 779 -178
rect 645 -212 661 -194
rect 585 -228 661 -212
rect 763 -212 779 -194
rect 823 -194 861 -178
rect 919 -178 1039 -140
rect 919 -194 957 -178
rect 823 -212 839 -194
rect 763 -228 839 -212
rect 941 -212 957 -194
rect 1001 -194 1039 -178
rect 1097 -178 1217 -140
rect 1097 -194 1135 -178
rect 1001 -212 1017 -194
rect 941 -228 1017 -212
rect 1119 -212 1135 -194
rect 1179 -194 1217 -178
rect 1275 -178 1395 -140
rect 1275 -194 1313 -178
rect 1179 -212 1195 -194
rect 1119 -228 1195 -212
rect 1297 -212 1313 -194
rect 1357 -194 1395 -178
rect 1453 -178 1573 -140
rect 1453 -194 1491 -178
rect 1357 -212 1373 -194
rect 1297 -228 1373 -212
rect 1475 -212 1491 -194
rect 1535 -194 1573 -178
rect 1631 -178 1751 -140
rect 1631 -194 1669 -178
rect 1535 -212 1551 -194
rect 1475 -228 1551 -212
rect 1653 -212 1669 -194
rect 1713 -194 1751 -178
rect 1809 -178 1929 -140
rect 1809 -194 1847 -178
rect 1713 -212 1729 -194
rect 1653 -228 1729 -212
rect 1831 -212 1847 -194
rect 1891 -194 1929 -178
rect 1987 -178 2107 -140
rect 1987 -194 2025 -178
rect 1891 -212 1907 -194
rect 1831 -228 1907 -212
rect 2009 -212 2025 -194
rect 2069 -194 2107 -178
rect 2165 -178 2285 -140
rect 2165 -194 2203 -178
rect 2069 -212 2085 -194
rect 2009 -228 2085 -212
rect 2187 -212 2203 -194
rect 2247 -194 2285 -178
rect 2343 -178 2463 -140
rect 2343 -194 2381 -178
rect 2247 -212 2263 -194
rect 2187 -228 2263 -212
rect 2365 -212 2381 -194
rect 2425 -194 2463 -178
rect 2521 -178 2641 -140
rect 2521 -194 2559 -178
rect 2425 -212 2441 -194
rect 2365 -228 2441 -212
rect 2543 -212 2559 -194
rect 2603 -194 2641 -178
rect 2699 -178 2819 -140
rect 2699 -194 2737 -178
rect 2603 -212 2619 -194
rect 2543 -228 2619 -212
rect 2721 -212 2737 -194
rect 2781 -194 2819 -178
rect 2877 -178 2997 -140
rect 2877 -194 2915 -178
rect 2781 -212 2797 -194
rect 2721 -228 2797 -212
rect 2899 -212 2915 -194
rect 2959 -194 2997 -178
rect 3055 -178 3175 -140
rect 3055 -194 3093 -178
rect 2959 -212 2975 -194
rect 2899 -228 2975 -212
rect 3077 -212 3093 -194
rect 3137 -194 3175 -178
rect 3233 -178 3353 -140
rect 3233 -194 3271 -178
rect 3137 -212 3153 -194
rect 3077 -228 3153 -212
rect 3255 -212 3271 -194
rect 3315 -194 3353 -178
rect 3411 -178 3531 -140
rect 3411 -194 3449 -178
rect 3315 -212 3331 -194
rect 3255 -228 3331 -212
rect 3433 -212 3449 -194
rect 3493 -194 3531 -178
rect 3493 -212 3509 -194
rect 3433 -228 3509 -212
<< polycont >>
rect -3493 178 -3449 212
rect -3315 178 -3271 212
rect -3137 178 -3093 212
rect -2959 178 -2915 212
rect -2781 178 -2737 212
rect -2603 178 -2559 212
rect -2425 178 -2381 212
rect -2247 178 -2203 212
rect -2069 178 -2025 212
rect -1891 178 -1847 212
rect -1713 178 -1669 212
rect -1535 178 -1491 212
rect -1357 178 -1313 212
rect -1179 178 -1135 212
rect -1001 178 -957 212
rect -823 178 -779 212
rect -645 178 -601 212
rect -467 178 -423 212
rect -289 178 -245 212
rect -111 178 -67 212
rect 67 178 111 212
rect 245 178 289 212
rect 423 178 467 212
rect 601 178 645 212
rect 779 178 823 212
rect 957 178 1001 212
rect 1135 178 1179 212
rect 1313 178 1357 212
rect 1491 178 1535 212
rect 1669 178 1713 212
rect 1847 178 1891 212
rect 2025 178 2069 212
rect 2203 178 2247 212
rect 2381 178 2425 212
rect 2559 178 2603 212
rect 2737 178 2781 212
rect 2915 178 2959 212
rect 3093 178 3137 212
rect 3271 178 3315 212
rect 3449 178 3493 212
rect -3493 -212 -3449 -178
rect -3315 -212 -3271 -178
rect -3137 -212 -3093 -178
rect -2959 -212 -2915 -178
rect -2781 -212 -2737 -178
rect -2603 -212 -2559 -178
rect -2425 -212 -2381 -178
rect -2247 -212 -2203 -178
rect -2069 -212 -2025 -178
rect -1891 -212 -1847 -178
rect -1713 -212 -1669 -178
rect -1535 -212 -1491 -178
rect -1357 -212 -1313 -178
rect -1179 -212 -1135 -178
rect -1001 -212 -957 -178
rect -823 -212 -779 -178
rect -645 -212 -601 -178
rect -467 -212 -423 -178
rect -289 -212 -245 -178
rect -111 -212 -67 -178
rect 67 -212 111 -178
rect 245 -212 289 -178
rect 423 -212 467 -178
rect 601 -212 645 -178
rect 779 -212 823 -178
rect 957 -212 1001 -178
rect 1135 -212 1179 -178
rect 1313 -212 1357 -178
rect 1491 -212 1535 -178
rect 1669 -212 1713 -178
rect 1847 -212 1891 -178
rect 2025 -212 2069 -178
rect 2203 -212 2247 -178
rect 2381 -212 2425 -178
rect 2559 -212 2603 -178
rect 2737 -212 2781 -178
rect 2915 -212 2959 -178
rect 3093 -212 3137 -178
rect 3271 -212 3315 -178
rect 3449 -212 3493 -178
<< locali >>
rect -3509 178 -3493 212
rect -3449 178 -3433 212
rect -3331 178 -3315 212
rect -3271 178 -3255 212
rect -3153 178 -3137 212
rect -3093 178 -3077 212
rect -2975 178 -2959 212
rect -2915 178 -2899 212
rect -2797 178 -2781 212
rect -2737 178 -2721 212
rect -2619 178 -2603 212
rect -2559 178 -2543 212
rect -2441 178 -2425 212
rect -2381 178 -2365 212
rect -2263 178 -2247 212
rect -2203 178 -2187 212
rect -2085 178 -2069 212
rect -2025 178 -2009 212
rect -1907 178 -1891 212
rect -1847 178 -1831 212
rect -1729 178 -1713 212
rect -1669 178 -1653 212
rect -1551 178 -1535 212
rect -1491 178 -1475 212
rect -1373 178 -1357 212
rect -1313 178 -1297 212
rect -1195 178 -1179 212
rect -1135 178 -1119 212
rect -1017 178 -1001 212
rect -957 178 -941 212
rect -839 178 -823 212
rect -779 178 -763 212
rect -661 178 -645 212
rect -601 178 -585 212
rect -483 178 -467 212
rect -423 178 -407 212
rect -305 178 -289 212
rect -245 178 -229 212
rect -127 178 -111 212
rect -67 178 -51 212
rect 51 178 67 212
rect 111 178 127 212
rect 229 178 245 212
rect 289 178 305 212
rect 407 178 423 212
rect 467 178 483 212
rect 585 178 601 212
rect 645 178 661 212
rect 763 178 779 212
rect 823 178 839 212
rect 941 178 957 212
rect 1001 178 1017 212
rect 1119 178 1135 212
rect 1179 178 1195 212
rect 1297 178 1313 212
rect 1357 178 1373 212
rect 1475 178 1491 212
rect 1535 178 1551 212
rect 1653 178 1669 212
rect 1713 178 1729 212
rect 1831 178 1847 212
rect 1891 178 1907 212
rect 2009 178 2025 212
rect 2069 178 2085 212
rect 2187 178 2203 212
rect 2247 178 2263 212
rect 2365 178 2381 212
rect 2425 178 2441 212
rect 2543 178 2559 212
rect 2603 178 2619 212
rect 2721 178 2737 212
rect 2781 178 2797 212
rect 2899 178 2915 212
rect 2959 178 2975 212
rect 3077 178 3093 212
rect 3137 178 3153 212
rect 3255 178 3271 212
rect 3315 178 3331 212
rect 3433 178 3449 212
rect 3493 178 3509 212
rect -3577 128 -3543 144
rect -3577 -144 -3543 -128
rect -3399 128 -3365 144
rect -3399 -144 -3365 -128
rect -3221 128 -3187 144
rect -3221 -144 -3187 -128
rect -3043 128 -3009 144
rect -3043 -144 -3009 -128
rect -2865 128 -2831 144
rect -2865 -144 -2831 -128
rect -2687 128 -2653 144
rect -2687 -144 -2653 -128
rect -2509 128 -2475 144
rect -2509 -144 -2475 -128
rect -2331 128 -2297 144
rect -2331 -144 -2297 -128
rect -2153 128 -2119 144
rect -2153 -144 -2119 -128
rect -1975 128 -1941 144
rect -1975 -144 -1941 -128
rect -1797 128 -1763 144
rect -1797 -144 -1763 -128
rect -1619 128 -1585 144
rect -1619 -144 -1585 -128
rect -1441 128 -1407 144
rect -1441 -144 -1407 -128
rect -1263 128 -1229 144
rect -1263 -144 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 144
rect 1229 -144 1263 -128
rect 1407 128 1441 144
rect 1407 -144 1441 -128
rect 1585 128 1619 144
rect 1585 -144 1619 -128
rect 1763 128 1797 144
rect 1763 -144 1797 -128
rect 1941 128 1975 144
rect 1941 -144 1975 -128
rect 2119 128 2153 144
rect 2119 -144 2153 -128
rect 2297 128 2331 144
rect 2297 -144 2331 -128
rect 2475 128 2509 144
rect 2475 -144 2509 -128
rect 2653 128 2687 144
rect 2653 -144 2687 -128
rect 2831 128 2865 144
rect 2831 -144 2865 -128
rect 3009 128 3043 144
rect 3009 -144 3043 -128
rect 3187 128 3221 144
rect 3187 -144 3221 -128
rect 3365 128 3399 144
rect 3365 -144 3399 -128
rect 3543 128 3577 144
rect 3543 -144 3577 -128
rect -3509 -212 -3493 -178
rect -3449 -212 -3433 -178
rect -3331 -212 -3315 -178
rect -3271 -212 -3255 -178
rect -3153 -212 -3137 -178
rect -3093 -212 -3077 -178
rect -2975 -212 -2959 -178
rect -2915 -212 -2899 -178
rect -2797 -212 -2781 -178
rect -2737 -212 -2721 -178
rect -2619 -212 -2603 -178
rect -2559 -212 -2543 -178
rect -2441 -212 -2425 -178
rect -2381 -212 -2365 -178
rect -2263 -212 -2247 -178
rect -2203 -212 -2187 -178
rect -2085 -212 -2069 -178
rect -2025 -212 -2009 -178
rect -1907 -212 -1891 -178
rect -1847 -212 -1831 -178
rect -1729 -212 -1713 -178
rect -1669 -212 -1653 -178
rect -1551 -212 -1535 -178
rect -1491 -212 -1475 -178
rect -1373 -212 -1357 -178
rect -1313 -212 -1297 -178
rect -1195 -212 -1179 -178
rect -1135 -212 -1119 -178
rect -1017 -212 -1001 -178
rect -957 -212 -941 -178
rect -839 -212 -823 -178
rect -779 -212 -763 -178
rect -661 -212 -645 -178
rect -601 -212 -585 -178
rect -483 -212 -467 -178
rect -423 -212 -407 -178
rect -305 -212 -289 -178
rect -245 -212 -229 -178
rect -127 -212 -111 -178
rect -67 -212 -51 -178
rect 51 -212 67 -178
rect 111 -212 127 -178
rect 229 -212 245 -178
rect 289 -212 305 -178
rect 407 -212 423 -178
rect 467 -212 483 -178
rect 585 -212 601 -178
rect 645 -212 661 -178
rect 763 -212 779 -178
rect 823 -212 839 -178
rect 941 -212 957 -178
rect 1001 -212 1017 -178
rect 1119 -212 1135 -178
rect 1179 -212 1195 -178
rect 1297 -212 1313 -178
rect 1357 -212 1373 -178
rect 1475 -212 1491 -178
rect 1535 -212 1551 -178
rect 1653 -212 1669 -178
rect 1713 -212 1729 -178
rect 1831 -212 1847 -178
rect 1891 -212 1907 -178
rect 2009 -212 2025 -178
rect 2069 -212 2085 -178
rect 2187 -212 2203 -178
rect 2247 -212 2263 -178
rect 2365 -212 2381 -178
rect 2425 -212 2441 -178
rect 2543 -212 2559 -178
rect 2603 -212 2619 -178
rect 2721 -212 2737 -178
rect 2781 -212 2797 -178
rect 2899 -212 2915 -178
rect 2959 -212 2975 -178
rect 3077 -212 3093 -178
rect 3137 -212 3153 -178
rect 3255 -212 3271 -178
rect 3315 -212 3331 -178
rect 3433 -212 3449 -178
rect 3493 -212 3509 -178
<< viali >>
rect -3493 178 -3449 212
rect -3315 178 -3271 212
rect -3137 178 -3093 212
rect -2959 178 -2915 212
rect -2781 178 -2737 212
rect -2603 178 -2559 212
rect -2425 178 -2381 212
rect -2247 178 -2203 212
rect -2069 178 -2025 212
rect -1891 178 -1847 212
rect -1713 178 -1669 212
rect -1535 178 -1491 212
rect -1357 178 -1313 212
rect -1179 178 -1135 212
rect -1001 178 -957 212
rect -823 178 -779 212
rect -645 178 -601 212
rect -467 178 -423 212
rect -289 178 -245 212
rect -111 178 -67 212
rect 67 178 111 212
rect 245 178 289 212
rect 423 178 467 212
rect 601 178 645 212
rect 779 178 823 212
rect 957 178 1001 212
rect 1135 178 1179 212
rect 1313 178 1357 212
rect 1491 178 1535 212
rect 1669 178 1713 212
rect 1847 178 1891 212
rect 2025 178 2069 212
rect 2203 178 2247 212
rect 2381 178 2425 212
rect 2559 178 2603 212
rect 2737 178 2781 212
rect 2915 178 2959 212
rect 3093 178 3137 212
rect 3271 178 3315 212
rect 3449 178 3493 212
rect -3577 -128 -3543 128
rect -3399 -128 -3365 128
rect -3221 -128 -3187 128
rect -3043 -128 -3009 128
rect -2865 -128 -2831 128
rect -2687 -128 -2653 128
rect -2509 -128 -2475 128
rect -2331 -128 -2297 128
rect -2153 -128 -2119 128
rect -1975 -128 -1941 128
rect -1797 -128 -1763 128
rect -1619 -128 -1585 128
rect -1441 -128 -1407 128
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
rect 1407 -128 1441 128
rect 1585 -128 1619 128
rect 1763 -128 1797 128
rect 1941 -128 1975 128
rect 2119 -128 2153 128
rect 2297 -128 2331 128
rect 2475 -128 2509 128
rect 2653 -128 2687 128
rect 2831 -128 2865 128
rect 3009 -128 3043 128
rect 3187 -128 3221 128
rect 3365 -128 3399 128
rect 3543 -128 3577 128
rect -3493 -212 -3449 -178
rect -3315 -212 -3271 -178
rect -3137 -212 -3093 -178
rect -2959 -212 -2915 -178
rect -2781 -212 -2737 -178
rect -2603 -212 -2559 -178
rect -2425 -212 -2381 -178
rect -2247 -212 -2203 -178
rect -2069 -212 -2025 -178
rect -1891 -212 -1847 -178
rect -1713 -212 -1669 -178
rect -1535 -212 -1491 -178
rect -1357 -212 -1313 -178
rect -1179 -212 -1135 -178
rect -1001 -212 -957 -178
rect -823 -212 -779 -178
rect -645 -212 -601 -178
rect -467 -212 -423 -178
rect -289 -212 -245 -178
rect -111 -212 -67 -178
rect 67 -212 111 -178
rect 245 -212 289 -178
rect 423 -212 467 -178
rect 601 -212 645 -178
rect 779 -212 823 -178
rect 957 -212 1001 -178
rect 1135 -212 1179 -178
rect 1313 -212 1357 -178
rect 1491 -212 1535 -178
rect 1669 -212 1713 -178
rect 1847 -212 1891 -178
rect 2025 -212 2069 -178
rect 2203 -212 2247 -178
rect 2381 -212 2425 -178
rect 2559 -212 2603 -178
rect 2737 -212 2781 -178
rect 2915 -212 2959 -178
rect 3093 -212 3137 -178
rect 3271 -212 3315 -178
rect 3449 -212 3493 -178
<< metal1 >>
rect -3509 212 -3433 228
rect -3509 178 -3493 212
rect -3449 178 -3433 212
rect -3509 172 -3433 178
rect -3331 212 -3255 228
rect -3331 178 -3315 212
rect -3271 178 -3255 212
rect -3331 172 -3255 178
rect -3153 212 -3077 228
rect -3153 178 -3137 212
rect -3093 178 -3077 212
rect -3153 172 -3077 178
rect -2975 212 -2899 228
rect -2975 178 -2959 212
rect -2915 178 -2899 212
rect -2975 172 -2899 178
rect -2797 212 -2721 228
rect -2797 178 -2781 212
rect -2737 178 -2721 212
rect -2797 172 -2721 178
rect -2619 212 -2543 228
rect -2619 178 -2603 212
rect -2559 178 -2543 212
rect -2619 172 -2543 178
rect -2441 212 -2365 228
rect -2441 178 -2425 212
rect -2381 178 -2365 212
rect -2441 172 -2365 178
rect -2263 212 -2187 228
rect -2263 178 -2247 212
rect -2203 178 -2187 212
rect -2263 172 -2187 178
rect -2085 212 -2009 228
rect -2085 178 -2069 212
rect -2025 178 -2009 212
rect -2085 172 -2009 178
rect -1907 212 -1831 228
rect -1907 178 -1891 212
rect -1847 178 -1831 212
rect -1907 172 -1831 178
rect -1729 212 -1653 228
rect -1729 178 -1713 212
rect -1669 178 -1653 212
rect -1729 172 -1653 178
rect -1551 212 -1475 228
rect -1551 178 -1535 212
rect -1491 178 -1475 212
rect -1551 172 -1475 178
rect -1373 212 -1297 228
rect -1373 178 -1357 212
rect -1313 178 -1297 212
rect -1373 172 -1297 178
rect -1195 212 -1119 228
rect -1195 178 -1179 212
rect -1135 178 -1119 212
rect -1195 172 -1119 178
rect -1017 212 -941 228
rect -1017 178 -1001 212
rect -957 178 -941 212
rect -1017 172 -941 178
rect -839 212 -763 228
rect -839 178 -823 212
rect -779 178 -763 212
rect -839 172 -763 178
rect -661 212 -585 228
rect -661 178 -645 212
rect -601 178 -585 212
rect -661 172 -585 178
rect -483 212 -407 228
rect -483 178 -467 212
rect -423 178 -407 212
rect -483 172 -407 178
rect -305 212 -229 228
rect -305 178 -289 212
rect -245 178 -229 212
rect -305 172 -229 178
rect -127 212 -51 228
rect -127 178 -111 212
rect -67 178 -51 212
rect -127 172 -51 178
rect 51 212 127 228
rect 51 178 67 212
rect 111 178 127 212
rect 51 172 127 178
rect 229 212 305 228
rect 229 178 245 212
rect 289 178 305 212
rect 229 172 305 178
rect 407 212 483 228
rect 407 178 423 212
rect 467 178 483 212
rect 407 172 483 178
rect 585 212 661 228
rect 585 178 601 212
rect 645 178 661 212
rect 585 172 661 178
rect 763 212 839 228
rect 763 178 779 212
rect 823 178 839 212
rect 763 172 839 178
rect 941 212 1017 228
rect 941 178 957 212
rect 1001 178 1017 212
rect 941 172 1017 178
rect 1119 212 1195 228
rect 1119 178 1135 212
rect 1179 178 1195 212
rect 1119 172 1195 178
rect 1297 212 1373 228
rect 1297 178 1313 212
rect 1357 178 1373 212
rect 1297 172 1373 178
rect 1475 212 1551 228
rect 1475 178 1491 212
rect 1535 178 1551 212
rect 1475 172 1551 178
rect 1653 212 1729 228
rect 1653 178 1669 212
rect 1713 178 1729 212
rect 1653 172 1729 178
rect 1831 212 1907 228
rect 1831 178 1847 212
rect 1891 178 1907 212
rect 1831 172 1907 178
rect 2009 212 2085 228
rect 2009 178 2025 212
rect 2069 178 2085 212
rect 2009 172 2085 178
rect 2187 212 2263 228
rect 2187 178 2203 212
rect 2247 178 2263 212
rect 2187 172 2263 178
rect 2365 212 2441 228
rect 2365 178 2381 212
rect 2425 178 2441 212
rect 2365 172 2441 178
rect 2543 212 2619 228
rect 2543 178 2559 212
rect 2603 178 2619 212
rect 2543 172 2619 178
rect 2721 212 2797 228
rect 2721 178 2737 212
rect 2781 178 2797 212
rect 2721 172 2797 178
rect 2899 212 2975 228
rect 2899 178 2915 212
rect 2959 178 2975 212
rect 2899 172 2975 178
rect 3077 212 3153 228
rect 3077 178 3093 212
rect 3137 178 3153 212
rect 3077 172 3153 178
rect 3255 212 3331 228
rect 3255 178 3271 212
rect 3315 178 3331 212
rect 3255 172 3331 178
rect 3433 212 3509 228
rect 3433 178 3449 212
rect 3493 178 3509 212
rect 3433 172 3509 178
rect -3583 128 -3537 140
rect -3583 -128 -3577 128
rect -3543 -128 -3537 128
rect -3583 -140 -3537 -128
rect -3405 128 -3359 140
rect -3405 -128 -3399 128
rect -3365 -128 -3359 128
rect -3405 -140 -3359 -128
rect -3227 128 -3181 140
rect -3227 -128 -3221 128
rect -3187 -128 -3181 128
rect -3227 -140 -3181 -128
rect -3049 128 -3003 140
rect -3049 -128 -3043 128
rect -3009 -128 -3003 128
rect -3049 -140 -3003 -128
rect -2871 128 -2825 140
rect -2871 -128 -2865 128
rect -2831 -128 -2825 128
rect -2871 -140 -2825 -128
rect -2693 128 -2647 140
rect -2693 -128 -2687 128
rect -2653 -128 -2647 128
rect -2693 -140 -2647 -128
rect -2515 128 -2469 140
rect -2515 -128 -2509 128
rect -2475 -128 -2469 128
rect -2515 -140 -2469 -128
rect -2337 128 -2291 140
rect -2337 -128 -2331 128
rect -2297 -128 -2291 128
rect -2337 -140 -2291 -128
rect -2159 128 -2113 140
rect -2159 -128 -2153 128
rect -2119 -128 -2113 128
rect -2159 -140 -2113 -128
rect -1981 128 -1935 140
rect -1981 -128 -1975 128
rect -1941 -128 -1935 128
rect -1981 -140 -1935 -128
rect -1803 128 -1757 140
rect -1803 -128 -1797 128
rect -1763 -128 -1757 128
rect -1803 -140 -1757 -128
rect -1625 128 -1579 140
rect -1625 -128 -1619 128
rect -1585 -128 -1579 128
rect -1625 -140 -1579 -128
rect -1447 128 -1401 140
rect -1447 -128 -1441 128
rect -1407 -128 -1401 128
rect -1447 -140 -1401 -128
rect -1269 128 -1223 140
rect -1269 -128 -1263 128
rect -1229 -128 -1223 128
rect -1269 -140 -1223 -128
rect -1091 128 -1045 140
rect -1091 -128 -1085 128
rect -1051 -128 -1045 128
rect -1091 -140 -1045 -128
rect -913 128 -867 140
rect -913 -128 -907 128
rect -873 -128 -867 128
rect -913 -140 -867 -128
rect -735 128 -689 140
rect -735 -128 -729 128
rect -695 -128 -689 128
rect -735 -140 -689 -128
rect -557 128 -511 140
rect -557 -128 -551 128
rect -517 -128 -511 128
rect -557 -140 -511 -128
rect -379 128 -333 140
rect -379 -128 -373 128
rect -339 -128 -333 128
rect -379 -140 -333 -128
rect -201 128 -155 140
rect -201 -128 -195 128
rect -161 -128 -155 128
rect -201 -140 -155 -128
rect -23 128 23 140
rect -23 -128 -17 128
rect 17 -128 23 128
rect -23 -140 23 -128
rect 155 128 201 140
rect 155 -128 161 128
rect 195 -128 201 128
rect 155 -140 201 -128
rect 333 128 379 140
rect 333 -128 339 128
rect 373 -128 379 128
rect 333 -140 379 -128
rect 511 128 557 140
rect 511 -128 517 128
rect 551 -128 557 128
rect 511 -140 557 -128
rect 689 128 735 140
rect 689 -128 695 128
rect 729 -128 735 128
rect 689 -140 735 -128
rect 867 128 913 140
rect 867 -128 873 128
rect 907 -128 913 128
rect 867 -140 913 -128
rect 1045 128 1091 140
rect 1045 -128 1051 128
rect 1085 -128 1091 128
rect 1045 -140 1091 -128
rect 1223 128 1269 140
rect 1223 -128 1229 128
rect 1263 -128 1269 128
rect 1223 -140 1269 -128
rect 1401 128 1447 140
rect 1401 -128 1407 128
rect 1441 -128 1447 128
rect 1401 -140 1447 -128
rect 1579 128 1625 140
rect 1579 -128 1585 128
rect 1619 -128 1625 128
rect 1579 -140 1625 -128
rect 1757 128 1803 140
rect 1757 -128 1763 128
rect 1797 -128 1803 128
rect 1757 -140 1803 -128
rect 1935 128 1981 140
rect 1935 -128 1941 128
rect 1975 -128 1981 128
rect 1935 -140 1981 -128
rect 2113 128 2159 140
rect 2113 -128 2119 128
rect 2153 -128 2159 128
rect 2113 -140 2159 -128
rect 2291 128 2337 140
rect 2291 -128 2297 128
rect 2331 -128 2337 128
rect 2291 -140 2337 -128
rect 2469 128 2515 140
rect 2469 -128 2475 128
rect 2509 -128 2515 128
rect 2469 -140 2515 -128
rect 2647 128 2693 140
rect 2647 -128 2653 128
rect 2687 -128 2693 128
rect 2647 -140 2693 -128
rect 2825 128 2871 140
rect 2825 -128 2831 128
rect 2865 -128 2871 128
rect 2825 -140 2871 -128
rect 3003 128 3049 140
rect 3003 -128 3009 128
rect 3043 -128 3049 128
rect 3003 -140 3049 -128
rect 3181 128 3227 140
rect 3181 -128 3187 128
rect 3221 -128 3227 128
rect 3181 -140 3227 -128
rect 3359 128 3405 140
rect 3359 -128 3365 128
rect 3399 -128 3405 128
rect 3359 -140 3405 -128
rect 3537 128 3583 140
rect 3537 -128 3543 128
rect 3577 -128 3583 128
rect 3537 -140 3583 -128
rect -3509 -178 -3433 -172
rect -3509 -212 -3493 -178
rect -3449 -212 -3433 -178
rect -3509 -228 -3433 -212
rect -3331 -178 -3255 -172
rect -3331 -212 -3315 -178
rect -3271 -212 -3255 -178
rect -3331 -228 -3255 -212
rect -3153 -178 -3077 -172
rect -3153 -212 -3137 -178
rect -3093 -212 -3077 -178
rect -3153 -228 -3077 -212
rect -2975 -178 -2899 -172
rect -2975 -212 -2959 -178
rect -2915 -212 -2899 -178
rect -2975 -228 -2899 -212
rect -2797 -178 -2721 -172
rect -2797 -212 -2781 -178
rect -2737 -212 -2721 -178
rect -2797 -228 -2721 -212
rect -2619 -178 -2543 -172
rect -2619 -212 -2603 -178
rect -2559 -212 -2543 -178
rect -2619 -228 -2543 -212
rect -2441 -178 -2365 -172
rect -2441 -212 -2425 -178
rect -2381 -212 -2365 -178
rect -2441 -228 -2365 -212
rect -2263 -178 -2187 -172
rect -2263 -212 -2247 -178
rect -2203 -212 -2187 -178
rect -2263 -228 -2187 -212
rect -2085 -178 -2009 -172
rect -2085 -212 -2069 -178
rect -2025 -212 -2009 -178
rect -2085 -228 -2009 -212
rect -1907 -178 -1831 -172
rect -1907 -212 -1891 -178
rect -1847 -212 -1831 -178
rect -1907 -228 -1831 -212
rect -1729 -178 -1653 -172
rect -1729 -212 -1713 -178
rect -1669 -212 -1653 -178
rect -1729 -228 -1653 -212
rect -1551 -178 -1475 -172
rect -1551 -212 -1535 -178
rect -1491 -212 -1475 -178
rect -1551 -228 -1475 -212
rect -1373 -178 -1297 -172
rect -1373 -212 -1357 -178
rect -1313 -212 -1297 -178
rect -1373 -228 -1297 -212
rect -1195 -178 -1119 -172
rect -1195 -212 -1179 -178
rect -1135 -212 -1119 -178
rect -1195 -228 -1119 -212
rect -1017 -178 -941 -172
rect -1017 -212 -1001 -178
rect -957 -212 -941 -178
rect -1017 -228 -941 -212
rect -839 -178 -763 -172
rect -839 -212 -823 -178
rect -779 -212 -763 -178
rect -839 -228 -763 -212
rect -661 -178 -585 -172
rect -661 -212 -645 -178
rect -601 -212 -585 -178
rect -661 -228 -585 -212
rect -483 -178 -407 -172
rect -483 -212 -467 -178
rect -423 -212 -407 -178
rect -483 -228 -407 -212
rect -305 -178 -229 -172
rect -305 -212 -289 -178
rect -245 -212 -229 -178
rect -305 -228 -229 -212
rect -127 -178 -51 -172
rect -127 -212 -111 -178
rect -67 -212 -51 -178
rect -127 -228 -51 -212
rect 51 -178 127 -172
rect 51 -212 67 -178
rect 111 -212 127 -178
rect 51 -228 127 -212
rect 229 -178 305 -172
rect 229 -212 245 -178
rect 289 -212 305 -178
rect 229 -228 305 -212
rect 407 -178 483 -172
rect 407 -212 423 -178
rect 467 -212 483 -178
rect 407 -228 483 -212
rect 585 -178 661 -172
rect 585 -212 601 -178
rect 645 -212 661 -178
rect 585 -228 661 -212
rect 763 -178 839 -172
rect 763 -212 779 -178
rect 823 -212 839 -178
rect 763 -228 839 -212
rect 941 -178 1017 -172
rect 941 -212 957 -178
rect 1001 -212 1017 -178
rect 941 -228 1017 -212
rect 1119 -178 1195 -172
rect 1119 -212 1135 -178
rect 1179 -212 1195 -178
rect 1119 -228 1195 -212
rect 1297 -178 1373 -172
rect 1297 -212 1313 -178
rect 1357 -212 1373 -178
rect 1297 -228 1373 -212
rect 1475 -178 1551 -172
rect 1475 -212 1491 -178
rect 1535 -212 1551 -178
rect 1475 -228 1551 -212
rect 1653 -178 1729 -172
rect 1653 -212 1669 -178
rect 1713 -212 1729 -178
rect 1653 -228 1729 -212
rect 1831 -178 1907 -172
rect 1831 -212 1847 -178
rect 1891 -212 1907 -178
rect 1831 -228 1907 -212
rect 2009 -178 2085 -172
rect 2009 -212 2025 -178
rect 2069 -212 2085 -178
rect 2009 -228 2085 -212
rect 2187 -178 2263 -172
rect 2187 -212 2203 -178
rect 2247 -212 2263 -178
rect 2187 -228 2263 -212
rect 2365 -178 2441 -172
rect 2365 -212 2381 -178
rect 2425 -212 2441 -178
rect 2365 -228 2441 -212
rect 2543 -178 2619 -172
rect 2543 -212 2559 -178
rect 2603 -212 2619 -178
rect 2543 -228 2619 -212
rect 2721 -178 2797 -172
rect 2721 -212 2737 -178
rect 2781 -212 2797 -178
rect 2721 -228 2797 -212
rect 2899 -178 2975 -172
rect 2899 -212 2915 -178
rect 2959 -212 2975 -178
rect 2899 -228 2975 -212
rect 3077 -178 3153 -172
rect 3077 -212 3093 -178
rect 3137 -212 3153 -178
rect 3077 -228 3153 -212
rect 3255 -178 3331 -172
rect 3255 -212 3271 -178
rect 3315 -212 3331 -178
rect 3255 -228 3331 -212
rect 3433 -178 3509 -172
rect 3433 -212 3449 -178
rect 3493 -212 3509 -178
rect 3433 -228 3509 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 40 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
