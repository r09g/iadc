* NGSPICE file created from analog_top.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_BRTJC6 a_n345_n500# a_1135_n588# a_n603_n588#
+ a_n1393_n588# a_n1609_n500# a_661_n588# a_n1135_n500# a_n977_n500# a_1293_n588#
+ a_n761_n588# a_n503_n500# a_n1551_n588# a_129_n500# a_n1293_n500# a_287_n500# a_n661_n500#
+ a_1451_n588# a_n1451_n500# a_919_n500# a_445_n500# a_1077_n500# a_29_n588# a_n129_n588#
+ a_603_n500# a_187_n588# a_1235_n500# a_n287_n588# a_761_n500# a_819_n588# a_345_n588#
+ a_n1077_n588# a_n29_n500# a_1393_n500# a_n919_n588# a_n1743_n722# a_n187_n500# a_977_n588#
+ a_n445_n588# a_503_n588# a_n1235_n588# a_1551_n500# a_n819_n500#
X0 a_n819_n500# a_n919_n588# a_n977_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n588# a_n819_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n588# a_761_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n588# a_n345_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n588# a_603_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n588# a_129_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n588# a_n1451_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n588# a_1235_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n588# a_n503_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n588# a_n29_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n588# a_287_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n588# a_n1609_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n588# a_1393_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n588# a_n1135_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_n503_n500# a_n603_n588# a_n661_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X15 a_1077_n500# a_977_n588# a_919_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n588# a_n187_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n588# a_445_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n588# a_n1293_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n588# a_1077_n500# a_n1743_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_n761_n588# a_503_n588# 0.01fF
C1 a_819_n588# a_977_n588# 0.12fF
C2 a_n445_n588# a_n1077_n588# 0.02fF
C3 a_n761_n588# a_n129_n588# 0.02fF
C4 a_661_n588# a_977_n588# 0.04fF
C5 a_n29_n500# a_1393_n500# 0.05fF
C6 a_n603_n588# a_n1077_n588# 0.02fF
C7 a_n761_n588# a_n287_n588# 0.02fF
C8 a_1235_n500# a_1551_n500# 0.24fF
C9 a_503_n588# a_977_n588# 0.02fF
C10 a_661_n588# a_819_n588# 0.12fF
C11 a_n345_n500# a_129_n500# 0.15fF
C12 a_503_n588# a_819_n588# 0.04fF
C13 a_445_n500# a_761_n500# 0.24fF
C14 a_287_n500# a_919_n500# 0.11fF
C15 a_129_n500# a_1077_n500# 0.07fF
C16 a_287_n500# a_n1135_n500# 0.05fF
C17 a_n1393_n588# a_n1077_n588# 0.04fF
C18 a_n129_n588# a_977_n588# 0.01fF
C19 a_503_n588# a_661_n588# 0.12fF
C20 a_n661_n500# a_287_n500# 0.07fF
C21 a_345_n588# a_n1077_n588# 0.01fF
C22 a_n129_n588# a_819_n588# 0.01fF
C23 a_n287_n588# a_977_n588# 0.01fF
C24 a_187_n588# a_n1077_n588# 0.01fF
C25 a_n1135_n500# a_n1609_n500# 0.15fF
C26 a_n287_n588# a_819_n588# 0.01fF
C27 a_n129_n588# a_661_n588# 0.01fF
C28 a_29_n588# a_n1077_n588# 0.01fF
C29 a_n819_n500# a_761_n500# 0.04fF
C30 a_n661_n500# a_n1609_n500# 0.07fF
C31 a_n287_n588# a_661_n588# 0.01fF
C32 a_n129_n588# a_503_n588# 0.02fF
C33 a_n29_n500# a_129_n500# 0.56fF
C34 a_n761_n588# a_n919_n588# 0.12fF
C35 a_n287_n588# a_503_n588# 0.01fF
C36 a_129_n500# a_1393_n500# 0.05fF
C37 a_n345_n500# a_287_n500# 0.11fF
C38 a_n1235_n588# a_n1077_n588# 0.12fF
C39 a_287_n500# a_1077_n500# 0.09fF
C40 a_445_n500# a_919_n500# 0.15fF
C41 a_603_n500# a_761_n500# 0.56fF
C42 a_445_n500# a_n1135_n500# 0.04fF
C43 a_n287_n588# a_n129_n588# 0.12fF
C44 a_n661_n500# a_445_n500# 0.06fF
C45 a_n603_n588# a_n445_n588# 0.12fF
C46 a_n503_n500# a_761_n500# 0.05fF
C47 a_n345_n500# a_n1609_n500# 0.05fF
C48 a_n1293_n500# a_n1135_n500# 0.56fF
C49 a_661_n588# a_n919_n588# 0.01fF
C50 a_n1393_n588# a_n445_n588# 0.01fF
C51 a_n819_n500# a_n1135_n500# 0.24fF
C52 a_n661_n500# a_n1293_n500# 0.11fF
C53 a_503_n588# a_n919_n588# 0.01fF
C54 a_n1393_n588# a_n603_n588# 0.01fF
C55 a_n445_n588# a_345_n588# 0.01fF
C56 a_n29_n500# a_287_n500# 0.24fF
C57 a_n819_n500# a_n661_n500# 0.56fF
C58 a_287_n500# a_1393_n500# 0.06fF
C59 a_n603_n588# a_345_n588# 0.01fF
C60 a_n445_n588# a_187_n588# 0.02fF
C61 a_n1551_n588# a_n1077_n588# 0.02fF
C62 a_n129_n588# a_n919_n588# 0.01fF
C63 a_n345_n500# a_445_n500# 0.09fF
C64 a_603_n500# a_919_n500# 0.24fF
C65 a_445_n500# a_1077_n500# 0.11fF
C66 a_n445_n588# a_29_n588# 0.02fF
C67 a_n603_n588# a_187_n588# 0.01fF
C68 a_n187_n500# a_761_n500# 0.07fF
C69 a_n29_n500# a_n1609_n500# 0.04fF
C70 a_n287_n588# a_n919_n588# 0.02fF
C71 a_761_n500# a_1235_n500# 0.15fF
C72 a_n1135_n500# a_n977_n500# 0.56fF
C73 a_n603_n588# a_29_n588# 0.02fF
C74 a_n661_n500# a_603_n500# 0.05fF
C75 a_n1393_n588# a_187_n588# 0.01fF
C76 a_n503_n500# a_919_n500# 0.05fF
C77 a_n345_n500# a_n1293_n500# 0.07fF
C78 a_n661_n500# a_n977_n500# 0.24fF
C79 a_n503_n500# a_n1135_n500# 0.11fF
C80 a_n1393_n588# a_29_n588# 0.01fF
C81 a_187_n588# a_345_n588# 0.12fF
C82 a_n661_n500# a_n503_n500# 0.56fF
C83 a_n819_n500# a_n345_n500# 0.15fF
C84 a_n445_n588# a_n1235_n588# 0.01fF
C85 a_29_n588# a_345_n588# 0.04fF
C86 a_n603_n588# a_n1235_n588# 0.02fF
C87 a_n29_n500# a_445_n500# 0.15fF
C88 a_129_n500# a_287_n500# 0.56fF
C89 a_29_n588# a_187_n588# 0.12fF
C90 a_445_n500# a_1393_n500# 0.07fF
C91 a_n1451_n500# a_n1135_n500# 0.24fF
C92 a_761_n500# a_1551_n500# 0.09fF
C93 a_n1393_n588# a_n1235_n588# 0.12fF
C94 a_n661_n500# a_n1451_n500# 0.09fF
C95 a_n345_n500# a_603_n500# 0.07fF
C96 a_603_n500# a_1077_n500# 0.15fF
C97 a_n187_n500# a_919_n500# 0.06fF
C98 a_n1235_n588# a_345_n588# 0.01fF
C99 a_n29_n500# a_n1293_n500# 0.05fF
C100 a_n187_n500# a_n1135_n500# 0.07fF
C101 a_n345_n500# a_n977_n500# 0.11fF
C102 a_919_n500# a_1235_n500# 0.24fF
C103 a_n1235_n588# a_187_n588# 0.01fF
C104 a_n445_n588# a_1135_n588# 0.01fF
C105 a_n661_n500# a_n187_n500# 0.15fF
C106 a_n503_n500# a_n345_n500# 0.56fF
C107 a_n819_n500# a_n29_n500# 0.09fF
C108 a_n503_n500# a_1077_n500# 0.04fF
C109 a_n1235_n588# a_29_n588# 0.01fF
C110 a_n1551_n588# a_n445_n588# 0.01fF
C111 a_1451_n588# a_345_n588# 0.01fF
C112 a_n1551_n588# a_n603_n588# 0.01fF
C113 a_1293_n588# a_345_n588# 0.01fF
C114 a_1451_n588# a_187_n588# 0.01fF
C115 a_n345_n500# a_n1451_n500# 0.06fF
C116 a_129_n500# a_445_n500# 0.24fF
C117 a_n29_n500# a_603_n500# 0.11fF
C118 a_n761_n588# a_n1077_n588# 0.04fF
C119 a_603_n500# a_1393_n500# 0.09fF
C120 a_n1551_n588# a_n1393_n588# 0.12fF
C121 a_1293_n588# a_187_n588# 0.01fF
C122 a_1451_n588# a_29_n588# 0.01fF
C123 a_1135_n588# a_345_n588# 0.01fF
C124 a_n29_n500# a_n977_n500# 0.07fF
C125 a_919_n500# a_1551_n500# 0.11fF
C126 a_1135_n588# a_187_n588# 0.01fF
C127 a_1293_n588# a_29_n588# 0.01fF
C128 a_n345_n500# a_n187_n500# 0.56fF
C129 a_n503_n500# a_n29_n500# 0.15fF
C130 a_n187_n500# a_1077_n500# 0.05fF
C131 a_n345_n500# a_1235_n500# 0.04fF
C132 a_129_n500# a_n1293_n500# 0.05fF
C133 a_1077_n500# a_1235_n500# 0.56fF
C134 a_1135_n588# a_29_n588# 0.01fF
C135 a_n819_n500# a_129_n500# 0.07fF
C136 a_n1551_n588# a_29_n588# 0.01fF
C137 a_n29_n500# a_n1451_n500# 0.05fF
C138 a_503_n588# a_n1077_n588# 0.01fF
C139 a_287_n500# a_445_n500# 0.56fF
C140 a_129_n500# a_603_n500# 0.15fF
C141 a_n1551_n588# a_n1235_n588# 0.04fF
C142 a_n187_n500# a_n29_n500# 0.56fF
C143 a_n187_n500# a_1393_n500# 0.04fF
C144 a_n29_n500# a_1235_n500# 0.05fF
C145 a_129_n500# a_n977_n500# 0.06fF
C146 a_1235_n500# a_1393_n500# 0.56fF
C147 a_1077_n500# a_1551_n500# 0.15fF
C148 a_1293_n588# a_1451_n588# 0.12fF
C149 a_n129_n588# a_n1077_n588# 0.01fF
C150 a_n503_n500# a_129_n500# 0.11fF
C151 a_1135_n588# a_1451_n588# 0.04fF
C152 a_287_n500# a_n1293_n500# 0.04fF
C153 a_n287_n588# a_n1077_n588# 0.01fF
C154 a_n445_n588# a_n761_n588# 0.04fF
C155 a_1135_n588# a_1293_n588# 0.12fF
C156 a_n819_n500# a_287_n500# 0.06fF
C157 a_n603_n588# a_n761_n588# 0.12fF
C158 a_n1293_n500# a_n1609_n500# 0.24fF
C159 a_129_n500# a_n1451_n500# 0.04fF
C160 a_n29_n500# a_1551_n500# 0.04fF
C161 a_n819_n500# a_n1609_n500# 0.09fF
C162 a_1393_n500# a_1551_n500# 0.56fF
C163 a_n1393_n588# a_n761_n588# 0.02fF
C164 a_n445_n588# a_977_n588# 0.01fF
C165 a_287_n500# a_603_n500# 0.24fF
C166 a_n187_n500# a_129_n500# 0.24fF
C167 a_n761_n588# a_345_n588# 0.01fF
C168 a_129_n500# a_1235_n500# 0.06fF
C169 a_n603_n588# a_977_n588# 0.01fF
C170 a_n445_n588# a_819_n588# 0.01fF
C171 a_287_n500# a_n977_n500# 0.05fF
C172 a_n761_n588# a_187_n588# 0.01fF
C173 a_n445_n588# a_661_n588# 0.01fF
C174 a_n603_n588# a_819_n588# 0.01fF
C175 a_n1077_n588# a_n919_n588# 0.12fF
C176 a_n503_n500# a_287_n500# 0.09fF
C177 a_n761_n588# a_29_n588# 0.01fF
C178 a_n445_n588# a_503_n588# 0.01fF
C179 a_n603_n588# a_661_n588# 0.01fF
C180 a_761_n500# a_919_n500# 0.56fF
C181 a_n977_n500# a_n1609_n500# 0.11fF
C182 a_n819_n500# a_445_n500# 0.05fF
C183 a_345_n588# a_977_n588# 0.02fF
C184 a_n603_n588# a_503_n588# 0.01fF
C185 a_n661_n500# a_761_n500# 0.05fF
C186 a_n503_n500# a_n1609_n500# 0.06fF
C187 a_345_n588# a_819_n588# 0.02fF
C188 a_187_n588# a_977_n588# 0.01fF
C189 a_n445_n588# a_n129_n588# 0.04fF
C190 a_345_n588# a_661_n588# 0.04fF
C191 a_29_n588# a_977_n588# 0.01fF
C192 a_187_n588# a_819_n588# 0.02fF
C193 a_129_n500# a_1551_n500# 0.05fF
C194 a_n445_n588# a_n287_n588# 0.12fF
C195 a_n1235_n588# a_n761_n588# 0.02fF
C196 a_n603_n588# a_n129_n588# 0.02fF
C197 a_n819_n500# a_n1293_n500# 0.15fF
C198 a_445_n500# a_603_n500# 0.56fF
C199 a_29_n588# a_819_n588# 0.01fF
C200 a_187_n588# a_661_n588# 0.02fF
C201 a_345_n588# a_503_n588# 0.12fF
C202 a_n603_n588# a_n287_n588# 0.04fF
C203 a_n187_n500# a_287_n500# 0.15fF
C204 a_287_n500# a_1235_n500# 0.07fF
C205 a_n1451_n500# a_n1609_n500# 0.56fF
C206 a_445_n500# a_n977_n500# 0.05fF
C207 a_n1393_n588# a_n129_n588# 0.01fF
C208 a_187_n588# a_503_n588# 0.04fF
C209 a_29_n588# a_661_n588# 0.02fF
C210 a_n503_n500# a_445_n500# 0.07fF
C211 a_n129_n588# a_345_n588# 0.02fF
C212 a_n1393_n588# a_n287_n588# 0.01fF
C213 a_29_n588# a_503_n588# 0.02fF
C214 a_n345_n500# a_761_n500# 0.06fF
C215 a_n187_n500# a_n1609_n500# 0.05fF
C216 a_761_n500# a_1077_n500# 0.24fF
C217 a_n287_n588# a_345_n588# 0.02fF
C218 a_n129_n588# a_187_n588# 0.04fF
C219 a_n1293_n500# a_n977_n500# 0.24fF
C220 a_n819_n500# a_603_n500# 0.05fF
C221 a_n129_n588# a_29_n588# 0.12fF
C222 a_n287_n588# a_187_n588# 0.02fF
C223 a_n661_n500# a_919_n500# 0.04fF
C224 a_n819_n500# a_n977_n500# 0.56fF
C225 a_n661_n500# a_n1135_n500# 0.15fF
C226 a_n503_n500# a_n1293_n500# 0.09fF
C227 a_n1551_n588# a_n761_n588# 0.01fF
C228 a_n287_n588# a_29_n588# 0.04fF
C229 a_1451_n588# a_977_n588# 0.02fF
C230 a_n445_n588# a_n919_n588# 0.02fF
C231 a_n819_n500# a_n503_n500# 0.24fF
C232 a_287_n500# a_1551_n500# 0.05fF
C233 a_1451_n588# a_819_n588# 0.02fF
C234 a_1293_n588# a_977_n588# 0.04fF
C235 a_n603_n588# a_n919_n588# 0.04fF
C236 a_n187_n500# a_445_n500# 0.11fF
C237 a_1135_n588# a_977_n588# 0.12fF
C238 a_1293_n588# a_819_n588# 0.02fF
C239 a_1451_n588# a_661_n588# 0.01fF
C240 a_445_n500# a_1235_n500# 0.09fF
C241 a_n1235_n588# a_n129_n588# 0.01fF
C242 a_n1451_n500# a_n1293_n500# 0.56fF
C243 a_603_n500# a_n977_n500# 0.04fF
C244 a_n29_n500# a_761_n500# 0.09fF
C245 a_761_n500# a_1393_n500# 0.11fF
C246 a_n1393_n588# a_n919_n588# 0.02fF
C247 a_1135_n588# a_819_n588# 0.04fF
C248 a_1451_n588# a_503_n588# 0.01fF
C249 a_1293_n588# a_661_n588# 0.02fF
C250 a_n1235_n588# a_n287_n588# 0.01fF
C251 a_n819_n500# a_n1451_n500# 0.11fF
C252 a_n503_n500# a_603_n500# 0.06fF
C253 a_345_n588# a_n919_n588# 0.01fF
C254 a_1135_n588# a_661_n588# 0.02fF
C255 a_1293_n588# a_503_n588# 0.01fF
C256 a_n345_n500# a_919_n500# 0.05fF
C257 a_n503_n500# a_n977_n500# 0.15fF
C258 a_n187_n500# a_n1293_n500# 0.06fF
C259 a_n345_n500# a_n1135_n500# 0.09fF
C260 a_919_n500# a_1077_n500# 0.56fF
C261 a_187_n588# a_n919_n588# 0.01fF
C262 a_n129_n588# a_1451_n588# 0.01fF
C263 a_1135_n588# a_503_n588# 0.02fF
C264 a_n819_n500# a_n187_n500# 0.11fF
C265 a_n661_n500# a_n345_n500# 0.24fF
C266 a_29_n588# a_n919_n588# 0.01fF
C267 a_n129_n588# a_1293_n588# 0.01fF
C268 a_n287_n588# a_1293_n588# 0.01fF
C269 a_n129_n588# a_1135_n588# 0.01fF
C270 a_445_n500# a_1551_n500# 0.06fF
C271 a_n1451_n500# a_n977_n500# 0.15fF
C272 a_n1551_n588# a_n129_n588# 0.01fF
C273 a_n287_n588# a_1135_n588# 0.01fF
C274 a_n503_n500# a_n1451_n500# 0.07fF
C275 a_n187_n500# a_603_n500# 0.09fF
C276 a_603_n500# a_1235_n500# 0.11fF
C277 a_n1551_n588# a_n287_n588# 0.01fF
C278 a_n1235_n588# a_n919_n588# 0.04fF
C279 a_129_n500# a_761_n500# 0.11fF
C280 a_n29_n500# a_919_n500# 0.07fF
C281 a_n187_n500# a_n977_n500# 0.09fF
C282 a_n29_n500# a_n1135_n500# 0.06fF
C283 a_919_n500# a_1393_n500# 0.15fF
C284 a_n661_n500# a_n29_n500# 0.11fF
C285 a_n503_n500# a_n187_n500# 0.24fF
C286 a_n345_n500# a_1077_n500# 0.05fF
C287 a_n187_n500# a_n1451_n500# 0.05fF
C288 a_603_n500# a_1551_n500# 0.07fF
C289 a_n1551_n588# a_n919_n588# 0.02fF
C290 a_n345_n500# a_n29_n500# 0.24fF
C291 a_n29_n500# a_1077_n500# 0.06fF
C292 a_n187_n500# a_1235_n500# 0.05fF
C293 a_287_n500# a_761_n500# 0.15fF
C294 a_129_n500# a_919_n500# 0.09fF
C295 a_129_n500# a_n1135_n500# 0.05fF
C296 a_n761_n588# a_819_n588# 0.01fF
C297 a_1077_n500# a_1393_n500# 0.24fF
C298 a_n661_n500# a_129_n500# 0.09fF
C299 a_n761_n588# a_661_n588# 0.01fF
C300 a_1551_n500# a_n1743_n722# 0.30fF
C301 a_1393_n500# a_n1743_n722# 0.13fF
C302 a_1235_n500# a_n1743_n722# 0.09fF
C303 a_1077_n500# a_n1743_n722# 0.07fF
C304 a_919_n500# a_n1743_n722# 0.06fF
C305 a_761_n500# a_n1743_n722# 0.05fF
C306 a_603_n500# a_n1743_n722# 0.05fF
C307 a_445_n500# a_n1743_n722# 0.04fF
C308 a_287_n500# a_n1743_n722# 0.04fF
C309 a_129_n500# a_n1743_n722# 0.04fF
C310 a_n29_n500# a_n1743_n722# 0.02fF
C311 a_n187_n500# a_n1743_n722# 0.04fF
C312 a_n345_n500# a_n1743_n722# 0.04fF
C313 a_n503_n500# a_n1743_n722# 0.04fF
C314 a_n661_n500# a_n1743_n722# 0.05fF
C315 a_n819_n500# a_n1743_n722# 0.05fF
C316 a_n977_n500# a_n1743_n722# 0.06fF
C317 a_n1135_n500# a_n1743_n722# 0.07fF
C318 a_n1293_n500# a_n1743_n722# 0.09fF
C319 a_n1451_n500# a_n1743_n722# 0.13fF
C320 a_n1609_n500# a_n1743_n722# 0.30fF
C321 a_1451_n588# a_n1743_n722# 0.28fF
C322 a_1293_n588# a_n1743_n722# 0.23fF
C323 a_1135_n588# a_n1743_n722# 0.24fF
C324 a_977_n588# a_n1743_n722# 0.25fF
C325 a_819_n588# a_n1743_n722# 0.26fF
C326 a_661_n588# a_n1743_n722# 0.26fF
C327 a_503_n588# a_n1743_n722# 0.27fF
C328 a_345_n588# a_n1743_n722# 0.28fF
C329 a_187_n588# a_n1743_n722# 0.28fF
C330 a_29_n588# a_n1743_n722# 0.28fF
C331 a_n129_n588# a_n1743_n722# 0.28fF
C332 a_n287_n588# a_n1743_n722# 0.28fF
C333 a_n445_n588# a_n1743_n722# 0.28fF
C334 a_n603_n588# a_n1743_n722# 0.28fF
C335 a_n761_n588# a_n1743_n722# 0.28fF
C336 a_n919_n588# a_n1743_n722# 0.28fF
C337 a_n1077_n588# a_n1743_n722# 0.28fF
C338 a_n1235_n588# a_n1743_n722# 0.29fF
C339 a_n1393_n588# a_n1743_n722# 0.29fF
C340 a_n1551_n588# a_n1743_n722# 0.34fF
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CADZ46 a_n345_n500# a_n1609_n500# a_n1135_n500#
+ a_29_n597# a_n977_n500# a_n129_n597# a_187_n597# a_n503_n500# a_129_n500# a_n1293_n500#
+ a_n287_n597# a_819_n597# a_n1077_n597# a_287_n500# a_n661_n500# a_345_n597# a_n919_n597#
+ a_n1451_n500# a_977_n597# a_n445_n597# a_919_n500# a_n1235_n597# a_445_n500# a_503_n597#
+ w_n1809_n797# a_n603_n597# a_1077_n500# a_1135_n597# a_661_n597# a_n1393_n597# a_603_n500#
+ a_1293_n597# a_n761_n597# a_1235_n500# a_n1551_n597# a_761_n500# a_n29_n500# a_1451_n597#
+ a_1393_n500# a_n187_n500# a_1551_n500# a_n819_n500# VSUBS
X0 a_n819_n500# a_n919_n597# a_n977_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X1 a_n661_n500# a_n761_n597# a_n819_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X2 a_919_n500# a_819_n597# a_761_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X3 a_n187_n500# a_n287_n597# a_n345_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X4 a_761_n500# a_661_n597# a_603_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X5 a_287_n500# a_187_n597# a_129_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X6 a_n1293_n500# a_n1393_n597# a_n1451_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X7 a_1393_n500# a_1293_n597# a_1235_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X8 a_n345_n500# a_n445_n597# a_n503_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X9 a_129_n500# a_29_n597# a_n29_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X10 a_445_n500# a_345_n597# a_287_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X11 a_n1451_n500# a_n1551_n597# a_n1609_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X12 a_1551_n500# a_1451_n597# a_1393_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X13 a_n977_n500# a_n1077_n597# a_n1135_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=500000u
X14 a_1077_n500# a_977_n597# a_919_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=500000u
X15 a_n503_n500# a_n603_n597# a_n661_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 a_n29_n500# a_n129_n597# a_n187_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X17 a_603_n500# a_503_n597# a_445_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X18 a_n1135_n500# a_n1235_n597# a_n1293_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X19 a_1235_n500# a_1135_n597# a_1077_n500# w_n1809_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
C0 a_345_n597# a_1293_n597# 0.01fF
C1 a_661_n597# a_n761_n597# 0.01fF
C2 a_n761_n597# a_n129_n597# 0.02fF
C3 a_n977_n500# a_n345_n500# 0.11fF
C4 a_661_n597# a_n919_n597# 0.01fF
C5 a_345_n597# a_503_n597# 0.12fF
C6 a_1451_n597# a_187_n597# 0.01fF
C7 a_n1293_n500# a_n345_n500# 0.07fF
C8 w_n1809_n797# a_1451_n597# 0.24fF
C9 a_n129_n597# a_n919_n597# 0.01fF
C10 a_445_n500# a_n345_n500# 0.09fF
C11 w_n1809_n797# a_n1451_n500# 0.13fF
C12 a_n1077_n597# a_503_n597# 0.01fF
C13 a_603_n500# a_1077_n500# 0.15fF
C14 a_761_n500# a_919_n500# 0.56fF
C15 a_n187_n500# a_n1609_n500# 0.05fF
C16 a_n1393_n597# a_n129_n597# 0.01fF
C17 w_n1809_n797# a_1235_n500# 0.09fF
C18 a_n661_n500# a_603_n500# 0.05fF
C19 a_n819_n500# a_n977_n500# 0.56fF
C20 a_n1135_n500# a_n1609_n500# 0.15fF
C21 w_n1809_n797# a_n503_n500# 0.04fF
C22 a_n1293_n500# a_n819_n500# 0.15fF
C23 a_n187_n500# a_761_n500# 0.07fF
C24 a_n819_n500# a_445_n500# 0.05fF
C25 a_287_n500# a_1235_n500# 0.07fF
C26 a_n287_n597# a_n603_n597# 0.04fF
C27 a_977_n597# a_819_n597# 0.12fF
C28 a_287_n500# a_n503_n500# 0.09fF
C29 a_n977_n500# a_n29_n500# 0.07fF
C30 a_919_n500# a_1551_n500# 0.11fF
C31 a_661_n597# a_187_n597# 0.02fF
C32 a_n761_n597# a_503_n597# 0.01fF
C33 a_977_n597# a_29_n597# 0.01fF
C34 a_n129_n597# a_187_n597# 0.04fF
C35 a_n919_n597# a_503_n597# 0.01fF
C36 w_n1809_n797# a_661_n597# 0.22fF
C37 a_n1293_n500# a_n29_n500# 0.05fF
C38 a_445_n500# a_n29_n500# 0.15fF
C39 w_n1809_n797# a_n129_n597# 0.24fF
C40 a_345_n597# a_977_n597# 0.02fF
C41 a_603_n500# a_1393_n500# 0.09fF
C42 a_n1235_n597# a_n287_n597# 0.01fF
C43 a_n661_n500# a_n1609_n500# 0.07fF
C44 a_761_n500# a_1077_n500# 0.24fF
C45 a_n977_n500# a_n1451_n500# 0.15fF
C46 a_n1293_n500# a_n1451_n500# 0.56fF
C47 a_n661_n500# a_761_n500# 0.05fF
C48 a_n819_n500# a_n345_n500# 0.15fF
C49 a_n187_n500# a_919_n500# 0.06fF
C50 a_1293_n597# a_187_n597# 0.01fF
C51 w_n1809_n797# a_1293_n597# 0.19fF
C52 a_503_n597# a_187_n597# 0.04fF
C53 a_445_n500# a_1235_n500# 0.09fF
C54 w_n1809_n797# a_503_n597# 0.23fF
C55 a_n287_n597# a_819_n597# 0.01fF
C56 a_129_n500# a_603_n500# 0.15fF
C57 a_n977_n500# a_n503_n500# 0.15fF
C58 a_n1293_n500# a_n503_n500# 0.09fF
C59 a_n345_n500# a_n29_n500# 0.24fF
C60 a_1077_n500# a_1551_n500# 0.15fF
C61 a_445_n500# a_n503_n500# 0.07fF
C62 a_n287_n597# a_29_n597# 0.04fF
C63 a_n1135_n500# a_n187_n500# 0.07fF
C64 a_345_n597# a_n287_n597# 0.02fF
C65 a_761_n500# a_1393_n500# 0.11fF
C66 a_n1077_n597# a_n287_n597# 0.01fF
C67 a_n1235_n597# a_n603_n597# 0.02fF
C68 a_n819_n500# a_n29_n500# 0.09fF
C69 a_919_n500# a_1077_n500# 0.56fF
C70 a_n345_n500# a_n1451_n500# 0.06fF
C71 w_n1809_n797# a_603_n500# 0.05fF
C72 a_n661_n500# a_919_n500# 0.04fF
C73 a_n187_n500# a_1077_n500# 0.05fF
C74 a_n345_n500# a_1235_n500# 0.04fF
C75 a_1393_n500# a_1551_n500# 0.56fF
C76 a_977_n597# a_187_n597# 0.01fF
C77 w_n1809_n797# a_977_n597# 0.20fF
C78 a_n603_n597# a_819_n597# 0.01fF
C79 a_287_n500# a_603_n500# 0.24fF
C80 a_129_n500# a_761_n500# 0.11fF
C81 a_n503_n500# a_n345_n500# 0.56fF
C82 a_n661_n500# a_n187_n500# 0.15fF
C83 a_n761_n597# a_n287_n597# 0.02fF
C84 a_n287_n597# a_n919_n597# 0.02fF
C85 a_n603_n597# a_29_n597# 0.02fF
C86 a_n819_n500# a_n1451_n500# 0.11fF
C87 a_n1135_n500# a_n661_n500# 0.15fF
C88 a_n1551_n597# a_n445_n597# 0.01fF
C89 a_345_n597# a_n603_n597# 0.01fF
C90 a_n1393_n597# a_n287_n597# 0.01fF
C91 a_919_n500# a_1393_n500# 0.15fF
C92 a_n1077_n597# a_n603_n597# 0.02fF
C93 a_n29_n500# a_n1451_n500# 0.05fF
C94 a_n819_n500# a_n503_n500# 0.24fF
C95 a_n445_n597# a_1135_n597# 0.01fF
C96 w_n1809_n797# a_n1609_n500# 0.30fF
C97 a_129_n500# a_1551_n500# 0.05fF
C98 a_n29_n500# a_1235_n500# 0.05fF
C99 a_n187_n500# a_1393_n500# 0.04fF
C100 a_n1235_n597# a_29_n597# 0.01fF
C101 a_1451_n597# a_1135_n597# 0.04fF
C102 w_n1809_n797# a_761_n500# 0.05fF
C103 a_n503_n500# a_n29_n500# 0.15fF
C104 a_n1235_n597# a_345_n597# 0.01fF
C105 a_n287_n597# a_187_n597# 0.02fF
C106 w_n1809_n797# a_n287_n597# 0.24fF
C107 a_n977_n500# a_603_n500# 0.04fF
C108 a_n1235_n597# a_n1077_n597# 0.12fF
C109 a_129_n500# a_919_n500# 0.09fF
C110 a_287_n500# a_761_n500# 0.15fF
C111 a_445_n500# a_603_n500# 0.56fF
C112 a_n761_n597# a_n603_n597# 0.12fF
C113 a_n603_n597# a_n919_n597# 0.04fF
C114 a_819_n597# a_29_n597# 0.01fF
C115 a_n1551_n597# a_n129_n597# 0.01fF
C116 w_n1809_n797# a_1551_n500# 0.30fF
C117 a_129_n500# a_n187_n500# 0.24fF
C118 a_345_n597# a_819_n597# 0.02fF
C119 a_n1393_n597# a_n603_n597# 0.01fF
C120 a_1077_n500# a_1393_n500# 0.24fF
C121 a_n503_n500# a_n1451_n500# 0.07fF
C122 a_661_n597# a_1135_n597# 0.02fF
C123 a_661_n597# a_n445_n597# 0.01fF
C124 a_n1135_n500# a_129_n500# 0.05fF
C125 a_345_n597# a_29_n597# 0.04fF
C126 a_1135_n597# a_n129_n597# 0.01fF
C127 a_n445_n597# a_n129_n597# 0.04fF
C128 a_287_n500# a_1551_n500# 0.05fF
C129 a_n1077_n597# a_29_n597# 0.01fF
C130 a_n1235_n597# a_n761_n597# 0.02fF
C131 a_1451_n597# a_661_n597# 0.01fF
C132 a_n1235_n597# a_n919_n597# 0.04fF
C133 a_1451_n597# a_n129_n597# 0.01fF
C134 a_n977_n500# a_n1609_n500# 0.11fF
C135 w_n1809_n797# a_919_n500# 0.06fF
C136 a_n1077_n597# a_345_n597# 0.01fF
C137 a_n1293_n500# a_n1609_n500# 0.24fF
C138 a_n1393_n597# a_n1235_n597# 0.12fF
C139 a_n603_n597# a_187_n597# 0.01fF
C140 w_n1809_n797# a_n603_n597# 0.24fF
C141 a_n345_n500# a_603_n500# 0.07fF
C142 w_n1809_n797# a_n187_n500# 0.04fF
C143 a_445_n500# a_761_n500# 0.24fF
C144 a_287_n500# a_919_n500# 0.11fF
C145 a_129_n500# a_1077_n500# 0.07fF
C146 a_n761_n597# a_819_n597# 0.01fF
C147 a_n1135_n500# w_n1809_n797# 0.07fF
C148 a_129_n500# a_n661_n500# 0.09fF
C149 a_1293_n597# a_1135_n597# 0.12fF
C150 a_n761_n597# a_29_n597# 0.01fF
C151 a_1135_n597# a_503_n597# 0.02fF
C152 a_287_n500# a_n187_n500# 0.15fF
C153 a_n445_n597# a_503_n597# 0.01fF
C154 a_29_n597# a_n919_n597# 0.01fF
C155 a_n819_n500# a_603_n500# 0.05fF
C156 a_345_n597# a_n761_n597# 0.01fF
C157 a_1451_n597# a_1293_n597# 0.12fF
C158 a_n1235_n597# a_187_n597# 0.01fF
C159 a_1451_n597# a_503_n597# 0.01fF
C160 a_661_n597# a_n129_n597# 0.01fF
C161 a_345_n597# a_n919_n597# 0.01fF
C162 a_n1235_n597# w_n1809_n797# 0.24fF
C163 a_n1135_n500# a_287_n500# 0.05fF
C164 a_n1393_n597# a_29_n597# 0.01fF
C165 a_445_n500# a_1551_n500# 0.06fF
C166 a_n1077_n597# a_n761_n597# 0.04fF
C167 a_n1077_n597# a_n919_n597# 0.12fF
C168 a_n29_n500# a_603_n500# 0.11fF
C169 a_n345_n500# a_n1609_n500# 0.05fF
C170 w_n1809_n797# a_1077_n500# 0.07fF
C171 a_129_n500# a_1393_n500# 0.05fF
C172 a_n1393_n597# a_n1077_n597# 0.04fF
C173 a_819_n597# a_187_n597# 0.02fF
C174 w_n1809_n797# a_n661_n500# 0.05fF
C175 w_n1809_n797# a_819_n597# 0.21fF
C176 a_n345_n500# a_761_n500# 0.06fF
C177 a_287_n500# a_1077_n500# 0.09fF
C178 a_445_n500# a_919_n500# 0.15fF
C179 a_29_n597# a_187_n597# 0.12fF
C180 w_n1809_n797# a_29_n597# 0.24fF
C181 a_n819_n500# a_n1609_n500# 0.09fF
C182 a_661_n597# a_1293_n597# 0.02fF
C183 a_287_n500# a_n661_n500# 0.07fF
C184 a_n977_n500# a_n187_n500# 0.09fF
C185 a_1293_n597# a_n129_n597# 0.01fF
C186 a_977_n597# a_1135_n597# 0.12fF
C187 a_661_n597# a_503_n597# 0.12fF
C188 a_n761_n597# a_n919_n597# 0.12fF
C189 a_345_n597# a_187_n597# 0.12fF
C190 a_977_n597# a_n445_n597# 0.01fF
C191 a_n129_n597# a_503_n597# 0.02fF
C192 a_n1293_n500# a_n187_n500# 0.06fF
C193 w_n1809_n797# a_345_n597# 0.23fF
C194 a_445_n500# a_n187_n500# 0.11fF
C195 a_n1077_n597# a_187_n597# 0.01fF
C196 a_n819_n500# a_761_n500# 0.04fF
C197 a_n1135_n500# a_n977_n500# 0.56fF
C198 a_1451_n597# a_977_n597# 0.02fF
C199 a_n1077_n597# w_n1809_n797# 0.24fF
C200 a_n1135_n500# a_n1293_n500# 0.56fF
C201 a_n1393_n597# a_n761_n597# 0.02fF
C202 a_n1135_n500# a_445_n500# 0.04fF
C203 a_603_n500# a_1235_n500# 0.11fF
C204 a_n29_n500# a_n1609_n500# 0.04fF
C205 a_n1393_n597# a_n919_n597# 0.02fF
C206 w_n1809_n797# a_1393_n500# 0.13fF
C207 a_n503_n500# a_603_n500# 0.06fF
C208 a_n29_n500# a_761_n500# 0.09fF
C209 a_287_n500# a_1393_n500# 0.06fF
C210 a_n345_n500# a_919_n500# 0.05fF
C211 a_n1551_n597# a_n287_n597# 0.01fF
C212 a_n761_n597# a_187_n597# 0.01fF
C213 a_1293_n597# a_503_n597# 0.01fF
C214 a_n919_n597# a_187_n597# 0.01fF
C215 w_n1809_n797# a_n761_n597# 0.24fF
C216 a_445_n500# a_1077_n500# 0.11fF
C217 w_n1809_n797# a_n919_n597# 0.24fF
C218 a_n1609_n500# a_n1451_n500# 0.56fF
C219 a_n977_n500# a_n661_n500# 0.24fF
C220 w_n1809_n797# a_129_n500# 0.04fF
C221 a_661_n597# a_977_n597# 0.04fF
C222 a_n1293_n500# a_n661_n500# 0.11fF
C223 a_n345_n500# a_n187_n500# 0.56fF
C224 a_445_n500# a_n661_n500# 0.06fF
C225 a_n29_n500# a_1551_n500# 0.04fF
C226 a_977_n597# a_n129_n597# 0.01fF
C227 a_n287_n597# a_1135_n597# 0.01fF
C228 a_n287_n597# a_n445_n597# 0.12fF
C229 a_n1393_n597# a_187_n597# 0.01fF
C230 a_n1393_n597# w_n1809_n797# 0.25fF
C231 a_n1135_n500# a_n345_n500# 0.09fF
C232 a_n503_n500# a_n1609_n500# 0.06fF
C233 a_129_n500# a_287_n500# 0.56fF
C234 a_761_n500# a_1235_n500# 0.15fF
C235 a_n819_n500# a_n187_n500# 0.11fF
C236 a_n503_n500# a_761_n500# 0.05fF
C237 a_n29_n500# a_919_n500# 0.07fF
C238 a_445_n500# a_1393_n500# 0.07fF
C239 a_n1135_n500# a_n819_n500# 0.24fF
C240 w_n1809_n797# a_187_n597# 0.24fF
C241 a_1293_n597# a_977_n597# 0.04fF
C242 a_n345_n500# a_1077_n500# 0.05fF
C243 a_n187_n500# a_n29_n500# 0.56fF
C244 a_n1551_n597# a_n603_n597# 0.01fF
C245 a_1235_n500# a_1551_n500# 0.24fF
C246 a_977_n597# a_503_n597# 0.02fF
C247 a_n661_n500# a_n345_n500# 0.24fF
C248 a_n1135_n500# a_n29_n500# 0.06fF
C249 w_n1809_n797# a_287_n500# 0.04fF
C250 a_661_n597# a_n287_n597# 0.01fF
C251 a_n287_n597# a_n129_n597# 0.12fF
C252 a_n603_n597# a_n445_n597# 0.12fF
C253 a_n977_n500# a_129_n500# 0.06fF
C254 a_n1293_n500# a_129_n500# 0.05fF
C255 a_129_n500# a_445_n500# 0.24fF
C256 a_919_n500# a_1235_n500# 0.24fF
C257 a_n1551_n597# a_n1235_n597# 0.04fF
C258 a_n187_n500# a_n1451_n500# 0.05fF
C259 a_n819_n500# a_n661_n500# 0.56fF
C260 a_n503_n500# a_919_n500# 0.05fF
C261 a_n187_n500# a_1235_n500# 0.05fF
C262 a_n29_n500# a_1077_n500# 0.06fF
C263 a_n1135_n500# a_n1451_n500# 0.24fF
C264 a_n1235_n597# a_n445_n597# 0.01fF
C265 a_n661_n500# a_n29_n500# 0.11fF
C266 a_n503_n500# a_n187_n500# 0.24fF
C267 a_1293_n597# a_n287_n597# 0.01fF
C268 a_n287_n597# a_503_n597# 0.01fF
C269 a_n1135_n500# a_n503_n500# 0.11fF
C270 w_n1809_n797# a_n977_n500# 0.06fF
C271 a_n1551_n597# a_29_n597# 0.01fF
C272 a_n1293_n500# w_n1809_n797# 0.09fF
C273 w_n1809_n797# a_445_n500# 0.04fF
C274 a_661_n597# a_n603_n597# 0.01fF
C275 a_n603_n597# a_n129_n597# 0.02fF
C276 a_819_n597# a_1135_n597# 0.04fF
C277 a_819_n597# a_n445_n597# 0.01fF
C278 a_29_n597# a_1135_n597# 0.01fF
C279 a_129_n500# a_n345_n500# 0.15fF
C280 a_n977_n500# a_287_n500# 0.05fF
C281 a_n445_n597# a_29_n597# 0.02fF
C282 a_1451_n597# a_819_n597# 0.02fF
C283 a_n1551_n597# a_n1077_n597# 0.02fF
C284 a_n1293_n500# a_287_n500# 0.04fF
C285 a_287_n500# a_445_n500# 0.56fF
C286 a_1077_n500# a_1235_n500# 0.56fF
C287 a_n29_n500# a_1393_n500# 0.05fF
C288 a_n661_n500# a_n1451_n500# 0.09fF
C289 a_345_n597# a_1135_n597# 0.01fF
C290 a_345_n597# a_n445_n597# 0.01fF
C291 a_1451_n597# a_29_n597# 0.01fF
C292 a_603_n500# a_761_n500# 0.56fF
C293 a_n503_n500# a_1077_n500# 0.04fF
C294 a_n1077_n597# a_n445_n597# 0.02fF
C295 a_1451_n597# a_345_n597# 0.01fF
C296 a_n1235_n597# a_n129_n597# 0.01fF
C297 a_n661_n500# a_n503_n500# 0.56fF
C298 a_n819_n500# a_129_n500# 0.07fF
C299 a_977_n597# a_n287_n597# 0.01fF
C300 a_n603_n597# a_503_n597# 0.01fF
C301 a_n1551_n597# a_n761_n597# 0.01fF
C302 a_603_n500# a_1551_n500# 0.07fF
C303 w_n1809_n797# a_n345_n500# 0.04fF
C304 a_n1551_n597# a_n919_n597# 0.02fF
C305 a_129_n500# a_n29_n500# 0.56fF
C306 a_661_n597# a_819_n597# 0.12fF
C307 a_819_n597# a_n129_n597# 0.01fF
C308 a_1235_n500# a_1393_n500# 0.56fF
C309 a_661_n597# a_29_n597# 0.02fF
C310 a_n761_n597# a_n445_n597# 0.04fF
C311 a_n1551_n597# a_n1393_n597# 0.12fF
C312 a_n445_n597# a_n919_n597# 0.02fF
C313 a_287_n500# a_n345_n500# 0.11fF
C314 a_n1293_n500# a_n977_n500# 0.24fF
C315 a_29_n597# a_n129_n597# 0.12fF
C316 a_n977_n500# a_445_n500# 0.05fF
C317 a_345_n597# a_661_n597# 0.04fF
C318 a_n819_n500# w_n1809_n797# 0.05fF
C319 a_345_n597# a_n129_n597# 0.02fF
C320 a_603_n500# a_919_n500# 0.24fF
C321 a_n1393_n597# a_n445_n597# 0.01fF
C322 a_n1077_n597# a_n129_n597# 0.01fF
C323 a_129_n500# a_n1451_n500# 0.04fF
C324 a_n819_n500# a_287_n500# 0.06fF
C325 a_n187_n500# a_603_n500# 0.09fF
C326 w_n1809_n797# a_n29_n500# 0.02fF
C327 a_129_n500# a_1235_n500# 0.06fF
C328 a_n1551_n597# w_n1809_n797# 0.30fF
C329 a_977_n597# a_n603_n597# 0.01fF
C330 a_1293_n597# a_819_n597# 0.02fF
C331 a_819_n597# a_503_n597# 0.04fF
C332 a_129_n500# a_n503_n500# 0.11fF
C333 a_761_n500# a_1551_n500# 0.09fF
C334 a_1293_n597# a_29_n597# 0.01fF
C335 a_1135_n597# a_187_n597# 0.01fF
C336 a_n445_n597# a_187_n597# 0.02fF
C337 a_287_n500# a_n29_n500# 0.24fF
C338 a_29_n597# a_503_n597# 0.02fF
C339 w_n1809_n797# a_1135_n597# 0.20fF
C340 w_n1809_n797# a_n445_n597# 0.24fF
C341 w_n1809_n797# VSUBS 17.30fF
.ends

.subckt esd_cell esd VSS VDD
Xsky130_fd_pr__nfet_g5v0d10v5_BRTJC6_0 VSS VSS VSS VSS VSS VSS esd VSS VSS VSS esd
+ VSS esd VSS VSS VSS VSS esd VSS esd esd VSS VSS VSS VSS VSS VSS esd VSS VSS VSS
+ VSS esd VSS VSS esd VSS VSS VSS VSS VSS esd sky130_fd_pr__nfet_g5v0d10v5_BRTJC6
Xsky130_fd_pr__pfet_g5v0d10v5_CADZ46_0 VDD VDD esd VDD VDD VDD VDD esd esd VDD VDD
+ VDD VDD VDD VDD VDD VDD esd VDD VDD VDD VDD esd VDD VDD VDD esd VDD VDD VDD VDD
+ VDD VDD VDD VDD esd VDD VDD esd esd VDD esd VSS sky130_fd_pr__pfet_g5v0d10v5_CADZ46
C0 esd VDD 7.39fF
C1 VDD VSS -181.47fF
C2 esd VSS 8.04fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CEWQ64 c1_n260_n210# m3_n360_n310# VSUBS
X0 c1_n260_n210# m3_n360_n310# sky130_fd_pr__cap_mim_m3_1 l=2.1e+06u w=2.1e+06u
C0 m3_n360_n310# c1_n260_n210# 0.73fF
C1 m3_n360_n310# VSUBS 0.63fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_CGPBWM m3_n1030_n980# c1_n930_n880# VSUBS
X0 c1_n930_n880# m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1 l=8.8e+06u w=8.8e+06u
C0 c1_n930_n880# m3_n1030_n980# 8.32fF
C1 m3_n1030_n980# VSUBS 2.84fF
.ends

.subckt sky130_fd_pr__pfet_01v8_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136# VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_352_n136# a_n416_n136# 0.02fF
C1 a_160_n136# a_448_n136# 0.07fF
C2 a_160_n136# a_n416_n136# 0.03fF
C3 a_n512_n234# a_n320_n136# 0.06fF
C4 a_n224_n136# a_n128_n136# 0.33fF
C5 a_n32_n136# a_352_n136# 0.05fF
C6 a_160_n136# a_n32_n136# 0.12fF
C7 a_64_n136# w_n646_n356# 0.05fF
C8 a_64_n136# a_n508_n136# 0.03fF
C9 a_352_n136# a_256_n136# 0.33fF
C10 a_n128_n136# a_n320_n136# 0.12fF
C11 a_160_n136# a_256_n136# 0.33fF
C12 a_448_n136# w_n646_n356# 0.13fF
C13 a_n508_n136# a_448_n136# 0.02fF
C14 w_n646_n356# a_n416_n136# 0.08fF
C15 a_n508_n136# a_n416_n136# 0.33fF
C16 a_n32_n136# w_n646_n356# 0.05fF
C17 a_n508_n136# a_n32_n136# 0.04fF
C18 w_n646_n356# a_256_n136# 0.06fF
C19 a_n224_n136# a_352_n136# 0.03fF
C20 a_n508_n136# a_256_n136# 0.02fF
C21 a_160_n136# a_n224_n136# 0.05fF
C22 a_n512_n234# a_n128_n136# 0.06fF
C23 a_352_n136# a_n320_n136# 0.03fF
C24 a_64_n136# a_448_n136# 0.05fF
C25 a_160_n136# a_n320_n136# 0.04fF
C26 a_64_n136# a_n416_n136# 0.04fF
C27 a_448_n136# a_n416_n136# 0.02fF
C28 a_n224_n136# w_n646_n356# 0.06fF
C29 a_64_n136# a_n32_n136# 0.33fF
C30 a_n508_n136# a_n224_n136# 0.07fF
C31 a_64_n136# a_256_n136# 0.12fF
C32 a_448_n136# a_n32_n136# 0.04fF
C33 w_n646_n356# a_n320_n136# 0.06fF
C34 a_n32_n136# a_n416_n136# 0.05fF
C35 a_n508_n136# a_n320_n136# 0.12fF
C36 a_448_n136# a_256_n136# 0.12fF
C37 a_256_n136# a_n416_n136# 0.03fF
C38 a_n32_n136# a_256_n136# 0.07fF
C39 a_n128_n136# a_352_n136# 0.04fF
C40 a_160_n136# a_n128_n136# 0.07fF
C41 a_64_n136# a_n224_n136# 0.07fF
C42 a_n512_n234# w_n646_n356# 1.13fF
C43 a_448_n136# a_n224_n136# 0.03fF
C44 a_n512_n234# a_n508_n136# 0.06fF
C45 a_n224_n136# a_n416_n136# 0.12fF
C46 a_64_n136# a_n320_n136# 0.05fF
C47 a_448_n136# a_n320_n136# 0.02fF
C48 a_n320_n136# a_n416_n136# 0.33fF
C49 a_n128_n136# w_n646_n356# 0.05fF
C50 a_n32_n136# a_n224_n136# 0.12fF
C51 a_n508_n136# a_n128_n136# 0.05fF
C52 a_n224_n136# a_256_n136# 0.04fF
C53 a_n32_n136# a_n320_n136# 0.07fF
C54 a_160_n136# a_352_n136# 0.12fF
C55 a_256_n136# a_n320_n136# 0.03fF
C56 a_64_n136# a_n512_n234# 0.06fF
C57 a_n512_n234# a_448_n136# 0.06fF
C58 a_64_n136# a_n128_n136# 0.12fF
C59 w_n646_n356# a_352_n136# 0.08fF
C60 a_n508_n136# a_352_n136# 0.02fF
C61 a_160_n136# w_n646_n356# 0.06fF
C62 a_n508_n136# a_160_n136# 0.03fF
C63 a_448_n136# a_n128_n136# 0.03fF
C64 a_n128_n136# a_n416_n136# 0.07fF
C65 a_n224_n136# a_n320_n136# 0.33fF
C66 a_n512_n234# a_256_n136# 0.06fF
C67 a_n32_n136# a_n128_n136# 0.33fF
C68 a_n508_n136# w_n646_n356# 0.13fF
C69 a_n128_n136# a_256_n136# 0.05fF
C70 a_64_n136# a_352_n136# 0.07fF
C71 a_64_n136# a_160_n136# 0.33fF
C72 a_448_n136# a_352_n136# 0.33fF
C73 w_n646_n356# VSUBS 2.52fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# w_n646_n262#
+ a_448_n52# a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52#
+ a_n320_n52# a_n508_n52# a_64_n52#
X0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_n416_n52# a_n128_n52# 0.03fF
C1 a_64_n52# a_n320_n52# 0.02fF
C2 a_n128_n52# a_n32_n52# 0.13fF
C3 a_n128_n52# a_256_n52# 0.02fF
C4 a_n416_n52# a_n320_n52# 0.13fF
C5 a_n128_n52# a_448_n52# 0.01fF
C6 a_n128_n52# a_n512_n140# 0.09fF
C7 a_n32_n52# a_n320_n52# 0.03fF
C8 a_256_n52# a_n320_n52# 0.01fF
C9 a_n508_n52# a_160_n52# 0.01fF
C10 a_352_n52# a_160_n52# 0.05fF
C11 a_448_n52# a_n320_n52# 0.01fF
C12 a_n512_n140# a_n320_n52# 0.09fF
C13 a_n224_n52# a_64_n52# 0.03fF
C14 a_n416_n52# a_n224_n52# 0.05fF
C15 a_352_n52# a_n508_n52# 0.01fF
C16 a_n224_n52# a_n32_n52# 0.05fF
C17 a_n128_n52# a_160_n52# 0.03fF
C18 a_n224_n52# a_256_n52# 0.02fF
C19 a_n416_n52# a_64_n52# 0.02fF
C20 a_n224_n52# a_448_n52# 0.01fF
C21 a_160_n52# a_n320_n52# 0.02fF
C22 a_64_n52# a_n32_n52# 0.13fF
C23 a_256_n52# a_64_n52# 0.05fF
C24 a_n128_n52# a_n508_n52# 0.02fF
C25 a_352_n52# a_n128_n52# 0.02fF
C26 a_n416_n52# a_n32_n52# 0.02fF
C27 a_n416_n52# a_256_n52# 0.01fF
C28 a_448_n52# a_64_n52# 0.02fF
C29 a_64_n52# a_n512_n140# 0.09fF
C30 a_n508_n52# a_n320_n52# 0.05fF
C31 a_352_n52# a_n320_n52# 0.01fF
C32 a_n416_n52# a_448_n52# 0.01fF
C33 a_256_n52# a_n32_n52# 0.03fF
C34 a_448_n52# a_n32_n52# 0.02fF
C35 a_256_n52# a_448_n52# 0.05fF
C36 a_256_n52# a_n512_n140# 0.09fF
C37 a_n224_n52# a_160_n52# 0.02fF
C38 a_448_n52# a_n512_n140# 0.09fF
C39 a_n128_n52# a_n320_n52# 0.05fF
C40 a_64_n52# a_160_n52# 0.13fF
C41 a_n224_n52# a_n508_n52# 0.03fF
C42 a_352_n52# a_n224_n52# 0.01fF
C43 a_n416_n52# a_160_n52# 0.01fF
C44 a_n508_n52# a_64_n52# 0.01fF
C45 a_160_n52# a_n32_n52# 0.05fF
C46 a_256_n52# a_160_n52# 0.13fF
C47 a_352_n52# a_64_n52# 0.03fF
C48 a_n416_n52# a_n508_n52# 0.13fF
C49 a_n416_n52# a_352_n52# 0.01fF
C50 a_n128_n52# a_n224_n52# 0.13fF
C51 a_448_n52# a_160_n52# 0.03fF
C52 a_n508_n52# a_n32_n52# 0.02fF
C53 a_n508_n52# a_256_n52# 0.01fF
C54 a_352_n52# a_n32_n52# 0.02fF
C55 a_352_n52# a_256_n52# 0.13fF
C56 a_n224_n52# a_n320_n52# 0.13fF
C57 a_n128_n52# a_64_n52# 0.05fF
C58 a_n508_n52# a_448_n52# 0.01fF
C59 a_n508_n52# a_n512_n140# 0.09fF
C60 a_352_n52# a_448_n52# 0.13fF
C61 a_448_n52# a_n610_n226# 0.07fF
C62 a_352_n52# a_n610_n226# 0.05fF
C63 a_256_n52# a_n610_n226# 0.04fF
C64 a_160_n52# a_n610_n226# 0.04fF
C65 a_64_n52# a_n610_n226# 0.04fF
C66 a_n32_n52# a_n610_n226# 0.04fF
C67 a_n128_n52# a_n610_n226# 0.04fF
C68 a_n224_n52# a_n610_n226# 0.04fF
C69 a_n320_n52# a_n610_n226# 0.04fF
C70 a_n416_n52# a_n610_n226# 0.05fF
C71 a_n508_n52# a_n610_n226# 0.07fF
C72 a_n512_n140# a_n610_n226# 1.45fF
.ends

.subckt transmission_gate en VDD sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# in
+ out VSS en_b
Xsky130_fd_pr__pfet_01v8_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ VSS sky130_fd_pr__pfet_01v8_UNG2NQ
Xsky130_fd_pr__nfet_01v8_6J4AMR_0 out in in sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ out in in VSS out en in out out out sky130_fd_pr__nfet_01v8_6J4AMR
C0 VDD out 0.40fF
C1 en_b out 0.03fF
C2 in en 1.30fF
C3 VDD en 0.05fF
C4 VDD in 0.92fF
C5 en_b en 0.14fF
C6 out en 0.05fF
C7 en_b in 1.18fF
C8 en_b VDD 0.10fF
C9 out in 0.71fF
C10 en VSS 1.66fF
C11 out VSS 1.04fF
C12 in VSS 1.15fF
C13 en_b VSS 0.24fF
C14 VDD VSS 3.18fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_II a_n207_n140# a_n1039_n205# a_1275_n205# a_29_n205#
+ a_327_n140# a_n1275_n140# a_n683_n205# a_741_n205# a_n29_n140# a_149_n140# a_n1097_n140#
+ a_1097_n205# a_1395_n140# a_n505_n205# a_n741_n140# a_563_n205# a_861_n140# a_919_n205#
+ a_n327_n205# a_n563_n140# a_385_n205# a_1217_n140# a_n1395_n205# a_683_n140# a_n919_n140#
+ a_n149_n205# w_n1489_n241# a_1039_n140# a_n385_n140# a_207_n205# a_n1217_n205# a_505_n140#
+ a_n1453_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1395_n140# a_1275_n205# a_1217_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_327_n140# a_207_n205# a_149_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_149_n140# a_29_n205# a_n29_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_861_n140# a_741_n205# a_683_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n207_n140# a_n327_n205# a_n385_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_1217_n140# a_1097_n205# a_1039_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n1275_n140# a_n1395_n205# a_n1453_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n205# a_n919_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1217_n205# a_n1275_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n205# a_505_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n205# a_861_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n29_n140# a_n149_n205# a_n207_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_n563_n140# a_n683_n205# a_n741_n140# w_n1489_n241# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_327_n140# a_n1275_n140# 0.01fF
C1 a_919_n205# a_1097_n205# 0.11fF
C2 a_n29_n140# a_n563_n140# 0.04fF
C3 a_861_n140# a_327_n140# 0.04fF
C4 a_n741_n140# w_n1489_n241# 0.02fF
C5 a_n1453_n140# a_n207_n140# 0.02fF
C6 a_1097_n205# w_n1489_n241# 0.18fF
C7 a_n1097_n140# a_n563_n140# 0.04fF
C8 a_1395_n140# a_1217_n140# 0.13fF
C9 a_149_n140# w_n1489_n241# 0.02fF
C10 a_n919_n140# w_n1489_n241# 0.02fF
C11 a_207_n205# a_n1395_n205# 0.01fF
C12 a_n861_n205# a_n505_n205# 0.03fF
C13 a_385_n205# a_n1039_n205# 0.01fF
C14 a_n1217_n205# a_207_n205# 0.01fF
C15 a_149_n140# a_1039_n140# 0.02fF
C16 a_n1453_n140# a_n563_n140# 0.02fF
C17 a_207_n205# a_29_n205# 0.11fF
C18 a_n149_n205# a_1275_n205# 0.01fF
C19 a_741_n205# a_n861_n205# 0.01fF
C20 a_1217_n140# a_n29_n140# 0.02fF
C21 a_n741_n140# a_n207_n140# 0.04fF
C22 a_385_n205# a_n149_n205# 0.02fF
C23 a_505_n140# w_n1489_n241# 0.02fF
C24 a_149_n140# a_n207_n140# 0.06fF
C25 a_n1275_n140# w_n1489_n241# 0.02fF
C26 a_861_n140# w_n1489_n241# 0.02fF
C27 a_n919_n140# a_n207_n140# 0.03fF
C28 a_n1395_n205# a_n327_n205# 0.01fF
C29 a_505_n140# a_1039_n140# 0.04fF
C30 a_n1217_n205# a_n327_n205# 0.01fF
C31 a_n741_n140# a_n563_n140# 0.13fF
C32 a_n327_n205# a_29_n205# 0.03fF
C33 a_n861_n205# a_n1039_n205# 0.11fF
C34 a_861_n140# a_1039_n140# 0.13fF
C35 a_149_n140# a_n563_n140# 0.03fF
C36 a_n919_n140# a_n563_n140# 0.06fF
C37 a_29_n205# a_563_n205# 0.02fF
C38 a_505_n140# a_n207_n140# 0.03fF
C39 a_n207_n140# a_n1275_n140# 0.02fF
C40 a_1097_n205# a_n505_n205# 0.01fF
C41 a_861_n140# a_n207_n140# 0.02fF
C42 a_n149_n205# a_n861_n205# 0.01fF
C43 a_741_n205# a_1097_n205# 0.03fF
C44 a_683_n140# a_n385_n140# 0.02fF
C45 a_385_n205# a_1275_n205# 0.01fF
C46 a_505_n140# a_n563_n140# 0.02fF
C47 a_n1275_n140# a_n563_n140# 0.03fF
C48 a_1217_n140# a_149_n140# 0.02fF
C49 a_861_n140# a_n563_n140# 0.01fF
C50 a_919_n205# a_29_n205# 0.01fF
C51 a_n1395_n205# w_n1489_n241# 0.31fF
C52 a_327_n140# a_n385_n140# 0.03fF
C53 a_n1217_n205# w_n1489_n241# 0.24fF
C54 w_n1489_n241# a_29_n205# 0.24fF
C55 a_207_n205# a_n327_n205# 0.02fF
C56 a_1217_n140# a_505_n140# 0.03fF
C57 a_1217_n140# a_861_n140# 0.06fF
C58 a_n149_n205# a_1097_n205# 0.01fF
C59 a_207_n205# a_563_n205# 0.03fF
C60 a_n683_n205# a_n1395_n205# 0.01fF
C61 a_n1217_n205# a_n683_n205# 0.02fF
C62 a_385_n205# a_n861_n205# 0.01fF
C63 a_n683_n205# a_29_n205# 0.01fF
C64 a_683_n140# a_327_n140# 0.06fF
C65 a_1395_n140# a_n29_n140# 0.01fF
C66 a_n385_n140# w_n1489_n241# 0.02fF
C67 a_n327_n205# a_563_n205# 0.01fF
C68 a_n385_n140# a_1039_n140# 0.01fF
C69 a_207_n205# a_919_n205# 0.01fF
C70 a_n1395_n205# a_n505_n205# 0.01fF
C71 a_n1217_n205# a_n505_n205# 0.01fF
C72 a_207_n205# w_n1489_n241# 0.23fF
C73 a_n505_n205# a_29_n205# 0.02fF
C74 a_1275_n205# a_1097_n205# 0.11fF
C75 a_n1097_n140# a_n29_n140# 0.02fF
C76 a_n385_n140# a_n207_n140# 0.13fF
C77 a_741_n205# a_29_n205# 0.01fF
C78 a_385_n205# a_1097_n205# 0.01fF
C79 a_683_n140# w_n1489_n241# 0.02fF
C80 a_n1453_n140# a_n29_n140# 0.01fF
C81 a_919_n205# a_n327_n205# 0.01fF
C82 a_n385_n140# a_n563_n140# 0.13fF
C83 a_207_n205# a_n683_n205# 0.01fF
C84 a_n1453_n140# a_n1097_n140# 0.06fF
C85 a_683_n140# a_1039_n140# 0.06fF
C86 a_n327_n205# w_n1489_n241# 0.24fF
C87 a_n1395_n205# a_n1039_n205# 0.03fF
C88 a_919_n205# a_563_n205# 0.03fF
C89 a_1395_n140# a_149_n140# 0.02fF
C90 a_n1217_n205# a_n1039_n205# 0.11fF
C91 a_327_n140# w_n1489_n241# 0.02fF
C92 a_29_n205# a_n1039_n205# 0.01fF
C93 w_n1489_n241# a_563_n205# 0.21fF
C94 a_683_n140# a_n207_n140# 0.02fF
C95 a_327_n140# a_1039_n140# 0.03fF
C96 a_n741_n140# a_n29_n140# 0.03fF
C97 a_n149_n205# a_n1395_n205# 0.01fF
C98 a_149_n140# a_n29_n140# 0.13fF
C99 a_n1217_n205# a_n149_n205# 0.01fF
C100 a_n741_n140# a_n1097_n140# 0.06fF
C101 a_n683_n205# a_n327_n205# 0.03fF
C102 a_1217_n140# a_n385_n140# 0.01fF
C103 a_n149_n205# a_29_n205# 0.11fF
C104 a_n919_n140# a_n29_n140# 0.02fF
C105 a_1395_n140# a_505_n140# 0.02fF
C106 a_n1097_n140# a_149_n140# 0.02fF
C107 a_683_n140# a_n563_n140# 0.02fF
C108 a_207_n205# a_n505_n205# 0.01fF
C109 a_327_n140# a_n207_n140# 0.04fF
C110 a_1395_n140# a_861_n140# 0.04fF
C111 a_n683_n205# a_563_n205# 0.01fF
C112 a_n919_n140# a_n1097_n140# 0.13fF
C113 a_n1453_n140# a_n741_n140# 0.03fF
C114 a_207_n205# a_741_n205# 0.02fF
C115 a_919_n205# w_n1489_n241# 0.19fF
C116 a_n1453_n140# a_149_n140# 0.01fF
C117 a_505_n140# a_n29_n140# 0.04fF
C118 a_327_n140# a_n563_n140# 0.02fF
C119 a_n919_n140# a_n1453_n140# 0.04fF
C120 a_n29_n140# a_n1275_n140# 0.02fF
C121 a_861_n140# a_n29_n140# 0.02fF
C122 a_n1097_n140# a_505_n140# 0.01fF
C123 a_1039_n140# w_n1489_n241# 0.02fF
C124 a_n1097_n140# a_n1275_n140# 0.13fF
C125 a_n327_n205# a_n505_n205# 0.11fF
C126 a_683_n140# a_1217_n140# 0.04fF
C127 a_919_n205# a_n683_n205# 0.01fF
C128 a_207_n205# a_n1039_n205# 0.01fF
C129 a_741_n205# a_n327_n205# 0.01fF
C130 a_1275_n205# a_29_n205# 0.01fF
C131 a_n741_n140# a_149_n140# 0.02fF
C132 a_n505_n205# a_563_n205# 0.01fF
C133 a_n683_n205# w_n1489_n241# 0.24fF
C134 a_n1453_n140# a_n1275_n140# 0.13fF
C135 a_n207_n140# w_n1489_n241# 0.02fF
C136 a_385_n205# a_n1217_n205# 0.01fF
C137 a_n919_n140# a_n741_n140# 0.13fF
C138 a_741_n205# a_563_n205# 0.11fF
C139 a_385_n205# a_29_n205# 0.03fF
C140 a_1217_n140# a_327_n140# 0.02fF
C141 a_207_n205# a_n149_n205# 0.03fF
C142 a_n919_n140# a_149_n140# 0.02fF
C143 a_1039_n140# a_n207_n140# 0.02fF
C144 w_n1489_n241# a_n563_n140# 0.02fF
C145 a_n327_n205# a_n1039_n205# 0.01fF
C146 a_n741_n140# a_505_n140# 0.02fF
C147 a_919_n205# a_n505_n205# 0.01fF
C148 a_n741_n140# a_n1275_n140# 0.04fF
C149 a_1039_n140# a_n563_n140# 0.01fF
C150 a_861_n140# a_n741_n140# 0.01fF
C151 a_149_n140# a_505_n140# 0.06fF
C152 a_n1039_n205# a_563_n205# 0.01fF
C153 a_149_n140# a_n1275_n140# 0.01fF
C154 a_n861_n205# a_n1395_n205# 0.02fF
C155 a_861_n140# a_149_n140# 0.03fF
C156 a_n505_n205# w_n1489_n241# 0.24fF
C157 a_919_n205# a_741_n205# 0.11fF
C158 a_n919_n140# a_505_n140# 0.01fF
C159 a_n1217_n205# a_n861_n205# 0.03fF
C160 a_n149_n205# a_n327_n205# 0.11fF
C161 a_n919_n140# a_n1275_n140# 0.06fF
C162 a_n861_n205# a_29_n205# 0.01fF
C163 a_741_n205# w_n1489_n241# 0.20fF
C164 a_n207_n140# a_n563_n140# 0.06fF
C165 a_1217_n140# w_n1489_n241# 0.02fF
C166 a_n149_n205# a_563_n205# 0.01fF
C167 a_207_n205# a_1275_n205# 0.01fF
C168 a_1217_n140# a_1039_n140# 0.13fF
C169 a_n683_n205# a_n505_n205# 0.11fF
C170 a_861_n140# a_505_n140# 0.06fF
C171 a_385_n205# a_207_n205# 0.11fF
C172 w_n1489_n241# a_n1039_n205# 0.24fF
C173 a_n683_n205# a_741_n205# 0.01fF
C174 a_1217_n140# a_n207_n140# 0.01fF
C175 a_n29_n140# a_n385_n140# 0.06fF
C176 a_919_n205# a_n149_n205# 0.01fF
C177 a_1275_n205# a_n327_n205# 0.01fF
C178 a_n1097_n140# a_n385_n140# 0.03fF
C179 a_n149_n205# w_n1489_n241# 0.24fF
C180 a_1097_n205# a_29_n205# 0.01fF
C181 a_385_n205# a_n327_n205# 0.01fF
C182 a_683_n140# a_1395_n140# 0.03fF
C183 a_1275_n205# a_563_n205# 0.01fF
C184 a_n683_n205# a_n1039_n205# 0.03fF
C185 a_207_n205# a_n861_n205# 0.01fF
C186 a_n1453_n140# a_n385_n140# 0.02fF
C187 a_385_n205# a_563_n205# 0.11fF
C188 a_741_n205# a_n505_n205# 0.01fF
C189 a_1395_n140# a_327_n140# 0.02fF
C190 a_n683_n205# a_n149_n205# 0.02fF
C191 a_683_n140# a_n29_n140# 0.03fF
C192 a_919_n205# a_1275_n205# 0.03fF
C193 a_n741_n140# a_n385_n140# 0.06fF
C194 a_n861_n205# a_n327_n205# 0.02fF
C195 a_n505_n205# a_n1039_n205# 0.02fF
C196 a_149_n140# a_n385_n140# 0.04fF
C197 a_1275_n205# w_n1489_n241# 0.24fF
C198 a_327_n140# a_n29_n140# 0.06fF
C199 a_385_n205# a_919_n205# 0.02fF
C200 a_n861_n205# a_563_n205# 0.01fF
C201 a_n919_n140# a_n385_n140# 0.04fF
C202 a_327_n140# a_n1097_n140# 0.01fF
C203 a_385_n205# w_n1489_n241# 0.22fF
C204 a_207_n205# a_1097_n205# 0.01fF
C205 a_n149_n205# a_n505_n205# 0.03fF
C206 a_1395_n140# w_n1489_n241# 0.02fF
C207 a_741_n205# a_n149_n205# 0.01fF
C208 a_505_n140# a_n385_n140# 0.02fF
C209 a_n385_n140# a_n1275_n140# 0.02fF
C210 a_683_n140# a_n741_n140# 0.01fF
C211 a_861_n140# a_n385_n140# 0.02fF
C212 a_1395_n140# a_1039_n140# 0.06fF
C213 a_385_n205# a_n683_n205# 0.01fF
C214 a_683_n140# a_149_n140# 0.04fF
C215 a_683_n140# a_n919_n140# 0.01fF
C216 a_n29_n140# w_n1489_n241# 0.02fF
C217 a_n327_n205# a_1097_n205# 0.01fF
C218 a_n1217_n205# a_n1395_n205# 0.11fF
C219 a_n861_n205# w_n1489_n241# 0.24fF
C220 a_n1395_n205# a_29_n205# 0.01fF
C221 a_327_n140# a_n741_n140# 0.02fF
C222 a_n1217_n205# a_29_n205# 0.01fF
C223 a_1395_n140# a_n207_n140# 0.01fF
C224 a_n1097_n140# w_n1489_n241# 0.02fF
C225 a_n149_n205# a_n1039_n205# 0.01fF
C226 a_n29_n140# a_1039_n140# 0.02fF
C227 a_327_n140# a_149_n140# 0.13fF
C228 a_1097_n205# a_563_n205# 0.02fF
C229 a_n919_n140# a_327_n140# 0.02fF
C230 a_683_n140# a_505_n140# 0.13fF
C231 a_n1453_n140# w_n1489_n241# 0.02fF
C232 a_683_n140# a_861_n140# 0.13fF
C233 a_n683_n205# a_n861_n205# 0.11fF
C234 a_741_n205# a_1275_n205# 0.02fF
C235 a_n29_n140# a_n207_n140# 0.13fF
C236 a_385_n205# a_n505_n205# 0.01fF
C237 a_n1097_n140# a_n207_n140# 0.02fF
C238 a_385_n205# a_741_n205# 0.03fF
C239 a_327_n140# a_505_n140# 0.13fF
C240 w_n1489_n241# VSUBS 4.31fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FF a_20_n120# a_n78_n120# a_n33_n208# VSUBS
X0 a_20_n120# a_n33_n208# a_n78_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
C0 a_n33_n208# a_20_n120# 0.02fF
C1 a_n78_n120# a_20_n120# 0.28fF
C2 a_n78_n120# a_n33_n208# 0.02fF
C3 a_20_n120# VSUBS 0.02fF
C4 a_n78_n120# VSUBS 0.02fF
C5 a_n33_n208# VSUBS 0.29fF
.ends

.subckt sky130_fd_pr__nfet_01v8_DD a_1751_n140# a_n149_n194# a_1987_n194# a_n2819_n194#
+ a_n207_n140# a_n1809_n140# a_n2877_n140# a_207_n194# a_n2285_n194# a_1453_n194#
+ a_n1217_n194# a_n3353_n194# a_327_n140# a_n1275_n140# a_n2343_n140# a_2521_n194#
+ a_n861_n194# a_1573_n140# a_n3411_n140# a_2641_n140# a_n2699_n140# a_2877_n194#
+ a_1809_n194# a_2997_n140# a_n29_n140# a_n1039_n194# a_n3175_n194# a_1929_n140# a_149_n140#
+ a_n1097_n140# a_2343_n194# a_1275_n194# a_29_n194# a_n2107_n194# a_n2165_n140# a_n3233_n140#
+ a_3411_n194# a_n683_n194# a_1395_n140# a_3531_n140# a_2463_n140# a_n741_n140# a_2699_n194#
+ a_741_n194# a_n3589_n140# a_n1751_n194# a_861_n140# a_1097_n194# a_2819_n140# a_3233_n194#
+ a_2165_n194# a_n3055_n140# a_n505_n194# a_2285_n140# a_n563_n140# a_563_n194# a_3353_n140#
+ a_1217_n140# a_n1573_n194# a_n2641_n194# a_683_n140# a_n919_n140# a_n1631_n140#
+ a_919_n194# a_3055_n194# a_n2997_n194# a_n1987_n140# a_n327_n194# a_n1929_n194#
+ a_3175_n140# a_1039_n140# a_n385_n140# a_385_n194# a_2107_n140# a_n1395_n194# a_n2463_n194#
+ a_n3531_n194# a_505_n140# a_n1453_n140# a_1631_n194# a_n2521_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2165_n140# a_n2285_n194# a_n2343_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_3175_n140# a_3055_n194# a_2997_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n3233_n140# a_n3353_n194# a_n3411_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_2997_n140# a_2877_n194# a_2819_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1987_n140# a_n2107_n194# a_n2165_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1809_n140# a_n1929_n194# a_n1987_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n1453_n140# a_n1573_n194# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2463_n140# a_2343_n194# a_2285_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n2521_n140# a_n2641_n194# a_n2699_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_3531_n140# a_3411_n194# a_3353_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1751_n140# a_1631_n194# a_1573_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n3055_n140# a_n3175_n194# a_n3233_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_2819_n140# a_2699_n194# a_2641_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n2877_n140# a_n2997_n194# a_n3055_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_2285_n140# a_2165_n194# a_2107_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_n2699_n140# a_n2819_n194# a_n2877_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n2343_n140# a_n2463_n194# a_n2521_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_2107_n140# a_1987_n194# a_1929_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X31 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_3353_n140# a_3233_n194# a_3175_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_n3411_n140# a_n3531_n194# a_n3589_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X36 a_1573_n140# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_1929_n140# a_1809_n194# a_1751_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_n1631_n140# a_n1751_n194# a_n1809_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_2641_n140# a_2521_n194# a_2463_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1395_n194# a_n2641_n194# 0.01fF
C1 a_n563_n140# a_149_n140# 0.03fF
C2 a_n1395_n194# a_n1573_n194# 0.10fF
C3 a_n3233_n140# a_n1809_n140# 0.01fF
C4 a_n3353_n194# a_n2819_n194# 0.02fF
C5 a_n207_n140# a_327_n140# 0.04fF
C6 a_n385_n140# a_505_n140# 0.02fF
C7 a_n29_n140# a_149_n140# 0.13fF
C8 a_n2107_n194# a_n1039_n194# 0.01fF
C9 a_n3411_n140# a_n3589_n140# 0.13fF
C10 a_n1929_n194# a_n3175_n194# 0.01fF
C11 a_n563_n140# a_n29_n140# 0.04fF
C12 a_n3589_n140# a_n2343_n140# 0.02fF
C13 a_1631_n194# a_2877_n194# 0.01fF
C14 a_n2285_n194# a_n2819_n194# 0.02fF
C15 a_n207_n140# a_149_n140# 0.06fF
C16 a_n385_n140# a_327_n140# 0.03fF
C17 a_n2463_n194# a_n1395_n194# 0.01fF
C18 a_2343_n194# a_2165_n194# 0.10fF
C19 a_n563_n140# a_n207_n140# 0.06fF
C20 a_n207_n140# a_n29_n140# 0.13fF
C21 a_n385_n140# a_149_n140# 0.04fF
C22 a_2877_n194# a_3055_n194# 0.10fF
C23 a_385_n194# a_29_n194# 0.03fF
C24 a_n683_n194# a_919_n194# 0.01fF
C25 a_n861_n194# a_563_n194# 0.01fF
C26 a_n563_n140# a_n385_n140# 0.13fF
C27 a_741_n194# a_n683_n194# 0.01fF
C28 a_n385_n140# a_n29_n140# 0.06fF
C29 a_n1929_n194# a_n2819_n194# 0.01fF
C30 a_n2521_n140# a_n919_n140# 0.01fF
C31 a_n1809_n140# a_n1631_n140# 0.13fF
C32 a_n2165_n140# a_n1275_n140# 0.02fF
C33 a_n2343_n140# a_n1097_n140# 0.02fF
C34 a_n1987_n140# a_n1453_n140# 0.04fF
C35 a_n683_n194# a_n505_n194# 0.10fF
C36 a_2343_n194# a_2521_n194# 0.10fF
C37 a_n327_n194# a_n1751_n194# 0.01fF
C38 a_n1217_n194# a_385_n194# 0.01fF
C39 a_n385_n140# a_n207_n140# 0.13fF
C40 a_n1395_n194# a_n2107_n194# 0.01fF
C41 a_n2641_n194# a_n3175_n194# 0.02fF
C42 a_n1217_n194# a_n2285_n194# 0.01fF
C43 a_n1573_n194# a_n3175_n194# 0.01fF
C44 a_1631_n194# a_919_n194# 0.01fF
C45 a_1809_n194# a_3233_n194# 0.01fF
C46 a_1631_n194# a_741_n194# 0.01fF
C47 a_n861_n194# a_n327_n194# 0.02fF
C48 a_1453_n194# a_1097_n194# 0.03fF
C49 a_n3531_n194# a_n3175_n194# 0.03fF
C50 a_n3589_n140# a_n1987_n140# 0.01fF
C51 a_1809_n194# a_1097_n194# 0.01fF
C52 a_n3055_n140# a_n2699_n140# 0.06fF
C53 a_n2463_n194# a_n3175_n194# 0.01fF
C54 a_2165_n194# a_3411_n194# 0.01fF
C55 a_919_n194# a_n149_n194# 0.01fF
C56 a_n1929_n194# a_n1217_n194# 0.01fF
C57 a_1631_n194# a_1275_n194# 0.03fF
C58 a_1453_n194# a_1987_n194# 0.02fF
C59 a_n3233_n140# a_n3589_n140# 0.06fF
C60 a_741_n194# a_n149_n194# 0.01fF
C61 a_n2641_n194# a_n2819_n194# 0.10fF
C62 a_n1573_n194# a_n2819_n194# 0.01fF
C63 a_n149_n194# a_n505_n194# 0.03fF
C64 a_385_n194# a_563_n194# 0.10fF
C65 a_1809_n194# a_1987_n194# 0.10fF
C66 a_n3531_n194# a_n2819_n194# 0.01fF
C67 a_n2343_n140# a_n741_n140# 0.01fF
C68 a_n1987_n140# a_n1097_n140# 0.02fF
C69 a_n1809_n140# a_n1275_n140# 0.04fF
C70 a_n1631_n140# a_n1453_n140# 0.13fF
C71 a_n2165_n140# a_n919_n140# 0.02fF
C72 a_2343_n194# a_2699_n194# 0.03fF
C73 a_n149_n194# a_1275_n194# 0.01fF
C74 a_3411_n194# a_2521_n194# 0.01fF
C75 a_2877_n194# a_3233_n194# 0.03fF
C76 a_n2463_n194# a_n2819_n194# 0.03fF
C77 a_207_n194# a_1453_n194# 0.01fF
C78 a_n505_n194# a_n1039_n194# 0.02fF
C79 a_n3175_n194# a_n2107_n194# 0.01fF
C80 a_1809_n194# a_207_n194# 0.01fF
C81 a_n1573_n194# a_29_n194# 0.01fF
C82 a_n327_n194# a_385_n194# 0.01fF
C83 a_n2641_n194# a_n1217_n194# 0.01fF
C84 a_n1217_n194# a_n1573_n194# 0.03fF
C85 a_n3411_n140# a_n3055_n140# 0.06fF
C86 a_n2877_n140# a_n2521_n140# 0.06fF
C87 a_n3055_n140# a_n2343_n140# 0.03fF
C88 a_2877_n194# a_1987_n194# 0.01fF
C89 a_n861_n194# a_n1751_n194# 0.01fF
C90 a_n2107_n194# a_n2819_n194# 0.01fF
C91 a_n2463_n194# a_n1217_n194# 0.01fF
C92 a_n1987_n140# a_n741_n140# 0.02fF
C93 a_n1631_n140# a_n1097_n140# 0.04fF
C94 a_n2165_n140# a_n563_n140# 0.01fF
C95 a_n1453_n140# a_n1275_n140# 0.13fF
C96 a_n1809_n140# a_n919_n140# 0.02fF
C97 a_n1929_n194# a_n327_n194# 0.01fF
C98 a_n1395_n194# a_n505_n194# 0.01fF
C99 a_3411_n194# a_2699_n194# 0.01fF
C100 a_919_n194# a_1097_n194# 0.10fF
C101 a_741_n194# a_1097_n194# 0.03fF
C102 a_1453_n194# a_29_n194# 0.01fF
C103 a_1097_n194# a_n505_n194# 0.01fF
C104 a_919_n194# a_1987_n194# 0.01fF
C105 a_741_n194# a_1987_n194# 0.01fF
C106 a_1275_n194# a_1097_n194# 0.10fF
C107 a_n683_n194# a_n149_n194# 0.02fF
C108 a_n1217_n194# a_n2107_n194# 0.01fF
C109 a_n3411_n140# a_n2699_n140# 0.03fF
C110 a_n2877_n140# a_n2165_n140# 0.03fF
C111 a_n3055_n140# a_n1987_n140# 0.02fF
C112 a_n2699_n140# a_n2343_n140# 0.06fF
C113 a_2165_n194# a_1453_n194# 0.01fF
C114 a_n1751_n194# a_n3353_n194# 0.01fF
C115 a_2165_n194# a_1809_n194# 0.03fF
C116 a_1275_n194# a_1987_n194# 0.01fF
C117 a_n327_n194# a_n1573_n194# 0.01fF
C118 a_n1751_n194# a_n2285_n194# 0.02fF
C119 a_n3233_n140# a_n3055_n140# 0.13fF
C120 a_n683_n194# a_n1039_n194# 0.03fF
C121 a_207_n194# a_919_n194# 0.01fF
C122 a_741_n194# a_207_n194# 0.02fF
C123 a_n1453_n140# a_n919_n140# 0.04fF
C124 a_n1275_n140# a_n1097_n140# 0.13fF
C125 a_n1631_n140# a_n741_n140# 0.02fF
C126 a_n1809_n140# a_n563_n140# 0.02fF
C127 a_1631_n194# a_3055_n194# 0.01fF
C128 a_n861_n194# a_385_n194# 0.01fF
C129 a_1453_n194# a_2521_n194# 0.01fF
C130 a_207_n194# a_n505_n194# 0.01fF
C131 a_1809_n194# a_2521_n194# 0.01fF
C132 a_n1395_n194# a_n2997_n194# 0.01fF
C133 a_n861_n194# a_n2285_n194# 0.01fF
C134 a_1453_n194# a_563_n194# 0.01fF
C135 a_207_n194# a_1275_n194# 0.01fF
C136 a_n1809_n140# a_n207_n140# 0.01fF
C137 a_n1929_n194# a_n1751_n194# 0.10fF
C138 a_1809_n194# a_563_n194# 0.01fF
C139 a_n1809_n140# a_n385_n140# 0.01fF
C140 a_2165_n194# a_2877_n194# 0.01fF
C141 a_n3411_n140# a_n2343_n140# 0.02fF
C142 a_n2877_n140# a_n1809_n140# 0.02fF
C143 a_n2699_n140# a_n1987_n140# 0.03fF
C144 a_n2521_n140# a_n2165_n140# 0.06fF
C145 a_n3055_n140# a_n1631_n140# 0.01fF
C146 a_n861_n194# a_n1929_n194# 0.01fF
C147 a_n149_n194# a_n1039_n194# 0.01fF
C148 a_n683_n194# a_n1395_n194# 0.01fF
C149 a_2343_n194# a_3411_n194# 0.01fF
C150 a_n1453_n140# a_149_n140# 0.01fF
C151 a_n3233_n140# a_n2699_n140# 0.04fF
C152 a_2877_n194# a_2521_n194# 0.03fF
C153 a_919_n194# a_29_n194# 0.01fF
C154 a_n1453_n140# a_n563_n140# 0.02fF
C155 a_n1097_n140# a_n919_n140# 0.13fF
C156 a_n1275_n140# a_n741_n140# 0.04fF
C157 a_741_n194# a_29_n194# 0.01fF
C158 a_1453_n194# a_2699_n194# 0.01fF
C159 a_n1453_n140# a_n29_n140# 0.01fF
C160 a_29_n194# a_n505_n194# 0.02fF
C161 a_n2641_n194# a_n1751_n194# 0.01fF
C162 a_n1751_n194# a_n1573_n194# 0.10fF
C163 a_1809_n194# a_2699_n194# 0.01fF
C164 a_n2285_n194# a_n3353_n194# 0.01fF
C165 a_n2997_n194# a_n3175_n194# 0.10fF
C166 a_n1453_n140# a_n207_n140# 0.02fF
C167 a_1631_n194# a_3233_n194# 0.01fF
C168 a_1275_n194# a_29_n194# 0.01fF
C169 a_2165_n194# a_919_n194# 0.01fF
C170 a_n1217_n194# a_n505_n194# 0.01fF
C171 a_741_n194# a_2165_n194# 0.01fF
C172 a_n861_n194# a_n1573_n194# 0.01fF
C173 a_n1097_n140# a_505_n140# 0.01fF
C174 a_n1453_n140# a_n385_n140# 0.02fF
C175 a_n2463_n194# a_n1751_n194# 0.01fF
C176 a_1631_n194# a_1097_n194# 0.02fF
C177 a_n3411_n140# a_n1987_n140# 0.01fF
C178 a_n1929_n194# a_n3353_n194# 0.01fF
C179 a_n1395_n194# a_n149_n194# 0.01fF
C180 a_n2699_n140# a_n1631_n140# 0.02fF
C181 a_n2877_n140# a_n1453_n140# 0.01fF
C182 a_n2521_n140# a_n1809_n140# 0.03fF
C183 a_n2343_n140# a_n1987_n140# 0.06fF
C184 a_3055_n194# a_3233_n194# 0.10fF
C185 a_n1097_n140# a_327_n140# 0.01fF
C186 a_2165_n194# a_1275_n194# 0.01fF
C187 a_n2997_n194# a_n2819_n194# 0.10fF
C188 a_919_n194# a_2521_n194# 0.01fF
C189 a_n683_n194# a_207_n194# 0.01fF
C190 a_n1929_n194# a_n2285_n194# 0.03fF
C191 a_n2463_n194# a_n861_n194# 0.01fF
C192 a_1631_n194# a_1987_n194# 0.03fF
C193 a_n149_n194# a_1097_n194# 0.01fF
C194 a_n3411_n140# a_n3233_n140# 0.13fF
C195 a_n1097_n140# a_149_n140# 0.02fF
C196 a_n3233_n140# a_n2343_n140# 0.02fF
C197 a_2877_n194# a_2699_n194# 0.10fF
C198 a_n1395_n194# a_n1039_n194# 0.03fF
C199 a_919_n194# a_563_n194# 0.03fF
C200 a_n919_n140# a_n741_n140# 0.13fF
C201 a_n1097_n140# a_n563_n140# 0.04fF
C202 a_741_n194# a_563_n194# 0.10fF
C203 a_n741_n140# a_861_n140# 0.01fF
C204 a_n3589_n140# a_n2877_n140# 0.03fF
C205 a_n1097_n140# a_n29_n140# 0.02fF
C206 a_n505_n194# a_563_n194# 0.01fF
C207 a_1987_n194# a_3055_n194# 0.01fF
C208 a_1275_n194# a_2521_n194# 0.01fF
C209 a_n1751_n194# a_n2107_n194# 0.03fF
C210 a_1631_n194# a_207_n194# 0.01fF
C211 a_n1097_n140# a_n207_n140# 0.02fF
C212 a_n741_n140# a_683_n140# 0.01fF
C213 a_1275_n194# a_563_n194# 0.01fF
C214 a_n2641_n194# a_n3353_n194# 0.01fF
C215 a_n741_n140# a_505_n140# 0.02fF
C216 a_n861_n194# a_n2107_n194# 0.01fF
C217 a_n1097_n140# a_n385_n140# 0.03fF
C218 a_n327_n194# a_919_n194# 0.01fF
C219 a_n3531_n194# a_n3353_n194# 0.10fF
C220 a_741_n194# a_n327_n194# 0.01fF
C221 a_207_n194# a_n149_n194# 0.03fF
C222 a_n2699_n140# a_n1275_n140# 0.01fF
C223 a_n2165_n140# a_n1809_n140# 0.06fF
C224 a_n2343_n140# a_n1631_n140# 0.03fF
C225 a_n2641_n194# a_n2285_n194# 0.03fF
C226 a_n2521_n140# a_n1453_n140# 0.02fF
C227 a_n2285_n194# a_n1573_n194# 0.01fF
C228 a_n327_n194# a_n505_n194# 0.10fF
C229 a_n741_n140# a_327_n140# 0.02fF
C230 a_n2463_n194# a_n3353_n194# 0.01fF
C231 a_2343_n194# a_1453_n194# 0.01fF
C232 a_n2285_n194# a_n3531_n194# 0.01fF
C233 a_n683_n194# a_29_n194# 0.01fF
C234 a_n741_n140# a_149_n140# 0.02fF
C235 a_n327_n194# a_1275_n194# 0.01fF
C236 a_n3233_n140# a_n1987_n140# 0.02fF
C237 a_2343_n194# a_1809_n194# 0.02fF
C238 a_3353_n140# a_3531_n140# 0.13fF
C239 a_207_n194# a_n1039_n194# 0.01fF
C240 a_n2463_n194# a_n2285_n194# 0.10fF
C241 a_n741_n140# a_n563_n140# 0.13fF
C242 a_n1929_n194# a_n2641_n194# 0.01fF
C243 a_n1929_n194# a_n1573_n194# 0.03fF
C244 a_n683_n194# a_n1217_n194# 0.02fF
C245 a_n3589_n140# a_n2521_n140# 0.02fF
C246 a_n741_n140# a_n29_n140# 0.03fF
C247 a_1275_n194# a_2699_n194# 0.01fF
C248 a_3175_n140# a_3531_n140# 0.06fF
C249 a_n1929_n194# a_n3531_n194# 0.01fF
C250 a_n741_n140# a_n207_n140# 0.04fF
C251 a_1631_n194# a_29_n194# 0.01fF
C252 a_3175_n140# a_3353_n140# 0.13fF
C253 a_2997_n140# a_3531_n140# 0.04fF
C254 a_385_n194# a_1453_n194# 0.01fF
C255 a_n2463_n194# a_n1929_n194# 0.02fF
C256 a_1987_n194# a_3233_n194# 0.01fF
C257 a_n3353_n194# a_n2107_n194# 0.01fF
C258 a_n741_n140# a_n385_n140# 0.06fF
C259 a_1809_n194# a_385_n194# 0.01fF
C260 a_2997_n140# a_3353_n140# 0.06fF
C261 a_2819_n140# a_3531_n140# 0.03fF
C262 a_n1987_n140# a_n1631_n140# 0.06fF
C263 a_n2521_n140# a_n1097_n140# 0.01fF
C264 a_n2343_n140# a_n1275_n140# 0.02fF
C265 a_n2165_n140# a_n1453_n140# 0.03fF
C266 a_1987_n194# a_1097_n194# 0.01fF
C267 a_n2285_n194# a_n2107_n194# 0.10fF
C268 a_n149_n194# a_29_n194# 0.10fF
C269 a_2343_n194# a_2877_n194# 0.02fF
C270 a_1631_n194# a_2165_n194# 0.02fF
C271 a_2997_n140# a_3175_n140# 0.13fF
C272 a_2641_n140# a_3531_n140# 0.02fF
C273 a_2819_n140# a_3353_n140# 0.04fF
C274 a_n1395_n194# a_207_n194# 0.01fF
C275 a_n683_n194# a_563_n194# 0.01fF
C276 a_n2641_n194# a_n1573_n194# 0.01fF
C277 a_n3233_n140# a_n1631_n140# 0.01fF
C278 a_n1217_n194# a_n149_n194# 0.01fF
C279 a_1809_n194# a_3411_n194# 0.01fF
C280 a_2819_n140# a_3175_n140# 0.06fF
C281 a_2641_n140# a_3353_n140# 0.03fF
C282 a_2463_n140# a_3531_n140# 0.02fF
C283 a_n1751_n194# a_n505_n194# 0.01fF
C284 a_n2641_n194# a_n3531_n194# 0.01fF
C285 a_29_n194# a_n1039_n194# 0.01fF
C286 a_2165_n194# a_3055_n194# 0.01fF
C287 a_n1929_n194# a_n2107_n194# 0.10fF
C288 a_207_n194# a_1097_n194# 0.01fF
C289 a_n3589_n140# a_n2165_n140# 0.01fF
C290 a_1631_n194# a_2521_n194# 0.01fF
C291 a_2463_n140# a_3353_n140# 0.02fF
C292 a_2285_n140# a_3531_n140# 0.02fF
C293 a_2641_n140# a_3175_n140# 0.04fF
C294 a_2819_n140# a_2997_n140# 0.13fF
C295 a_n861_n194# a_741_n194# 0.01fF
C296 a_n2463_n194# a_n2641_n194# 0.10fF
C297 a_n3055_n140# a_n2877_n140# 0.13fF
C298 a_n2463_n194# a_n1573_n194# 0.01fF
C299 a_n1217_n194# a_n1039_n194# 0.10fF
C300 a_n861_n194# a_n505_n194# 0.03fF
C301 a_1631_n194# a_563_n194# 0.01fF
C302 a_2285_n140# a_3353_n140# 0.02fF
C303 a_2641_n140# a_2997_n140# 0.06fF
C304 a_2107_n140# a_3531_n140# 0.01fF
C305 a_2463_n140# a_3175_n140# 0.03fF
C306 a_n683_n194# a_n327_n194# 0.03fF
C307 a_n2463_n194# a_n3531_n194# 0.01fF
C308 a_n1395_n194# a_n2819_n194# 0.01fF
C309 a_3055_n194# a_2521_n194# 0.02fF
C310 a_2343_n194# a_919_n194# 0.01fF
C311 a_2107_n140# a_3353_n140# 0.02fF
C312 a_2641_n140# a_2819_n140# 0.13fF
C313 a_2343_n194# a_741_n194# 0.01fF
C314 a_2463_n140# a_2997_n140# 0.04fF
C315 a_2285_n140# a_3175_n140# 0.02fF
C316 a_1929_n140# a_3531_n140# 0.01fF
C317 a_n2343_n140# a_n919_n140# 0.01fF
C318 a_n2165_n140# a_n1097_n140# 0.02fF
C319 a_n1987_n140# a_n1275_n140# 0.03fF
C320 a_n1809_n140# a_n1453_n140# 0.06fF
C321 a_n149_n194# a_563_n194# 0.01fF
C322 a_3411_n194# a_2877_n194# 0.02fF
C323 a_1929_n140# a_3353_n140# 0.01fF
C324 a_2463_n140# a_2819_n140# 0.06fF
C325 a_2285_n140# a_2997_n140# 0.03fF
C326 a_2107_n140# a_3175_n140# 0.02fF
C327 a_2343_n194# a_1275_n194# 0.01fF
C328 a_n1395_n194# a_29_n194# 0.01fF
C329 a_n2641_n194# a_n2107_n194# 0.02fF
C330 a_n1573_n194# a_n2107_n194# 0.02fF
C331 a_2285_n140# a_2819_n140# 0.04fF
C332 a_2107_n140# a_2997_n140# 0.02fF
C333 a_2463_n140# a_2641_n140# 0.13fF
C334 a_1751_n140# a_3353_n140# 0.01fF
C335 a_1929_n140# a_3175_n140# 0.02fF
C336 a_563_n194# a_n1039_n194# 0.01fF
C337 a_n3531_n194# a_n2107_n194# 0.01fF
C338 a_n1751_n194# a_n2997_n194# 0.01fF
C339 a_1631_n194# a_2699_n194# 0.01fF
C340 a_385_n194# a_919_n194# 0.02fF
C341 a_29_n194# a_1097_n194# 0.01fF
C342 a_n1395_n194# a_n1217_n194# 0.10fF
C343 a_2285_n140# a_2641_n140# 0.06fF
C344 a_1929_n140# a_2997_n140# 0.02fF
C345 a_1751_n140# a_3175_n140# 0.01fF
C346 a_2107_n140# a_2819_n140# 0.03fF
C347 a_741_n194# a_385_n194# 0.03fF
C348 a_n327_n194# a_n149_n194# 0.10fF
C349 a_n2877_n140# a_n2699_n140# 0.13fF
C350 a_n3055_n140# a_n2521_n140# 0.04fF
C351 a_n2463_n194# a_n2107_n194# 0.03fF
C352 a_385_n194# a_n505_n194# 0.01fF
C353 a_2165_n194# a_3233_n194# 0.01fF
C354 a_1573_n140# a_3175_n140# 0.01fF
C355 a_1929_n140# a_2819_n140# 0.02fF
C356 a_2285_n140# a_2463_n140# 0.13fF
C357 a_2107_n140# a_2641_n140# 0.04fF
C358 a_1751_n140# a_2997_n140# 0.02fF
C359 a_3055_n194# a_2699_n194# 0.03fF
C360 a_n3175_n194# a_n2819_n194# 0.03fF
C361 a_385_n194# a_1275_n194# 0.01fF
C362 a_2165_n194# a_1097_n194# 0.01fF
C363 a_2107_n140# a_2463_n140# 0.06fF
C364 a_1751_n140# a_2819_n140# 0.02fF
C365 a_1573_n140# a_2997_n140# 0.01fF
C366 a_1929_n140# a_2641_n140# 0.03fF
C367 a_n327_n194# a_n1039_n194# 0.01fF
C368 a_n1631_n140# a_n1275_n140# 0.06fF
C369 a_n1809_n140# a_n1097_n140# 0.03fF
C370 a_n2165_n140# a_n741_n140# 0.01fF
C371 a_n1987_n140# a_n919_n140# 0.02fF
C372 a_n683_n194# a_n1751_n194# 0.01fF
C373 a_3233_n194# a_2521_n194# 0.01fF
C374 a_1929_n140# a_2463_n140# 0.04fF
C375 a_1751_n140# a_2641_n140# 0.02fF
C376 a_1395_n140# a_2997_n140# 0.01fF
C377 a_2107_n140# a_2285_n140# 0.13fF
C378 a_1573_n140# a_2819_n140# 0.02fF
C379 a_2165_n194# a_1987_n194# 0.10fF
C380 a_n1929_n194# a_n505_n194# 0.01fF
C381 a_207_n194# a_29_n194# 0.10fF
C382 a_1809_n194# a_1453_n194# 0.03fF
C383 a_1097_n194# a_2521_n194# 0.01fF
C384 a_1929_n140# a_2285_n140# 0.06fF
C385 a_1395_n140# a_2819_n140# 0.01fF
C386 a_1751_n140# a_2463_n140# 0.03fF
C387 a_1573_n140# a_2641_n140# 0.02fF
C388 a_n861_n194# a_n683_n194# 0.10fF
C389 a_1097_n194# a_563_n194# 0.02fF
C390 a_207_n194# a_n1217_n194# 0.01fF
C391 a_1929_n140# a_2107_n140# 0.13fF
C392 a_1751_n140# a_2285_n140# 0.04fF
C393 a_1573_n140# a_2463_n140# 0.02fF
C394 a_1395_n140# a_2641_n140# 0.02fF
C395 a_1217_n140# a_2819_n140# 0.01fF
C396 a_n3411_n140# a_n2877_n140# 0.04fF
C397 a_n2877_n140# a_n2343_n140# 0.04fF
C398 a_n2699_n140# a_n2521_n140# 0.13fF
C399 a_1987_n194# a_2521_n194# 0.02fF
C400 a_n3055_n140# a_n2165_n140# 0.02fF
C401 a_1395_n140# a_2463_n140# 0.02fF
C402 a_n3353_n194# a_n2997_n194# 0.03fF
C403 a_1751_n140# a_2107_n140# 0.06fF
C404 a_1573_n140# a_2285_n140# 0.03fF
C405 a_1217_n140# a_2641_n140# 0.01fF
C406 a_n1395_n194# a_n327_n194# 0.01fF
C407 a_1987_n194# a_563_n194# 0.01fF
C408 a_n1751_n194# a_n149_n194# 0.01fF
C409 a_1573_n140# a_2107_n140# 0.04fF
C410 a_1217_n140# a_2463_n140# 0.02fF
C411 a_1039_n140# a_2641_n140# 0.01fF
C412 a_1395_n140# a_2285_n140# 0.02fF
C413 a_1751_n140# a_1929_n140# 0.13fF
C414 a_n2285_n194# a_n2997_n194# 0.01fF
C415 a_n1809_n140# a_n741_n140# 0.02fF
C416 a_n1631_n140# a_n919_n140# 0.03fF
C417 a_n1453_n140# a_n1097_n140# 0.06fF
C418 a_n1987_n140# a_n563_n140# 0.01fF
C419 a_1453_n194# a_2877_n194# 0.01fF
C420 a_n327_n194# a_1097_n194# 0.01fF
C421 a_n1217_n194# a_n2819_n194# 0.01fF
C422 a_n1573_n194# a_n505_n194# 0.01fF
C423 a_3233_n194# a_2699_n194# 0.02fF
C424 a_1395_n140# a_2107_n140# 0.03fF
C425 a_1573_n140# a_1929_n140# 0.06fF
C426 a_1039_n140# a_2463_n140# 0.01fF
C427 a_1217_n140# a_2285_n140# 0.02fF
C428 a_1809_n194# a_2877_n194# 0.01fF
C429 a_n861_n194# a_n149_n194# 0.01fF
C430 a_1631_n194# a_2343_n194# 0.01fF
C431 a_n1751_n194# a_n1039_n194# 0.01fF
C432 a_207_n194# a_563_n194# 0.03fF
C433 a_1097_n194# a_2699_n194# 0.01fF
C434 a_1039_n140# a_2285_n140# 0.02fF
C435 a_1217_n140# a_2107_n140# 0.02fF
C436 a_1573_n140# a_1751_n140# 0.13fF
C437 a_861_n140# a_2463_n140# 0.01fF
C438 a_1395_n140# a_1929_n140# 0.04fF
C439 a_n683_n194# a_385_n194# 0.01fF
C440 a_n1929_n194# a_n2997_n194# 0.01fF
C441 a_n1987_n140# a_n385_n140# 0.01fF
C442 a_n683_n194# a_n2285_n194# 0.01fF
C443 a_2343_n194# a_3055_n194# 0.01fF
C444 a_n861_n194# a_n1039_n194# 0.10fF
C445 a_1217_n140# a_1929_n140# 0.03fF
C446 a_861_n140# a_2285_n140# 0.01fF
C447 a_1395_n140# a_1751_n140# 0.06fF
C448 a_n1217_n194# a_29_n194# 0.01fF
C449 a_1039_n140# a_2107_n140# 0.02fF
C450 a_n3411_n140# a_n2521_n140# 0.02fF
C451 a_n2877_n140# a_n1987_n140# 0.02fF
C452 a_n3055_n140# a_n1809_n140# 0.02fF
C453 a_1987_n194# a_2699_n194# 0.01fF
C454 a_n2699_n140# a_n2165_n140# 0.04fF
C455 a_n2521_n140# a_n2343_n140# 0.13fF
C456 a_1395_n140# a_1573_n140# 0.13fF
C457 a_683_n140# a_2285_n140# 0.01fF
C458 a_1039_n140# a_1929_n140# 0.02fF
C459 a_861_n140# a_2107_n140# 0.02fF
C460 a_1217_n140# a_1751_n140# 0.04fF
C461 a_207_n194# a_n327_n194# 0.02fF
C462 a_1631_n194# a_385_n194# 0.01fF
C463 a_919_n194# a_1453_n194# 0.02fF
C464 a_n3233_n140# a_n2877_n140# 0.06fF
C465 a_741_n194# a_1453_n194# 0.01fF
C466 a_n1929_n194# a_n683_n194# 0.01fF
C467 a_1039_n140# a_1751_n140# 0.03fF
C468 a_1217_n140# a_1573_n140# 0.06fF
C469 a_861_n140# a_1929_n140# 0.02fF
C470 a_683_n140# a_2107_n140# 0.01fF
C471 a_n1453_n140# a_n741_n140# 0.03fF
C472 a_n1631_n140# a_n563_n140# 0.02fF
C473 a_n1275_n140# a_n919_n140# 0.06fF
C474 a_1809_n194# a_919_n194# 0.01fF
C475 a_741_n194# a_1809_n194# 0.01fF
C476 a_n1631_n140# a_n29_n140# 0.01fF
C477 a_n1395_n194# a_n1751_n194# 0.03fF
C478 a_n2107_n194# a_n505_n194# 0.01fF
C479 a_1039_n140# a_1573_n140# 0.04fF
C480 a_1217_n140# a_1395_n140# 0.13fF
C481 a_861_n140# a_1751_n140# 0.02fF
C482 a_683_n140# a_1929_n140# 0.02fF
C483 a_505_n140# a_2107_n140# 0.01fF
C484 a_n2641_n194# a_n2997_n194# 0.03fF
C485 a_385_n194# a_n149_n194# 0.02fF
C486 a_n2997_n194# a_n1573_n194# 0.01fF
C487 a_1453_n194# a_1275_n194# 0.10fF
C488 a_n1631_n140# a_n207_n140# 0.01fF
C489 a_29_n194# a_563_n194# 0.02fF
C490 a_n3531_n194# a_n2997_n194# 0.02fF
C491 a_861_n140# a_1573_n140# 0.03fF
C492 a_683_n140# a_1751_n140# 0.02fF
C493 a_505_n140# a_1929_n140# 0.01fF
C494 a_1039_n140# a_1395_n140# 0.06fF
C495 a_1809_n194# a_1275_n194# 0.02fF
C496 a_n861_n194# a_n1395_n194# 0.02fF
C497 a_n1631_n140# a_n385_n140# 0.02fF
C498 a_2165_n194# a_2521_n194# 0.03fF
C499 a_327_n140# a_1929_n140# 0.01fF
C500 a_683_n140# a_1573_n140# 0.02fF
C501 a_1039_n140# a_1217_n140# 0.13fF
C502 a_505_n140# a_1751_n140# 0.02fF
C503 a_385_n194# a_n1039_n194# 0.01fF
C504 a_n2463_n194# a_n2997_n194# 0.02fF
C505 a_861_n140# a_1395_n140# 0.04fF
C506 a_3411_n194# a_3055_n194# 0.03fF
C507 a_n3411_n140# a_n2165_n140# 0.02fF
C508 a_n3055_n140# a_n1453_n140# 0.01fF
C509 a_n2699_n140# a_n1809_n140# 0.02fF
C510 a_n2521_n140# a_n1987_n140# 0.04fF
C511 a_n2343_n140# a_n2165_n140# 0.13fF
C512 a_n2877_n140# a_n1631_n140# 0.02fF
C513 a_n1275_n140# a_327_n140# 0.01fF
C514 a_2165_n194# a_563_n194# 0.01fF
C515 a_n2285_n194# a_n1039_n194# 0.01fF
C516 a_861_n140# a_1217_n140# 0.06fF
C517 a_327_n140# a_1751_n140# 0.01fF
C518 a_683_n140# a_1395_n140# 0.03fF
C519 a_505_n140# a_1573_n140# 0.02fF
C520 a_n683_n194# a_n1573_n194# 0.01fF
C521 a_2343_n194# a_3233_n194# 0.01fF
C522 a_n327_n194# a_29_n194# 0.03fF
C523 a_n1275_n140# a_149_n140# 0.01fF
C524 a_n3233_n140# a_n2521_n140# 0.03fF
C525 a_683_n140# a_1217_n140# 0.04fF
C526 a_149_n140# a_1751_n140# 0.01fF
C527 a_327_n140# a_1573_n140# 0.02fF
C528 a_861_n140# a_1039_n140# 0.13fF
C529 a_505_n140# a_1395_n140# 0.02fF
C530 a_n1275_n140# a_n563_n140# 0.03fF
C531 a_n1097_n140# a_n741_n140# 0.06fF
C532 a_2343_n194# a_1097_n194# 0.01fF
C533 a_n1275_n140# a_n29_n140# 0.02fF
C534 a_n3589_n140# a_n3055_n140# 0.04fF
C535 a_n1217_n194# a_n327_n194# 0.01fF
C536 a_1275_n194# a_2877_n194# 0.01fF
C537 a_n1929_n194# a_n1039_n194# 0.01fF
C538 a_327_n140# a_1395_n140# 0.02fF
C539 a_n1751_n194# a_n3175_n194# 0.01fF
C540 a_505_n140# a_1217_n140# 0.03fF
C541 a_683_n140# a_1039_n140# 0.06fF
C542 a_149_n140# a_1573_n140# 0.01fF
C543 a_n2997_n194# a_n2107_n194# 0.01fF
C544 a_n1275_n140# a_n207_n140# 0.02fF
C545 a_n919_n140# a_683_n140# 0.01fF
C546 a_2343_n194# a_1987_n194# 0.03fF
C547 a_n29_n140# a_1573_n140# 0.01fF
C548 a_327_n140# a_1217_n140# 0.02fF
C549 a_505_n140# a_1039_n140# 0.04fF
C550 a_149_n140# a_1395_n140# 0.02fF
C551 a_683_n140# a_861_n140# 0.13fF
C552 a_n861_n194# a_207_n194# 0.01fF
C553 a_n919_n140# a_505_n140# 0.01fF
C554 a_n1275_n140# a_n385_n140# 0.02fF
C555 a_2165_n194# a_2699_n194# 0.02fF
C556 a_n29_n140# a_1395_n140# 0.01fF
C557 a_505_n140# a_861_n140# 0.06fF
C558 a_327_n140# a_1039_n140# 0.03fF
C559 a_149_n140# a_1217_n140# 0.02fF
C560 a_n3411_n140# a_n1809_n140# 0.01fF
C561 a_n2877_n140# a_n1275_n140# 0.01fF
C562 a_n1395_n194# a_n2285_n194# 0.01fF
C563 a_n2165_n140# a_n1987_n140# 0.13fF
C564 a_n2521_n140# a_n1631_n140# 0.02fF
C565 a_n2343_n140# a_n1809_n140# 0.04fF
C566 a_n2699_n140# a_n1453_n140# 0.02fF
C567 a_741_n194# a_919_n194# 0.10fF
C568 a_n149_n194# a_n1573_n194# 0.01fF
C569 a_n1751_n194# a_n2819_n194# 0.01fF
C570 a_385_n194# a_1097_n194# 0.01fF
C571 a_n919_n140# a_327_n140# 0.02fF
C572 a_919_n194# a_n505_n194# 0.01fF
C573 a_n207_n140# a_1395_n140# 0.01fF
C574 a_149_n140# a_1039_n140# 0.02fF
C575 a_n29_n140# a_1217_n140# 0.02fF
C576 a_505_n140# a_683_n140# 0.13fF
C577 a_327_n140# a_861_n140# 0.04fF
C578 a_n683_n194# a_n2107_n194# 0.01fF
C579 a_741_n194# a_n505_n194# 0.01fF
C580 a_n327_n194# a_563_n194# 0.01fF
C581 a_n919_n140# a_149_n140# 0.02fF
C582 a_n563_n140# a_1039_n140# 0.01fF
C583 a_3411_n194# a_3233_n194# 0.10fF
C584 a_n3233_n140# a_n2165_n140# 0.02fF
C585 a_2521_n194# a_2699_n194# 0.10fF
C586 a_149_n140# a_861_n140# 0.03fF
C587 a_n207_n140# a_1217_n140# 0.01fF
C588 a_327_n140# a_683_n140# 0.06fF
C589 a_n2641_n194# a_n1039_n194# 0.01fF
C590 a_n29_n140# a_1039_n140# 0.02fF
C591 a_385_n194# a_1987_n194# 0.01fF
C592 a_919_n194# a_1275_n194# 0.03fF
C593 a_n919_n140# a_n563_n140# 0.06fF
C594 a_n1929_n194# a_n1395_n194# 0.02fF
C595 a_n1573_n194# a_n1039_n194# 0.02fF
C596 a_741_n194# a_1275_n194# 0.02fF
C597 a_n563_n140# a_861_n140# 0.01fF
C598 a_n3589_n140# a_n2699_n140# 0.02fF
C599 a_n919_n140# a_n29_n140# 0.02fF
C600 a_n207_n140# a_1039_n140# 0.02fF
C601 a_n385_n140# a_1217_n140# 0.01fF
C602 a_149_n140# a_683_n140# 0.04fF
C603 a_327_n140# a_505_n140# 0.13fF
C604 a_n29_n140# a_861_n140# 0.02fF
C605 a_1631_n194# a_1453_n194# 0.10fF
C606 a_n919_n140# a_n207_n140# 0.03fF
C607 a_n563_n140# a_683_n140# 0.02fF
C608 a_n2463_n194# a_n1039_n194# 0.01fF
C609 a_n29_n140# a_683_n140# 0.03fF
C610 a_n207_n140# a_861_n140# 0.02fF
C611 a_149_n140# a_505_n140# 0.06fF
C612 a_n385_n140# a_1039_n140# 0.01fF
C613 a_1631_n194# a_1809_n194# 0.10fF
C614 a_3411_n194# a_1987_n194# 0.01fF
C615 a_207_n194# a_385_n194# 0.10fF
C616 a_n1217_n194# a_n1751_n194# 0.02fF
C617 a_n3353_n194# a_n3175_n194# 0.10fF
C618 a_n563_n140# a_505_n140# 0.02fF
C619 a_n861_n194# a_29_n194# 0.01fF
C620 a_n919_n140# a_n385_n140# 0.04fF
C621 a_1453_n194# a_3055_n194# 0.01fF
C622 a_n207_n140# a_683_n140# 0.02fF
C623 a_n149_n194# a_1453_n194# 0.01fF
C624 a_149_n140# a_327_n140# 0.13fF
C625 a_n385_n140# a_861_n140# 0.02fF
C626 a_n29_n140# a_505_n140# 0.04fF
C627 a_n2343_n140# a_n1453_n140# 0.02fF
C628 a_n2165_n140# a_n1631_n140# 0.04fF
C629 a_n2699_n140# a_n1097_n140# 0.01fF
C630 a_n1987_n140# a_n1809_n140# 0.13fF
C631 a_n2521_n140# a_n1275_n140# 0.02fF
C632 a_n2285_n194# a_n3175_n194# 0.01fF
C633 a_n563_n140# a_327_n140# 0.02fF
C634 a_1809_n194# a_3055_n194# 0.01fF
C635 a_n861_n194# a_n1217_n194# 0.03fF
C636 a_n207_n140# a_505_n140# 0.03fF
C637 a_n29_n140# a_327_n140# 0.06fF
C638 a_n385_n140# a_683_n140# 0.02fF
C639 a_3531_n140# VSUBS 0.02fF
C640 a_3353_n140# VSUBS 0.02fF
C641 a_3175_n140# VSUBS 0.02fF
C642 a_2997_n140# VSUBS 0.02fF
C643 a_2819_n140# VSUBS 0.02fF
C644 a_2641_n140# VSUBS 0.02fF
C645 a_2463_n140# VSUBS 0.02fF
C646 a_2285_n140# VSUBS 0.02fF
C647 a_2107_n140# VSUBS 0.02fF
C648 a_1929_n140# VSUBS 0.02fF
C649 a_1751_n140# VSUBS 0.02fF
C650 a_1573_n140# VSUBS 0.02fF
C651 a_1395_n140# VSUBS 0.02fF
C652 a_1217_n140# VSUBS 0.02fF
C653 a_1039_n140# VSUBS 0.02fF
C654 a_861_n140# VSUBS 0.02fF
C655 a_683_n140# VSUBS 0.02fF
C656 a_505_n140# VSUBS 0.02fF
C657 a_327_n140# VSUBS 0.02fF
C658 a_149_n140# VSUBS 0.02fF
C659 a_n29_n140# VSUBS 0.02fF
C660 a_n207_n140# VSUBS 0.02fF
C661 a_n385_n140# VSUBS 0.02fF
C662 a_n563_n140# VSUBS 0.02fF
C663 a_n741_n140# VSUBS 0.02fF
C664 a_n919_n140# VSUBS 0.02fF
C665 a_n1097_n140# VSUBS 0.02fF
C666 a_n1275_n140# VSUBS 0.02fF
C667 a_n1453_n140# VSUBS 0.02fF
C668 a_n1631_n140# VSUBS 0.02fF
C669 a_n1809_n140# VSUBS 0.02fF
C670 a_n1987_n140# VSUBS 0.02fF
C671 a_n2165_n140# VSUBS 0.02fF
C672 a_n2343_n140# VSUBS 0.02fF
C673 a_n2521_n140# VSUBS 0.02fF
C674 a_n2699_n140# VSUBS 0.02fF
C675 a_n2877_n140# VSUBS 0.02fF
C676 a_n3055_n140# VSUBS 0.02fF
C677 a_n3233_n140# VSUBS 0.02fF
C678 a_n3411_n140# VSUBS 0.02fF
C679 a_n3589_n140# VSUBS 0.02fF
C680 a_3411_n194# VSUBS 0.29fF
C681 a_3233_n194# VSUBS 0.23fF
C682 a_3055_n194# VSUBS 0.24fF
C683 a_2877_n194# VSUBS 0.25fF
C684 a_2699_n194# VSUBS 0.26fF
C685 a_2521_n194# VSUBS 0.27fF
C686 a_2343_n194# VSUBS 0.28fF
C687 a_2165_n194# VSUBS 0.28fF
C688 a_1987_n194# VSUBS 0.29fF
C689 a_1809_n194# VSUBS 0.29fF
C690 a_1631_n194# VSUBS 0.29fF
C691 a_1453_n194# VSUBS 0.29fF
C692 a_1275_n194# VSUBS 0.29fF
C693 a_1097_n194# VSUBS 0.29fF
C694 a_919_n194# VSUBS 0.29fF
C695 a_741_n194# VSUBS 0.29fF
C696 a_563_n194# VSUBS 0.29fF
C697 a_385_n194# VSUBS 0.29fF
C698 a_207_n194# VSUBS 0.29fF
C699 a_29_n194# VSUBS 0.29fF
C700 a_n149_n194# VSUBS 0.29fF
C701 a_n327_n194# VSUBS 0.29fF
C702 a_n505_n194# VSUBS 0.29fF
C703 a_n683_n194# VSUBS 0.29fF
C704 a_n861_n194# VSUBS 0.29fF
C705 a_n1039_n194# VSUBS 0.29fF
C706 a_n1217_n194# VSUBS 0.29fF
C707 a_n1395_n194# VSUBS 0.29fF
C708 a_n1573_n194# VSUBS 0.29fF
C709 a_n1751_n194# VSUBS 0.29fF
C710 a_n1929_n194# VSUBS 0.29fF
C711 a_n2107_n194# VSUBS 0.29fF
C712 a_n2285_n194# VSUBS 0.29fF
C713 a_n2463_n194# VSUBS 0.29fF
C714 a_n2641_n194# VSUBS 0.29fF
C715 a_n2819_n194# VSUBS 0.29fF
C716 a_n2997_n194# VSUBS 0.29fF
C717 a_n3175_n194# VSUBS 0.29fF
C718 a_n3353_n194# VSUBS 0.29fF
C719 a_n3531_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CC a_n1008_n140# a_2374_n140# a_1306_n140# a_n652_n140#
+ a_652_n194# a_n1662_n194# a_772_n140# a_n2730_n194# a_n1720_n140# a_n60_n194# a_2076_n194#
+ a_1008_n194# a_2196_n140# a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194#
+ a_n2552_n194# a_594_n140# a_n1542_n140# a_n2610_n140# a_1720_n194# a_1840_n140#
+ a_n238_n194# a_n2908_n194# a_3086_n140# a_n296_n140# a_n1898_n140# a_n2966_n140#
+ a_296_n194# a_2018_n140# a_60_n140# a_n1306_n194# a_n2374_n194# a_n1364_n140# a_1542_n194#
+ a_416_n140# a_n2432_n140# a_2610_n194# a_n950_n194# a_1662_n140# a_2730_n140# a_2966_n194#
+ a_1898_n194# a_n2788_n140# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194#
+ a_238_n140# a_n1186_n140# a_n2254_n140# a_2432_n194# a_1364_n194# a_n772_n194# a_2552_n140#
+ a_1484_n140# a_n830_n140# a_2788_n194# a_830_n194# a_n1840_n194# a_950_n140# a_n3086_n194#
+ a_2908_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_n3144_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2374_n140# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2788_n140# a_n2908_n194# a_n2966_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n2432_n140# a_n2552_n194# a_n2610_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2966_n140# a_n3086_n194# a_n3144_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_2730_n140# a_2610_n194# a_2552_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n2610_n140# a_n2730_n194# a_n2788_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n2254_n140# a_n2374_n194# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_3086_n140# a_2966_n194# a_2908_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_2552_n140# a_2432_n194# a_2374_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_2908_n140# a_2788_n194# a_2730_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_1186_n194# a_2432_n194# 0.01fF
C1 a_60_n140# a_1662_n140# 0.01fF
C2 a_1186_n194# a_1364_n194# 0.10fF
C3 a_772_n140# a_2374_n140# 0.01fF
C4 a_n474_n140# a_60_n140# 0.04fF
C5 a_n1720_n140# a_n118_n140# 0.01fF
C6 a_n1364_n140# a_n1898_n140# 0.04fF
C7 a_416_n140# a_238_n140# 0.13fF
C8 a_1898_n194# a_830_n194# 0.01fF
C9 a_n652_n140# a_n1542_n140# 0.02fF
C10 a_1720_n194# a_2966_n194# 0.01fF
C11 a_n652_n140# a_416_n140# 0.02fF
C12 a_2076_n194# a_2610_n194# 0.02fF
C13 a_2254_n194# a_1186_n194# 0.01fF
C14 a_950_n140# a_2018_n140# 0.02fF
C15 a_n2432_n140# a_n2610_n140# 0.13fF
C16 a_n3144_n140# a_n1542_n140# 0.01fF
C17 a_594_n140# a_1484_n140# 0.02fF
C18 a_1662_n140# a_3086_n140# 0.01fF
C19 a_1840_n140# a_2908_n140# 0.02fF
C20 a_n1364_n140# a_n1186_n140# 0.13fF
C21 a_474_n194# a_n1128_n194# 0.01fF
C22 a_n594_n194# a_n238_n194# 0.03fF
C23 a_652_n194# a_n772_n194# 0.01fF
C24 a_n950_n194# a_474_n194# 0.01fF
C25 a_1306_n140# a_1484_n140# 0.13fF
C26 a_1128_n140# a_1662_n140# 0.04fF
C27 a_1720_n194# a_2610_n194# 0.01fF
C28 a_n2374_n194# a_n2908_n194# 0.02fF
C29 a_474_n194# a_296_n194# 0.10fF
C30 a_n474_n140# a_1128_n140# 0.01fF
C31 a_n2432_n140# a_n1720_n140# 0.03fF
C32 a_n1840_n194# a_n2908_n194# 0.01fF
C33 a_60_n140# a_1128_n140# 0.02fF
C34 a_n830_n140# a_n1542_n140# 0.03fF
C35 a_n2788_n140# a_n1364_n140# 0.01fF
C36 a_118_n194# a_1542_n194# 0.01fF
C37 a_1008_n194# a_n594_n194# 0.01fF
C38 a_n830_n140# a_416_n140# 0.02fF
C39 a_772_n140# a_1840_n140# 0.02fF
C40 a_n1008_n140# a_n2254_n140# 0.02fF
C41 a_n2610_n140# a_n3144_n140# 0.04fF
C42 a_2432_n194# a_2966_n194# 0.02fF
C43 a_1186_n194# a_1898_n194# 0.01fF
C44 a_1008_n194# a_2076_n194# 0.01fF
C45 a_n1128_n194# a_n2374_n194# 0.01fF
C46 a_1364_n194# a_2966_n194# 0.01fF
C47 a_n1840_n194# a_n1128_n194# 0.01fF
C48 a_n474_n140# a_n118_n140# 0.06fF
C49 a_n950_n194# a_n2374_n194# 0.01fF
C50 a_60_n140# a_n118_n140# 0.13fF
C51 a_n2076_n140# a_n1898_n140# 0.13fF
C52 a_n1840_n194# a_n950_n194# 0.01fF
C53 a_950_n140# a_1484_n140# 0.04fF
C54 a_652_n194# a_118_n194# 0.02fF
C55 a_n652_n140# a_n1720_n140# 0.02fF
C56 a_n1662_n194# a_n1306_n194# 0.03fF
C57 a_n2018_n194# a_n1306_n194# 0.01fF
C58 a_n1662_n194# a_n2730_n194# 0.01fF
C59 a_1306_n140# a_2908_n140# 0.01fF
C60 a_n3144_n140# a_n1720_n140# 0.01fF
C61 a_2254_n194# a_2966_n194# 0.01fF
C62 a_594_n140# a_772_n140# 0.13fF
C63 a_n1484_n194# a_n2374_n194# 0.01fF
C64 a_n1128_n194# a_n60_n194# 0.01fF
C65 a_n1840_n194# a_n1484_n194# 0.03fF
C66 a_1720_n194# a_1008_n194# 0.01fF
C67 a_n2018_n194# a_n2730_n194# 0.01fF
C68 a_n1662_n194# a_n2196_n194# 0.02fF
C69 a_n296_n140# a_n1542_n140# 0.02fF
C70 a_n950_n194# a_n60_n194# 0.01fF
C71 a_2432_n194# a_2610_n194# 0.10fF
C72 a_n296_n140# a_416_n140# 0.03fF
C73 a_1364_n194# a_2610_n194# 0.01fF
C74 a_n60_n194# a_296_n194# 0.03fF
C75 a_n1186_n140# a_n2076_n140# 0.02fF
C76 a_n594_n194# a_n772_n194# 0.10fF
C77 a_n2018_n194# a_n2196_n194# 0.10fF
C78 a_2552_n140# a_2730_n140# 0.13fF
C79 a_772_n140# a_1306_n140# 0.04fF
C80 a_n2552_n194# a_n3086_n194# 0.02fF
C81 a_n118_n140# a_1128_n140# 0.02fF
C82 a_n830_n140# a_n1720_n140# 0.02fF
C83 a_n60_n194# a_n1484_n194# 0.01fF
C84 a_n2788_n140# a_n2076_n140# 0.03fF
C85 a_n1364_n140# a_n1008_n140# 0.06fF
C86 a_2254_n194# a_2610_n194# 0.03fF
C87 a_n416_n194# a_n1662_n194# 0.01fF
C88 a_296_n194# a_830_n194# 0.02fF
C89 a_n2966_n140# a_n1542_n140# 0.01fF
C90 a_238_n140# a_1662_n140# 0.01fF
C91 a_n2018_n194# a_n416_n194# 0.01fF
C92 a_1364_n194# a_n238_n194# 0.01fF
C93 a_2966_n194# a_1898_n194# 0.01fF
C94 a_n474_n140# a_238_n140# 0.03fF
C95 a_60_n140# a_238_n140# 0.13fF
C96 a_118_n194# a_n594_n194# 0.01fF
C97 a_n652_n140# a_n474_n140# 0.13fF
C98 a_772_n140# a_950_n140# 0.13fF
C99 a_416_n140# a_2018_n140# 0.01fF
C100 a_n652_n140# a_60_n140# 0.03fF
C101 a_2432_n194# a_1008_n194# 0.01fF
C102 a_1008_n194# a_1364_n194# 0.03fF
C103 a_2196_n140# a_2552_n140# 0.06fF
C104 a_652_n194# a_1542_n194# 0.01fF
C105 a_2018_n140# a_2730_n140# 0.03fF
C106 a_n296_n140# a_n1720_n140# 0.01fF
C107 a_1898_n194# a_2610_n194# 0.01fF
C108 a_n2610_n140# a_n2966_n140# 0.06fF
C109 a_n1306_n194# a_n2908_n194# 0.01fF
C110 a_2254_n194# a_1008_n194# 0.01fF
C111 a_n1542_n140# a_n2254_n140# 0.03fF
C112 a_n2730_n194# a_n2908_n194# 0.10fF
C113 a_1720_n194# a_118_n194# 0.01fF
C114 a_n830_n140# a_n474_n140# 0.06fF
C115 a_238_n140# a_1128_n140# 0.02fF
C116 a_1186_n194# a_296_n194# 0.01fF
C117 a_n830_n140# a_60_n140# 0.02fF
C118 a_n1128_n194# a_n1306_n194# 0.10fF
C119 a_n2196_n194# a_n2908_n194# 0.01fF
C120 a_n1008_n140# a_n2076_n140# 0.02fF
C121 a_n950_n194# a_n1306_n194# 0.03fF
C122 a_n1662_n194# a_n238_n194# 0.01fF
C123 a_n2966_n140# a_n1720_n140# 0.02fF
C124 a_416_n140# a_1484_n140# 0.02fF
C125 a_n1128_n194# a_n2730_n194# 0.01fF
C126 a_n1306_n194# a_296_n194# 0.01fF
C127 a_n118_n140# a_238_n140# 0.06fF
C128 a_n1128_n194# a_n2196_n194# 0.01fF
C129 a_n652_n140# a_n118_n140# 0.04fF
C130 a_1484_n140# a_2730_n140# 0.02fF
C131 a_1840_n140# a_2374_n140# 0.04fF
C132 a_1662_n140# a_2552_n140# 0.02fF
C133 a_2018_n140# a_2196_n140# 0.13fF
C134 a_n1484_n194# a_n1306_n194# 0.10fF
C135 a_n950_n194# a_n2196_n194# 0.01fF
C136 a_474_n194# a_n60_n194# 0.02fF
C137 a_n2610_n140# a_n2254_n140# 0.06fF
C138 a_1008_n194# a_1898_n194# 0.01fF
C139 a_n1840_n194# a_n2374_n194# 0.02fF
C140 a_n1484_n194# a_n2730_n194# 0.01fF
C141 a_n296_n140# a_n474_n140# 0.13fF
C142 a_n296_n140# a_60_n140# 0.06fF
C143 a_n1484_n194# a_n2196_n194# 0.01fF
C144 a_n1186_n140# a_n1898_n140# 0.03fF
C145 a_118_n194# a_1364_n194# 0.01fF
C146 a_1542_n194# a_2076_n194# 0.02fF
C147 a_474_n194# a_830_n194# 0.03fF
C148 a_n416_n194# a_n1128_n194# 0.01fF
C149 a_n1542_n140# a_n1364_n140# 0.13fF
C150 a_n1720_n140# a_n2254_n140# 0.04fF
C151 a_n950_n194# a_n416_n194# 0.02fF
C152 a_652_n194# a_n594_n194# 0.01fF
C153 a_n416_n194# a_296_n194# 0.01fF
C154 a_n2788_n140# a_n1898_n140# 0.02fF
C155 a_n830_n140# a_n118_n140# 0.03fF
C156 a_1186_n194# a_2788_n194# 0.01fF
C157 a_2730_n140# a_2908_n140# 0.13fF
C158 a_2552_n140# a_3086_n140# 0.04fF
C159 a_652_n194# a_2076_n194# 0.01fF
C160 a_n1662_n194# a_n772_n194# 0.01fF
C161 a_416_n140# a_772_n140# 0.06fF
C162 a_n416_n194# a_n1484_n194# 0.01fF
C163 a_1720_n194# a_1542_n194# 0.10fF
C164 a_1662_n140# a_2018_n140# 0.06fF
C165 a_1128_n140# a_2552_n140# 0.01fF
C166 a_1484_n140# a_2196_n140# 0.03fF
C167 a_1306_n140# a_2374_n140# 0.02fF
C168 a_n2432_n140# a_n3144_n140# 0.03fF
C169 a_n2018_n194# a_n772_n194# 0.01fF
C170 a_n296_n140# a_1128_n140# 0.01fF
C171 a_n652_n140# a_238_n140# 0.02fF
C172 a_n2610_n140# a_n1364_n140# 0.02fF
C173 a_n1662_n194# a_n3086_n194# 0.01fF
C174 a_n2788_n140# a_n1186_n140# 0.01fF
C175 a_652_n194# a_1720_n194# 0.01fF
C176 a_n2018_n194# a_n3086_n194# 0.01fF
C177 a_n60_n194# a_830_n194# 0.01fF
C178 a_474_n194# a_1186_n194# 0.01fF
C179 a_n296_n140# a_n118_n140# 0.13fF
C180 a_n2432_n140# a_n830_n140# 0.01fF
C181 a_950_n140# a_2374_n140# 0.01fF
C182 a_594_n140# a_1840_n140# 0.02fF
C183 a_n1364_n140# a_n1720_n140# 0.06fF
C184 a_n1128_n194# a_n238_n194# 0.01fF
C185 a_n1542_n140# a_n2076_n140# 0.04fF
C186 a_2018_n140# a_3086_n140# 0.02fF
C187 a_2196_n140# a_2908_n140# 0.03fF
C188 a_n950_n194# a_n238_n194# 0.01fF
C189 a_n830_n140# a_238_n140# 0.02fF
C190 a_n238_n194# a_296_n194# 0.02fF
C191 a_2432_n194# a_1542_n194# 0.01fF
C192 a_1128_n140# a_2018_n140# 0.02fF
C193 a_1306_n140# a_1840_n140# 0.04fF
C194 a_1484_n140# a_1662_n140# 0.13fF
C195 a_n1008_n140# a_n1898_n140# 0.02fF
C196 a_1542_n194# a_1364_n194# 0.10fF
C197 a_n830_n140# a_n652_n140# 0.13fF
C198 a_2788_n194# a_2966_n194# 0.10fF
C199 a_60_n140# a_1484_n140# 0.01fF
C200 a_772_n140# a_2196_n140# 0.01fF
C201 a_n1484_n194# a_n238_n194# 0.01fF
C202 a_1008_n194# a_296_n194# 0.01fF
C203 a_n1306_n194# a_n2374_n194# 0.01fF
C204 a_652_n194# a_1364_n194# 0.01fF
C205 a_2254_n194# a_1542_n194# 0.01fF
C206 a_n1840_n194# a_n1306_n194# 0.02fF
C207 a_n2610_n140# a_n2076_n140# 0.04fF
C208 a_1186_n194# a_n60_n194# 0.01fF
C209 a_n2374_n194# a_n2730_n194# 0.03fF
C210 a_n1186_n140# a_n1008_n140# 0.13fF
C211 a_950_n140# a_1840_n140# 0.02fF
C212 a_n1840_n194# a_n2730_n194# 0.01fF
C213 a_594_n140# a_1306_n140# 0.03fF
C214 a_2788_n194# a_2610_n194# 0.10fF
C215 a_474_n194# a_n416_n194# 0.01fF
C216 a_n2196_n194# a_n2374_n194# 0.10fF
C217 a_n296_n140# a_238_n140# 0.04fF
C218 a_1720_n194# a_2076_n194# 0.03fF
C219 a_2254_n194# a_652_n194# 0.01fF
C220 a_n1840_n194# a_n2196_n194# 0.03fF
C221 a_1662_n140# a_2908_n140# 0.02fF
C222 a_1484_n140# a_3086_n140# 0.01fF
C223 a_n60_n194# a_n1306_n194# 0.01fF
C224 a_n652_n140# a_n296_n140# 0.06fF
C225 a_n1364_n140# a_n474_n140# 0.02fF
C226 a_1128_n140# a_1484_n140# 0.06fF
C227 a_n1128_n194# a_n772_n194# 0.03fF
C228 a_n2432_n140# a_n2966_n140# 0.04fF
C229 a_1186_n194# a_830_n194# 0.03fF
C230 a_n1720_n140# a_n2076_n140# 0.06fF
C231 a_n1364_n140# a_60_n140# 0.01fF
C232 a_n2908_n194# a_n3086_n194# 0.10fF
C233 a_n950_n194# a_n772_n194# 0.10fF
C234 a_296_n194# a_n772_n194# 0.01fF
C235 a_772_n140# a_1662_n140# 0.02fF
C236 a_n1008_n140# a_594_n140# 0.01fF
C237 a_594_n140# a_950_n140# 0.06fF
C238 a_1542_n194# a_1898_n194# 0.03fF
C239 a_n474_n140# a_772_n140# 0.02fF
C240 a_n1840_n194# a_n416_n194# 0.01fF
C241 a_60_n140# a_772_n140# 0.03fF
C242 a_n118_n140# a_1484_n140# 0.01fF
C243 a_n1484_n194# a_n772_n194# 0.01fF
C244 a_950_n140# a_1306_n140# 0.06fF
C245 a_652_n194# a_1898_n194# 0.01fF
C246 a_2908_n140# a_3086_n140# 0.13fF
C247 a_118_n194# a_n1128_n194# 0.01fF
C248 a_n830_n140# a_n296_n140# 0.04fF
C249 a_n2966_n140# a_n3144_n140# 0.13fF
C250 a_n950_n194# a_118_n194# 0.01fF
C251 a_2432_n194# a_2076_n194# 0.03fF
C252 a_n416_n194# a_n60_n194# 0.03fF
C253 a_2076_n194# a_1364_n194# 0.01fF
C254 a_n1484_n194# a_n3086_n194# 0.01fF
C255 a_118_n194# a_296_n194# 0.10fF
C256 a_n2432_n140# a_n2254_n140# 0.13fF
C257 a_474_n194# a_n238_n194# 0.01fF
C258 a_118_n194# a_n1484_n194# 0.01fF
C259 a_2374_n140# a_2730_n140# 0.06fF
C260 a_772_n140# a_1128_n140# 0.06fF
C261 a_n416_n194# a_830_n194# 0.01fF
C262 a_n474_n140# a_n2076_n140# 0.01fF
C263 a_n1364_n140# a_n118_n140# 0.02fF
C264 a_n1542_n140# a_n1898_n140# 0.06fF
C265 a_2254_n194# a_2076_n194# 0.10fF
C266 a_1720_n194# a_2432_n194# 0.01fF
C267 a_1720_n194# a_1364_n194# 0.03fF
C268 a_474_n194# a_1008_n194# 0.02fF
C269 a_n652_n140# a_n2254_n140# 0.01fF
C270 a_n1662_n194# a_n2552_n194# 0.01fF
C271 a_n118_n140# a_772_n140# 0.02fF
C272 a_238_n140# a_1484_n140# 0.02fF
C273 a_n3144_n140# a_n2254_n140# 0.02fF
C274 a_n1840_n194# a_n238_n194# 0.01fF
C275 a_n2018_n194# a_n2552_n194# 0.02fF
C276 a_2254_n194# a_1720_n194# 0.02fF
C277 a_n594_n194# a_n1662_n194# 0.01fF
C278 a_n1542_n140# a_n1186_n140# 0.06fF
C279 a_n1306_n194# a_n2730_n194# 0.01fF
C280 a_416_n140# a_1840_n140# 0.01fF
C281 a_n1186_n140# a_416_n140# 0.01fF
C282 a_n2018_n194# a_n594_n194# 0.01fF
C283 a_n2610_n140# a_n1898_n140# 0.03fF
C284 a_n2196_n194# a_n1306_n194# 0.01fF
C285 a_n2432_n140# a_n1364_n140# 0.02fF
C286 a_n60_n194# a_n238_n194# 0.10fF
C287 a_2076_n194# a_1898_n194# 0.10fF
C288 a_n2788_n140# a_n1542_n140# 0.02fF
C289 a_2196_n140# a_2374_n140# 0.13fF
C290 a_1840_n140# a_2730_n140# 0.02fF
C291 a_2018_n140# a_2552_n140# 0.04fF
C292 a_n830_n140# a_n2254_n140# 0.01fF
C293 a_n2196_n194# a_n2730_n194# 0.02fF
C294 a_1186_n194# a_n416_n194# 0.01fF
C295 a_474_n194# a_n772_n194# 0.01fF
C296 a_2432_n194# a_1364_n194# 0.01fF
C297 a_1008_n194# a_n60_n194# 0.01fF
C298 a_1542_n194# a_296_n194# 0.01fF
C299 a_n1720_n140# a_n1898_n140# 0.13fF
C300 a_n1364_n140# a_238_n140# 0.01fF
C301 a_416_n140# a_594_n140# 0.13fF
C302 a_n238_n194# a_830_n194# 0.01fF
C303 a_n2610_n140# a_n1186_n140# 0.01fF
C304 a_n652_n140# a_n1364_n140# 0.03fF
C305 a_1720_n194# a_1898_n194# 0.10fF
C306 a_n416_n194# a_n1306_n194# 0.01fF
C307 a_652_n194# a_n950_n194# 0.01fF
C308 a_2254_n194# a_2432_n194# 0.10fF
C309 a_2254_n194# a_1364_n194# 0.01fF
C310 a_238_n140# a_772_n140# 0.04fF
C311 a_1008_n194# a_830_n194# 0.10fF
C312 a_n772_n194# a_n2374_n194# 0.01fF
C313 a_416_n140# a_1306_n140# 0.02fF
C314 a_652_n194# a_296_n194# 0.03fF
C315 a_n2610_n140# a_n2788_n140# 0.13fF
C316 a_n1840_n194# a_n772_n194# 0.01fF
C317 a_n652_n140# a_772_n140# 0.01fF
C318 a_474_n194# a_118_n194# 0.03fF
C319 a_1186_n194# a_2610_n194# 0.01fF
C320 a_n1186_n140# a_n1720_n140# 0.04fF
C321 a_1306_n140# a_2730_n140# 0.01fF
C322 a_1840_n140# a_2196_n140# 0.06fF
C323 a_1662_n140# a_2374_n140# 0.03fF
C324 a_1484_n140# a_2552_n140# 0.02fF
C325 a_n2374_n194# a_n3086_n194# 0.01fF
C326 a_n2552_n194# a_n2908_n194# 0.03fF
C327 a_n1840_n194# a_n3086_n194# 0.01fF
C328 a_n60_n194# a_n772_n194# 0.01fF
C329 a_n2788_n140# a_n1720_n140# 0.02fF
C330 a_n2432_n140# a_n2076_n140# 0.06fF
C331 a_n830_n140# a_n1364_n140# 0.04fF
C332 a_n1542_n140# a_n1008_n140# 0.04fF
C333 a_416_n140# a_950_n140# 0.04fF
C334 a_n1008_n140# a_416_n140# 0.01fF
C335 a_2432_n194# a_1898_n194# 0.02fF
C336 a_1186_n194# a_n238_n194# 0.01fF
C337 a_n2966_n140# a_n2254_n140# 0.03fF
C338 a_n1128_n194# a_n2552_n194# 0.01fF
C339 a_1364_n194# a_1898_n194# 0.02fF
C340 a_n474_n140# a_n1898_n140# 0.01fF
C341 a_n950_n194# a_n2552_n194# 0.01fF
C342 a_n830_n140# a_772_n140# 0.01fF
C343 a_n772_n194# a_830_n194# 0.01fF
C344 a_594_n140# a_2196_n140# 0.01fF
C345 a_n652_n140# a_n2076_n140# 0.01fF
C346 a_1542_n194# a_2788_n194# 0.01fF
C347 a_n594_n194# a_n1128_n194# 0.02fF
C348 a_1186_n194# a_1008_n194# 0.10fF
C349 a_n238_n194# a_n1306_n194# 0.01fF
C350 a_n950_n194# a_n594_n194# 0.03fF
C351 a_2374_n140# a_3086_n140# 0.03fF
C352 a_2552_n140# a_2908_n140# 0.06fF
C353 a_118_n194# a_n60_n194# 0.10fF
C354 a_2254_n194# a_1898_n194# 0.03fF
C355 a_n594_n194# a_296_n194# 0.01fF
C356 a_n1484_n194# a_n2552_n194# 0.01fF
C357 a_n3144_n140# a_n2076_n140# 0.02fF
C358 a_1306_n140# a_2196_n140# 0.02fF
C359 a_n2610_n140# a_n1008_n140# 0.01fF
C360 a_1662_n140# a_1840_n140# 0.13fF
C361 a_1128_n140# a_2374_n140# 0.02fF
C362 a_1484_n140# a_2018_n140# 0.04fF
C363 a_n296_n140# a_n1364_n140# 0.02fF
C364 a_n1186_n140# a_n474_n140# 0.03fF
C365 a_2966_n194# a_2610_n194# 0.03fF
C366 a_n1186_n140# a_60_n140# 0.02fF
C367 a_n594_n194# a_n1484_n194# 0.01fF
C368 a_118_n194# a_830_n194# 0.01fF
C369 a_n296_n140# a_772_n140# 0.02fF
C370 a_474_n194# a_1542_n194# 0.01fF
C371 a_n830_n140# a_n2076_n140# 0.02fF
C372 a_n1008_n140# a_n1720_n140# 0.03fF
C373 a_950_n140# a_2196_n140# 0.02fF
C374 a_n2966_n140# a_n1364_n140# 0.01fF
C375 a_1720_n194# a_296_n194# 0.01fF
C376 a_594_n140# a_1662_n140# 0.02fF
C377 a_n416_n194# a_n238_n194# 0.10fF
C378 a_n2018_n194# a_n1662_n194# 0.03fF
C379 a_n474_n140# a_594_n140# 0.02fF
C380 a_652_n194# a_474_n194# 0.10fF
C381 a_60_n140# a_594_n140# 0.04fF
C382 a_1840_n140# a_3086_n140# 0.02fF
C383 a_2018_n140# a_2908_n140# 0.02fF
C384 a_n1306_n194# a_n772_n194# 0.02fF
C385 a_1306_n140# a_1662_n140# 0.06fF
C386 a_n416_n194# a_1008_n194# 0.01fF
C387 a_1128_n140# a_1840_n140# 0.03fF
C388 a_60_n140# a_1306_n140# 0.02fF
C389 a_772_n140# a_2018_n140# 0.02fF
C390 a_1186_n194# a_118_n194# 0.01fF
C391 a_n2196_n194# a_n772_n194# 0.01fF
C392 a_n1186_n140# a_n118_n140# 0.02fF
C393 a_1542_n194# a_n60_n194# 0.01fF
C394 a_2076_n194# a_2788_n194# 0.01fF
C395 a_n1364_n140# a_n2254_n140# 0.02fF
C396 a_n2730_n194# a_n3086_n194# 0.03fF
C397 a_950_n140# a_1662_n140# 0.03fF
C398 a_1008_n194# a_2610_n194# 0.01fF
C399 a_118_n194# a_n1306_n194# 0.01fF
C400 a_594_n140# a_1128_n140# 0.04fF
C401 a_n2432_n140# a_n1898_n140# 0.04fF
C402 a_n474_n140# a_950_n140# 0.01fF
C403 a_1364_n194# a_296_n194# 0.01fF
C404 a_n1008_n140# a_n474_n140# 0.04fF
C405 a_n2196_n194# a_n3086_n194# 0.01fF
C406 a_n1008_n140# a_60_n140# 0.02fF
C407 a_60_n140# a_950_n140# 0.02fF
C408 a_1484_n140# a_2908_n140# 0.01fF
C409 a_652_n194# a_n60_n194# 0.01fF
C410 a_1542_n194# a_830_n194# 0.01fF
C411 a_n416_n194# a_n772_n194# 0.03fF
C412 a_n2966_n140# a_n2076_n140# 0.02fF
C413 a_1128_n140# a_1306_n140# 0.13fF
C414 a_474_n194# a_n594_n194# 0.01fF
C415 a_1720_n194# a_2788_n194# 0.01fF
C416 a_n118_n140# a_594_n140# 0.03fF
C417 a_n652_n140# a_n1898_n140# 0.02fF
C418 a_n2610_n140# a_n1542_n140# 0.02fF
C419 a_772_n140# a_1484_n140# 0.03fF
C420 a_n2432_n140# a_n1186_n140# 0.02fF
C421 a_474_n194# a_2076_n194# 0.01fF
C422 a_1008_n194# a_n238_n194# 0.01fF
C423 a_652_n194# a_830_n194# 0.10fF
C424 a_n1662_n194# a_n2908_n194# 0.01fF
C425 a_n2374_n194# a_n2552_n194# 0.10fF
C426 a_n1840_n194# a_n2552_n194# 0.01fF
C427 a_n118_n140# a_1306_n140# 0.01fF
C428 a_n3144_n140# a_n1898_n140# 0.02fF
C429 a_n2018_n194# a_n2908_n194# 0.01fF
C430 a_n2432_n140# a_n2788_n140# 0.06fF
C431 a_n416_n194# a_118_n194# 0.02fF
C432 a_950_n140# a_1128_n140# 0.13fF
C433 a_n1840_n194# a_n594_n194# 0.01fF
C434 a_238_n140# a_1840_n140# 0.01fF
C435 a_n1186_n140# a_238_n140# 0.01fF
C436 a_n1128_n194# a_n1662_n194# 0.02fF
C437 a_n1542_n140# a_n1720_n140# 0.13fF
C438 a_n652_n140# a_n1186_n140# 0.04fF
C439 a_n950_n194# a_n1662_n194# 0.01fF
C440 a_1720_n194# a_474_n194# 0.01fF
C441 a_n2018_n194# a_n1128_n194# 0.01fF
C442 a_n2254_n140# a_n2076_n140# 0.13fF
C443 a_n950_n194# a_n2018_n194# 0.01fF
C444 a_1186_n194# a_1542_n194# 0.03fF
C445 a_n830_n140# a_n1898_n140# 0.02fF
C446 a_1898_n194# a_296_n194# 0.01fF
C447 a_n1008_n140# a_n118_n140# 0.02fF
C448 a_n118_n140# a_950_n140# 0.02fF
C449 a_2432_n194# a_2788_n194# 0.03fF
C450 a_n594_n194# a_n60_n194# 0.02fF
C451 a_2788_n194# a_1364_n194# 0.01fF
C452 a_n1662_n194# a_n1484_n194# 0.10fF
C453 a_2374_n140# a_2552_n140# 0.13fF
C454 a_2196_n140# a_2730_n140# 0.04fF
C455 a_n238_n194# a_n772_n194# 0.02fF
C456 a_238_n140# a_594_n140# 0.06fF
C457 a_n2788_n140# a_n3144_n140# 0.06fF
C458 a_n2018_n194# a_n1484_n194# 0.02fF
C459 a_652_n194# a_1186_n194# 0.02fF
C460 a_n652_n140# a_594_n140# 0.02fF
C461 a_n2610_n140# a_n1720_n140# 0.02fF
C462 a_n594_n194# a_830_n194# 0.01fF
C463 a_2254_n194# a_2788_n194# 0.02fF
C464 a_n830_n140# a_n1186_n140# 0.06fF
C465 a_238_n140# a_1306_n140# 0.02fF
C466 a_2076_n194# a_830_n194# 0.01fF
C467 a_n296_n140# a_n1898_n140# 0.01fF
C468 a_474_n194# a_1364_n194# 0.01fF
C469 a_n2432_n140# a_n1008_n140# 0.01fF
C470 a_416_n140# a_1662_n140# 0.02fF
C471 a_118_n194# a_n238_n194# 0.03fF
C472 a_n1542_n140# a_n474_n140# 0.02fF
C473 a_n474_n140# a_416_n140# 0.02fF
C474 a_n1364_n140# a_n2076_n140# 0.03fF
C475 a_n1542_n140# a_60_n140# 0.01fF
C476 a_416_n140# a_60_n140# 0.06fF
C477 a_n830_n140# a_594_n140# 0.01fF
C478 a_1840_n140# a_2552_n140# 0.03fF
C479 a_1008_n194# a_118_n194# 0.01fF
C480 a_2018_n140# a_2374_n140# 0.06fF
C481 a_1662_n140# a_2730_n140# 0.02fF
C482 a_n1008_n140# a_238_n140# 0.02fF
C483 a_1720_n194# a_830_n194# 0.01fF
C484 a_1542_n194# a_2966_n194# 0.01fF
C485 a_238_n140# a_950_n140# 0.03fF
C486 a_2788_n194# a_1898_n194# 0.01fF
C487 a_n296_n140# a_n1186_n140# 0.02fF
C488 a_n652_n140# a_n1008_n140# 0.06fF
C489 a_n652_n140# a_950_n140# 0.01fF
C490 a_n2966_n140# a_n1898_n140# 0.02fF
C491 a_652_n194# a_n416_n194# 0.01fF
C492 a_n1306_n194# a_n2552_n194# 0.01fF
C493 a_n2552_n194# a_n2730_n194# 0.10fF
C494 a_1186_n194# a_2076_n194# 0.01fF
C495 a_n950_n194# a_n1128_n194# 0.10fF
C496 a_n60_n194# a_1364_n194# 0.01fF
C497 a_416_n140# a_1128_n140# 0.03fF
C498 a_n594_n194# a_n1306_n194# 0.01fF
C499 a_n1484_n194# a_n2908_n194# 0.01fF
C500 a_1542_n194# a_2610_n194# 0.01fF
C501 a_n1128_n194# a_296_n194# 0.01fF
C502 a_n2196_n194# a_n2552_n194# 0.03fF
C503 a_n296_n140# a_594_n140# 0.02fF
C504 a_2730_n140# a_3086_n140# 0.06fF
C505 a_474_n194# a_1898_n194# 0.01fF
C506 a_n950_n194# a_296_n194# 0.01fF
C507 a_118_n194# a_n772_n194# 0.01fF
C508 a_n830_n140# a_n1008_n140# 0.13fF
C509 a_n1720_n140# a_n474_n140# 0.02fF
C510 a_1484_n140# a_2374_n140# 0.02fF
C511 a_1306_n140# a_2552_n140# 0.02fF
C512 a_1128_n140# a_2730_n140# 0.01fF
C513 a_1840_n140# a_2018_n140# 0.13fF
C514 a_1662_n140# a_2196_n140# 0.04fF
C515 a_2432_n194# a_830_n194# 0.01fF
C516 a_n1128_n194# a_n1484_n194# 0.03fF
C517 a_n594_n194# a_n2196_n194# 0.01fF
C518 a_n1542_n140# a_n118_n140# 0.01fF
C519 a_n2788_n140# a_n2966_n140# 0.13fF
C520 a_n2254_n140# a_n1898_n140# 0.06fF
C521 a_416_n140# a_n118_n140# 0.04fF
C522 a_1720_n194# a_1186_n194# 0.02fF
C523 a_1364_n194# a_830_n194# 0.02fF
C524 a_n950_n194# a_n1484_n194# 0.02fF
C525 a_n296_n140# a_1306_n140# 0.01fF
C526 a_n1662_n194# a_n2374_n194# 0.01fF
C527 a_n1840_n194# a_n1662_n194# 0.10fF
C528 a_n2018_n194# a_n2374_n194# 0.03fF
C529 a_2254_n194# a_830_n194# 0.01fF
C530 a_n1840_n194# a_n2018_n194# 0.10fF
C531 a_950_n140# a_2552_n140# 0.01fF
C532 a_n416_n194# a_n594_n194# 0.10fF
C533 a_1008_n194# a_1542_n194# 0.02fF
C534 a_594_n140# a_2018_n140# 0.01fF
C535 a_n1186_n140# a_n2254_n140# 0.02fF
C536 a_652_n194# a_n238_n194# 0.01fF
C537 a_n296_n140# a_n1008_n140# 0.03fF
C538 a_n296_n140# a_950_n140# 0.02fF
C539 a_n60_n194# a_n1662_n194# 0.01fF
C540 a_2374_n140# a_2908_n140# 0.04fF
C541 a_2196_n140# a_3086_n140# 0.02fF
C542 a_n2432_n140# a_n1542_n140# 0.02fF
C543 a_2076_n194# a_2966_n194# 0.01fF
C544 a_1128_n140# a_2196_n140# 0.02fF
C545 a_1484_n140# a_1840_n140# 0.06fF
C546 a_n2788_n140# a_n2254_n140# 0.04fF
C547 a_1306_n140# a_2018_n140# 0.03fF
C548 a_652_n194# a_1008_n194# 0.03fF
C549 a_3086_n140# VSUBS 0.02fF
C550 a_2908_n140# VSUBS 0.02fF
C551 a_2730_n140# VSUBS 0.02fF
C552 a_2552_n140# VSUBS 0.02fF
C553 a_2374_n140# VSUBS 0.02fF
C554 a_2196_n140# VSUBS 0.02fF
C555 a_2018_n140# VSUBS 0.02fF
C556 a_1840_n140# VSUBS 0.02fF
C557 a_1662_n140# VSUBS 0.02fF
C558 a_1484_n140# VSUBS 0.02fF
C559 a_1306_n140# VSUBS 0.02fF
C560 a_1128_n140# VSUBS 0.02fF
C561 a_950_n140# VSUBS 0.02fF
C562 a_772_n140# VSUBS 0.02fF
C563 a_594_n140# VSUBS 0.02fF
C564 a_416_n140# VSUBS 0.02fF
C565 a_238_n140# VSUBS 0.02fF
C566 a_60_n140# VSUBS 0.02fF
C567 a_n118_n140# VSUBS 0.02fF
C568 a_n296_n140# VSUBS 0.02fF
C569 a_n474_n140# VSUBS 0.02fF
C570 a_n652_n140# VSUBS 0.02fF
C571 a_n830_n140# VSUBS 0.02fF
C572 a_n1008_n140# VSUBS 0.02fF
C573 a_n1186_n140# VSUBS 0.02fF
C574 a_n1364_n140# VSUBS 0.02fF
C575 a_n1542_n140# VSUBS 0.02fF
C576 a_n1720_n140# VSUBS 0.02fF
C577 a_n1898_n140# VSUBS 0.02fF
C578 a_n2076_n140# VSUBS 0.02fF
C579 a_n2254_n140# VSUBS 0.02fF
C580 a_n2432_n140# VSUBS 0.02fF
C581 a_n2610_n140# VSUBS 0.02fF
C582 a_n2788_n140# VSUBS 0.02fF
C583 a_n2966_n140# VSUBS 0.02fF
C584 a_n3144_n140# VSUBS 0.02fF
C585 a_2966_n194# VSUBS 0.29fF
C586 a_2788_n194# VSUBS 0.23fF
C587 a_2610_n194# VSUBS 0.24fF
C588 a_2432_n194# VSUBS 0.25fF
C589 a_2254_n194# VSUBS 0.26fF
C590 a_2076_n194# VSUBS 0.27fF
C591 a_1898_n194# VSUBS 0.28fF
C592 a_1720_n194# VSUBS 0.28fF
C593 a_1542_n194# VSUBS 0.29fF
C594 a_1364_n194# VSUBS 0.29fF
C595 a_1186_n194# VSUBS 0.29fF
C596 a_1008_n194# VSUBS 0.29fF
C597 a_830_n194# VSUBS 0.29fF
C598 a_652_n194# VSUBS 0.29fF
C599 a_474_n194# VSUBS 0.29fF
C600 a_296_n194# VSUBS 0.29fF
C601 a_118_n194# VSUBS 0.29fF
C602 a_n60_n194# VSUBS 0.29fF
C603 a_n238_n194# VSUBS 0.29fF
C604 a_n416_n194# VSUBS 0.29fF
C605 a_n594_n194# VSUBS 0.29fF
C606 a_n772_n194# VSUBS 0.29fF
C607 a_n950_n194# VSUBS 0.29fF
C608 a_n1128_n194# VSUBS 0.29fF
C609 a_n1306_n194# VSUBS 0.29fF
C610 a_n1484_n194# VSUBS 0.29fF
C611 a_n1662_n194# VSUBS 0.29fF
C612 a_n1840_n194# VSUBS 0.29fF
C613 a_n2018_n194# VSUBS 0.29fF
C614 a_n2196_n194# VSUBS 0.29fF
C615 a_n2374_n194# VSUBS 0.29fF
C616 a_n2552_n194# VSUBS 0.29fF
C617 a_n2730_n194# VSUBS 0.29fF
C618 a_n2908_n194# VSUBS 0.29fF
C619 a_n3086_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BB a_n1008_n140# a_n652_n140# a_652_n194# a_772_n140#
+ a_n60_n194# a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140#
+ a_296_n194# a_60_n140# a_416_n140# a_n950_n194# a_n118_n140# a_118_n194# a_238_n140#
+ a_n772_n194# a_n830_n140# a_830_n194# a_950_n140# a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n474_n140# a_n652_n140# 0.13fF
C1 a_n772_n194# a_830_n194# 0.01fF
C2 a_n416_n194# a_118_n194# 0.02fF
C3 a_652_n194# a_118_n194# 0.02fF
C4 a_238_n140# a_416_n140# 0.13fF
C5 a_594_n140# a_n830_n140# 0.01fF
C6 a_296_n194# a_n238_n194# 0.02fF
C7 a_60_n140# a_594_n140# 0.04fF
C8 a_n594_n194# a_n238_n194# 0.03fF
C9 a_474_n194# a_n238_n194# 0.01fF
C10 a_n1008_n140# a_n296_n140# 0.03fF
C11 a_296_n194# a_118_n194# 0.10fF
C12 a_772_n140# a_416_n140# 0.06fF
C13 a_n594_n194# a_118_n194# 0.01fF
C14 a_474_n194# a_118_n194# 0.03fF
C15 a_416_n140# a_n118_n140# 0.04fF
C16 a_n652_n140# a_950_n140# 0.01fF
C17 a_n238_n194# a_830_n194# 0.01fF
C18 a_n296_n140# a_n652_n140# 0.06fF
C19 a_60_n140# a_n830_n140# 0.02fF
C20 a_830_n194# a_118_n194# 0.01fF
C21 a_n1008_n140# a_594_n140# 0.01fF
C22 a_n474_n140# a_416_n140# 0.02fF
C23 a_n772_n194# a_n60_n194# 0.01fF
C24 a_238_n140# a_772_n140# 0.04fF
C25 a_594_n140# a_n652_n140# 0.02fF
C26 a_238_n140# a_n118_n140# 0.06fF
C27 a_n1008_n140# a_n830_n140# 0.13fF
C28 a_n950_n194# a_n416_n194# 0.02fF
C29 a_n950_n194# a_652_n194# 0.01fF
C30 a_60_n140# a_n1008_n140# 0.02fF
C31 a_772_n140# a_n118_n140# 0.02fF
C32 a_238_n140# a_n474_n140# 0.03fF
C33 a_950_n140# a_416_n140# 0.04fF
C34 a_652_n194# a_n416_n194# 0.01fF
C35 a_n830_n140# a_n652_n140# 0.13fF
C36 a_n60_n194# a_n238_n194# 0.10fF
C37 a_n296_n140# a_416_n140# 0.03fF
C38 a_60_n140# a_n652_n140# 0.03fF
C39 a_n474_n140# a_772_n140# 0.02fF
C40 a_n60_n194# a_118_n194# 0.10fF
C41 a_n950_n194# a_296_n194# 0.01fF
C42 a_n474_n140# a_n118_n140# 0.06fF
C43 a_n950_n194# a_n594_n194# 0.03fF
C44 a_474_n194# a_n950_n194# 0.01fF
C45 a_296_n194# a_n416_n194# 0.01fF
C46 a_n594_n194# a_n416_n194# 0.10fF
C47 a_296_n194# a_652_n194# 0.03fF
C48 a_594_n140# a_416_n140# 0.13fF
C49 a_474_n194# a_n416_n194# 0.01fF
C50 a_652_n194# a_n594_n194# 0.01fF
C51 a_238_n140# a_950_n140# 0.03fF
C52 a_n772_n194# a_n238_n194# 0.02fF
C53 a_474_n194# a_652_n194# 0.10fF
C54 a_238_n140# a_n296_n140# 0.04fF
C55 a_n1008_n140# a_n652_n140# 0.06fF
C56 a_n772_n194# a_118_n194# 0.01fF
C57 a_n416_n194# a_830_n194# 0.01fF
C58 a_652_n194# a_830_n194# 0.10fF
C59 a_772_n140# a_950_n140# 0.13fF
C60 a_n296_n140# a_772_n140# 0.02fF
C61 a_n830_n140# a_416_n140# 0.02fF
C62 a_296_n194# a_n594_n194# 0.01fF
C63 a_950_n140# a_n118_n140# 0.02fF
C64 a_474_n194# a_296_n194# 0.10fF
C65 a_n296_n140# a_n118_n140# 0.13fF
C66 a_60_n140# a_416_n140# 0.06fF
C67 a_474_n194# a_n594_n194# 0.01fF
C68 a_238_n140# a_594_n140# 0.06fF
C69 a_n474_n140# a_950_n140# 0.01fF
C70 a_296_n194# a_830_n194# 0.02fF
C71 a_n594_n194# a_830_n194# 0.01fF
C72 a_n474_n140# a_n296_n140# 0.13fF
C73 a_594_n140# a_772_n140# 0.13fF
C74 a_474_n194# a_830_n194# 0.03fF
C75 a_n238_n194# a_118_n194# 0.03fF
C76 a_594_n140# a_n118_n140# 0.03fF
C77 a_238_n140# a_n830_n140# 0.02fF
C78 a_n950_n194# a_n60_n194# 0.01fF
C79 a_n1008_n140# a_416_n140# 0.01fF
C80 a_60_n140# a_238_n140# 0.13fF
C81 a_n416_n194# a_n60_n194# 0.03fF
C82 a_n474_n140# a_594_n140# 0.02fF
C83 a_n830_n140# a_772_n140# 0.01fF
C84 a_652_n194# a_n60_n194# 0.01fF
C85 a_n652_n140# a_416_n140# 0.02fF
C86 a_60_n140# a_772_n140# 0.03fF
C87 a_n830_n140# a_n118_n140# 0.03fF
C88 a_n296_n140# a_950_n140# 0.02fF
C89 a_60_n140# a_n118_n140# 0.13fF
C90 a_n950_n194# a_n772_n194# 0.10fF
C91 a_n1008_n140# a_238_n140# 0.02fF
C92 a_n474_n140# a_n830_n140# 0.06fF
C93 a_296_n194# a_n60_n194# 0.03fF
C94 a_n594_n194# a_n60_n194# 0.02fF
C95 a_n772_n194# a_n416_n194# 0.03fF
C96 a_60_n140# a_n474_n140# 0.04fF
C97 a_474_n194# a_n60_n194# 0.02fF
C98 a_n772_n194# a_652_n194# 0.01fF
C99 a_238_n140# a_n652_n140# 0.02fF
C100 a_594_n140# a_950_n140# 0.06fF
C101 a_n296_n140# a_594_n140# 0.02fF
C102 a_n1008_n140# a_n118_n140# 0.02fF
C103 a_n60_n194# a_830_n194# 0.01fF
C104 a_772_n140# a_n652_n140# 0.01fF
C105 a_n772_n194# a_296_n194# 0.01fF
C106 a_n950_n194# a_n238_n194# 0.01fF
C107 a_n772_n194# a_n594_n194# 0.10fF
C108 a_n652_n140# a_n118_n140# 0.04fF
C109 a_n1008_n140# a_n474_n140# 0.04fF
C110 a_474_n194# a_n772_n194# 0.01fF
C111 a_n950_n194# a_118_n194# 0.01fF
C112 a_n296_n140# a_n830_n140# 0.04fF
C113 a_n416_n194# a_n238_n194# 0.10fF
C114 a_60_n140# a_950_n140# 0.02fF
C115 a_652_n194# a_n238_n194# 0.01fF
C116 a_60_n140# a_n296_n140# 0.06fF
C117 a_950_n140# VSUBS 0.02fF
C118 a_772_n140# VSUBS 0.02fF
C119 a_594_n140# VSUBS 0.02fF
C120 a_416_n140# VSUBS 0.02fF
C121 a_238_n140# VSUBS 0.02fF
C122 a_60_n140# VSUBS 0.02fF
C123 a_n118_n140# VSUBS 0.02fF
C124 a_n296_n140# VSUBS 0.02fF
C125 a_n474_n140# VSUBS 0.02fF
C126 a_n652_n140# VSUBS 0.02fF
C127 a_n830_n140# VSUBS 0.02fF
C128 a_n1008_n140# VSUBS 0.02fF
C129 a_830_n194# VSUBS 0.29fF
C130 a_652_n194# VSUBS 0.23fF
C131 a_474_n194# VSUBS 0.24fF
C132 a_296_n194# VSUBS 0.25fF
C133 a_118_n194# VSUBS 0.26fF
C134 a_n60_n194# VSUBS 0.27fF
C135 a_n238_n194# VSUBS 0.28fF
C136 a_n416_n194# VSUBS 0.28fF
C137 a_n594_n194# VSUBS 0.29fF
C138 a_n772_n194# VSUBS 0.29fF
C139 a_n950_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_HH a_n1008_n140# a_n416_n205# a_1306_n140# a_n652_n140#
+ a_474_n205# a_n1484_n205# a_772_n140# a_n1720_n140# a_1720_n205# a_n238_n205# a_n474_n140#
+ a_296_n205# a_1128_n140# a_594_n140# a_1542_n205# a_n1306_n205# w_n2112_n240# a_n1542_n140#
+ a_n950_n205# a_1840_n140# a_1898_n205# a_n296_n140# a_n1898_n140# a_2018_n140# a_60_n140#
+ a_118_n205# a_n1128_n205# a_n1364_n140# a_1364_n205# a_416_n140# a_n772_n205# a_1662_n140#
+ a_830_n205# a_n1840_n205# a_n118_n140# a_1186_n205# a_n2018_n205# a_238_n140# a_n1186_n140#
+ a_n594_n205# a_1484_n140# a_n830_n140# a_652_n205# a_n1662_n205# a_950_n140# a_n60_n205#
+ a_n2076_n140# a_1008_n205# VSUBS
X0 a_1662_n140# a_1542_n205# a_1484_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n205# a_n296_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n205# a_n830_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_2018_n140# a_1898_n205# a_1840_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1008_n140# a_n1128_n205# a_n1186_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_594_n140# a_474_n205# a_416_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_60_n140# a_n60_n205# a_n118_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1484_n140# a_1364_n205# a_1306_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1542_n140# a_n1662_n205# a_n1720_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_950_n140# a_830_n205# a_772_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n830_n140# a_n950_n205# a_n1008_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n474_n140# a_n594_n205# a_n652_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_1840_n140# a_1720_n205# a_1662_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_416_n140# a_296_n205# a_238_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1898_n140# a_n2018_n205# a_n2076_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n296_n140# a_n416_n205# a_n474_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n1720_n140# a_n1840_n205# a_n1898_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1306_n140# a_1186_n205# a_1128_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1364_n140# a_n1484_n205# a_n1542_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_238_n140# a_118_n205# a_60_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_1128_n140# a_1008_n205# a_950_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_n1186_n140# a_n1306_n205# a_n1364_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_772_n140# a_652_n205# a_594_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n2076_n140# a_n830_n140# 0.02fF
C1 a_238_n140# a_n1364_n140# 0.01fF
C2 a_n2076_n140# a_n1898_n140# 0.13fF
C3 a_950_n140# a_594_n140# 0.06fF
C4 a_n118_n140# a_n652_n140# 0.04fF
C5 a_n1542_n140# a_n296_n140# 0.02fF
C6 a_n1186_n140# a_n652_n140# 0.04fF
C7 a_1364_n205# a_n60_n205# 0.01fF
C8 a_n1720_n140# w_n2112_n240# 0.02fF
C9 a_n1008_n140# a_n2076_n140# 0.02fF
C10 a_416_n140# a_2018_n140# 0.01fF
C11 a_416_n140# a_772_n140# 0.06fF
C12 a_652_n205# a_n416_n205# 0.01fF
C13 a_238_n140# a_1840_n140# 0.01fF
C14 a_1542_n205# w_n2112_n240# 0.19fF
C15 a_n1542_n140# a_n652_n140# 0.02fF
C16 a_n594_n205# a_n60_n205# 0.02fF
C17 a_1364_n205# a_1186_n205# 0.11fF
C18 a_n1128_n205# a_n60_n205# 0.01fF
C19 a_238_n140# a_594_n140# 0.06fF
C20 a_1542_n205# a_118_n205# 0.01fF
C21 a_772_n140# a_n118_n140# 0.02fF
C22 a_416_n140# w_n2112_n240# 0.02fF
C23 a_n830_n140# a_n296_n140# 0.04fF
C24 a_n2076_n140# a_n1364_n140# 0.03fF
C25 a_n1840_n205# a_n594_n205# 0.01fF
C26 a_n1898_n140# a_n296_n140# 0.01fF
C27 a_n1128_n205# a_n1840_n205# 0.01fF
C28 a_n2018_n205# a_n594_n205# 0.01fF
C29 a_830_n205# a_n60_n205# 0.01fF
C30 a_1840_n140# a_1128_n140# 0.03fF
C31 a_n1128_n205# a_n2018_n205# 0.01fF
C32 a_1542_n205# a_1008_n205# 0.02fF
C33 a_60_n140# a_n296_n140# 0.06fF
C34 a_416_n140# a_1662_n140# 0.02fF
C35 a_n1306_n205# a_n1662_n205# 0.03fF
C36 a_1364_n205# a_296_n205# 0.01fF
C37 a_n950_n205# a_n1662_n205# 0.01fF
C38 a_n1306_n205# a_n238_n205# 0.01fF
C39 a_n1008_n140# a_n296_n140# 0.03fF
C40 w_n2112_n240# a_n416_n205# 0.24fF
C41 a_n1484_n205# a_n594_n205# 0.01fF
C42 a_n950_n205# a_n238_n205# 0.01fF
C43 a_n1128_n205# a_n1484_n205# 0.03fF
C44 a_n1306_n205# a_n772_n205# 0.02fF
C45 a_n830_n140# a_n652_n140# 0.13fF
C46 a_594_n140# a_1128_n140# 0.04fF
C47 a_n1898_n140# a_n652_n140# 0.02fF
C48 a_830_n205# a_1186_n205# 0.03fF
C49 a_n118_n140# w_n2112_n240# 0.02fF
C50 a_n950_n205# a_n772_n205# 0.11fF
C51 a_60_n140# a_n652_n140# 0.03fF
C52 a_n594_n205# a_296_n205# 0.01fF
C53 a_n416_n205# a_118_n205# 0.02fF
C54 a_n1128_n205# a_296_n205# 0.01fF
C55 a_n1186_n140# w_n2112_n240# 0.02fF
C56 a_n1008_n140# a_n652_n140# 0.06fF
C57 a_1186_n205# a_1720_n205# 0.02fF
C58 a_1008_n205# a_n416_n205# 0.01fF
C59 a_416_n140# a_1306_n140# 0.02fF
C60 a_n950_n205# a_474_n205# 0.01fF
C61 a_n296_n140# a_n1364_n140# 0.02fF
C62 a_830_n205# a_296_n205# 0.02fF
C63 a_n474_n140# a_950_n140# 0.01fF
C64 a_n1542_n140# w_n2112_n240# 0.02fF
C65 a_950_n140# a_1484_n140# 0.04fF
C66 a_772_n140# a_n830_n140# 0.01fF
C67 a_1720_n205# a_296_n205# 0.01fF
C68 a_n1364_n140# a_n652_n140# 0.03fF
C69 a_772_n140# a_60_n140# 0.03fF
C70 a_n118_n140# a_1306_n140# 0.01fF
C71 a_n1662_n205# a_n60_n205# 0.01fF
C72 a_n238_n205# a_n60_n205# 0.11fF
C73 a_n296_n140# a_594_n140# 0.02fF
C74 a_n772_n205# a_n60_n205# 0.01fF
C75 a_n1840_n205# a_n1662_n205# 0.11fF
C76 a_238_n140# a_n474_n140# 0.03fF
C77 a_n2018_n205# a_n1662_n205# 0.03fF
C78 a_n830_n140# w_n2112_n240# 0.02fF
C79 a_238_n140# a_1484_n140# 0.02fF
C80 a_n1840_n205# a_n238_n205# 0.01fF
C81 a_n1898_n140# w_n2112_n240# 0.02fF
C82 a_n950_n205# a_652_n205# 0.01fF
C83 a_1186_n205# a_n238_n205# 0.01fF
C84 a_60_n140# w_n2112_n240# 0.02fF
C85 a_n1840_n205# a_n772_n205# 0.01fF
C86 a_n2018_n205# a_n772_n205# 0.01fF
C87 a_n1484_n205# a_n1662_n205# 0.11fF
C88 a_1364_n205# a_830_n205# 0.02fF
C89 a_474_n205# a_n60_n205# 0.02fF
C90 a_n652_n140# a_594_n140# 0.02fF
C91 a_60_n140# a_1662_n140# 0.01fF
C92 a_n1008_n140# w_n2112_n240# 0.02fF
C93 a_n1128_n205# a_n594_n205# 0.02fF
C94 a_n1484_n205# a_n238_n205# 0.01fF
C95 a_n1720_n140# a_n118_n140# 0.01fF
C96 a_n1484_n205# a_n772_n205# 0.01fF
C97 a_n1720_n140# a_n1186_n140# 0.04fF
C98 a_1364_n205# a_1720_n205# 0.03fF
C99 a_n474_n140# a_1128_n140# 0.01fF
C100 a_n238_n205# a_296_n205# 0.02fF
C101 a_1484_n140# a_1128_n140# 0.06fF
C102 a_830_n205# a_n594_n205# 0.01fF
C103 a_474_n205# a_1186_n205# 0.01fF
C104 a_238_n140# a_950_n140# 0.03fF
C105 a_1840_n140# a_2018_n140# 0.13fF
C106 a_772_n140# a_1840_n140# 0.02fF
C107 a_n772_n205# a_296_n205# 0.01fF
C108 a_n2076_n140# a_n474_n140# 0.01fF
C109 a_n1306_n205# w_n2112_n240# 0.24fF
C110 a_n1542_n140# a_n1720_n140# 0.13fF
C111 a_n1364_n140# w_n2112_n240# 0.02fF
C112 a_416_n140# a_n118_n140# 0.04fF
C113 a_n950_n205# w_n2112_n240# 0.24fF
C114 a_60_n140# a_1306_n140# 0.02fF
C115 a_2018_n140# a_594_n140# 0.01fF
C116 a_772_n140# a_594_n140# 0.13fF
C117 a_n1306_n205# a_118_n205# 0.01fF
C118 a_416_n140# a_n1186_n140# 0.01fF
C119 a_474_n205# a_296_n205# 0.11fF
C120 a_652_n205# a_n60_n205# 0.01fF
C121 a_n950_n205# a_118_n205# 0.01fF
C122 w_n2112_n240# a_1840_n140# 0.02fF
C123 a_830_n205# a_1720_n205# 0.01fF
C124 a_950_n140# a_1128_n140# 0.13fF
C125 a_1840_n140# a_1662_n140# 0.13fF
C126 w_n2112_n240# a_594_n140# 0.02fF
C127 a_n830_n140# a_n1720_n140# 0.02fF
C128 a_652_n205# a_1186_n205# 0.02fF
C129 a_1364_n205# a_n238_n205# 0.01fF
C130 a_n1186_n140# a_n118_n140# 0.02fF
C131 a_n1720_n140# a_n1898_n140# 0.13fF
C132 a_n474_n140# a_n296_n140# 0.13fF
C133 a_1662_n140# a_594_n140# 0.02fF
C134 a_1898_n205# a_1186_n205# 0.01fF
C135 a_n1662_n205# a_n594_n205# 0.01fF
C136 a_n1008_n140# a_n1720_n140# 0.03fF
C137 a_n1128_n205# a_n1662_n205# 0.02fF
C138 a_238_n140# a_1128_n140# 0.02fF
C139 a_n1542_n140# a_n118_n140# 0.01fF
C140 a_n594_n205# a_n238_n205# 0.03fF
C141 a_n1128_n205# a_n238_n205# 0.01fF
C142 a_652_n205# a_296_n205# 0.03fF
C143 w_n2112_n240# a_n60_n205# 0.24fF
C144 a_n474_n140# a_n652_n140# 0.13fF
C145 a_1840_n140# a_1306_n140# 0.04fF
C146 a_1364_n205# a_474_n205# 0.01fF
C147 a_n772_n205# a_n594_n205# 0.11fF
C148 a_n1542_n140# a_n1186_n140# 0.06fF
C149 a_416_n140# a_n830_n140# 0.02fF
C150 a_n1128_n205# a_n772_n205# 0.03fF
C151 a_1898_n205# a_296_n205# 0.01fF
C152 a_416_n140# a_60_n140# 0.06fF
C153 a_n1840_n205# w_n2112_n240# 0.24fF
C154 a_n60_n205# a_118_n205# 0.11fF
C155 a_830_n205# a_n238_n205# 0.01fF
C156 a_n2018_n205# w_n2112_n240# 0.31fF
C157 a_1306_n140# a_594_n140# 0.03fF
C158 a_n296_n140# a_950_n140# 0.02fF
C159 a_1186_n205# w_n2112_n240# 0.21fF
C160 a_n1008_n140# a_416_n140# 0.01fF
C161 a_830_n205# a_n772_n205# 0.01fF
C162 a_n1720_n140# a_n1364_n140# 0.06fF
C163 a_1008_n205# a_n60_n205# 0.01fF
C164 a_474_n205# a_n594_n205# 0.01fF
C165 a_n1128_n205# a_474_n205# 0.01fF
C166 a_n1484_n205# w_n2112_n240# 0.24fF
C167 a_n830_n140# a_n118_n140# 0.03fF
C168 a_1186_n205# a_118_n205# 0.01fF
C169 a_60_n140# a_n118_n140# 0.13fF
C170 a_n830_n140# a_n1186_n140# 0.06fF
C171 a_474_n205# a_830_n205# 0.03fF
C172 a_n652_n140# a_950_n140# 0.01fF
C173 a_772_n140# a_n474_n140# 0.02fF
C174 w_n2112_n240# a_296_n205# 0.24fF
C175 a_n1186_n140# a_n1898_n140# 0.03fF
C176 a_1008_n205# a_1186_n205# 0.11fF
C177 a_n1484_n205# a_118_n205# 0.01fF
C178 a_2018_n140# a_1484_n140# 0.04fF
C179 a_772_n140# a_1484_n140# 0.03fF
C180 a_n1008_n140# a_n118_n140# 0.02fF
C181 a_n1186_n140# a_60_n140# 0.02fF
C182 a_1364_n205# a_652_n205# 0.01fF
C183 a_238_n140# a_n296_n140# 0.04fF
C184 a_474_n205# a_1720_n205# 0.01fF
C185 a_n1008_n140# a_n1186_n140# 0.13fF
C186 a_118_n205# a_296_n205# 0.11fF
C187 a_n1542_n140# a_n830_n140# 0.03fF
C188 a_n1542_n140# a_n1898_n140# 0.06fF
C189 a_1364_n205# a_1898_n205# 0.02fF
C190 a_n1306_n205# a_n416_n205# 0.01fF
C191 a_1008_n205# a_296_n205# 0.01fF
C192 a_n1542_n140# a_60_n140# 0.01fF
C193 a_416_n140# a_1840_n140# 0.01fF
C194 a_n474_n140# w_n2112_n240# 0.02fF
C195 a_652_n205# a_n594_n205# 0.01fF
C196 w_n2112_n240# a_1484_n140# 0.02fF
C197 a_n950_n205# a_n416_n205# 0.02fF
C198 a_238_n140# a_n652_n140# 0.02fF
C199 a_n1008_n140# a_n1542_n140# 0.04fF
C200 a_n118_n140# a_n1364_n140# 0.02fF
C201 a_n1662_n205# a_n238_n205# 0.01fF
C202 a_1662_n140# a_1484_n140# 0.13fF
C203 a_950_n140# a_2018_n140# 0.02fF
C204 a_772_n140# a_950_n140# 0.13fF
C205 a_n296_n140# a_1128_n140# 0.01fF
C206 a_n772_n205# a_n1662_n205# 0.01fF
C207 a_416_n140# a_594_n140# 0.13fF
C208 a_n1186_n140# a_n1364_n140# 0.13fF
C209 a_830_n205# a_652_n205# 0.11fF
C210 a_n772_n205# a_n238_n205# 0.02fF
C211 a_1542_n205# a_n60_n205# 0.01fF
C212 a_1364_n205# w_n2112_n240# 0.20fF
C213 a_n830_n140# a_n1898_n140# 0.02fF
C214 a_1898_n205# a_830_n205# 0.01fF
C215 a_n830_n140# a_60_n140# 0.02fF
C216 a_652_n205# a_1720_n205# 0.01fF
C217 a_n1542_n140# a_n1364_n140# 0.13fF
C218 w_n2112_n240# a_950_n140# 0.02fF
C219 a_1364_n205# a_118_n205# 0.01fF
C220 a_n1008_n140# a_n830_n140# 0.13fF
C221 a_474_n205# a_n238_n205# 0.01fF
C222 a_n118_n140# a_594_n140# 0.03fF
C223 a_n1008_n140# a_n1898_n140# 0.02fF
C224 a_1898_n205# a_1720_n205# 0.11fF
C225 w_n2112_n240# a_n594_n205# 0.24fF
C226 a_772_n140# a_238_n140# 0.04fF
C227 a_1542_n205# a_1186_n205# 0.03fF
C228 a_n1128_n205# w_n2112_n240# 0.24fF
C229 a_1306_n140# a_1484_n140# 0.13fF
C230 a_1662_n140# a_950_n140# 0.03fF
C231 a_1364_n205# a_1008_n205# 0.03fF
C232 a_n1008_n140# a_60_n140# 0.02fF
C233 a_n2076_n140# a_n652_n140# 0.01fF
C234 a_474_n205# a_n772_n205# 0.01fF
C235 a_n416_n205# a_n60_n205# 0.03fF
C236 a_n594_n205# a_118_n205# 0.01fF
C237 a_n1128_n205# a_118_n205# 0.01fF
C238 a_830_n205# w_n2112_n240# 0.23fF
C239 a_1542_n205# a_296_n205# 0.01fF
C240 a_1008_n205# a_n594_n205# 0.01fF
C241 a_n830_n140# a_n1364_n140# 0.04fF
C242 a_238_n140# w_n2112_n240# 0.02fF
C243 a_n1840_n205# a_n416_n205# 0.01fF
C244 a_n1898_n140# a_n1364_n140# 0.04fF
C245 a_n2018_n205# a_n416_n205# 0.01fF
C246 a_830_n205# a_118_n205# 0.01fF
C247 a_2018_n140# a_1128_n140# 0.02fF
C248 a_772_n140# a_1128_n140# 0.06fF
C249 w_n2112_n240# a_1720_n205# 0.18fF
C250 a_60_n140# a_n1364_n140# 0.01fF
C251 a_1186_n205# a_n416_n205# 0.01fF
C252 a_238_n140# a_1662_n140# 0.01fF
C253 a_n1720_n140# a_n474_n140# 0.02fF
C254 a_1306_n140# a_950_n140# 0.06fF
C255 a_1008_n205# a_830_n205# 0.11fF
C256 a_n1008_n140# a_n1364_n140# 0.06fF
C257 a_652_n205# a_n238_n205# 0.01fF
C258 a_n1484_n205# a_n416_n205# 0.01fF
C259 a_1720_n205# a_118_n205# 0.01fF
C260 a_n296_n140# a_n652_n140# 0.06fF
C261 a_n772_n205# a_652_n205# 0.01fF
C262 a_1008_n205# a_1720_n205# 0.01fF
C263 a_n416_n205# a_296_n205# 0.01fF
C264 w_n2112_n240# a_1128_n140# 0.02fF
C265 a_n830_n140# a_594_n140# 0.01fF
C266 a_416_n140# a_n474_n140# 0.02fF
C267 a_1662_n140# a_1128_n140# 0.04fF
C268 a_416_n140# a_1484_n140# 0.02fF
C269 a_60_n140# a_594_n140# 0.04fF
C270 a_474_n205# a_652_n205# 0.11fF
C271 a_238_n140# a_1306_n140# 0.02fF
C272 a_n2076_n140# w_n2112_n240# 0.02fF
C273 a_n950_n205# a_n1306_n205# 0.03fF
C274 a_1542_n205# a_1364_n205# 0.11fF
C275 a_n1008_n140# a_594_n140# 0.01fF
C276 a_n1662_n205# w_n2112_n240# 0.24fF
C277 a_474_n205# a_1898_n205# 0.01fF
C278 w_n2112_n240# a_n238_n205# 0.24fF
C279 a_772_n140# a_n296_n140# 0.02fF
C280 a_n118_n140# a_n474_n140# 0.06fF
C281 a_n118_n140# a_1484_n140# 0.01fF
C282 a_n772_n205# w_n2112_n240# 0.24fF
C283 a_n1186_n140# a_n474_n140# 0.03fF
C284 a_n238_n205# a_118_n205# 0.03fF
C285 a_1306_n140# a_1128_n140# 0.13fF
C286 a_416_n140# a_950_n140# 0.04fF
C287 a_n772_n205# a_118_n205# 0.01fF
C288 a_1542_n205# a_830_n205# 0.01fF
C289 a_772_n140# a_n652_n140# 0.01fF
C290 a_1008_n205# a_n238_n205# 0.01fF
C291 a_474_n205# w_n2112_n240# 0.24fF
C292 a_n296_n140# w_n2112_n240# 0.02fF
C293 a_n1542_n140# a_n474_n140# 0.02fF
C294 a_1840_n140# a_594_n140# 0.02fF
C295 a_1542_n205# a_1720_n205# 0.11fF
C296 a_1898_n205# a_652_n205# 0.01fF
C297 a_n1306_n205# a_n60_n205# 0.01fF
C298 a_474_n205# a_118_n205# 0.03fF
C299 a_n594_n205# a_n416_n205# 0.11fF
C300 a_n118_n140# a_950_n140# 0.02fF
C301 a_n1128_n205# a_n416_n205# 0.01fF
C302 a_n950_n205# a_n60_n205# 0.01fF
C303 a_416_n140# a_238_n140# 0.13fF
C304 a_474_n205# a_1008_n205# 0.02fF
C305 a_n652_n140# w_n2112_n240# 0.02fF
C306 a_n1840_n205# a_n1306_n205# 0.02fF
C307 a_n2018_n205# a_n1306_n205# 0.01fF
C308 a_n950_n205# a_n1840_n205# 0.01fF
C309 a_830_n205# a_n416_n205# 0.01fF
C310 a_n2018_n205# a_n950_n205# 0.01fF
C311 a_n2076_n140# a_n1720_n140# 0.06fF
C312 a_772_n140# a_2018_n140# 0.02fF
C313 a_n830_n140# a_n474_n140# 0.06fF
C314 a_n474_n140# a_n1898_n140# 0.01fF
C315 a_n1306_n205# a_n1484_n205# 0.11fF
C316 a_n296_n140# a_1306_n140# 0.01fF
C317 a_652_n205# w_n2112_n240# 0.24fF
C318 a_60_n140# a_n474_n140# 0.04fF
C319 a_238_n140# a_n118_n140# 0.06fF
C320 a_n950_n205# a_n1484_n205# 0.02fF
C321 a_60_n140# a_1484_n140# 0.01fF
C322 a_416_n140# a_1128_n140# 0.03fF
C323 a_n1008_n140# a_n474_n140# 0.04fF
C324 a_1898_n205# w_n2112_n240# 0.24fF
C325 a_n1306_n205# a_296_n205# 0.01fF
C326 a_238_n140# a_n1186_n140# 0.01fF
C327 a_652_n205# a_118_n205# 0.02fF
C328 a_n950_n205# a_296_n205# 0.01fF
C329 a_772_n140# w_n2112_n240# 0.02fF
C330 w_n2112_n240# a_2018_n140# 0.02fF
C331 a_1008_n205# a_652_n205# 0.03fF
C332 a_1662_n140# a_2018_n140# 0.06fF
C333 a_772_n140# a_1662_n140# 0.02fF
C334 a_1898_n205# a_1008_n205# 0.01fF
C335 a_n118_n140# a_1128_n140# 0.02fF
C336 a_n1720_n140# a_n296_n140# 0.01fF
C337 a_n474_n140# a_n1364_n140# 0.02fF
C338 a_60_n140# a_950_n140# 0.02fF
C339 a_1542_n205# a_474_n205# 0.01fF
C340 a_1186_n205# a_n60_n205# 0.01fF
C341 a_n1662_n205# a_n416_n205# 0.01fF
C342 w_n2112_n240# a_1662_n140# 0.02fF
C343 a_n2076_n140# a_n1186_n140# 0.02fF
C344 a_n416_n205# a_n238_n205# 0.11fF
C345 w_n2112_n240# a_118_n205# 0.24fF
C346 a_n2018_n205# a_n1840_n205# 0.11fF
C347 a_n1720_n140# a_n652_n140# 0.02fF
C348 a_n1484_n205# a_n60_n205# 0.01fF
C349 a_1840_n140# a_1484_n140# 0.06fF
C350 a_1306_n140# a_2018_n140# 0.03fF
C351 a_772_n140# a_1306_n140# 0.04fF
C352 a_n772_n205# a_n416_n205# 0.03fF
C353 a_238_n140# a_n830_n140# 0.02fF
C354 a_416_n140# a_n296_n140# 0.03fF
C355 a_1008_n205# w_n2112_n240# 0.22fF
C356 a_n1840_n205# a_n1484_n205# 0.03fF
C357 a_n60_n205# a_296_n205# 0.03fF
C358 a_238_n140# a_60_n140# 0.13fF
C359 a_n474_n140# a_594_n140# 0.02fF
C360 a_n1542_n140# a_n2076_n140# 0.04fF
C361 a_n2018_n205# a_n1484_n205# 0.02fF
C362 a_1484_n140# a_594_n140# 0.02fF
C363 a_n1306_n205# a_n594_n205# 0.01fF
C364 a_n1008_n140# a_238_n140# 0.02fF
C365 a_1008_n205# a_118_n205# 0.01fF
C366 a_474_n205# a_n416_n205# 0.01fF
C367 a_n1128_n205# a_n1306_n205# 0.11fF
C368 w_n2112_n240# a_1306_n140# 0.02fF
C369 a_n950_n205# a_n594_n205# 0.03fF
C370 a_416_n140# a_n652_n140# 0.02fF
C371 a_n1128_n205# a_n950_n205# 0.11fF
C372 a_n118_n140# a_n296_n140# 0.13fF
C373 a_1186_n205# a_296_n205# 0.01fF
C374 a_1542_n205# a_652_n205# 0.01fF
C375 a_1306_n140# a_1662_n140# 0.06fF
C376 a_1840_n140# a_950_n140# 0.02fF
C377 a_n1186_n140# a_n296_n140# 0.02fF
C378 a_1542_n205# a_1898_n205# 0.03fF
C379 a_60_n140# a_1128_n140# 0.02fF
C380 w_n2112_n240# VSUBS 6.08fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_GG a_n652_n140# a_652_n194# a_772_n140# a_n60_n194#
+ a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140# a_296_n194#
+ a_60_n140# a_416_n140# a_n118_n140# a_118_n194# a_238_n140# a_n772_n194# a_n830_n140#
+ a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n830_n140# a_n296_n140# 0.04fF
C1 a_594_n140# a_n652_n140# 0.02fF
C2 a_238_n140# a_n296_n140# 0.04fF
C3 a_474_n194# a_n772_n194# 0.01fF
C4 a_594_n140# a_n296_n140# 0.02fF
C5 a_474_n194# a_118_n194# 0.03fF
C6 a_n118_n140# a_n652_n140# 0.04fF
C7 a_n772_n194# a_n60_n194# 0.01fF
C8 a_296_n194# a_n594_n194# 0.01fF
C9 a_60_n140# a_n652_n140# 0.03fF
C10 a_n118_n140# a_n296_n140# 0.13fF
C11 a_118_n194# a_n60_n194# 0.10fF
C12 a_60_n140# a_n296_n140# 0.06fF
C13 a_296_n194# a_n238_n194# 0.02fF
C14 a_n652_n140# a_416_n140# 0.02fF
C15 a_416_n140# a_n296_n140# 0.03fF
C16 a_474_n194# a_n416_n194# 0.01fF
C17 a_652_n194# a_n594_n194# 0.01fF
C18 a_772_n140# a_n830_n140# 0.01fF
C19 a_772_n140# a_238_n140# 0.04fF
C20 a_n416_n194# a_n60_n194# 0.03fF
C21 a_594_n140# a_772_n140# 0.13fF
C22 a_652_n194# a_n238_n194# 0.01fF
C23 a_n772_n194# a_n594_n194# 0.10fF
C24 a_n118_n140# a_772_n140# 0.02fF
C25 a_238_n140# a_n830_n140# 0.02fF
C26 a_n474_n140# a_n652_n140# 0.13fF
C27 a_n594_n194# a_118_n194# 0.01fF
C28 a_60_n140# a_772_n140# 0.03fF
C29 a_474_n194# a_n60_n194# 0.02fF
C30 a_594_n140# a_n830_n140# 0.01fF
C31 a_n772_n194# a_n238_n194# 0.02fF
C32 a_n474_n140# a_n296_n140# 0.13fF
C33 a_594_n140# a_238_n140# 0.06fF
C34 a_296_n194# a_652_n194# 0.03fF
C35 a_n238_n194# a_118_n194# 0.03fF
C36 a_772_n140# a_416_n140# 0.06fF
C37 a_n118_n140# a_n830_n140# 0.03fF
C38 a_n118_n140# a_238_n140# 0.06fF
C39 a_60_n140# a_n830_n140# 0.02fF
C40 a_60_n140# a_238_n140# 0.13fF
C41 a_594_n140# a_n118_n140# 0.03fF
C42 a_296_n194# a_n772_n194# 0.01fF
C43 a_60_n140# a_594_n140# 0.04fF
C44 a_n830_n140# a_416_n140# 0.02fF
C45 a_n594_n194# a_n416_n194# 0.10fF
C46 a_296_n194# a_118_n194# 0.10fF
C47 a_238_n140# a_416_n140# 0.13fF
C48 a_594_n140# a_416_n140# 0.13fF
C49 a_60_n140# a_n118_n140# 0.13fF
C50 a_n238_n194# a_n416_n194# 0.10fF
C51 a_n118_n140# a_416_n140# 0.04fF
C52 a_474_n194# a_n594_n194# 0.01fF
C53 a_772_n140# a_n474_n140# 0.02fF
C54 a_60_n140# a_416_n140# 0.06fF
C55 a_n652_n140# a_n296_n140# 0.06fF
C56 a_652_n194# a_n772_n194# 0.01fF
C57 a_n594_n194# a_n60_n194# 0.02fF
C58 a_652_n194# a_118_n194# 0.02fF
C59 a_296_n194# a_n416_n194# 0.01fF
C60 a_474_n194# a_n238_n194# 0.01fF
C61 a_n830_n140# a_n474_n140# 0.06fF
C62 a_238_n140# a_n474_n140# 0.03fF
C63 a_n238_n194# a_n60_n194# 0.10fF
C64 a_594_n140# a_n474_n140# 0.02fF
C65 a_n772_n194# a_118_n194# 0.01fF
C66 a_296_n194# a_474_n194# 0.10fF
C67 a_n118_n140# a_n474_n140# 0.06fF
C68 a_652_n194# a_n416_n194# 0.01fF
C69 a_296_n194# a_n60_n194# 0.03fF
C70 a_60_n140# a_n474_n140# 0.04fF
C71 a_772_n140# a_n652_n140# 0.01fF
C72 a_n474_n140# a_416_n140# 0.02fF
C73 a_772_n140# a_n296_n140# 0.02fF
C74 a_n772_n194# a_n416_n194# 0.03fF
C75 a_474_n194# a_652_n194# 0.10fF
C76 a_n416_n194# a_118_n194# 0.02fF
C77 a_n830_n140# a_n652_n140# 0.13fF
C78 a_n238_n194# a_n594_n194# 0.03fF
C79 a_238_n140# a_n652_n140# 0.02fF
C80 a_652_n194# a_n60_n194# 0.01fF
C81 a_772_n140# VSUBS 0.02fF
C82 a_594_n140# VSUBS 0.02fF
C83 a_416_n140# VSUBS 0.02fF
C84 a_238_n140# VSUBS 0.02fF
C85 a_60_n140# VSUBS 0.02fF
C86 a_n118_n140# VSUBS 0.02fF
C87 a_n296_n140# VSUBS 0.02fF
C88 a_n474_n140# VSUBS 0.02fF
C89 a_n652_n140# VSUBS 0.02fF
C90 a_n830_n140# VSUBS 0.02fF
C91 a_652_n194# VSUBS 0.29fF
C92 a_474_n194# VSUBS 0.23fF
C93 a_296_n194# VSUBS 0.24fF
C94 a_118_n194# VSUBS 0.25fF
C95 a_n60_n194# VSUBS 0.26fF
C96 a_n238_n194# VSUBS 0.27fF
C97 a_n416_n194# VSUBS 0.28fF
C98 a_n594_n194# VSUBS 0.28fF
C99 a_n772_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_AA a_n149_n194# a_n207_n140# a_207_n194# a_n1217_n194#
+ a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140# a_n1097_n140#
+ a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194# a_861_n140#
+ a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140# a_n919_n140#
+ a_919_n194# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194# a_n1395_n194# a_505_n140#
+ a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n29_n140# a_1395_n140# 0.01fF
C1 a_149_n140# a_n741_n140# 0.02fF
C2 a_n861_n194# a_563_n194# 0.01fF
C3 a_861_n140# a_1395_n140# 0.04fF
C4 a_327_n140# a_n207_n140# 0.04fF
C5 a_n149_n194# a_919_n194# 0.01fF
C6 a_505_n140# a_1395_n140# 0.02fF
C7 a_1097_n194# a_563_n194# 0.02fF
C8 a_n861_n194# a_n683_n194# 0.10fF
C9 a_n1039_n194# a_385_n194# 0.01fF
C10 a_n1275_n140# a_n563_n140# 0.03fF
C11 a_n327_n194# a_563_n194# 0.01fF
C12 a_n1275_n140# a_n385_n140# 0.02fF
C13 a_n1039_n194# a_n505_n194# 0.02fF
C14 a_n1097_n140# a_n741_n140# 0.06fF
C15 a_683_n140# a_n741_n140# 0.01fF
C16 a_n861_n194# a_207_n194# 0.01fF
C17 a_n1453_n140# a_n741_n140# 0.03fF
C18 a_n1275_n140# a_n919_n140# 0.06fF
C19 a_1217_n140# a_1395_n140# 0.13fF
C20 a_149_n140# a_1395_n140# 0.02fF
C21 a_n327_n194# a_n683_n194# 0.03fF
C22 a_n29_n140# a_n207_n140# 0.13fF
C23 a_1097_n194# a_207_n194# 0.01fF
C24 a_919_n194# a_385_n194# 0.02fF
C25 a_861_n140# a_n207_n140# 0.02fF
C26 a_1039_n140# a_1395_n140# 0.06fF
C27 a_n683_n194# a_n1217_n194# 0.02fF
C28 a_n505_n194# a_919_n194# 0.01fF
C29 a_n327_n194# a_207_n194# 0.02fF
C30 a_505_n140# a_n207_n140# 0.03fF
C31 a_n1217_n194# a_207_n194# 0.01fF
C32 a_683_n140# a_1395_n140# 0.03fF
C33 a_741_n194# a_563_n194# 0.10fF
C34 a_1275_n194# a_563_n194# 0.01fF
C35 a_n563_n140# a_n741_n140# 0.13fF
C36 a_n385_n140# a_n741_n140# 0.06fF
C37 a_1217_n140# a_n207_n140# 0.01fF
C38 a_149_n140# a_n207_n140# 0.06fF
C39 a_n683_n194# a_741_n194# 0.01fF
C40 a_n919_n140# a_n741_n140# 0.13fF
C41 a_n861_n194# a_n327_n194# 0.02fF
C42 a_29_n194# a_563_n194# 0.02fF
C43 a_1039_n140# a_n207_n140# 0.02fF
C44 a_327_n140# a_n29_n140# 0.06fF
C45 a_327_n140# a_861_n140# 0.04fF
C46 a_n861_n194# a_n1217_n194# 0.03fF
C47 a_741_n194# a_207_n194# 0.02fF
C48 a_n327_n194# a_1097_n194# 0.01fF
C49 a_29_n194# a_n683_n194# 0.01fF
C50 a_1275_n194# a_207_n194# 0.01fF
C51 a_n1097_n140# a_n207_n140# 0.02fF
C52 a_505_n140# a_327_n140# 0.13fF
C53 a_683_n140# a_n207_n140# 0.02fF
C54 a_n1453_n140# a_n207_n140# 0.02fF
C55 a_29_n194# a_207_n194# 0.10fF
C56 a_n149_n194# a_563_n194# 0.01fF
C57 a_n327_n194# a_n1217_n194# 0.01fF
C58 a_1217_n140# a_327_n140# 0.02fF
C59 a_n149_n194# a_n683_n194# 0.02fF
C60 a_n861_n194# a_741_n194# 0.01fF
C61 a_327_n140# a_149_n140# 0.13fF
C62 a_n29_n140# a_861_n140# 0.02fF
C63 a_n1395_n194# a_n683_n194# 0.01fF
C64 a_1039_n140# a_327_n140# 0.03fF
C65 a_n1275_n140# a_n741_n140# 0.04fF
C66 a_1097_n194# a_741_n194# 0.03fF
C67 a_505_n140# a_n29_n140# 0.04fF
C68 a_n149_n194# a_207_n194# 0.03fF
C69 a_n861_n194# a_29_n194# 0.01fF
C70 a_1275_n194# a_1097_n194# 0.10fF
C71 a_505_n140# a_861_n140# 0.06fF
C72 a_n1395_n194# a_207_n194# 0.01fF
C73 a_n563_n140# a_n207_n140# 0.06fF
C74 a_563_n194# a_385_n194# 0.10fF
C75 a_n327_n194# a_741_n194# 0.01fF
C76 a_n385_n140# a_n207_n140# 0.13fF
C77 a_327_n140# a_n1097_n140# 0.01fF
C78 a_n327_n194# a_1275_n194# 0.01fF
C79 a_327_n140# a_683_n140# 0.06fF
C80 a_n505_n194# a_563_n194# 0.01fF
C81 a_29_n194# a_1097_n194# 0.01fF
C82 a_n919_n140# a_n207_n140# 0.03fF
C83 a_1217_n140# a_n29_n140# 0.02fF
C84 a_n683_n194# a_385_n194# 0.01fF
C85 a_n29_n140# a_149_n140# 0.13fF
C86 a_1217_n140# a_861_n140# 0.06fF
C87 a_29_n194# a_n327_n194# 0.03fF
C88 a_861_n140# a_149_n140# 0.03fF
C89 a_n505_n194# a_n683_n194# 0.10fF
C90 a_1039_n140# a_n29_n140# 0.02fF
C91 a_n861_n194# a_n149_n194# 0.01fF
C92 a_29_n194# a_n1217_n194# 0.01fF
C93 a_1039_n140# a_861_n140# 0.13fF
C94 a_385_n194# a_207_n194# 0.10fF
C95 a_505_n140# a_1217_n140# 0.03fF
C96 a_n861_n194# a_n1395_n194# 0.02fF
C97 a_505_n140# a_149_n140# 0.06fF
C98 a_n505_n194# a_207_n194# 0.01fF
C99 a_n149_n194# a_1097_n194# 0.01fF
C100 a_1039_n140# a_505_n140# 0.04fF
C101 a_n29_n140# a_n1097_n140# 0.02fF
C102 a_n29_n140# a_683_n140# 0.03fF
C103 a_n1453_n140# a_n29_n140# 0.01fF
C104 a_861_n140# a_683_n140# 0.13fF
C105 a_n327_n194# a_n149_n194# 0.10fF
C106 a_1275_n194# a_741_n194# 0.02fF
C107 a_n1039_n194# a_563_n194# 0.01fF
C108 a_327_n140# a_n563_n140# 0.02fF
C109 a_1217_n140# a_149_n140# 0.02fF
C110 a_n385_n140# a_327_n140# 0.03fF
C111 a_n1395_n194# a_n327_n194# 0.01fF
C112 a_505_n140# a_n1097_n140# 0.01fF
C113 a_n149_n194# a_n1217_n194# 0.01fF
C114 a_505_n140# a_683_n140# 0.13fF
C115 a_n861_n194# a_385_n194# 0.01fF
C116 a_327_n140# a_n919_n140# 0.02fF
C117 a_1039_n140# a_1217_n140# 0.13fF
C118 a_29_n194# a_741_n194# 0.01fF
C119 a_1039_n140# a_149_n140# 0.02fF
C120 a_n1395_n194# a_n1217_n194# 0.10fF
C121 a_n1039_n194# a_n683_n194# 0.03fF
C122 a_n1275_n140# a_n207_n140# 0.02fF
C123 a_n861_n194# a_n505_n194# 0.03fF
C124 a_29_n194# a_1275_n194# 0.01fF
C125 a_919_n194# a_563_n194# 0.03fF
C126 a_1097_n194# a_385_n194# 0.01fF
C127 a_n1039_n194# a_207_n194# 0.01fF
C128 a_n505_n194# a_1097_n194# 0.01fF
C129 a_n1097_n140# a_149_n140# 0.02fF
C130 a_1217_n140# a_683_n140# 0.04fF
C131 a_149_n140# a_683_n140# 0.04fF
C132 a_n1453_n140# a_149_n140# 0.01fF
C133 a_n327_n194# a_385_n194# 0.01fF
C134 a_n683_n194# a_919_n194# 0.01fF
C135 a_n29_n140# a_n563_n140# 0.04fF
C136 a_n385_n140# a_n29_n140# 0.06fF
C137 a_n505_n194# a_n327_n194# 0.10fF
C138 a_1039_n140# a_683_n140# 0.06fF
C139 a_n149_n194# a_741_n194# 0.01fF
C140 a_n563_n140# a_861_n140# 0.01fF
C141 a_n1217_n194# a_385_n194# 0.01fF
C142 a_n385_n140# a_861_n140# 0.02fF
C143 a_1275_n194# a_n149_n194# 0.01fF
C144 a_n29_n140# a_n919_n140# 0.02fF
C145 a_n505_n194# a_n1217_n194# 0.01fF
C146 a_919_n194# a_207_n194# 0.01fF
C147 a_505_n140# a_n563_n140# 0.02fF
C148 a_505_n140# a_n385_n140# 0.02fF
C149 a_29_n194# a_n149_n194# 0.10fF
C150 a_n1453_n140# a_n1097_n140# 0.06fF
C151 a_n1039_n194# a_n861_n194# 0.10fF
C152 a_505_n140# a_n919_n140# 0.01fF
C153 a_29_n194# a_n1395_n194# 0.01fF
C154 a_n741_n140# a_n207_n140# 0.04fF
C155 a_n1275_n140# a_327_n140# 0.01fF
C156 a_n563_n140# a_149_n140# 0.03fF
C157 a_n385_n140# a_1217_n140# 0.01fF
C158 a_741_n194# a_385_n194# 0.03fF
C159 a_n385_n140# a_149_n140# 0.04fF
C160 a_1275_n194# a_385_n194# 0.01fF
C161 a_n505_n194# a_741_n194# 0.01fF
C162 a_n1039_n194# a_n327_n194# 0.01fF
C163 a_1039_n140# a_n563_n140# 0.01fF
C164 a_n919_n140# a_149_n140# 0.02fF
C165 a_1039_n140# a_n385_n140# 0.01fF
C166 a_n1395_n194# a_n149_n194# 0.01fF
C167 a_n1039_n194# a_n1217_n194# 0.10fF
C168 a_29_n194# a_385_n194# 0.03fF
C169 a_1097_n194# a_919_n194# 0.10fF
C170 a_29_n194# a_n505_n194# 0.02fF
C171 a_1395_n140# a_n207_n140# 0.01fF
C172 a_n1275_n140# a_n29_n140# 0.02fF
C173 a_n563_n140# a_n1097_n140# 0.04fF
C174 a_n385_n140# a_n1097_n140# 0.03fF
C175 a_n563_n140# a_683_n140# 0.02fF
C176 a_n1453_n140# a_n563_n140# 0.02fF
C177 a_n327_n194# a_919_n194# 0.01fF
C178 a_n385_n140# a_683_n140# 0.02fF
C179 a_n385_n140# a_n1453_n140# 0.02fF
C180 a_n1097_n140# a_n919_n140# 0.13fF
C181 a_n919_n140# a_683_n140# 0.01fF
C182 a_327_n140# a_n741_n140# 0.02fF
C183 a_n1453_n140# a_n919_n140# 0.04fF
C184 a_n149_n194# a_385_n194# 0.02fF
C185 a_n505_n194# a_n149_n194# 0.03fF
C186 a_n1395_n194# a_n505_n194# 0.01fF
C187 a_n1275_n140# a_149_n140# 0.01fF
C188 a_n1039_n194# a_29_n194# 0.01fF
C189 a_n683_n194# a_563_n194# 0.01fF
C190 a_919_n194# a_741_n194# 0.10fF
C191 a_n385_n140# a_n563_n140# 0.13fF
C192 a_327_n140# a_1395_n140# 0.02fF
C193 a_n29_n140# a_n741_n140# 0.03fF
C194 a_1275_n194# a_919_n194# 0.03fF
C195 a_861_n140# a_n741_n140# 0.01fF
C196 a_n563_n140# a_n919_n140# 0.06fF
C197 a_563_n194# a_207_n194# 0.03fF
C198 a_n385_n140# a_n919_n140# 0.04fF
C199 a_n505_n194# a_385_n194# 0.01fF
C200 a_29_n194# a_919_n194# 0.01fF
C201 a_n1275_n140# a_n1097_n140# 0.13fF
C202 a_505_n140# a_n741_n140# 0.02fF
C203 a_n1275_n140# a_n1453_n140# 0.13fF
C204 a_n683_n194# a_207_n194# 0.01fF
C205 a_n1039_n194# a_n149_n194# 0.01fF
C206 a_n1039_n194# a_n1395_n194# 0.03fF
C207 a_1395_n140# VSUBS 0.02fF
C208 a_1217_n140# VSUBS 0.02fF
C209 a_1039_n140# VSUBS 0.02fF
C210 a_861_n140# VSUBS 0.02fF
C211 a_683_n140# VSUBS 0.02fF
C212 a_505_n140# VSUBS 0.02fF
C213 a_327_n140# VSUBS 0.02fF
C214 a_149_n140# VSUBS 0.02fF
C215 a_n29_n140# VSUBS 0.02fF
C216 a_n207_n140# VSUBS 0.02fF
C217 a_n385_n140# VSUBS 0.02fF
C218 a_n563_n140# VSUBS 0.02fF
C219 a_n741_n140# VSUBS 0.02fF
C220 a_n919_n140# VSUBS 0.02fF
C221 a_n1097_n140# VSUBS 0.02fF
C222 a_n1275_n140# VSUBS 0.02fF
C223 a_n1453_n140# VSUBS 0.02fF
C224 a_1275_n194# VSUBS 0.29fF
C225 a_1097_n194# VSUBS 0.23fF
C226 a_919_n194# VSUBS 0.24fF
C227 a_741_n194# VSUBS 0.25fF
C228 a_563_n194# VSUBS 0.26fF
C229 a_385_n194# VSUBS 0.27fF
C230 a_207_n194# VSUBS 0.28fF
C231 a_29_n194# VSUBS 0.28fF
C232 a_n149_n194# VSUBS 0.29fF
C233 a_n327_n194# VSUBS 0.29fF
C234 a_n505_n194# VSUBS 0.29fF
C235 a_n683_n194# VSUBS 0.29fF
C236 a_n861_n194# VSUBS 0.29fF
C237 a_n1039_n194# VSUBS 0.29fF
C238 a_n1217_n194# VSUBS 0.29fF
C239 a_n1395_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_EE a_n352_n194# a_n60_n194# a_n644_n194# a_n936_n194#
+ a_n410_n140# a_n994_n140# a_n702_n140# a_n232_n140# a_n524_n140# a_524_n194# a_232_n194#
+ a_n816_n140# a_816_n194# a_644_n140# a_352_n140# a_936_n140# a_60_n140# a_174_n140#
+ a_466_n140# a_758_n140# a_n118_n140# VSUBS
X0 a_n232_n140# a_n352_n194# a_n410_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n524_n140# a_n644_n194# a_n702_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n816_n140# a_n936_n194# a_n994_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_352_n140# a_232_n194# a_174_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_644_n140# a_524_n194# a_466_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_936_n140# a_816_n194# a_758_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_936_n140# a_n232_n140# 0.02fF
C1 a_466_n140# a_n410_n140# 0.02fF
C2 a_174_n140# a_n232_n140# 0.05fF
C3 a_644_n140# a_n994_n140# 0.01fF
C4 a_466_n140# a_n232_n140# 0.03fF
C5 a_n644_n194# a_n60_n194# 0.02fF
C6 a_936_n140# a_n702_n140# 0.01fF
C7 a_n118_n140# a_n410_n140# 0.07fF
C8 a_758_n140# a_n410_n140# 0.02fF
C9 a_174_n140# a_n702_n140# 0.02fF
C10 a_60_n140# a_n410_n140# 0.04fF
C11 a_n118_n140# a_n232_n140# 0.25fF
C12 a_n60_n194# a_232_n194# 0.04fF
C13 a_758_n140# a_n232_n140# 0.02fF
C14 a_466_n140# a_n702_n140# 0.02fF
C15 a_60_n140# a_n232_n140# 0.07fF
C16 a_174_n140# a_n994_n140# 0.02fF
C17 a_n352_n194# a_524_n194# 0.01fF
C18 a_n410_n140# a_352_n140# 0.03fF
C19 a_n118_n140# a_n702_n140# 0.03fF
C20 a_466_n140# a_n994_n140# 0.01fF
C21 a_758_n140# a_n702_n140# 0.01fF
C22 a_n410_n140# a_n816_n140# 0.05fF
C23 a_352_n140# a_n232_n140# 0.03fF
C24 a_60_n140# a_n702_n140# 0.03fF
C25 a_n232_n140# a_n816_n140# 0.03fF
C26 a_n644_n194# a_816_n194# 0.01fF
C27 a_n118_n140# a_n994_n140# 0.02fF
C28 a_644_n140# a_936_n140# 0.07fF
C29 a_352_n140# a_n702_n140# 0.02fF
C30 a_60_n140# a_n994_n140# 0.02fF
C31 a_644_n140# a_174_n140# 0.04fF
C32 a_816_n194# a_232_n194# 0.02fF
C33 a_n816_n140# a_n702_n140# 0.25fF
C34 a_466_n140# a_644_n140# 0.13fF
C35 a_n936_n194# a_524_n194# 0.01fF
C36 a_352_n140# a_n994_n140# 0.01fF
C37 a_n816_n140# a_n994_n140# 0.13fF
C38 a_n118_n140# a_644_n140# 0.03fF
C39 a_644_n140# a_758_n140# 0.25fF
C40 a_936_n140# a_174_n140# 0.03fF
C41 a_n524_n140# a_n410_n140# 0.25fF
C42 a_60_n140# a_644_n140# 0.03fF
C43 a_n644_n194# a_232_n194# 0.01fF
C44 a_466_n140# a_936_n140# 0.04fF
C45 a_n524_n140# a_n232_n140# 0.07fF
C46 a_466_n140# a_174_n140# 0.07fF
C47 a_n352_n194# a_n936_n194# 0.02fF
C48 a_524_n194# a_n60_n194# 0.02fF
C49 a_644_n140# a_352_n140# 0.07fF
C50 a_n118_n140# a_936_n140# 0.02fF
C51 a_936_n140# a_758_n140# 0.13fF
C52 a_644_n140# a_n816_n140# 0.01fF
C53 a_n118_n140# a_174_n140# 0.07fF
C54 a_n524_n140# a_n702_n140# 0.13fF
C55 a_174_n140# a_758_n140# 0.03fF
C56 a_60_n140# a_936_n140# 0.02fF
C57 a_60_n140# a_174_n140# 0.25fF
C58 a_466_n140# a_n118_n140# 0.03fF
C59 a_466_n140# a_758_n140# 0.07fF
C60 a_60_n140# a_466_n140# 0.05fF
C61 a_n524_n140# a_n994_n140# 0.04fF
C62 a_936_n140# a_352_n140# 0.03fF
C63 a_n352_n194# a_n60_n194# 0.04fF
C64 a_174_n140# a_352_n140# 0.13fF
C65 a_n118_n140# a_758_n140# 0.02fF
C66 a_174_n140# a_n816_n140# 0.02fF
C67 a_466_n140# a_352_n140# 0.25fF
C68 a_60_n140# a_n118_n140# 0.13fF
C69 a_60_n140# a_758_n140# 0.03fF
C70 a_524_n194# a_816_n194# 0.04fF
C71 a_466_n140# a_n816_n140# 0.01fF
C72 a_n118_n140# a_352_n140# 0.04fF
C73 a_758_n140# a_352_n140# 0.05fF
C74 a_644_n140# a_n524_n140# 0.02fF
C75 a_60_n140# a_352_n140# 0.07fF
C76 a_n118_n140# a_n816_n140# 0.03fF
C77 a_758_n140# a_n816_n140# 0.01fF
C78 a_n410_n140# a_n232_n140# 0.13fF
C79 a_60_n140# a_n816_n140# 0.02fF
C80 a_n352_n194# a_816_n194# 0.01fF
C81 a_n936_n194# a_n60_n194# 0.01fF
C82 a_n644_n194# a_524_n194# 0.01fF
C83 a_n410_n140# a_n702_n140# 0.07fF
C84 a_352_n140# a_n816_n140# 0.02fF
C85 a_936_n140# a_n524_n140# 0.01fF
C86 a_174_n140# a_n524_n140# 0.03fF
C87 a_524_n194# a_232_n194# 0.04fF
C88 a_n232_n140# a_n702_n140# 0.04fF
C89 a_466_n140# a_n524_n140# 0.02fF
C90 a_n410_n140# a_n994_n140# 0.03fF
C91 a_n352_n194# a_n644_n194# 0.04fF
C92 a_n232_n140# a_n994_n140# 0.03fF
C93 a_n118_n140# a_n524_n140# 0.05fF
C94 a_n524_n140# a_758_n140# 0.01fF
C95 a_n352_n194# a_232_n194# 0.02fF
C96 a_60_n140# a_n524_n140# 0.03fF
C97 a_n994_n140# a_n702_n140# 0.07fF
C98 a_644_n140# a_n410_n140# 0.02fF
C99 a_n524_n140# a_352_n140# 0.02fF
C100 a_n524_n140# a_n816_n140# 0.07fF
C101 a_644_n140# a_n232_n140# 0.02fF
C102 a_n644_n194# a_n936_n194# 0.04fF
C103 a_816_n194# a_n60_n194# 0.01fF
C104 a_936_n140# a_n410_n140# 0.01fF
C105 a_644_n140# a_n702_n140# 0.01fF
C106 a_174_n140# a_n410_n140# 0.03fF
C107 a_n936_n194# a_232_n194# 0.01fF
C108 a_936_n140# VSUBS 0.02fF
C109 a_758_n140# VSUBS 0.02fF
C110 a_644_n140# VSUBS 0.02fF
C111 a_466_n140# VSUBS 0.02fF
C112 a_352_n140# VSUBS 0.02fF
C113 a_174_n140# VSUBS 0.02fF
C114 a_60_n140# VSUBS 0.02fF
C115 a_n118_n140# VSUBS 0.02fF
C116 a_n232_n140# VSUBS 0.02fF
C117 a_n410_n140# VSUBS 0.02fF
C118 a_n524_n140# VSUBS 0.02fF
C119 a_n702_n140# VSUBS 0.02fF
C120 a_n816_n140# VSUBS 0.02fF
C121 a_n994_n140# VSUBS 0.02fF
C122 a_816_n194# VSUBS 0.29fF
C123 a_524_n194# VSUBS 0.24fF
C124 a_232_n194# VSUBS 0.26fF
C125 a_n60_n194# VSUBS 0.27fF
C126 a_n352_n194# VSUBS 0.29fF
C127 a_n644_n194# VSUBS 0.29fF
C128 a_n936_n194# VSUBS 0.35fF
.ends

.subckt unit_cap_mim_m3m4 c1_n530_n480# m3_n630_n580# VSUBS
X0 c1_n530_n480# m3_n630_n580# sky130_fd_pr__cap_mim_m3_1 l=4.8e+06u w=4.8e+06u
C0 m3_n630_n580# c1_n530_n480# 2.88fF
C1 m3_n630_n580# VSUBS 1.37fF
.ends

.subckt sc_cmfb unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_26/c1_n530_n480#
+ unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580#
+ unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_20/m3_n630_n580#
+ unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480#
+ unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580#
+ unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580#
+ unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ transmission_gate_4/out unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480#
+ unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480#
+ unit_cap_mim_m3m4_34/c1_n530_n480# bias_a unit_cap_mim_m3m4_24/m3_n630_n580# p2_b
+ unit_cap_mim_m3m4_25/c1_n530_n480# p1 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_16/c1_n530_n480#
+ unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_28/c1_n530_n480# p2 VDD unit_cap_mim_m3m4_32/c1_n530_n480#
+ unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580# transmission_gate_3/out
+ transmission_gate_6/in cmc unit_cap_mim_m3m4_19/c1_n530_n480# on transmission_gate_8/in
+ unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_7/in
+ cm transmission_gate_9/in unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480#
+ p1_b VSS op
Xtransmission_gate_10 p1 VDD transmission_gate_10/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_3/out on VSS p1_b transmission_gate
Xtransmission_gate_11 p1 VDD transmission_gate_11/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_4/out op VSS p1_b transmission_gate
Xtransmission_gate_0 p1 VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ cm transmission_gate_7/in VSS p1_b transmission_gate
Xtransmission_gate_1 p1 VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ cm transmission_gate_6/in VSS p1_b transmission_gate
Xtransmission_gate_2 p1 VDD transmission_gate_2/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ bias_a transmission_gate_8/in VSS p1_b transmission_gate
Xtransmission_gate_3 p2 VDD transmission_gate_3/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ cm transmission_gate_3/out VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_0 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xtransmission_gate_4 p2 VDD transmission_gate_4/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ cm transmission_gate_4/out VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_1 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_5 p2 VDD transmission_gate_5/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ bias_a transmission_gate_9/in VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_2 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_30 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_6 p2 VDD transmission_gate_6/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_6/in op VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_20 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_20/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_3 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_31 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xtransmission_gate_7 p2 VDD transmission_gate_7/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_7/in on VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_10 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_21 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_21/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_4 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_32 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_12 transmission_gate_4/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_11 on cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_8 p2 VDD transmission_gate_8/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_8/in cmc VSS p2_b transmission_gate
Xunit_cap_mim_m3m4_5 transmission_gate_6/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_22 unit_cap_mim_m3m4_22/c1_n530_n480# unit_cap_mim_m3m4_22/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_23 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_34 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_33 unit_cap_mim_m3m4_33/c1_n530_n480# unit_cap_mim_m3m4_33/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_24 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_13 on cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_6 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_7 op cmc VSS unit_cap_mim_m3m4
Xtransmission_gate_9 p1 VDD transmission_gate_9/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_9/in cmc VSS p1_b transmission_gate
Xunit_cap_mim_m3m4_35 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_25 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_25/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_14 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_8 op cmc VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_26 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_26/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_15 transmission_gate_7/in transmission_gate_8/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_9 transmission_gate_3/out transmission_gate_9/in VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_27 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_27/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_16 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_16/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_28 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_28/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_17 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_17/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_29 unit_cap_mim_m3m4_29/c1_n530_n480# unit_cap_mim_m3m4_29/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_18 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_18/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
Xunit_cap_mim_m3m4_19 unit_cap_mim_m3m4_19/c1_n530_n480# unit_cap_mim_m3m4_19/m3_n630_n580#
+ VSS unit_cap_mim_m3m4
C0 transmission_gate_6/in p2_b 0.02fF
C1 p2_b unit_cap_mim_m3m4_17/m3_n630_n580# -0.46fF
C2 p2_b unit_cap_mim_m3m4_16/c1_n530_n480# -0.07fF
C3 p1 p2 0.01fF
C4 bias_a VDD -0.01fF
C5 op unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C6 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C7 cmc transmission_gate_9/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# 0.00fF
C8 on p2 0.28fF
C9 transmission_gate_4/out VDD 0.20fF
C10 cm unit_cap_mim_m3m4_18/c1_n530_n480# -0.22fF
C11 transmission_gate_8/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.17fF
C12 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_24/m3_n630_n580# -0.24fF
C13 transmission_gate_3/out unit_cap_mim_m3m4_23/m3_n630_n580# 0.61fF
C14 transmission_gate_7/in transmission_gate_9/in 0.02fF
C15 transmission_gate_6/in op 0.68fF
C16 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.17fF
C17 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_25/m3_n630_n580# 0.17fF
C18 cmc unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C19 p1 transmission_gate_9/in 0.01fF
C20 p1_b cm 0.27fF
C21 transmission_gate_8/in unit_cap_mim_m3m4_21/m3_n630_n580# 0.59fF
C22 on transmission_gate_9/in 0.79fF
C23 transmission_gate_8/in cmc 8.00fF
C24 transmission_gate_4/out unit_cap_mim_m3m4_16/m3_n630_n580# 0.62fF
C25 transmission_gate_7/in unit_cap_mim_m3m4_19/m3_n630_n580# 0.63fF
C26 unit_cap_mim_m3m4_18/c1_n530_n480# unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C27 transmission_gate_6/in VDD 0.31fF
C28 VDD unit_cap_mim_m3m4_17/m3_n630_n580# -0.16fF
C29 VDD unit_cap_mim_m3m4_16/c1_n530_n480# -0.06fF
C30 op unit_cap_mim_m3m4_30/m3_n630_n580# 0.31fF
C31 p1_b transmission_gate_3/out 0.08fF
C32 p1 unit_cap_mim_m3m4_19/m3_n630_n580# -0.29fF
C33 p1_b p2_b 0.01fF
C34 p1_b unit_cap_mim_m3m4_22/m3_n630_n580# -0.63fF
C35 VDD unit_cap_mim_m3m4_30/m3_n630_n580# 0.28fF
C36 p1_b unit_cap_mim_m3m4_19/c1_n530_n480# 0.07fF
C37 transmission_gate_7/in cmc 0.07fF
C38 p2 transmission_gate_9/in 0.02fF
C39 VDD unit_cap_mim_m3m4_23/m3_n630_n580# 0.33fF
C40 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_17/m3_n630_n580# 0.10fF
C41 unit_cap_mim_m3m4_16/m3_n630_n580# unit_cap_mim_m3m4_16/c1_n530_n480# -0.35fF
C42 on unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C43 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_26/c1_n530_n480# -0.20fF
C44 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_32/m3_n630_n580# -0.15fF
C45 transmission_gate_8/in unit_cap_mim_m3m4_34/m3_n630_n580# 0.56fF
C46 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.12fF
C47 bias_a transmission_gate_8/in 0.04fF
C48 p1 cmc 0.03fF
C49 VDD unit_cap_mim_m3m4_18/c1_n530_n480# -0.06fF
C50 p2_b unit_cap_mim_m3m4_24/c1_n530_n480# -0.07fF
C51 p1_b op 0.10fF
C52 transmission_gate_8/in transmission_gate_4/out 0.26fF
C53 on cmc 2.26fF
C54 cmc unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C55 bias_a unit_cap_mim_m3m4_35/c1_n530_n480# -0.22fF
C56 p2_b unit_cap_mim_m3m4_24/m3_n630_n580# -0.55fF
C57 p1_b VDD 0.07fF
C58 unit_cap_mim_m3m4_20/m3_n630_n580# p2_b -0.65fF
C59 bias_a transmission_gate_7/in 0.09fF
C60 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C61 transmission_gate_6/in unit_cap_mim_m3m4_18/m3_n630_n580# 0.62fF
C62 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C63 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_18/m3_n630_n580# 0.17fF
C64 unit_cap_mim_m3m4_17/m3_n630_n580# unit_cap_mim_m3m4_17/c1_n530_n480# -0.15fF
C65 unit_cap_mim_m3m4_16/c1_n530_n480# unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C66 unit_cap_mim_m3m4_21/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C67 transmission_gate_4/out transmission_gate_7/in 0.61fF
C68 unit_cap_mim_m3m4_21/m3_n630_n580# p2 -1.16fF
C69 p2 cmc 0.61fF
C70 transmission_gate_8/in transmission_gate_6/in -0.10fF
C71 bias_a p1 0.06fF
C72 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_25/c1_n530_n480# -0.19fF
C73 VDD unit_cap_mim_m3m4_35/m3_n630_n580# -0.40fF
C74 unit_cap_mim_m3m4_26/c1_n530_n480# unit_cap_mim_m3m4_27/c1_n530_n480# 0.06fF
C75 transmission_gate_4/out p1 0.01fF
C76 op unit_cap_mim_m3m4_27/m3_n630_n580# 0.28fF
C77 VDD unit_cap_mim_m3m4_24/c1_n530_n480# -0.06fF
C78 unit_cap_mim_m3m4_30/c1_n530_n480# op 0.05fF
C79 on transmission_gate_4/out 3.14fF
C80 transmission_gate_3/out cm 0.19fF
C81 p2_b unit_cap_mim_m3m4_29/m3_n630_n580# -0.58fF
C82 cm p2_b 0.16fF
C83 transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# cm 0.00fF
C84 VDD unit_cap_mim_m3m4_24/m3_n630_n580# -0.50fF
C85 transmission_gate_6/in transmission_gate_7/in 0.44fF
C86 unit_cap_mim_m3m4_18/m3_n630_n580# unit_cap_mim_m3m4_18/c1_n530_n480# -0.15fF
C87 unit_cap_mim_m3m4_17/c1_n530_n480# unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C88 transmission_gate_9/in cmc 6.71fF
C89 cm unit_cap_mim_m3m4_19/c1_n530_n480# -0.22fF
C90 VDD unit_cap_mim_m3m4_20/m3_n630_n580# 0.33fF
C91 bias_a p2 0.05fF
C92 transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# transmission_gate_3/out 0.00fF
C93 op unit_cap_mim_m3m4_31/m3_n630_n580# 0.02fF
C94 unit_cap_mim_m3m4_33/m3_n630_n580# cmc 0.10fF
C95 transmission_gate_4/out p2 0.02fF
C96 op unit_cap_mim_m3m4_29/m3_n630_n580# 0.42fF
C97 op unit_cap_mim_m3m4_28/c1_n530_n480# 0.17fF
C98 on transmission_gate_6/in 0.40fF
C99 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_31/m3_n630_n580# 0.17fF
C100 p1_b unit_cap_mim_m3m4_18/m3_n630_n580# -0.41fF
C101 unit_cap_mim_m3m4_24/m3_n630_n580# unit_cap_mim_m3m4_16/m3_n630_n580# 0.12fF
C102 transmission_gate_8/in p1_b 0.02fF
C103 p1 unit_cap_mim_m3m4_30/m3_n630_n580# -0.67fF
C104 on unit_cap_mim_m3m4_21/c1_n530_n480# 0.06fF
C105 transmission_gate_3/out op 0.42fF
C106 VDD unit_cap_mim_m3m4_29/m3_n630_n580# 0.35fF
C107 bias_a transmission_gate_9/in 0.02fF
C108 p1 unit_cap_mim_m3m4_23/m3_n630_n580# -0.71fF
C109 VDD cm 0.00fF
C110 p1_b unit_cap_mim_m3m4_35/c1_n530_n480# -0.07fF
C111 op p2_b 0.17fF
C112 transmission_gate_4/out transmission_gate_9/in 3.03fF
C113 transmission_gate_6/in p2 0.00fF
C114 unit_cap_mim_m3m4_21/m3_n630_n580# cmc 0.58fF
C115 p1 unit_cap_mim_m3m4_18/c1_n530_n480# -0.30fF
C116 p2 unit_cap_mim_m3m4_17/m3_n630_n580# -0.56fF
C117 p2 unit_cap_mim_m3m4_16/c1_n530_n480# -0.30fF
C118 on unit_cap_mim_m3m4_23/m3_n630_n580# 0.02fF
C119 transmission_gate_8/in unit_cap_mim_m3m4_35/m3_n630_n580# 0.58fF
C120 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C121 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_20/c1_n530_n480# -0.20fF
C122 transmission_gate_3/out VDD 0.27fF
C123 on unit_cap_mim_m3m4_18/c1_n530_n480# 0.06fF
C124 p1_b transmission_gate_7/in 0.03fF
C125 transmission_gate_4/out unit_cap_mim_m3m4_31/c1_n530_n480# 0.06fF
C126 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_35/m3_n630_n580# -0.33fF
C127 VDD p2_b 0.27fF
C128 unit_cap_mim_m3m4_21/c1_n530_n480# p2 0.03fF
C129 on unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C130 VDD unit_cap_mim_m3m4_22/m3_n630_n580# 0.33fF
C131 transmission_gate_6/in unit_cap_mim_m3m4_28/m3_n630_n580# -1.01fF
C132 transmission_gate_6/in unit_cap_mim_m3m4_27/c1_n530_n480# -0.04fF
C133 transmission_gate_4/out unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C134 p1_b p1 2.54fF
C135 cm unit_cap_mim_m3m4_16/m3_n630_n580# 0.36fF
C136 VDD unit_cap_mim_m3m4_19/c1_n530_n480# -0.06fF
C137 unit_cap_mim_m3m4_33/m3_n630_n580# unit_cap_mim_m3m4_33/c1_n530_n480# -0.20fF
C138 transmission_gate_6/in transmission_gate_9/in 0.09fF
C139 on p1_b 0.12fF
C140 transmission_gate_8/in unit_cap_mim_m3m4_20/m3_n630_n580# 0.17fF
C141 p1 unit_cap_mim_m3m4_35/m3_n630_n580# -0.25fF
C142 VDD op 0.19fF
C143 p2_b unit_cap_mim_m3m4_16/m3_n630_n580# -0.37fF
C144 transmission_gate_4/out cmc 0.10fF
C145 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_35/c1_n530_n480# 0.06fF
C146 p1_b p2 0.29fF
C147 unit_cap_mim_m3m4_23/m3_n630_n580# transmission_gate_9/in 0.17fF
C148 cm unit_cap_mim_m3m4_18/m3_n630_n580# 0.39fF
C149 cm unit_cap_mim_m3m4_17/c1_n530_n480# -0.22fF
C150 transmission_gate_7/in unit_cap_mim_m3m4_20/m3_n630_n580# 0.64fF
C151 transmission_gate_8/in cm 0.03fF
C152 unit_cap_mim_m3m4_25/m3_n630_n580# unit_cap_mim_m3m4_26/m3_n630_n580# 0.12fF
C153 unit_cap_mim_m3m4_22/m3_n630_n580# unit_cap_mim_m3m4_22/c1_n530_n480# -0.20fF
C154 transmission_gate_7/in unit_cap_mim_m3m4_34/c1_n530_n480# 0.06fF
C155 transmission_gate_3/out unit_cap_mim_m3m4_17/c1_n530_n480# -0.03fF
C156 unit_cap_mim_m3m4_26/m3_n630_n580# unit_cap_mim_m3m4_27/m3_n630_n580# 0.12fF
C157 transmission_gate_6/in cmc 0.92fF
C158 cmc unit_cap_mim_m3m4_17/m3_n630_n580# 0.17fF
C159 on unit_cap_mim_m3m4_20/m3_n630_n580# 0.40fF
C160 p2_b unit_cap_mim_m3m4_17/c1_n530_n480# -0.07fF
C161 transmission_gate_8/in transmission_gate_3/out 0.24fF
C162 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_23/m3_n630_n580# -0.20fF
C163 unit_cap_mim_m3m4_24/c1_n530_n480# p2 -0.30fF
C164 bias_a transmission_gate_4/out 0.09fF
C165 transmission_gate_8/in p2_b -0.02fF
C166 p1_b transmission_gate_9/in 0.00fF
C167 VDD unit_cap_mim_m3m4_16/m3_n630_n580# -0.43fF
C168 transmission_gate_7/in unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C169 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_32/c1_n530_n480# 0.06fF
C170 op unit_cap_mim_m3m4_22/c1_n530_n480# 0.07fF
C171 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_21/c1_n530_n480# -0.20fF
C172 transmission_gate_7/in cm 0.11fF
C173 p2 unit_cap_mim_m3m4_24/m3_n630_n580# -0.47fF
C174 cm p1 0.12fF
C175 unit_cap_mim_m3m4_20/m3_n630_n580# p2 -0.71fF
C176 op unit_cap_mim_m3m4_17/c1_n530_n480# 0.06fF
C177 transmission_gate_3/out transmission_gate_7/in 0.28fF
C178 unit_cap_mim_m3m4_35/c1_n530_n480# unit_cap_mim_m3m4_19/c1_n530_n480# 0.06fF
C179 p1_b unit_cap_mim_m3m4_19/m3_n630_n580# -0.65fF
C180 p1_b unit_cap_mim_m3m4_23/c1_n530_n480# 0.13fF
C181 unit_cap_mim_m3m4_24/c1_n530_n480# transmission_gate_9/in -0.01fF
C182 transmission_gate_8/in op 0.88fF
C183 transmission_gate_7/in p2_b 0.00fF
C184 bias_a transmission_gate_6/in 0.05fF
C185 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_28/m3_n630_n580# 0.17fF
C186 unit_cap_mim_m3m4_27/m3_n630_n580# unit_cap_mim_m3m4_27/c1_n530_n480# -0.13fF
C187 transmission_gate_3/out p1 -0.00fF
C188 transmission_gate_4/out transmission_gate_6/in 0.46fF
C189 transmission_gate_4/out unit_cap_mim_m3m4_16/c1_n530_n480# 0.03fF
C190 transmission_gate_7/in unit_cap_mim_m3m4_19/c1_n530_n480# 0.03fF
C191 VDD unit_cap_mim_m3m4_18/m3_n630_n580# -0.26fF
C192 VDD unit_cap_mim_m3m4_17/c1_n530_n480# -0.06fF
C193 transmission_gate_9/in unit_cap_mim_m3m4_25/m3_n630_n580# 0.43fF
C194 on transmission_gate_3/out 0.48fF
C195 unit_cap_mim_m3m4_35/m3_n630_n580# unit_cap_mim_m3m4_19/m3_n630_n580# 0.10fF
C196 p1 unit_cap_mim_m3m4_22/m3_n630_n580# -0.76fF
C197 unit_cap_mim_m3m4_24/m3_n630_n580# transmission_gate_9/in 0.58fF
C198 transmission_gate_8/in VDD 0.21fF
C199 on p2_b 0.11fF
C200 p1_b cmc 0.31fF
C201 p2 unit_cap_mim_m3m4_29/m3_n630_n580# -0.78fF
C202 p1 unit_cap_mim_m3m4_19/c1_n530_n480# -0.30fF
C203 cm p2 0.21fF
C204 transmission_gate_4/out unit_cap_mim_m3m4_30/m3_n630_n580# 0.57fF
C205 transmission_gate_7/in op 2.64fF
C206 VDD unit_cap_mim_m3m4_35/c1_n530_n480# -0.06fF
C207 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C208 p1 op 0.10fF
C209 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_29/m3_n630_n580# 0.17fF
C210 unit_cap_mim_m3m4_28/m3_n630_n580# unit_cap_mim_m3m4_28/c1_n530_n480# -0.17fF
C211 transmission_gate_3/out p2 0.02fF
C212 unit_cap_mim_m3m4_27/c1_n530_n480# unit_cap_mim_m3m4_28/c1_n530_n480# 0.06fF
C213 VDD transmission_gate_7/in 0.25fF
C214 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C215 on op 1.88fF
C216 unit_cap_mim_m3m4_31/m3_n630_n580# transmission_gate_9/in 0.10fF
C217 p2_b p2 2.48fF
C218 transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# p2 0.00fF
C219 cm transmission_gate_9/in 0.04fF
C220 VDD p1 0.08fF
C221 bias_a p1_b 0.04fF
C222 transmission_gate_8/in transmission_gate_9/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# 0.00fF
C223 unit_cap_mim_m3m4_31/c1_n530_n480# unit_cap_mim_m3m4_31/m3_n630_n580# -0.49fF
C224 cmc unit_cap_mim_m3m4_27/m3_n630_n580# 0.12fF
C225 on VDD 0.45fF
C226 p1_b transmission_gate_4/out -0.01fF
C227 unit_cap_mim_m3m4_32/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C228 unit_cap_mim_m3m4_20/m3_n630_n580# unit_cap_mim_m3m4_21/m3_n630_n580# 0.10fF
C229 transmission_gate_3/out transmission_gate_9/in 2.49fF
C230 op p2 0.04fF
C231 transmission_gate_6/in unit_cap_mim_m3m4_18/c1_n530_n480# -0.03fF
C232 unit_cap_mim_m3m4_29/m3_n630_n580# unit_cap_mim_m3m4_29/c1_n530_n480# -0.13fF
C233 unit_cap_mim_m3m4_28/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C234 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_35/m3_n630_n580# 0.17fF
C235 bias_a unit_cap_mim_m3m4_35/m3_n630_n580# 0.33fF
C236 p2_b transmission_gate_9/in 0.03fF
C237 cm unit_cap_mim_m3m4_19/m3_n630_n580# 0.38fF
C238 unit_cap_mim_m3m4_22/m3_n630_n580# transmission_gate_9/in 0.59fF
C239 bias_a unit_cap_mim_m3m4_24/c1_n530_n480# -0.22fF
C240 unit_cap_mim_m3m4_30/m3_n630_n580# unit_cap_mim_m3m4_23/m3_n630_n580# 0.10fF
C241 op unit_cap_mim_m3m4_28/m3_n630_n580# 0.66fF
C242 op unit_cap_mim_m3m4_27/c1_n530_n480# -0.09fF
C243 VDD p2 0.15fF
C244 transmission_gate_7/in unit_cap_mim_m3m4_20/c1_n530_n480# 0.07fF
C245 p1_b transmission_gate_6/in 0.04fF
C246 bias_a unit_cap_mim_m3m4_24/m3_n630_n580# 0.35fF
C247 transmission_gate_8/in unit_cap_mim_m3m4_35/c1_n530_n480# -0.01fF
C248 op transmission_gate_9/in 0.68fF
C249 unit_cap_mim_m3m4_19/m3_n630_n580# unit_cap_mim_m3m4_19/c1_n530_n480# -0.34fF
C250 p1_b unit_cap_mim_m3m4_30/m3_n630_n580# -0.72fF
C251 transmission_gate_3/out cmc 0.79fF
C252 unit_cap_mim_m3m4_34/m3_n630_n580# unit_cap_mim_m3m4_34/c1_n530_n480# -0.19fF
C253 unit_cap_mim_m3m4_31/c1_n530_n480# op 0.05fF
C254 transmission_gate_8/in transmission_gate_7/in -0.06fF
C255 p1 unit_cap_mim_m3m4_18/m3_n630_n580# -0.55fF
C256 p2 unit_cap_mim_m3m4_16/m3_n630_n580# -0.29fF
C257 unit_cap_mim_m3m4_24/c1_n530_n480# unit_cap_mim_m3m4_16/c1_n530_n480# 0.06fF
C258 VDD transmission_gate_9/in 0.21fF
C259 p2_b cmc 0.03fF
C260 unit_cap_mim_m3m4_21/m3_n630_n580# p2_b -0.72fF
C261 unit_cap_mim_m3m4_32/m3_n630_n580# unit_cap_mim_m3m4_33/m3_n630_n580# 0.12fF
C262 p1_b unit_cap_mim_m3m4_23/m3_n630_n580# -1.03fF
C263 unit_cap_mim_m3m4_21/m3_n630_n580# unit_cap_mim_m3m4_22/m3_n630_n580# 0.17fF
C264 unit_cap_mim_m3m4_22/m3_n630_n580# cmc 0.60fF
C265 op unit_cap_mim_m3m4_23/c1_n530_n480# 0.13fF
C266 transmission_gate_8/in p1 0.02fF
C267 p1_b unit_cap_mim_m3m4_18/c1_n530_n480# -0.07fF
C268 p2 transmission_gate_9/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# 0.00fF
C269 transmission_gate_4/out unit_cap_mim_m3m4_31/m3_n630_n580# 0.53fF
C270 transmission_gate_8/in on 0.83fF
C271 unit_cap_mim_m3m4_25/c1_n530_n480# unit_cap_mim_m3m4_26/c1_n530_n480# 0.06fF
C272 unit_cap_mim_m3m4_34/c1_n530_n480# unit_cap_mim_m3m4_33/c1_n530_n480# 0.06fF
C273 transmission_gate_6/in unit_cap_mim_m3m4_27/m3_n630_n580# 0.21fF
C274 bias_a cm 0.91fF
C275 p1 unit_cap_mim_m3m4_35/c1_n530_n480# -0.30fF
C276 VDD unit_cap_mim_m3m4_19/m3_n630_n580# -0.52fF
C277 transmission_gate_4/out cm 0.08fF
C278 op cmc 4.31fF
C279 transmission_gate_9/in unit_cap_mim_m3m4_16/m3_n630_n580# 0.17fF
C280 bias_a transmission_gate_3/out 0.05fF
C281 transmission_gate_7/in p1 0.02fF
C282 p2 unit_cap_mim_m3m4_17/c1_n530_n480# -0.25fF
C283 unit_cap_mim_m3m4_32/m3_n630_n580# cmc 0.10fF
C284 transmission_gate_3/out transmission_gate_4/out 0.37fF
C285 bias_a p2_b 0.06fF
C286 unit_cap_mim_m3m4_30/c1_n530_n480# unit_cap_mim_m3m4_30/m3_n630_n580# -0.13fF
C287 on transmission_gate_7/in 3.18fF
C288 transmission_gate_8/in p2 -0.01fF
C289 VDD unit_cap_mim_m3m4_21/m3_n630_n580# 0.33fF
C290 VDD cmc 0.66fF
C291 transmission_gate_4/out p2_b 0.03fF
C292 p1_b unit_cap_mim_m3m4_35/m3_n630_n580# -0.40fF
C293 transmission_gate_6/in unit_cap_mim_m3m4_29/m3_n630_n580# 0.63fF
C294 transmission_gate_6/in unit_cap_mim_m3m4_28/c1_n530_n480# -0.32fF
C295 on p1 0.22fF
C296 transmission_gate_6/in cm 0.19fF
C297 cm unit_cap_mim_m3m4_17/m3_n630_n580# 0.41fF
C298 cm unit_cap_mim_m3m4_16/c1_n530_n480# -0.22fF
C299 transmission_gate_8/in unit_cap_mim_m3m4_28/m3_n630_n580# 0.12fF
C300 unit_cap_mim_m3m4_31/m3_n630_n580# unit_cap_mim_m3m4_30/m3_n630_n580# 0.17fF
C301 transmission_gate_7/in p2 -0.01fF
C302 transmission_gate_3/out transmission_gate_6/in 0.76fF
C303 transmission_gate_3/out unit_cap_mim_m3m4_17/m3_n630_n580# 0.62fF
C304 unit_cap_mim_m3m4_20/c1_n530_n480# unit_cap_mim_m3m4_29/c1_n530_n480# 0.06fF
C305 transmission_gate_4/out unit_cap_mim_m3m4_25/c1_n530_n480# 0.06fF
C306 transmission_gate_4/out op 1.08fF
C307 transmission_gate_8/in transmission_gate_9/in 3.34fF
C308 unit_cap_mim_m3m4_23/c1_n530_n480# unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C309 unit_cap_mim_m3m4_19/c1_n530_n480# VSS -0.06fF
C310 unit_cap_mim_m3m4_19/m3_n630_n580# VSS 0.87fF
C311 unit_cap_mim_m3m4_18/c1_n530_n480# VSS -0.06fF
C312 unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.14fF
C313 unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.64fF
C314 unit_cap_mim_m3m4_17/c1_n530_n480# VSS -0.06fF
C315 unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.05fF
C316 unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C317 unit_cap_mim_m3m4_16/c1_n530_n480# VSS -0.06fF
C318 unit_cap_mim_m3m4_16/m3_n630_n580# VSS 0.87fF
C319 unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C320 unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C321 unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C322 unit_cap_mim_m3m4_35/c1_n530_n480# VSS -0.06fF
C323 unit_cap_mim_m3m4_35/m3_n630_n580# VSS 0.94fF
C324 cmc VSS -12.07fF
C325 transmission_gate_9/in VSS -27.53fF
C326 unit_cap_mim_m3m4_24/c1_n530_n480# VSS -0.06fF
C327 unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.10fF
C328 unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C329 unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C330 unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.62fF
C331 unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.64fF
C332 p2 VSS 9.29fF
C333 p2_b VSS 1.84fF
C334 unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C335 unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.63fF
C336 unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C337 unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.62fF
C338 unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.61fF
C339 transmission_gate_8/in VSS -0.19fF
C340 bias_a VSS 7.51fF
C341 transmission_gate_6/in VSS 2.86fF
C342 transmission_gate_7/in VSS 2.35fF
C343 cm VSS 0.43fF
C344 p1 VSS 10.10fF
C345 op VSS 11.93fF
C346 transmission_gate_4/out VSS 1.26fF
C347 p1_b VSS 2.50fF
C348 VDD VSS 16.22fF
C349 on VSS -9.15fF
C350 transmission_gate_3/out VSS -4.23fF
.ends

.subckt ota_w_test sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# m1_12118_n9704# m1_12410_n9718#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# m1_11356_n10481# m1_11063_n10490# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# m1_11940_n10482# m1_12232_n10488# sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580#
+ m1_11825_n9711# m1_11534_n9706# m1_11242_n9716# m1_n6302_n3889# on sc_cmfb_0/transmission_gate_8/in
+ sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# p2_b m1_11648_n10486# sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_6/in ip sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# m1_2462_n3318# m1_n208_n2883# cm in
+ m1_2463_n5585# sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# m1_n1659_n11581# sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580#
+ m1_6690_n8907# sc_cmfb_0/transmission_gate_9/in p1_b sc_cmfb_0/transmission_gate_4/out
+ m1_n2176_n12171# i_bias sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ bias_b sc_cmfb_0/transmission_gate_7/in VDD bias_a m1_1038_n2886# op p2 VSS sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580#
+ m1_n5574_n13620# m1_n947_n12836# p1 cmc bias_c bias_d
Xsky130_fd_pr__pfet_01v8_lvt_II_2 m1_n6302_n3889# bias_b m1_n6302_n3889# bias_b VDD
+ m1_n6302_n3889# bias_b bias_b VDD m1_n6302_n3889# VDD bias_b m1_n6302_n3889# bias_b
+ VDD bias_b m1_n208_n2883# bias_b bias_b m1_1038_n2886# bias_b m1_n6302_n3889# m1_n6302_n3889#
+ VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b bias_b m1_1038_n2886# m1_n6302_n3889#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_lvt_FF_9 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_DD_2 m1_n947_n12836# bias_d VSS bias_d bias_a m1_n1659_n11581#
+ m1_n947_n12836# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# op on bias_d
+ bias_d on on op on bias_d VSS op m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n1659_n11581#
+ bias_d bias_d bias_d VSS m1_n947_n12836# m1_n947_n12836# op VSS m1_n947_n12836#
+ op m1_n1659_n11581# m1_n1659_n11581# bias_d bias_d on bias_d on bias_d m1_n1659_n11581#
+ bias_d bias_d on VSS op VSS VSS op on bias_d bias_d m1_n947_n12836# op op bias_d
+ bias_d bias_d VSS bias_d VSS m1_n1659_n11581# m1_n947_n12836# m1_n2176_n12171# VSS
+ m1_n1659_n11581# bias_d bias_d on VSS m1_n1659_n11581# bias_d m1_n947_n12836# VSS
+ sky130_fd_pr__nfet_01v8_DD
Xsky130_fd_pr__pfet_01v8_lvt_II_3 m1_2462_n3318# bias_b m1_2463_n5585# bias_b VDD
+ m1_2462_n3318# bias_b bias_b VDD m1_2463_n5585# VDD bias_b m1_2463_n5585# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2463_n5585# m1_2462_n3318#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2462_n3318#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__pfet_01v8_lvt_II_4 m1_1038_n2886# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_n208_n2883# VDD VDD VDD bias_b VDD bias_b m1_n208_n2883# bias_b bias_b
+ m1_n208_n2883# bias_b VDD VDD VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b VDD m1_1038_n2886#
+ VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_CC_4 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a
+ VSS cmc VSS cmc cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc VSS cmc cmc VSS VSS m1_n5574_n13620# m1_n5574_n13620#
+ bias_a m1_n5574_n13620# VSS bias_a cmc VSS cmc VSS VSS bias_a bias_a m1_n5574_n13620#
+ m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620# m1_n5574_n13620#
+ m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a bias_a bias_a m1_n5574_n13620#
+ m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620# cmc cmc VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_5 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS
+ bias_a VSS VSS bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS VSS bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS VSS VSS cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS m1_n5574_n13620# bias_a
+ bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_6 VSS VSS VSS VSS bias_a bias_a m1_n947_n12836# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n1659_n11581# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n947_n12836# bias_a m1_n1659_n11581# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n1659_n11581# m1_n947_n12836# bias_a bias_a bias_a
+ m1_n1659_n11581# m1_n2176_n12171# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_10 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS
+ bias_a VSS cmc cmc bias_a VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS cmc bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_7 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n947_n12836# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n1659_n11581# m1_n2176_n12171# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n2176_n12171# m1_n1659_n11581# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_0 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias i_bias
+ i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__nfet_01v8_CC_11 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a
+ VSS cmc VSS bias_a bias_a cmc VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc VSS bias_a cmc VSS VSS m1_n5574_n13620# m1_n5574_n13620#
+ bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620# bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ cmc bias_a m1_n5574_n13620# m1_n5574_n13620# VSS cmc bias_a VSS m1_n5574_n13620#
+ bias_a cmc VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_CC_8 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n947_n12836# m1_n947_n12836# bias_a m1_n1659_n11581# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n1659_n11581# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n1659_n11581# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n1659_n11581# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n947_n12836# m1_n2176_n12171# m1_n947_n12836# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_1 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__nfet_01v8_CC_9 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a
+ VSS cmc VSS VSS cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc VSS VSS cmc VSS VSS m1_n5574_n13620# m1_n5574_n13620#
+ bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# VSS cmc VSS VSS VSS bias_a cmc m1_n5574_n13620# m1_n5574_n13620#
+ m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a bias_a bias_a m1_n5574_n13620#
+ m1_n5574_n13620# VSS bias_a bias_a VSS m1_n5574_n13620# cmc cmc VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_2 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias bias_c
+ i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__nfet_01v8_CC_12 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS
+ bias_a VSS bias_a bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS bias_a bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS cmc bias_a VSS bias_a VSS VSS cmc cmc
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620# bias_a bias_a
+ cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS
+ m1_n5574_n13620# cmc cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc bias_a VSS
+ m1_n5574_n13620# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_CC
Xsky130_fd_pr__nfet_01v8_BB_3 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias i_bias
+ i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS i_bias
+ VSS sky130_fd_pr__nfet_01v8_BB
Xsky130_fd_pr__pfet_01v8_HH_0 VDD bias_c m1_6690_n8907# op bias_c bias_c m1_1038_n2886#
+ bias_b bias_c VDD m1_n208_n2883# bias_c VDD on bias_c VDD VDD m1_2463_n5585# VDD
+ m1_2462_n3318# m1_2462_n3318# op m1_2463_n5585# m1_2462_n3318# VDD VDD VDD bias_b
+ bias_c m1_1038_n2886# bias_c m1_6690_n8907# VDD bias_c VDD VDD m1_2463_n5585# on
+ VDD bias_c m1_2462_n3318# m1_n208_n2883# bias_c bias_c VDD VDD m1_2463_n5585# VDD
+ VSS sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__nfet_01v8_lvt_GG_0 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_10 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__pfet_01v8_HH_1 op VDD on op VDD bias_c m1_1038_n2886# op bias_c bias_c
+ VDD VDD m1_1038_n2886# on bias_c bias_c VDD m1_n208_n2883# bias_c m1_1038_n2886#
+ m1_1038_n2886# m1_n6302_n3889# m1_n208_n2883# m1_1038_n2886# m1_n6302_n3889# bias_c
+ bias_c op bias_c VDD bias_c on bias_c bias_c cm bias_c m1_n208_n2883# cm m1_n208_n2883#
+ VDD m1_1038_n2886# m1_n208_n2883# bias_c bias_c on bias_c m1_n208_n2883# bias_c
+ VSS sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__nfet_01v8_AA_0 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_lvt_GG_1 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_11 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__pfet_01v8_HH_3 VDD bias_c bias_b on bias_c bias_c m1_n208_n2883# m1_6690_n8907#
+ bias_c VDD m1_1038_n2886# bias_c VDD op bias_c VDD VDD m1_2462_n3318# VDD m1_2463_n5585#
+ m1_2463_n5585# on m1_2462_n3318# m1_2463_n5585# VDD VDD VDD m1_6690_n8907# bias_c
+ m1_n208_n2883# bias_c bias_b VDD bias_c VDD VDD m1_2462_n3318# op VDD bias_c m1_2463_n5585#
+ m1_1038_n2886# bias_c bias_c VDD VDD m1_2462_n3318# VDD VSS sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__pfet_01v8_HH_2 on VDD op on VDD bias_c m1_n208_n2883# on bias_c bias_c
+ VDD VDD m1_n208_n2883# op bias_c bias_c VDD m1_1038_n2886# bias_c m1_n208_n2883#
+ m1_n208_n2883# m1_n6302_n3889# m1_1038_n2886# m1_n208_n2883# m1_n6302_n3889# bias_c
+ bias_c on bias_c VDD bias_c op bias_c bias_c cm bias_c m1_1038_n2886# cm m1_1038_n2886#
+ VDD m1_n208_n2883# m1_1038_n2886# bias_c bias_c op bias_c m1_1038_n2886# bias_c
+ VSS sky130_fd_pr__pfet_01v8_HH
Xsky130_fd_pr__nfet_01v8_lvt_GG_2 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_AA_1 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d bias_a m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_a m1_6690_n8907# bias_a VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_AA_2 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_a
+ m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_lvt_FF_12 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_GG_3 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_AA_3 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d
+ m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_AA
Xsky130_fd_pr__nfet_01v8_lvt_FF_13 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_GG_4 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_14 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_15 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_GG_5 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_EE_0 cm cm cm cm cm cm cm m1_11534_n9706# m1_11242_n9716#
+ cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# cm cm cm cm VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_GG_6 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_EE_1 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490# m1_11534_n9706#
+ m1_11242_n9716# cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# m1_11940_n10482#
+ m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_GG_7 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_GG
Xsky130_fd_pr__nfet_01v8_lvt_FF_0 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_EE_2 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490# m1_11534_n11258#
+ m1_11244_n11260# cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260#
+ m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_FF_1 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_EE_3 cm cm cm cm VSS cm VSS m1_11534_n11258# m1_11244_n11260#
+ cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260# VSS VSS cm VSS
+ VSS sky130_fd_pr__nfet_01v8_EE
Xsky130_fd_pr__nfet_01v8_lvt_FF_2 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsc_cmfb_0 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480#
+ bias_a sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# p2_b sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480#
+ p1 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480#
+ p2 VDD sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_6/in
+ cmc sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# on sc_cmfb_0/transmission_gate_8/in
+ sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_7/in cm sc_cmfb_0/transmission_gate_9/in sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# p1_b VSS op sc_cmfb
Xsky130_fd_pr__nfet_01v8_lvt_FF_3 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_4 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_5 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_lvt_FF_6 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__pfet_01v8_lvt_II_0 m1_n208_n2883# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_1038_n2886# VDD VDD VDD bias_b VDD bias_b m1_1038_n2886# bias_b bias_b
+ m1_1038_n2886# bias_b VDD VDD VDD m1_n208_n2883# bias_b VDD VDD VDD bias_b VDD m1_n208_n2883#
+ VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_lvt_FF_7 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_DD_0 m1_n1659_n11581# bias_d VSS bias_d bias_a m1_n947_n12836#
+ m1_n1659_n11581# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# on op bias_d
+ bias_d op op on op bias_d VSS on m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n947_n12836#
+ bias_d bias_d bias_d VSS m1_n1659_n11581# m1_n1659_n11581# on VSS m1_n1659_n11581#
+ on m1_n947_n12836# m1_n947_n12836# bias_d bias_d op bias_d op bias_d m1_n947_n12836#
+ bias_d bias_d op VSS on VSS VSS on op bias_d bias_d m1_n1659_n11581# on on bias_d
+ bias_d bias_d VSS bias_d VSS m1_n947_n12836# m1_n1659_n11581# m1_n2176_n12171# VSS
+ m1_n947_n12836# bias_d bias_d op VSS m1_n947_n12836# bias_d m1_n1659_n11581# VSS
+ sky130_fd_pr__nfet_01v8_DD
Xsky130_fd_pr__pfet_01v8_lvt_II_1 m1_2463_n5585# bias_b m1_2462_n3318# bias_b VDD
+ m1_2463_n5585# bias_b bias_b VDD m1_2462_n3318# VDD bias_b m1_2462_n3318# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2462_n3318# m1_2463_n5585#
+ VDD m1_1038_n2886# bias_b VDD VDD VDD bias_b bias_b m1_n208_n2883# m1_2463_n5585#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_II
Xsky130_fd_pr__nfet_01v8_lvt_FF_8 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886# VSS
+ sky130_fd_pr__nfet_01v8_lvt_FF
Xsky130_fd_pr__nfet_01v8_DD_1 m1_n947_n12836# bias_d bias_d bias_d op m1_n947_n12836#
+ m1_n2176_n12171# bias_d VSS bias_d VSS bias_d m1_n1659_n11581# on VSS bias_d bias_d
+ on bias_a bias_a bias_a bias_d bias_d bias_a m1_n1659_n11581# VSS bias_d on op VSS
+ VSS bias_d bias_d bias_d m1_n947_n12836# m1_n2176_n12171# bias_a bias_d m1_n947_n12836#
+ bias_a m1_n2176_n12171# m1_n1659_n11581# bias_d bias_d bias_a bias_d op VSS m1_n2176_n12171#
+ bias_d VSS bias_a bias_d VSS op bias_d bias_a on bias_d bias_d m1_n1659_n11581#
+ op on VSS bias_d bias_d on bias_d bias_d m1_n2176_n12171# VSS m1_n1659_n11581# bias_d
+ m1_n947_n12836# bias_d VSS bias_a op m1_n947_n12836# bias_d m1_n2176_n12171# VSS
+ sky130_fd_pr__nfet_01v8_DD
C0 m1_2462_n3318# bias_b 3.43fF
C1 bias_a m1_2462_n3318# 0.11fF
C2 cmc op 1.20fF
C3 m1_2463_n5585# VDD 7.63fF
C4 VSS m1_6690_n8907# 0.22fF
C5 m1_11242_n9716# m1_11244_n11260# 0.01fF
C6 m1_12410_n9718# m1_12410_n11263# 0.01fF
C7 m1_11534_n9706# m1_11825_n9711# 0.07fF
C8 m1_11940_n10482# m1_12232_n10488# 0.07fF
C9 on cm 1.01fF
C10 m1_12410_n9718# cm 0.64fF
C11 m1_12118_n11263# m1_12410_n11263# 0.07fF
C12 VSS m1_11825_n9711# 0.00fF
C13 m1_11940_n10482# cm 0.59fF
C14 op bias_d 12.45fF
C15 m1_12118_n11263# cm 0.57fF
C16 op m1_1038_n2886# 0.78fF
C17 cm sc_cmfb_0/transmission_gate_8/in 0.04fF
C18 VSS m1_2462_n3318# 0.00fF
C19 m1_2462_n3318# m1_6690_n8907# 2.72fF
C20 bias_b m1_n208_n2883# 9.15fF
C21 bias_c op 5.30fF
C22 bias_a m1_n208_n2883# 0.04fF
C23 m1_n6302_n3889# cm 2.61fF
C24 m1_n947_n12836# cmc 0.37fF
C25 m1_11063_n10490# m1_11940_n10482# 0.02fF
C26 cmc bias_a 12.12fF
C27 m1_n5574_n13620# cm 0.02fF
C28 VSS m1_11244_n11260# -0.00fF
C29 m1_n5574_n13620# ip 1.01fF
C30 cmc p1_b 0.04fF
C31 m1_2463_n5585# op 0.25fF
C32 on VDD 5.69fF
C33 m1_n947_n12836# bias_d 16.58fF
C34 bias_a bias_d 8.20fF
C35 m1_11242_n9716# m1_12118_n9704# 0.02fF
C36 bias_b m1_1038_n2886# 10.79fF
C37 bias_a m1_1038_n2886# 0.07fF
C38 VSS m1_n208_n2883# 0.03fF
C39 m1_6690_n8907# m1_n208_n2883# 0.10fF
C40 m1_11356_n10481# m1_11940_n10482# 0.03fF
C41 on m1_n2176_n12171# 8.63fF
C42 cmc VSS 32.86fF
C43 m1_11534_n9706# m1_11534_n11258# 0.01fF
C44 bias_c bias_b 25.24fF
C45 bias_a bias_c 0.00fF
C46 cmc m1_6690_n8907# 0.46fF
C47 sc_cmfb_0/transmission_gate_3/out op 0.00fF
C48 m1_n6302_n3889# VDD 3.85fF
C49 in ip 3.13fF
C50 VSS m1_11534_n11258# 0.00fF
C51 m1_n5574_n13620# VDD 0.03fF
C52 m1_n1659_n11581# on 1.52fF
C53 m1_n5574_n13620# m1_n2176_n12171# 0.57fF
C54 VSS bias_d 1.08fF
C55 m1_2462_n3318# m1_n208_n2883# 3.03fF
C56 m1_11534_n9706# m1_12118_n9704# 0.03fF
C57 m1_6690_n8907# bias_d 35.87fF
C58 m1_2463_n5585# bias_b 6.62fF
C59 VSS m1_1038_n2886# 0.20fF
C60 m1_6690_n8907# m1_1038_n2886# 0.28fF
C61 on p1 0.01fF
C62 m1_11648_n10486# m1_11940_n10482# 0.07fF
C63 m1_n1659_n11581# m1_n5574_n13620# 0.14fF
C64 VSS bias_c 3.39fF
C65 cm sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.01fF
C66 VSS m1_12118_n9704# 0.01fF
C67 m1_12232_n10488# cm 0.57fF
C68 bias_c m1_6690_n8907# 1.61fF
C69 m1_12410_n11263# cm 0.58fF
C70 i_bias VSS 13.74fF
C71 VSS m1_11826_n11260# -0.00fF
C72 on op 7.65fF
C73 m1_11063_n10490# m1_12232_n10488# 0.02fF
C74 cmc p2_b 0.01fF
C75 m1_2462_n3318# m1_1038_n2886# 4.36fF
C76 m1_11063_n10490# cm 0.61fF
C77 m1_11825_n9711# m1_12118_n9704# 0.07fF
C78 m1_11244_n11260# m1_11534_n11258# 0.07fF
C79 m1_2463_n5585# VSS 0.00fF
C80 m1_2463_n5585# m1_6690_n8907# 0.36fF
C81 bias_c m1_2462_n3318# 4.04fF
C82 m1_11825_n9711# m1_11826_n11260# 0.01fF
C83 m1_n6302_n3889# op 0.17fF
C84 VSS sc_cmfb_0/transmission_gate_7/in 0.01fF
C85 cmc m1_n208_n2883# 0.14fF
C86 m1_n5574_n13620# op 0.17fF
C87 m1_11242_n9716# m1_12410_n9718# 0.02fF
C88 m1_n947_n12836# on 8.70fF
C89 m1_11356_n10481# m1_12232_n10488# 0.02fF
C90 cm VDD 3.69fF
C91 bias_b on 0.07fF
C92 bias_a on 4.51fF
C93 m1_2463_n5585# m1_2462_n3318# 4.55fF
C94 m1_11356_n10481# cm 0.58fF
C95 m1_11244_n11260# m1_11826_n11260# 0.03fF
C96 m1_n208_n2883# m1_1038_n2886# 17.20fF
C97 cmc bias_d 0.03fF
C98 bias_a sc_cmfb_0/transmission_gate_8/in 0.02fF
C99 cmc m1_1038_n2886# 0.17fF
C100 sc_cmfb_0/transmission_gate_4/out VDD 0.01fF
C101 bias_c m1_n208_n2883# 8.21fF
C102 m1_n6302_n3889# bias_b 2.49fF
C103 m1_n947_n12836# m1_n5574_n13620# 0.12fF
C104 i_bias m1_n208_n2883# 0.24fF
C105 cmc bias_c 0.07fF
C106 m1_11063_n10490# m1_11356_n10481# 0.07fF
C107 m1_n5574_n13620# bias_b 0.11fF
C108 bias_a m1_n5574_n13620# 21.14fF
C109 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.08fF
C110 m1_11534_n9706# m1_12410_n9718# 0.02fF
C111 m1_11648_n10486# m1_12232_n10488# 0.03fF
C112 VSS on 0.66fF
C113 p1 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.00fF
C114 VSS m1_12410_n9718# 0.01fF
C115 m1_6690_n8907# on 1.68fF
C116 m1_11648_n10486# cm 0.59fF
C117 m1_11534_n11258# m1_11826_n11260# 0.07fF
C118 VSS m1_11940_n10482# 0.01fF
C119 VSS m1_12118_n11263# 0.01fF
C120 cm p1 0.17fF
C121 m1_2463_n5585# m1_n208_n2883# 3.39fF
C122 VSS sc_cmfb_0/transmission_gate_8/in 0.06fF
C123 bias_c m1_1038_n2886# 7.06fF
C124 i_bias m1_1038_n2886# 0.27fF
C125 bias_b in 0.09fF
C126 m1_11063_n10490# m1_11648_n10486# 0.03fF
C127 m1_n5574_n13620# VSS 19.74fF
C128 m1_11825_n9711# m1_12410_n9718# 0.03fF
C129 m1_n5574_n13620# m1_6690_n8907# 0.08fF
C130 sc_cmfb_0/transmission_gate_4/out p1 -0.00fF
C131 op cm 0.76fF
C132 i_bias bias_c 12.15fF
C133 m1_2462_n3318# on 0.27fF
C134 sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.00fF
C135 m1_2463_n5585# m1_1038_n2886# 3.88fF
C136 m1_n1659_n11581# m1_n2176_n12171# 10.31fF
C137 m1_2463_n5585# bias_c 2.57fF
C138 m1_n6302_n3889# m1_2462_n3318# 0.57fF
C139 VSS in 0.01fF
C140 m1_11356_n10481# m1_11648_n10486# 0.07fF
C141 m1_11242_n9716# cm 0.68fF
C142 VDD sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.02fF
C143 m1_11244_n11260# m1_12118_n11263# 0.02fF
C144 bias_b cm 0.36fF
C145 bias_a cm 0.62fF
C146 op VDD 5.61fF
C147 on m1_n208_n2883# 0.40fF
C148 cmc on 0.96fF
C149 bias_b ip 0.07fF
C150 p1_b cm 0.09fF
C151 op m1_n2176_n12171# 1.95fF
C152 m1_n6302_n3889# m1_n208_n2883# 3.54fF
C153 m1_11534_n9706# cm 0.65fF
C154 m1_11534_n11258# m1_12118_n11263# 0.03fF
C155 VSS m1_12232_n10488# 0.02fF
C156 m1_n5574_n13620# m1_n208_n2883# 2.49fF
C157 m1_n1659_n11581# op 8.09fF
C158 VSS m1_12410_n11263# 0.01fF
C159 cmc m1_n5574_n13620# 54.64fF
C160 on bias_d 13.96fF
C161 VSS cm 0.57fF
C162 p2_b p2 0.00fF
C163 p1 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.00fF
C164 m1_6690_n8907# cm 4.14fF
C165 on m1_1038_n2886# 3.37fF
C166 bias_b VDD 41.24fF
C167 bias_a VDD 0.11fF
C168 bias_c on 4.92fF
C169 VSS ip 0.00fF
C170 m1_12118_n9704# m1_12410_n9718# 0.07fF
C171 op p1 0.00fF
C172 VSS m1_11063_n10490# 0.01fF
C173 cmc p2 0.00fF
C174 VSS sc_cmfb_0/transmission_gate_4/out 0.03fF
C175 op sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.00fF
C176 m1_12118_n9704# m1_12118_n11263# 0.01fF
C177 m1_6690_n8907# sc_cmfb_0/transmission_gate_4/out 0.01fF
C178 m1_n947_n12836# m1_n2176_n12171# 10.60fF
C179 m1_n6302_n3889# m1_1038_n2886# 2.81fF
C180 bias_a m1_n2176_n12171# 23.78fF
C181 p1_b VDD -0.01fF
C182 m1_11825_n9711# cm 0.65fF
C183 in m1_n208_n2883# 3.17fF
C184 m1_n5574_n13620# m1_1038_n2886# 2.45fF
C185 m1_11826_n11260# m1_12118_n11263# 0.07fF
C186 cmc in 0.04fF
C187 m1_n6302_n3889# bias_c 3.58fF
C188 m1_2462_n3318# cm 1.44fF
C189 m1_n1659_n11581# m1_n947_n12836# 9.35fF
C190 m1_n5574_n13620# bias_c 0.50fF
C191 m1_n1659_n11581# bias_a 20.90fF
C192 m1_2463_n5585# on 0.09fF
C193 m1_n5574_n13620# i_bias 0.12fF
C194 VSS VDD 0.10fF
C195 m1_11244_n11260# m1_12410_n11263# 0.02fF
C196 m1_6690_n8907# VDD 3.64fF
C197 VSS m1_11356_n10481# 0.01fF
C198 m1_11244_n11260# cm 0.55fF
C199 bias_a p1 0.04fF
C200 m1_n6302_n3889# m1_2463_n5585# 0.56fF
C201 VSS m1_n2176_n12171# 4.39fF
C202 in m1_1038_n2886# 1.58fF
C203 m1_6690_n8907# m1_n2176_n12171# 0.00fF
C204 bias_c in 0.44fF
C205 p1 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.00fF
C206 p1_b p1 -0.00fF
C207 m1_n1659_n11581# VSS 5.68fF
C208 m1_n947_n12836# op 1.19fF
C209 i_bias in 0.29fF
C210 cm m1_n208_n2883# 0.17fF
C211 bias_b op 0.14fF
C212 bias_a op 2.42fF
C213 cmc cm 0.85fF
C214 m1_2462_n3318# VDD 7.01fF
C215 m1_11534_n11258# m1_12410_n11263# 0.02fF
C216 ip m1_n208_n2883# 1.08fF
C217 VSS m1_11648_n10486# 0.01fF
C218 m1_11534_n11258# cm 0.58fF
C219 VSS p1 0.04fF
C220 VSS sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.02fF
C221 cm bias_d 0.08fF
C222 VDD p2_b 0.00fF
C223 cm m1_1038_n2886# 1.34fF
C224 VSS op 0.86fF
C225 m1_6690_n8907# op 2.49fF
C226 m1_n947_n12836# bias_a 21.86fF
C227 bias_c cm 3.39fF
C228 m1_12118_n9704# cm 0.64fF
C229 m1_11826_n11260# m1_12410_n11263# 0.03fF
C230 VDD m1_n208_n2883# 15.19fF
C231 ip m1_1038_n2886# 1.68fF
C232 m1_n6302_n3889# on 0.08fF
C233 m1_11826_n11260# cm 0.58fF
C234 cmc VDD 0.08fF
C235 m1_n5574_n13620# on 0.06fF
C236 bias_c ip 0.11fF
C237 bias_a sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.05fF
C238 bias_a p1_b 0.01fF
C239 m1_n2176_n12171# m1_n208_n2883# 0.09fF
C240 i_bias ip 0.17fF
C241 m1_11242_n9716# m1_11534_n9706# 0.07fF
C242 cmc m1_n2176_n12171# 1.14fF
C243 sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.02fF
C244 VSS m1_11242_n9716# 0.00fF
C245 m1_2462_n3318# op 0.28fF
C246 m1_2463_n5585# cm 0.52fF
C247 m1_n1659_n11581# cmc 0.44fF
C248 m1_n947_n12836# VSS 7.60fF
C249 cm sc_cmfb_0/transmission_gate_7/in 0.04fF
C250 VSS bias_b 0.23fF
C251 bias_a VSS 70.68fF
C252 VDD m1_1038_n2886# 15.36fF
C253 m1_6690_n8907# bias_b 0.39fF
C254 bias_a m1_6690_n8907# 2.54fF
C255 bias_c VDD 10.55fF
C256 bias_d m1_n2176_n12171# 8.59fF
C257 m1_n2176_n12171# m1_1038_n2886# 0.11fF
C258 VSS p1_b 0.01fF
C259 m1_11242_n9716# m1_11825_n9711# 0.03fF
C260 cmc p1 0.00fF
C261 bias_c m1_n2176_n12171# 0.02fF
C262 m1_n1659_n11581# bias_d 12.63fF
C263 on sc_cmfb_0/transmission_gate_9/in 0.00fF
C264 VSS m1_11534_n9706# 0.00fF
C265 m1_n5574_n13620# in 2.04fF
C266 op m1_n208_n2883# 3.85fF
C267 m1_1038_n2886# 0 -76.00fF
C268 m1_n208_n2883# 0 -83.42fF
C269 m1_n2176_n12171# 0 12.82fF
C270 bias_d 0 119.38fF
C271 ip 0 2.31fF
C272 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0 1.37fF
C273 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# 0 1.37fF
C274 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0 1.37fF
C275 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# 0 1.37fF
C276 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# 0 1.37fF
C277 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0 1.37fF
C278 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# 0 1.37fF
C279 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# 0 1.37fF
C280 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# 0 1.37fF
C281 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0 1.37fF
C282 sc_cmfb_0/transmission_gate_9/in 0 -27.99fF
C283 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# 0 1.37fF
C284 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# 0 1.37fF
C285 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# 0 1.37fF
C286 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0 1.37fF
C287 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0 1.37fF
C288 p2 0 9.44fF
C289 p2_b 0 3.15fF
C290 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# 0 1.37fF
C291 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0 1.37fF
C292 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# 0 1.37fF
C293 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0 1.37fF
C294 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0 1.37fF
C295 sc_cmfb_0/transmission_gate_8/in 0 -0.42fF
C296 sc_cmfb_0/transmission_gate_6/in 0 2.41fF
C297 sc_cmfb_0/transmission_gate_7/in 0 1.91fF
C298 cm 0 -13.24fF
C299 p1 0 9.87fF
C300 op 0 -12.21fF
C301 sc_cmfb_0/transmission_gate_4/out 0 0.84fF
C302 p1_b 0 1.48fF
C303 VDD 0 364.20fF
C304 on 0 -77.28fF
C305 sc_cmfb_0/transmission_gate_3/out 0 -4.68fF
C306 in 0 2.38fF
C307 m1_12410_n11263# 0 0.16fF
C308 m1_12118_n11263# 0 0.30fF
C309 m1_11826_n11260# 0 0.32fF
C310 m1_11534_n11258# 0 0.23fF
C311 m1_11244_n11260# 0 0.24fF
C312 m1_12232_n10488# 0 0.22fF
C313 m1_11940_n10482# 0 0.34fF
C314 m1_11648_n10486# 0 0.25fF
C315 m1_11356_n10481# 0 0.26fF
C316 m1_11063_n10490# 0 0.26fF
C317 bias_b 0 12.75fF
C318 m1_12410_n9718# 0 0.16fF
C319 m1_12118_n9704# 0 0.27fF
C320 m1_11825_n9711# 0 0.29fF
C321 m1_11534_n9706# 0 0.22fF
C322 m1_11242_n9716# 0 0.23fF
C323 m1_6690_n8907# 0 -73.84fF
C324 m1_2462_n3318# 0 -13.18fF
C325 bias_c 0 43.28fF
C326 VSS 0 179.48fF
C327 i_bias 0 21.00fF
C328 m1_n5574_n13620# 0 183.14fF
C329 bias_a 0 -298.49fF
C330 cmc 0 0.86fF
C331 m1_2463_n5585# 0 0.31fF
C332 m1_n1659_n11581# 0 3.21fF
C333 m1_n947_n12836# 0 7.99fF
C334 m1_n6302_n3889# 0 10.46fF
.ends

.subckt sky130_fd_sc_hd__clkinv_16 A VGND VPWR Y VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.0605e+12p pd=1.261e+07u as=1.0059e+12p ps=1.151e+07u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.515e+12p pd=3.103e+07u as=3.655e+12p ps=3.331e+07u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 VPWR VGND 0.34fF
C1 A VGND 0.66fF
C2 Y VPB 0.09fF
C3 VPWR Y 4.41fF
C4 VPWR VPB 0.89fF
C5 A Y 1.32fF
C6 Y VGND 1.58fF
C7 A VPB 1.26fF
C8 VPWR A 0.64fF
C9 VGND VNB 1.26fF
C10 Y VNB 0.13fF
C11 VPWR VNB 0.47fF
C12 A VNB 1.70fF
C13 VPB VNB 2.20fF
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y w_82_21# VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=8.4e+11p pd=7.68e+06u as=1.21e+12p ps=1.042e+07u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=4.221e+11p pd=4.53e+06u as=2.352e+11p ps=2.8e+06u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 A VPB 0.21fF
C1 A VPWR 0.13fF
C2 Y A 0.88fF
C3 VGND VPWR 0.10fF
C4 VGND Y 0.56fF
C5 VGND A 0.13fF
C6 VPWR VPB 0.34fF
C7 Y VPB 0.05fF
C8 Y VPWR 1.13fF
C9 VGND VNB 0.40fF
C10 Y VNB 0.10fF
C11 VPWR VNB 0.14fF
C12 A VNB 0.47fF
C13 VPB VNB 0.69fF
.ends

.subckt onebit_dac VDD v v_b out v_lo v_hi VSS
Xtransmission_gate_0 v VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ v_hi out VSS v_b transmission_gate
Xtransmission_gate_1 v_b VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ v_lo out VSS v transmission_gate
C0 v_b out 0.47fF
C1 VDD v -0.13fF
C2 v_b v_hi 0.45fF
C3 VDD out 1.01fF
C4 v_b v_lo 0.45fF
C5 out v 0.19fF
C6 VDD v_hi 0.16fF
C7 VDD v_lo 0.04fF
C8 v v_hi 0.19fF
C9 out v_hi 0.20fF
C10 v_lo v 0.13fF
C11 out v_lo 0.29fF
C12 v_lo v_hi 0.50fF
C13 VDD v_b 0.15fF
C14 v_b v 0.62fF
C15 v_b VSS 1.48fF
C16 out VSS 3.17fF
C17 v_lo VSS 1.71fF
C18 v VSS 1.88fF
C19 VDD VSS 7.43fF
C20 v_hi VSS 1.27fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_VU7MNH a_n652_n140# a_652_n194# a_772_n140# a_n60_n194#
+ a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140# a_296_n194#
+ a_60_n140# a_416_n140# a_n118_n140# a_118_n194# a_238_n140# a_n772_n194# a_n830_n140#
+ a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X4 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n772_n194# a_n60_n194# 0.01fF
C1 a_n118_n140# a_416_n140# 0.04fF
C2 a_60_n140# a_772_n140# 0.03fF
C3 a_238_n140# a_772_n140# 0.04fF
C4 a_n652_n140# a_594_n140# 0.02fF
C5 a_n238_n194# a_474_n194# 0.01fF
C6 a_474_n194# a_296_n194# 0.10fF
C7 a_n652_n140# a_416_n140# 0.02fF
C8 a_n830_n140# a_n474_n140# 0.06fF
C9 a_n238_n194# a_n416_n194# 0.10fF
C10 a_n118_n140# a_n474_n140# 0.06fF
C11 a_296_n194# a_n416_n194# 0.01fF
C12 a_594_n140# a_n296_n140# 0.02fF
C13 a_416_n140# a_n296_n140# 0.03fF
C14 a_n772_n194# a_474_n194# 0.01fF
C15 a_118_n194# a_n594_n194# 0.01fF
C16 a_n238_n194# a_652_n194# 0.01fF
C17 a_n772_n194# a_n416_n194# 0.03fF
C18 a_296_n194# a_652_n194# 0.03fF
C19 a_n652_n140# a_n474_n140# 0.13fF
C20 a_n60_n194# a_n594_n194# 0.02fF
C21 a_594_n140# a_416_n140# 0.13fF
C22 a_60_n140# a_n830_n140# 0.02fF
C23 a_60_n140# a_n118_n140# 0.13fF
C24 a_n772_n194# a_652_n194# 0.01fF
C25 a_238_n140# a_n830_n140# 0.02fF
C26 a_n296_n140# a_n474_n140# 0.13fF
C27 a_238_n140# a_n118_n140# 0.06fF
C28 a_594_n140# a_n474_n140# 0.02fF
C29 a_n652_n140# a_60_n140# 0.03fF
C30 a_416_n140# a_n474_n140# 0.02fF
C31 a_474_n194# a_n594_n194# 0.01fF
C32 a_n238_n194# a_296_n194# 0.02fF
C33 a_238_n140# a_n652_n140# 0.02fF
C34 a_n416_n194# a_n594_n194# 0.10fF
C35 a_60_n140# a_n296_n140# 0.06fF
C36 a_238_n140# a_n296_n140# 0.04fF
C37 a_n772_n194# a_n238_n194# 0.02fF
C38 a_n772_n194# a_296_n194# 0.01fF
C39 a_652_n194# a_n594_n194# 0.01fF
C40 a_60_n140# a_594_n140# 0.04fF
C41 a_238_n140# a_594_n140# 0.06fF
C42 a_60_n140# a_416_n140# 0.06fF
C43 a_238_n140# a_416_n140# 0.13fF
C44 a_n60_n194# a_118_n194# 0.10fF
C45 a_60_n140# a_n474_n140# 0.04fF
C46 a_772_n140# a_n830_n140# 0.01fF
C47 a_238_n140# a_n474_n140# 0.03fF
C48 a_n118_n140# a_772_n140# 0.02fF
C49 a_n238_n194# a_n594_n194# 0.03fF
C50 a_296_n194# a_n594_n194# 0.01fF
C51 a_474_n194# a_118_n194# 0.03fF
C52 a_n772_n194# a_n594_n194# 0.10fF
C53 a_n652_n140# a_772_n140# 0.01fF
C54 a_n60_n194# a_474_n194# 0.02fF
C55 a_118_n194# a_n416_n194# 0.02fF
C56 a_238_n140# a_60_n140# 0.13fF
C57 a_n60_n194# a_n416_n194# 0.03fF
C58 a_772_n140# a_n296_n140# 0.02fF
C59 a_652_n194# a_118_n194# 0.02fF
C60 a_n118_n140# a_n830_n140# 0.03fF
C61 a_n60_n194# a_652_n194# 0.01fF
C62 a_772_n140# a_594_n140# 0.13fF
C63 a_772_n140# a_416_n140# 0.06fF
C64 a_n652_n140# a_n830_n140# 0.13fF
C65 a_474_n194# a_n416_n194# 0.01fF
C66 a_n652_n140# a_n118_n140# 0.04fF
C67 a_n830_n140# a_n296_n140# 0.04fF
C68 a_772_n140# a_n474_n140# 0.02fF
C69 a_n238_n194# a_118_n194# 0.03fF
C70 a_474_n194# a_652_n194# 0.10fF
C71 a_296_n194# a_118_n194# 0.10fF
C72 a_n118_n140# a_n296_n140# 0.13fF
C73 a_n60_n194# a_n238_n194# 0.10fF
C74 a_652_n194# a_n416_n194# 0.01fF
C75 a_n60_n194# a_296_n194# 0.03fF
C76 a_n830_n140# a_594_n140# 0.01fF
C77 a_n772_n194# a_118_n194# 0.01fF
C78 a_n118_n140# a_594_n140# 0.03fF
C79 a_n830_n140# a_416_n140# 0.02fF
C80 a_n652_n140# a_n296_n140# 0.06fF
C81 a_772_n140# VSUBS 0.02fF
C82 a_594_n140# VSUBS 0.02fF
C83 a_416_n140# VSUBS 0.02fF
C84 a_238_n140# VSUBS 0.02fF
C85 a_60_n140# VSUBS 0.02fF
C86 a_n118_n140# VSUBS 0.02fF
C87 a_n296_n140# VSUBS 0.02fF
C88 a_n474_n140# VSUBS 0.02fF
C89 a_n652_n140# VSUBS 0.02fF
C90 a_n830_n140# VSUBS 0.02fF
C91 a_652_n194# VSUBS 0.29fF
C92 a_474_n194# VSUBS 0.23fF
C93 a_296_n194# VSUBS 0.24fF
C94 a_118_n194# VSUBS 0.25fF
C95 a_n60_n194# VSUBS 0.26fF
C96 a_n238_n194# VSUBS 0.27fF
C97 a_n416_n194# VSUBS 0.28fF
C98 a_n594_n194# VSUBS 0.28fF
C99 a_n772_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_TRAZV8 a_20_n120# a_n78_n120# a_n33_n208# VSUBS
X0 a_20_n120# a_n33_n208# a_n78_n120# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=3.48e+11p pd=2.98e+06u as=3.48e+11p ps=2.98e+06u w=1.2e+06u l=200000u
C0 a_n78_n120# a_n33_n208# 0.02fF
C1 a_20_n120# a_n33_n208# 0.02fF
C2 a_n78_n120# a_20_n120# 0.28fF
C3 a_20_n120# VSUBS 0.02fF
C4 a_n78_n120# VSUBS 0.02fF
C5 a_n33_n208# VSUBS 0.29fF
.ends

.subckt sky130_fd_pr__nfet_01v8_BASQVB a_n1008_n140# a_n652_n140# a_652_n194# a_772_n140#
+ a_n60_n194# a_n474_n140# a_n416_n194# a_474_n194# a_594_n140# a_n238_n194# a_n296_n140#
+ a_296_n194# a_60_n140# a_416_n140# a_n950_n194# a_n118_n140# a_118_n194# a_238_n140#
+ a_n772_n194# a_n830_n140# a_830_n194# a_950_n140# a_n594_n194# VSUBS
X0 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X6 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_416_n140# a_238_n140# 0.13fF
C1 a_652_n194# a_n60_n194# 0.01fF
C2 a_296_n194# a_n594_n194# 0.01fF
C3 a_772_n140# a_950_n140# 0.13fF
C4 a_594_n140# a_60_n140# 0.04fF
C5 a_772_n140# a_n474_n140# 0.02fF
C6 a_474_n194# a_830_n194# 0.03fF
C7 a_118_n194# a_n60_n194# 0.10fF
C8 a_n830_n140# a_n652_n140# 0.13fF
C9 a_594_n140# a_n118_n140# 0.03fF
C10 a_n296_n140# a_238_n140# 0.04fF
C11 a_n652_n140# a_n1008_n140# 0.06fF
C12 a_296_n194# a_n238_n194# 0.02fF
C13 a_652_n194# a_n772_n194# 0.01fF
C14 a_416_n140# a_950_n140# 0.04fF
C15 a_n474_n140# a_416_n140# 0.02fF
C16 a_n830_n140# a_60_n140# 0.02fF
C17 a_118_n194# a_n772_n194# 0.01fF
C18 a_60_n140# a_n1008_n140# 0.02fF
C19 a_n830_n140# a_n118_n140# 0.03fF
C20 a_n416_n194# a_n594_n194# 0.10fF
C21 a_652_n194# a_n950_n194# 0.01fF
C22 a_n118_n140# a_n1008_n140# 0.02fF
C23 a_772_n140# a_n652_n140# 0.01fF
C24 a_n296_n140# a_950_n140# 0.02fF
C25 a_118_n194# a_n950_n194# 0.01fF
C26 a_474_n194# a_652_n194# 0.10fF
C27 a_n474_n140# a_n296_n140# 0.13fF
C28 a_296_n194# a_n60_n194# 0.03fF
C29 a_474_n194# a_118_n194# 0.03fF
C30 a_n238_n194# a_n416_n194# 0.10fF
C31 a_594_n140# a_n830_n140# 0.01fF
C32 a_772_n140# a_60_n140# 0.03fF
C33 a_594_n140# a_n1008_n140# 0.01fF
C34 a_416_n140# a_n652_n140# 0.02fF
C35 a_772_n140# a_n118_n140# 0.02fF
C36 a_n238_n194# a_n594_n194# 0.03fF
C37 a_296_n194# a_n772_n194# 0.01fF
C38 a_416_n140# a_60_n140# 0.06fF
C39 a_n60_n194# a_n416_n194# 0.03fF
C40 a_n830_n140# a_n1008_n140# 0.13fF
C41 a_n296_n140# a_n652_n140# 0.06fF
C42 a_652_n194# a_830_n194# 0.10fF
C43 a_594_n140# a_772_n140# 0.13fF
C44 a_296_n194# a_n950_n194# 0.01fF
C45 a_n118_n140# a_416_n140# 0.04fF
C46 a_118_n194# a_830_n194# 0.01fF
C47 a_474_n194# a_296_n194# 0.10fF
C48 a_n60_n194# a_n594_n194# 0.02fF
C49 a_n296_n140# a_60_n140# 0.06fF
C50 a_950_n140# a_238_n140# 0.03fF
C51 a_n474_n140# a_238_n140# 0.03fF
C52 a_n416_n194# a_n772_n194# 0.03fF
C53 a_594_n140# a_416_n140# 0.13fF
C54 a_n118_n140# a_n296_n140# 0.13fF
C55 a_772_n140# a_n830_n140# 0.01fF
C56 a_n60_n194# a_n238_n194# 0.10fF
C57 a_n594_n194# a_n772_n194# 0.10fF
C58 a_n416_n194# a_n950_n194# 0.02fF
C59 a_594_n140# a_n296_n140# 0.02fF
C60 a_474_n194# a_n416_n194# 0.01fF
C61 a_652_n194# a_118_n194# 0.02fF
C62 a_296_n194# a_830_n194# 0.02fF
C63 a_n830_n140# a_416_n140# 0.02fF
C64 a_n474_n140# a_950_n140# 0.01fF
C65 a_416_n140# a_n1008_n140# 0.01fF
C66 a_n594_n194# a_n950_n194# 0.03fF
C67 a_n238_n194# a_n772_n194# 0.02fF
C68 a_n652_n140# a_238_n140# 0.02fF
C69 a_474_n194# a_n594_n194# 0.01fF
C70 a_n830_n140# a_n296_n140# 0.04fF
C71 a_n238_n194# a_n950_n194# 0.01fF
C72 a_n296_n140# a_n1008_n140# 0.03fF
C73 a_60_n140# a_238_n140# 0.13fF
C74 a_474_n194# a_n238_n194# 0.01fF
C75 a_772_n140# a_416_n140# 0.06fF
C76 a_n416_n194# a_830_n194# 0.01fF
C77 a_n118_n140# a_238_n140# 0.06fF
C78 a_n60_n194# a_n772_n194# 0.01fF
C79 a_652_n194# a_296_n194# 0.03fF
C80 a_950_n140# a_n652_n140# 0.01fF
C81 a_n474_n140# a_n652_n140# 0.13fF
C82 a_118_n194# a_296_n194# 0.10fF
C83 a_772_n140# a_n296_n140# 0.02fF
C84 a_n594_n194# a_830_n194# 0.01fF
C85 a_n60_n194# a_n950_n194# 0.01fF
C86 a_594_n140# a_238_n140# 0.06fF
C87 a_60_n140# a_950_n140# 0.02fF
C88 a_n474_n140# a_60_n140# 0.04fF
C89 a_474_n194# a_n60_n194# 0.02fF
C90 a_n118_n140# a_950_n140# 0.02fF
C91 a_n474_n140# a_n118_n140# 0.06fF
C92 a_n238_n194# a_830_n194# 0.01fF
C93 a_n296_n140# a_416_n140# 0.03fF
C94 a_652_n194# a_n416_n194# 0.01fF
C95 a_n772_n194# a_n950_n194# 0.10fF
C96 a_n830_n140# a_238_n140# 0.02fF
C97 a_118_n194# a_n416_n194# 0.02fF
C98 a_474_n194# a_n772_n194# 0.01fF
C99 a_n1008_n140# a_238_n140# 0.02fF
C100 a_594_n140# a_950_n140# 0.06fF
C101 a_594_n140# a_n474_n140# 0.02fF
C102 a_652_n194# a_n594_n194# 0.01fF
C103 a_118_n194# a_n594_n194# 0.01fF
C104 a_60_n140# a_n652_n140# 0.03fF
C105 a_n60_n194# a_830_n194# 0.01fF
C106 a_474_n194# a_n950_n194# 0.01fF
C107 a_n118_n140# a_n652_n140# 0.04fF
C108 a_652_n194# a_n238_n194# 0.01fF
C109 a_772_n140# a_238_n140# 0.04fF
C110 a_n830_n140# a_n474_n140# 0.06fF
C111 a_118_n194# a_n238_n194# 0.03fF
C112 a_n474_n140# a_n1008_n140# 0.04fF
C113 a_n772_n194# a_830_n194# 0.01fF
C114 a_n118_n140# a_60_n140# 0.13fF
C115 a_296_n194# a_n416_n194# 0.01fF
C116 a_594_n140# a_n652_n140# 0.02fF
C117 a_950_n140# VSUBS 0.02fF
C118 a_772_n140# VSUBS 0.02fF
C119 a_594_n140# VSUBS 0.02fF
C120 a_416_n140# VSUBS 0.02fF
C121 a_238_n140# VSUBS 0.02fF
C122 a_60_n140# VSUBS 0.02fF
C123 a_n118_n140# VSUBS 0.02fF
C124 a_n296_n140# VSUBS 0.02fF
C125 a_n474_n140# VSUBS 0.02fF
C126 a_n652_n140# VSUBS 0.02fF
C127 a_n830_n140# VSUBS 0.02fF
C128 a_n1008_n140# VSUBS 0.02fF
C129 a_830_n194# VSUBS 0.29fF
C130 a_652_n194# VSUBS 0.23fF
C131 a_474_n194# VSUBS 0.24fF
C132 a_296_n194# VSUBS 0.25fF
C133 a_118_n194# VSUBS 0.26fF
C134 a_n60_n194# VSUBS 0.27fF
C135 a_n238_n194# VSUBS 0.28fF
C136 a_n416_n194# VSUBS 0.28fF
C137 a_n594_n194# VSUBS 0.29fF
C138 a_n772_n194# VSUBS 0.29fF
C139 a_n950_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_UFQYRB a_1751_n140# a_n149_n194# a_1987_n194# a_n2819_n194#
+ a_n207_n140# a_n1809_n140# a_n2877_n140# a_207_n194# a_n2285_n194# a_1453_n194#
+ a_n1217_n194# a_n3353_n194# a_327_n140# a_n1275_n140# a_n2343_n140# a_2521_n194#
+ a_n861_n194# a_1573_n140# a_n3411_n140# a_2641_n140# a_n2699_n140# a_2877_n194#
+ a_1809_n194# a_2997_n140# a_n29_n140# a_n1039_n194# a_n3175_n194# a_1929_n140# a_149_n140#
+ a_n1097_n140# a_2343_n194# a_1275_n194# a_29_n194# a_n2107_n194# a_n2165_n140# a_n3233_n140#
+ a_3411_n194# a_n683_n194# a_1395_n140# a_3531_n140# a_2463_n140# a_n741_n140# a_2699_n194#
+ a_741_n194# a_n3589_n140# a_n1751_n194# a_861_n140# a_1097_n194# a_2819_n140# a_3233_n194#
+ a_2165_n194# a_n3055_n140# a_n505_n194# a_2285_n140# a_n563_n140# a_563_n194# a_3353_n140#
+ a_1217_n140# a_n1573_n194# a_n2641_n194# a_683_n140# a_n919_n140# a_n1631_n140#
+ a_919_n194# a_3055_n194# a_n2997_n194# a_n1987_n140# a_n327_n194# a_n1929_n194#
+ a_3175_n140# a_1039_n140# a_n385_n140# a_385_n194# a_2107_n140# a_n1395_n194# a_n2463_n194#
+ a_n3531_n194# a_505_n140# a_n1453_n140# a_1631_n194# a_n2521_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2165_n140# a_n2285_n194# a_n2343_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_3175_n140# a_3055_n194# a_2997_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_n3233_n140# a_n3353_n194# a_n3411_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_2997_n140# a_2877_n194# a_2819_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1987_n140# a_n2107_n194# a_n2165_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X9 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1809_n140# a_n1929_n194# a_n1987_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n1453_n140# a_n1573_n194# a_n1631_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X13 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2463_n140# a_2343_n194# a_2285_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n2521_n140# a_n2641_n194# a_n2699_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X16 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_3531_n140# a_3411_n194# a_3353_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1751_n140# a_1631_n194# a_1573_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n3055_n140# a_n3175_n194# a_n3233_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_2819_n140# a_2699_n194# a_2641_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X22 a_n2877_n140# a_n2997_n194# a_n3055_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X25 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_2285_n140# a_2165_n194# a_2107_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X27 a_n2699_n140# a_n2819_n194# a_n2877_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X28 a_n2343_n140# a_n2463_n194# a_n2521_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_2107_n140# a_1987_n194# a_1929_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X31 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_3353_n140# a_3233_n194# a_3175_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X35 a_n3411_n140# a_n3531_n194# a_n3589_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X36 a_1573_n140# a_1453_n194# a_1395_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X37 a_1929_n140# a_1809_n194# a_1751_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X38 a_n1631_n140# a_n1751_n194# a_n1809_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X39 a_2641_n140# a_2521_n194# a_2463_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1631_n140# a_n2165_n140# 0.04fF
C1 a_1631_n194# a_3233_n194# 0.01fF
C2 a_n1453_n140# a_n29_n140# 0.01fF
C3 a_683_n140# a_1751_n140# 0.02fF
C4 a_n1039_n194# a_n327_n194# 0.01fF
C5 a_n1453_n140# a_n2521_n140# 0.02fF
C6 a_1751_n140# a_2463_n140# 0.03fF
C7 a_n385_n140# a_n563_n140# 0.13fF
C8 a_327_n140# a_n29_n140# 0.06fF
C9 a_2285_n140# a_2641_n140# 0.06fF
C10 a_1453_n194# a_207_n194# 0.01fF
C11 a_2107_n140# a_861_n140# 0.02fF
C12 a_683_n140# a_1217_n140# 0.04fF
C13 a_n505_n194# a_385_n194# 0.01fF
C14 a_n563_n140# a_149_n140# 0.03fF
C15 a_n505_n194# a_563_n194# 0.01fF
C16 a_n683_n194# a_n505_n194# 0.10fF
C17 a_2997_n140# a_3531_n140# 0.04fF
C18 a_1217_n140# a_2463_n140# 0.02fF
C19 a_n2285_n194# a_n861_n194# 0.01fF
C20 a_1987_n194# a_385_n194# 0.01fF
C21 a_n2819_n194# a_n3175_n194# 0.03fF
C22 a_29_n194# a_385_n194# 0.03fF
C23 a_1987_n194# a_563_n194# 0.01fF
C24 a_1929_n140# a_3531_n140# 0.01fF
C25 a_207_n194# a_n861_n194# 0.01fF
C26 a_2343_n194# a_3055_n194# 0.01fF
C27 a_n683_n194# a_29_n194# 0.01fF
C28 a_29_n194# a_563_n194# 0.02fF
C29 a_n1987_n140# a_n3411_n140# 0.01fF
C30 a_n919_n140# a_n1275_n140# 0.06fF
C31 a_n2107_n194# a_n1929_n194# 0.10fF
C32 a_n2521_n140# a_n1987_n140# 0.04fF
C33 a_n1809_n140# a_n1275_n140# 0.04fF
C34 a_n1275_n140# a_n2343_n140# 0.02fF
C35 a_1573_n140# a_861_n140# 0.03fF
C36 a_3175_n140# a_2463_n140# 0.03fF
C37 a_n741_n140# a_n919_n140# 0.13fF
C38 a_n1809_n140# a_n2877_n140# 0.02fF
C39 a_n2877_n140# a_n2343_n140# 0.04fF
C40 a_n505_n194# a_741_n194# 0.01fF
C41 a_n741_n140# a_n1809_n140# 0.02fF
C42 a_n2699_n140# a_n2165_n140# 0.04fF
C43 a_n741_n140# a_n2343_n140# 0.01fF
C44 a_1751_n140# a_1217_n140# 0.04fF
C45 a_2107_n140# a_2819_n140# 0.03fF
C46 a_1987_n194# a_741_n194# 0.01fF
C47 a_n563_n140# a_n2165_n140# 0.01fF
C48 a_29_n194# a_741_n194# 0.01fF
C49 a_1453_n194# a_2343_n194# 0.01fF
C50 a_2641_n140# a_3531_n140# 0.02fF
C51 a_n2521_n140# a_n3411_n140# 0.02fF
C52 a_n1395_n194# a_n1217_n194# 0.10fF
C53 a_3411_n194# a_2165_n194# 0.01fF
C54 a_1453_n194# a_919_n194# 0.02fF
C55 a_1751_n140# a_3175_n140# 0.01fF
C56 a_3353_n140# a_2463_n140# 0.02fF
C57 a_n207_n140# a_861_n140# 0.02fF
C58 a_1631_n194# a_3055_n194# 0.01fF
C59 a_n385_n140# a_n919_n140# 0.04fF
C60 a_n2641_n194# a_n1573_n194# 0.01fF
C61 a_n385_n140# a_n1809_n140# 0.01fF
C62 a_1573_n140# a_2819_n140# 0.02fF
C63 a_1809_n194# a_3411_n194# 0.01fF
C64 a_n919_n140# a_149_n140# 0.02fF
C65 a_n207_n140# a_n1097_n140# 0.02fF
C66 a_n149_n194# a_385_n194# 0.02fF
C67 a_n3175_n194# a_n3531_n194# 0.03fF
C68 a_1751_n140# a_3353_n140# 0.01fF
C69 a_n149_n194# a_563_n194# 0.01fF
C70 a_n683_n194# a_n149_n194# 0.02fF
C71 a_1453_n194# a_1631_n194# 0.10fF
C72 a_n505_n194# a_n1751_n194# 0.01fF
C73 a_1275_n194# a_2165_n194# 0.01fF
C74 a_1039_n140# a_1395_n140# 0.06fF
C75 a_n2877_n140# a_n3233_n140# 0.06fF
C76 a_n2819_n194# a_n2107_n194# 0.01fF
C77 a_1097_n194# a_1453_n194# 0.03fF
C78 a_n861_n194# a_n1395_n194# 0.02fF
C79 a_1275_n194# a_1809_n194# 0.02fF
C80 a_683_n140# a_505_n140# 0.13fF
C81 a_n149_n194# a_741_n194# 0.01fF
C82 a_n919_n140# a_n2165_n140# 0.02fF
C83 a_2877_n194# a_3411_n194# 0.02fF
C84 a_n2165_n140# a_n2343_n140# 0.13fF
C85 a_n1809_n140# a_n2165_n140# 0.06fF
C86 a_3353_n140# a_3175_n140# 0.13fF
C87 a_327_n140# a_1573_n140# 0.02fF
C88 a_3233_n194# a_2165_n194# 0.01fF
C89 a_n2107_n194# a_n683_n194# 0.01fF
C90 a_n3175_n194# a_n1751_n194# 0.01fF
C91 a_n1039_n194# a_n2641_n194# 0.01fF
C92 a_n2819_n194# a_n1929_n194# 0.01fF
C93 a_n385_n140# a_1039_n140# 0.01fF
C94 a_683_n140# a_1929_n140# 0.02fF
C95 a_1809_n194# a_3233_n194# 0.01fF
C96 a_2285_n140# a_1039_n140# 0.02fF
C97 a_1751_n140# a_505_n140# 0.02fF
C98 a_2463_n140# a_2997_n140# 0.04fF
C99 a_1039_n140# a_149_n140# 0.02fF
C100 a_n207_n140# a_n1453_n140# 0.02fF
C101 a_n505_n194# a_207_n194# 0.01fF
C102 a_1275_n194# a_2877_n194# 0.01fF
C103 a_1929_n140# a_2463_n140# 0.04fF
C104 a_n1573_n194# a_n1217_n194# 0.03fF
C105 a_327_n140# a_n207_n140# 0.04fF
C106 a_29_n194# a_207_n194# 0.10fF
C107 a_n2107_n194# a_n3531_n194# 0.01fF
C108 a_1217_n140# a_505_n140# 0.03fF
C109 a_n149_n194# a_n1751_n194# 0.01fF
C110 a_n1631_n140# a_n3055_n140# 0.01fF
C111 a_n683_n194# a_n1929_n194# 0.01fF
C112 a_1751_n140# a_2997_n140# 0.02fF
C113 a_683_n140# a_n563_n140# 0.02fF
C114 a_1929_n140# a_1751_n140# 0.13fF
C115 a_n2463_n194# a_n2641_n194# 0.10fF
C116 a_2641_n140# a_2463_n140# 0.13fF
C117 a_1573_n140# a_n29_n140# 0.01fF
C118 a_n3233_n140# a_n2165_n140# 0.02fF
C119 a_n2285_n194# a_n3175_n194# 0.01fF
C120 a_n3175_n194# a_n2997_n194# 0.10fF
C121 a_2877_n194# a_3233_n194# 0.03fF
C122 a_1275_n194# a_n327_n194# 0.01fF
C123 a_1929_n140# a_1217_n140# 0.03fF
C124 a_861_n140# a_1395_n140# 0.04fF
C125 a_n505_n194# a_919_n194# 0.01fF
C126 a_n3531_n194# a_n1929_n194# 0.01fF
C127 a_3055_n194# a_2165_n194# 0.01fF
C128 a_n861_n194# a_n1573_n194# 0.01fF
C129 a_1987_n194# a_2343_n194# 0.03fF
C130 a_3175_n140# a_2997_n140# 0.13fF
C131 a_1751_n140# a_2641_n140# 0.02fF
C132 a_n741_n140# a_861_n140# 0.01fF
C133 a_1929_n140# a_3175_n140# 0.02fF
C134 a_n207_n140# a_n29_n140# 0.13fF
C135 a_1987_n194# a_919_n194# 0.01fF
C136 a_n2107_n194# a_n1751_n194# 0.03fF
C137 a_29_n194# a_919_n194# 0.01fF
C138 a_1809_n194# a_3055_n194# 0.01fF
C139 a_n1275_n140# a_n1097_n140# 0.13fF
C140 a_n2699_n140# a_n3055_n140# 0.06fF
C141 a_n149_n194# a_207_n194# 0.03fF
C142 a_n1039_n194# a_n1217_n194# 0.10fF
C143 a_1217_n140# a_2641_n140# 0.01fF
C144 a_n741_n140# a_n1097_n140# 0.06fF
C145 a_n505_n194# a_n1395_n194# 0.01fF
C146 a_1453_n194# a_2165_n194# 0.01fF
C147 a_2699_n194# a_2343_n194# 0.03fF
C148 a_3353_n140# a_2997_n140# 0.06fF
C149 a_1929_n140# a_3353_n140# 0.01fF
C150 a_683_n140# a_n919_n140# 0.01fF
C151 a_2819_n140# a_1395_n140# 0.01fF
C152 a_29_n194# a_n1395_n194# 0.01fF
C153 a_n3353_n194# a_n3175_n194# 0.10fF
C154 a_1809_n194# a_1453_n194# 0.03fF
C155 a_3175_n140# a_2641_n140# 0.04fF
C156 a_1987_n194# a_1631_n194# 0.03fF
C157 a_861_n140# a_n385_n140# 0.02fF
C158 a_29_n194# a_1631_n194# 0.01fF
C159 a_1097_n194# a_n505_n194# 0.01fF
C160 a_861_n140# a_2285_n140# 0.01fF
C161 a_861_n140# a_149_n140# 0.03fF
C162 a_n1929_n194# a_n1751_n194# 0.10fF
C163 a_1097_n194# a_1987_n194# 0.01fF
C164 a_n2877_n140# a_n3589_n140# 0.03fF
C165 a_1097_n194# a_29_n194# 0.01fF
C166 a_n385_n140# a_n1097_n140# 0.03fF
C167 a_2877_n194# a_3055_n194# 0.10fF
C168 a_n2285_n194# a_n2107_n194# 0.10fF
C169 a_2699_n194# a_1631_n194# 0.01fF
C170 a_n2463_n194# a_n1217_n194# 0.01fF
C171 a_n2107_n194# a_n2997_n194# 0.01fF
C172 a_3353_n140# a_2641_n140# 0.03fF
C173 a_385_n194# a_563_n194# 0.10fF
C174 a_n1097_n140# a_149_n140# 0.02fF
C175 a_n1039_n194# a_n861_n194# 0.10fF
C176 a_n683_n194# a_385_n194# 0.01fF
C177 a_n2819_n194# a_n3531_n194# 0.01fF
C178 a_n683_n194# a_563_n194# 0.01fF
C179 a_n149_n194# a_919_n194# 0.01fF
C180 a_1097_n194# a_2699_n194# 0.01fF
C181 a_2107_n140# a_1573_n140# 0.04fF
C182 a_2285_n140# a_2819_n140# 0.04fF
C183 a_1453_n194# a_2877_n194# 0.01fF
C184 a_n1453_n140# a_n1275_n140# 0.13fF
C185 a_385_n194# a_741_n194# 0.03fF
C186 a_n1453_n140# a_n2877_n140# 0.01fF
C187 a_n741_n140# a_n1453_n140# 0.03fF
C188 a_563_n194# a_741_n194# 0.10fF
C189 a_1929_n140# a_505_n140# 0.01fF
C190 a_n683_n194# a_741_n194# 0.01fF
C191 a_327_n140# a_1395_n140# 0.02fF
C192 a_n149_n194# a_n1395_n194# 0.01fF
C193 a_n327_n194# a_n1217_n194# 0.01fF
C194 a_327_n140# a_n1275_n140# 0.01fF
C195 a_n2285_n194# a_n1929_n194# 0.03fF
C196 a_n1809_n140# a_n3055_n140# 0.02fF
C197 a_n3055_n140# a_n2343_n140# 0.03fF
C198 a_n1929_n194# a_n2997_n194# 0.01fF
C199 a_n741_n140# a_327_n140# 0.02fF
C200 a_n2165_n140# a_n1097_n140# 0.02fF
C201 a_683_n140# a_1039_n140# 0.06fF
C202 a_n2463_n194# a_n861_n194# 0.01fF
C203 a_3233_n194# a_3411_n194# 0.10fF
C204 a_n3353_n194# a_n2107_n194# 0.01fF
C205 a_1097_n194# a_n149_n194# 0.01fF
C206 a_n1631_n140# a_n2699_n140# 0.02fF
C207 a_n2819_n194# a_n1751_n194# 0.01fF
C208 a_2463_n140# a_1039_n140# 0.01fF
C209 a_1929_n140# a_2997_n140# 0.02fF
C210 a_n505_n194# a_n1573_n194# 0.01fF
C211 a_n563_n140# a_505_n140# 0.02fF
C212 a_n1453_n140# a_n385_n140# 0.02fF
C213 a_n1987_n140# a_n1275_n140# 0.03fF
C214 a_n563_n140# a_n1631_n140# 0.02fF
C215 a_n1987_n140# a_n2877_n140# 0.02fF
C216 a_2521_n194# a_2343_n194# 0.10fF
C217 a_2819_n140# a_3531_n140# 0.03fF
C218 a_n741_n140# a_n1987_n140# 0.02fF
C219 a_n1453_n140# a_149_n140# 0.01fF
C220 a_327_n140# a_n385_n140# 0.03fF
C221 a_2521_n194# a_919_n194# 0.01fF
C222 a_29_n194# a_n1573_n194# 0.01fF
C223 a_n2165_n140# a_n3589_n140# 0.01fF
C224 a_n327_n194# a_n861_n194# 0.02fF
C225 a_n2107_n194# a_n1395_n194# 0.01fF
C226 a_1751_n140# a_1039_n140# 0.03fF
C227 a_327_n140# a_149_n140# 0.13fF
C228 a_n29_n140# a_1395_n140# 0.01fF
C229 a_2641_n140# a_2997_n140# 0.06fF
C230 a_n29_n140# a_n1275_n140# 0.02fF
C231 a_n683_n194# a_n1751_n194# 0.01fF
C232 a_n2877_n140# a_n3411_n140# 0.04fF
C233 a_n2521_n140# a_n1275_n140# 0.02fF
C234 a_n3353_n194# a_n1929_n194# 0.01fF
C235 a_n741_n140# a_n29_n140# 0.03fF
C236 a_n2521_n140# a_n2877_n140# 0.06fF
C237 a_1929_n140# a_2641_n140# 0.03fF
C238 a_1217_n140# a_1039_n140# 0.13fF
C239 a_n3055_n140# a_n3233_n140# 0.13fF
C240 a_n385_n140# a_n1987_n140# 0.01fF
C241 a_2521_n194# a_1631_n194# 0.01fF
C242 a_n3175_n194# a_n1573_n194# 0.01fF
C243 a_n2819_n194# a_n2285_n194# 0.02fF
C244 a_n2819_n194# a_n2997_n194# 0.10fF
C245 a_n1453_n140# a_n2165_n140# 0.03fF
C246 a_1987_n194# a_2165_n194# 0.10fF
C247 a_1097_n194# a_2521_n194# 0.01fF
C248 a_n1929_n194# a_n1395_n194# 0.02fF
C249 a_3055_n194# a_3411_n194# 0.03fF
C250 a_n385_n140# a_n29_n140# 0.06fF
C251 a_n919_n140# a_505_n140# 0.01fF
C252 a_n1039_n194# a_n505_n194# 0.02fF
C253 a_1987_n194# a_1809_n194# 0.10fF
C254 a_n1631_n140# a_n919_n140# 0.03fF
C255 a_n1631_n140# a_n1809_n140# 0.13fF
C256 a_n1631_n140# a_n2343_n140# 0.03fF
C257 a_n29_n140# a_149_n140# 0.13fF
C258 a_n149_n194# a_n1573_n194# 0.01fF
C259 a_n2285_n194# a_n683_n194# 0.01fF
C260 a_385_n194# a_207_n194# 0.10fF
C261 a_n1039_n194# a_29_n194# 0.01fF
C262 a_2699_n194# a_2165_n194# 0.02fF
C263 a_207_n194# a_563_n194# 0.03fF
C264 a_n683_n194# a_207_n194# 0.01fF
C265 a_n1987_n140# a_n2165_n140# 0.13fF
C266 a_683_n140# a_861_n140# 0.13fF
C267 a_2699_n194# a_1809_n194# 0.01fF
C268 a_n3353_n194# a_n2819_n194# 0.02fF
C269 a_861_n140# a_2463_n140# 0.01fF
C270 a_207_n194# a_741_n194# 0.02fF
C271 a_n2285_n194# a_n3531_n194# 0.01fF
C272 a_n3531_n194# a_n2997_n194# 0.02fF
C273 a_n2165_n140# a_n3411_n140# 0.02fF
C274 a_1987_n194# a_2877_n194# 0.01fF
C275 a_n2521_n140# a_n2165_n140# 0.06fF
C276 a_n2641_n194# a_n1217_n194# 0.01fF
C277 a_n2107_n194# a_n1573_n194# 0.02fF
C278 a_1275_n194# a_1453_n194# 0.10fF
C279 a_1751_n140# a_861_n140# 0.02fF
C280 a_n1809_n140# a_n2699_n140# 0.02fF
C281 a_n2699_n140# a_n2343_n140# 0.06fF
C282 a_2107_n140# a_1395_n140# 0.03fF
C283 a_n2819_n194# a_n1395_n194# 0.01fF
C284 a_385_n194# a_919_n194# 0.02fF
C285 a_n563_n140# a_n919_n140# 0.06fF
C286 a_563_n194# a_919_n194# 0.03fF
C287 a_n683_n194# a_919_n194# 0.01fF
C288 a_n563_n140# a_n1809_n140# 0.02fF
C289 a_n1631_n140# a_n3233_n140# 0.01fF
C290 a_2463_n140# a_2819_n140# 0.06fF
C291 a_3055_n194# a_3233_n194# 0.10fF
C292 a_2699_n194# a_2877_n194# 0.10fF
C293 a_1039_n140# a_505_n140# 0.04fF
C294 a_n1039_n194# a_n149_n194# 0.01fF
C295 a_861_n140# a_1217_n140# 0.06fF
C296 a_n327_n194# a_n505_n194# 0.10fF
C297 a_2343_n194# a_741_n194# 0.01fF
C298 a_n3175_n194# a_n2463_n194# 0.01fF
C299 a_1573_n140# a_1395_n140# 0.13fF
C300 a_n327_n194# a_29_n194# 0.03fF
C301 a_n2285_n194# a_n1751_n194# 0.02fF
C302 a_919_n194# a_741_n194# 0.10fF
C303 a_1631_n194# a_385_n194# 0.01fF
C304 a_n683_n194# a_n1395_n194# 0.01fF
C305 a_n1751_n194# a_n2997_n194# 0.01fF
C306 a_n1929_n194# a_n1573_n194# 0.03fF
C307 a_1751_n140# a_2819_n140# 0.02fF
C308 a_n3353_n194# a_n3531_n194# 0.10fF
C309 a_1631_n194# a_563_n194# 0.01fF
C310 a_2107_n140# a_2285_n140# 0.13fF
C311 a_1929_n140# a_1039_n140# 0.02fF
C312 a_1097_n194# a_385_n194# 0.01fF
C313 a_1097_n194# a_563_n194# 0.02fF
C314 a_1217_n140# a_2819_n140# 0.01fF
C315 a_n207_n140# a_1395_n140# 0.01fF
C316 a_2521_n194# a_2165_n194# 0.03fF
C317 a_683_n140# a_327_n140# 0.06fF
C318 a_n207_n140# a_n1275_n140# 0.02fF
C319 a_n1039_n194# a_n2107_n194# 0.01fF
C320 a_1631_n194# a_741_n194# 0.01fF
C321 a_n2699_n140# a_n3233_n140# 0.04fF
C322 a_n741_n140# a_n207_n140# 0.04fF
C323 a_3175_n140# a_2819_n140# 0.06fF
C324 a_2521_n194# a_1809_n194# 0.01fF
C325 a_1573_n140# a_2285_n140# 0.03fF
C326 a_n3055_n140# a_n3589_n140# 0.04fF
C327 a_n919_n140# a_n1809_n140# 0.02fF
C328 a_1573_n140# a_149_n140# 0.01fF
C329 a_n919_n140# a_n2343_n140# 0.01fF
C330 a_2641_n140# a_1039_n140# 0.01fF
C331 a_1097_n194# a_741_n194# 0.03fF
C332 a_n1809_n140# a_n2343_n140# 0.04fF
C333 a_n563_n140# a_1039_n140# 0.01fF
C334 a_n2285_n194# a_n2997_n194# 0.01fF
C335 a_n3353_n194# a_n1751_n194# 0.01fF
C336 a_n149_n194# a_n327_n194# 0.10fF
C337 a_327_n140# a_1751_n140# 0.01fF
C338 a_2107_n140# a_3531_n140# 0.01fF
C339 a_3353_n140# a_2819_n140# 0.04fF
C340 a_n207_n140# a_n385_n140# 0.13fF
C341 a_n1039_n194# a_n1929_n194# 0.01fF
C342 a_n2819_n194# a_n1573_n194# 0.01fF
C343 a_n2107_n194# a_n2463_n194# 0.03fF
C344 a_n207_n140# a_149_n140# 0.06fF
C345 a_n1453_n140# a_n3055_n140# 0.01fF
C346 a_1453_n194# a_3055_n194# 0.01fF
C347 a_683_n140# a_n29_n140# 0.03fF
C348 a_327_n140# a_1217_n140# 0.02fF
C349 a_2521_n194# a_2877_n194# 0.03fF
C350 a_n1751_n194# a_n1395_n194# 0.03fF
C351 a_861_n140# a_505_n140# 0.06fF
C352 a_1987_n194# a_3411_n194# 0.01fF
C353 a_n861_n194# a_n1217_n194# 0.03fF
C354 a_505_n140# a_n1097_n140# 0.01fF
C355 a_n683_n194# a_n1573_n194# 0.01fF
C356 a_n3353_n194# a_n2285_n194# 0.01fF
C357 a_n1631_n140# a_n1097_n140# 0.04fF
C358 a_n3353_n194# a_n2997_n194# 0.03fF
C359 a_n2463_n194# a_n1929_n194# 0.02fF
C360 a_2699_n194# a_3411_n194# 0.01fF
C361 a_n3233_n140# a_n2343_n140# 0.02fF
C362 a_n1809_n140# a_n3233_n140# 0.01fF
C363 a_207_n194# a_919_n194# 0.01fF
C364 a_n1987_n140# a_n3055_n140# 0.02fF
C365 a_1929_n140# a_861_n140# 0.02fF
C366 a_1275_n194# a_1987_n194# 0.01fF
C367 a_1275_n194# a_29_n194# 0.01fF
C368 a_n2285_n194# a_n1395_n194# 0.01fF
C369 a_1217_n140# a_n29_n140# 0.02fF
C370 a_n3055_n140# a_n3411_n140# 0.06fF
C371 a_n2997_n194# a_n1395_n194# 0.01fF
C372 a_207_n194# a_n1395_n194# 0.01fF
C373 a_n2521_n140# a_n3055_n140# 0.04fF
C374 a_1631_n194# a_207_n194# 0.01fF
C375 a_n327_n194# a_n1929_n194# 0.01fF
C376 a_1275_n194# a_2699_n194# 0.01fF
C377 a_563_n194# a_2165_n194# 0.01fF
C378 a_861_n140# a_n563_n140# 0.01fF
C379 a_2819_n140# a_2997_n140# 0.13fF
C380 a_1929_n140# a_2819_n140# 0.02fF
C381 a_1809_n194# a_385_n194# 0.01fF
C382 a_n2699_n140# a_n1097_n140# 0.01fF
C383 a_1987_n194# a_3233_n194# 0.01fF
C384 a_1097_n194# a_207_n194# 0.01fF
C385 a_2343_n194# a_919_n194# 0.01fF
C386 a_1809_n194# a_563_n194# 0.01fF
C387 a_n1039_n194# a_385_n194# 0.01fF
C388 a_n1039_n194# a_n683_n194# 0.03fF
C389 a_n1039_n194# a_563_n194# 0.01fF
C390 a_n563_n140# a_n1097_n140# 0.04fF
C391 a_2165_n194# a_741_n194# 0.01fF
C392 a_n1453_n140# a_n1631_n140# 0.13fF
C393 a_n3175_n194# a_n2641_n194# 0.02fF
C394 a_n1275_n140# a_n2877_n140# 0.01fF
C395 a_n741_n140# a_n1275_n140# 0.04fF
C396 a_n2819_n194# a_n2463_n194# 0.03fF
C397 a_327_n140# a_505_n140# 0.13fF
C398 a_1275_n194# a_n149_n194# 0.01fF
C399 a_2107_n140# a_683_n140# 0.01fF
C400 a_2699_n194# a_3233_n194# 0.02fF
C401 a_1809_n194# a_741_n194# 0.01fF
C402 a_n1751_n194# a_n1573_n194# 0.10fF
C403 a_2641_n140# a_2819_n140# 0.13fF
C404 a_1631_n194# a_2343_n194# 0.01fF
C405 a_n2699_n140# a_n3589_n140# 0.02fF
C406 a_2107_n140# a_2463_n140# 0.06fF
C407 a_1631_n194# a_919_n194# 0.01fF
C408 a_1097_n194# a_2343_n194# 0.01fF
C409 a_n385_n140# a_n1275_n140# 0.02fF
C410 a_2285_n140# a_1395_n140# 0.02fF
C411 a_683_n140# a_1573_n140# 0.02fF
C412 a_1097_n194# a_919_n194# 0.10fF
C413 a_n1631_n140# a_n1987_n140# 0.06fF
C414 a_1395_n140# a_149_n140# 0.02fF
C415 a_n741_n140# a_n385_n140# 0.06fF
C416 a_2521_n194# a_3411_n194# 0.01fF
C417 a_1929_n140# a_327_n140# 0.01fF
C418 a_n1275_n140# a_149_n140# 0.01fF
C419 a_1573_n140# a_2463_n140# 0.02fF
C420 a_2107_n140# a_1751_n140# 0.06fF
C421 a_n505_n194# a_n1217_n194# 0.01fF
C422 a_n741_n140# a_149_n140# 0.02fF
C423 a_n1453_n140# a_n2699_n140# 0.02fF
C424 a_29_n194# a_n1217_n194# 0.01fF
C425 a_1987_n194# a_3055_n194# 0.01fF
C426 a_n29_n140# a_505_n140# 0.04fF
C427 a_n919_n140# a_n1097_n140# 0.13fF
C428 a_n1631_n140# a_n29_n140# 0.01fF
C429 a_n2285_n194# a_n1573_n194# 0.01fF
C430 a_n1453_n140# a_n563_n140# 0.02fF
C431 a_2107_n140# a_1217_n140# 0.02fF
C432 a_n1809_n140# a_n1097_n140# 0.03fF
C433 a_n2343_n140# a_n1097_n140# 0.02fF
C434 a_683_n140# a_n207_n140# 0.02fF
C435 a_n2997_n194# a_n1573_n194# 0.01fF
C436 a_n1631_n140# a_n2521_n140# 0.02fF
C437 a_1097_n194# a_1631_n194# 0.02fF
C438 a_n3531_n194# a_n2463_n194# 0.01fF
C439 a_n327_n194# a_385_n194# 0.01fF
C440 a_1573_n140# a_1751_n140# 0.13fF
C441 a_n683_n194# a_n327_n194# 0.03fF
C442 a_n327_n194# a_563_n194# 0.01fF
C443 a_1275_n194# a_2521_n194# 0.01fF
C444 a_327_n140# a_n563_n140# 0.02fF
C445 a_n1039_n194# a_n1751_n194# 0.01fF
C446 a_n2107_n194# a_n2641_n194# 0.02fF
C447 a_2107_n140# a_3175_n140# 0.02fF
C448 a_n385_n140# a_149_n140# 0.04fF
C449 a_n1275_n140# a_n2165_n140# 0.02fF
C450 a_1987_n194# a_1453_n194# 0.02fF
C451 a_2699_n194# a_3055_n194# 0.03fF
C452 a_n2877_n140# a_n2165_n140# 0.03fF
C453 a_29_n194# a_1453_n194# 0.01fF
C454 a_n741_n140# a_n2165_n140# 0.01fF
C455 a_1573_n140# a_1217_n140# 0.06fF
C456 a_n1987_n140# a_n2699_n140# 0.03fF
C457 a_n505_n194# a_n861_n194# 0.03fF
C458 a_n2343_n140# a_n3589_n140# 0.02fF
C459 a_n327_n194# a_741_n194# 0.01fF
C460 a_n563_n140# a_n1987_n140# 0.01fF
C461 a_29_n194# a_n861_n194# 0.01fF
C462 a_1573_n140# a_3175_n140# 0.01fF
C463 a_2107_n140# a_3353_n140# 0.02fF
C464 a_2699_n194# a_1453_n194# 0.01fF
C465 a_2521_n194# a_3233_n194# 0.01fF
C466 a_n2699_n140# a_n3411_n140# 0.03fF
C467 a_861_n140# a_1039_n140# 0.13fF
C468 a_n2641_n194# a_n1929_n194# 0.01fF
C469 a_n2521_n140# a_n2699_n140# 0.13fF
C470 a_n2463_n194# a_n1751_n194# 0.01fF
C471 a_n149_n194# a_n1217_n194# 0.01fF
C472 a_n207_n140# a_1217_n140# 0.01fF
C473 a_1809_n194# a_207_n194# 0.01fF
C474 a_n563_n140# a_n29_n140# 0.04fF
C475 a_n2285_n194# a_n1039_n194# 0.01fF
C476 a_n1453_n140# a_n919_n140# 0.04fF
C477 a_2285_n140# a_3531_n140# 0.02fF
C478 a_n1453_n140# a_n1809_n140# 0.06fF
C479 a_n1039_n194# a_207_n194# 0.01fF
C480 a_n1453_n140# a_n2343_n140# 0.02fF
C481 a_327_n140# a_n919_n140# 0.02fF
C482 a_n1573_n194# a_n1395_n194# 0.10fF
C483 a_n149_n194# a_1453_n194# 0.01fF
C484 a_n327_n194# a_n1751_n194# 0.01fF
C485 a_2343_n194# a_2165_n194# 0.10fF
C486 a_n3233_n140# a_n3589_n140# 0.06fF
C487 a_2107_n140# a_505_n140# 0.01fF
C488 a_n149_n194# a_n861_n194# 0.01fF
C489 a_919_n194# a_2165_n194# 0.01fF
C490 a_n2107_n194# a_n1217_n194# 0.01fF
C491 a_n919_n140# a_n1987_n140# 0.02fF
C492 a_1809_n194# a_2343_n194# 0.02fF
C493 a_n2285_n194# a_n2463_n194# 0.10fF
C494 a_n1809_n140# a_n1987_n140# 0.13fF
C495 a_n1987_n140# a_n2343_n140# 0.06fF
C496 a_n2463_n194# a_n2997_n194# 0.02fF
C497 a_1809_n194# a_919_n194# 0.01fF
C498 a_2521_n194# a_3055_n194# 0.02fF
C499 a_n2819_n194# a_n2641_n194# 0.10fF
C500 a_1573_n140# a_505_n140# 0.02fF
C501 a_2107_n140# a_2997_n140# 0.02fF
C502 a_n919_n140# a_n29_n140# 0.02fF
C503 a_n1809_n140# a_n3411_n140# 0.01fF
C504 a_1275_n194# a_385_n194# 0.01fF
C505 a_1631_n194# a_2165_n194# 0.02fF
C506 a_n2343_n140# a_n3411_n140# 0.02fF
C507 a_n919_n140# a_n2521_n140# 0.01fF
C508 a_1275_n194# a_563_n194# 0.01fF
C509 a_2107_n140# a_1929_n140# 0.13fF
C510 a_n1809_n140# a_n2521_n140# 0.03fF
C511 a_n2521_n140# a_n2343_n140# 0.13fF
C512 a_683_n140# a_1395_n140# 0.03fF
C513 a_n1929_n194# a_n1217_n194# 0.01fF
C514 a_1809_n194# a_1631_n194# 0.10fF
C515 a_1097_n194# a_2165_n194# 0.01fF
C516 a_2521_n194# a_1453_n194# 0.01fF
C517 a_n327_n194# a_207_n194# 0.02fF
C518 a_n1039_n194# a_n1395_n194# 0.03fF
C519 a_n741_n140# a_683_n140# 0.01fF
C520 a_n2107_n194# a_n861_n194# 0.01fF
C521 a_327_n140# a_1039_n140# 0.03fF
C522 a_2343_n194# a_2877_n194# 0.02fF
C523 a_2463_n140# a_1395_n140# 0.02fF
C524 a_1573_n140# a_2997_n140# 0.01fF
C525 a_n207_n140# a_505_n140# 0.03fF
C526 a_1097_n194# a_1809_n194# 0.01fF
C527 a_1275_n194# a_741_n194# 0.02fF
C528 a_n207_n140# a_n1631_n140# 0.01fF
C529 a_1929_n140# a_1573_n140# 0.06fF
C530 a_n3353_n194# a_n2463_n194# 0.01fF
C531 a_2107_n140# a_2641_n140# 0.04fF
C532 a_29_n194# a_n505_n194# 0.02fF
C533 a_n1987_n140# a_n3233_n140# 0.02fF
C534 a_1751_n140# a_1395_n140# 0.06fF
C535 a_683_n140# a_n385_n140# 0.02fF
C536 a_n3531_n194# a_n2641_n194# 0.01fF
C537 a_683_n140# a_2285_n140# 0.01fF
C538 a_1631_n194# a_2877_n194# 0.01fF
C539 a_n861_n194# a_n1929_n194# 0.01fF
C540 a_1573_n140# a_2641_n140# 0.02fF
C541 a_683_n140# a_149_n140# 0.04fF
C542 a_n2463_n194# a_n1395_n194# 0.01fF
C543 a_1217_n140# a_1395_n140# 0.13fF
C544 a_n3233_n140# a_n3411_n140# 0.13fF
C545 a_2285_n140# a_2463_n140# 0.13fF
C546 a_n327_n194# a_919_n194# 0.01fF
C547 a_2699_n194# a_1987_n194# 0.01fF
C548 a_n2521_n140# a_n3233_n140# 0.03fF
C549 a_1039_n140# a_n29_n140# 0.02fF
C550 a_n2877_n140# a_n3055_n140# 0.13fF
C551 a_n2819_n194# a_n1217_n194# 0.01fF
C552 a_1751_n140# a_2285_n140# 0.04fF
C553 a_n207_n140# a_n563_n140# 0.06fF
C554 a_n327_n194# a_n1395_n194# 0.01fF
C555 a_1751_n140# a_149_n140# 0.01fF
C556 a_n149_n194# a_n505_n194# 0.03fF
C557 a_n2641_n194# a_n1751_n194# 0.01fF
C558 a_1217_n140# a_n385_n140# 0.01fF
C559 a_n149_n194# a_29_n194# 0.10fF
C560 a_385_n194# a_n1217_n194# 0.01fF
C561 a_1217_n140# a_2285_n140# 0.02fF
C562 a_1097_n194# a_n327_n194# 0.01fF
C563 a_n683_n194# a_n1217_n194# 0.02fF
C564 a_1217_n140# a_149_n140# 0.02fF
C565 a_2463_n140# a_3531_n140# 0.02fF
C566 a_n1039_n194# a_n1573_n194# 0.02fF
C567 a_327_n140# a_861_n140# 0.04fF
C568 a_3175_n140# a_2285_n140# 0.02fF
C569 a_n1453_n140# a_n1097_n140# 0.06fF
C570 a_1453_n194# a_385_n194# 0.01fF
C571 a_1453_n194# a_563_n194# 0.01fF
C572 a_327_n140# a_n1097_n140# 0.01fF
C573 a_1275_n194# a_207_n194# 0.01fF
C574 a_n2107_n194# a_n505_n194# 0.01fF
C575 a_2343_n194# a_3411_n194# 0.01fF
C576 a_3353_n140# a_2285_n140# 0.02fF
C577 a_1809_n194# a_2165_n194# 0.03fF
C578 a_n2285_n194# a_n2641_n194# 0.03fF
C579 a_385_n194# a_n861_n194# 0.01fF
C580 a_n207_n140# a_n919_n140# 0.03fF
C581 a_n861_n194# a_563_n194# 0.01fF
C582 a_n683_n194# a_n861_n194# 0.10fF
C583 a_n3055_n140# a_n2165_n140# 0.02fF
C584 a_n2641_n194# a_n2997_n194# 0.03fF
C585 a_n2463_n194# a_n1573_n194# 0.01fF
C586 a_n207_n140# a_n1809_n140# 0.01fF
C587 a_1453_n194# a_741_n194# 0.01fF
C588 a_1395_n140# a_505_n140# 0.02fF
C589 a_n1987_n140# a_n1097_n140# 0.02fF
C590 a_n1631_n140# a_n1275_n140# 0.06fF
C591 a_2521_n194# a_1987_n194# 0.02fF
C592 a_n1631_n140# a_n2877_n140# 0.02fF
C593 a_861_n140# a_n29_n140# 0.02fF
C594 a_n741_n140# a_505_n140# 0.02fF
C595 a_3175_n140# a_3531_n140# 0.06fF
C596 a_2107_n140# a_1039_n140# 0.02fF
C597 a_n741_n140# a_n1631_n140# 0.02fF
C598 a_n861_n194# a_741_n194# 0.01fF
C599 a_n505_n194# a_n1929_n194# 0.01fF
C600 a_1275_n194# a_2343_n194# 0.01fF
C601 a_n3175_n194# a_n2107_n194# 0.01fF
C602 a_n29_n140# a_n1097_n140# 0.02fF
C603 a_n1751_n194# a_n1217_n194# 0.02fF
C604 a_1275_n194# a_919_n194# 0.03fF
C605 a_2997_n140# a_1395_n140# 0.01fF
C606 a_n2521_n140# a_n1097_n140# 0.01fF
C607 a_2699_n194# a_2521_n194# 0.10fF
C608 a_n327_n194# a_n1573_n194# 0.01fF
C609 a_1929_n140# a_1395_n140# 0.04fF
C610 a_2877_n194# a_2165_n194# 0.01fF
C611 a_n1987_n140# a_n3589_n140# 0.01fF
C612 a_1573_n140# a_1039_n140# 0.04fF
C613 a_3353_n140# a_3531_n140# 0.13fF
C614 a_n385_n140# a_505_n140# 0.02fF
C615 a_n385_n140# a_n1631_n140# 0.02fF
C616 a_n3353_n194# a_n2641_n194# 0.01fF
C617 a_1809_n194# a_2877_n194# 0.01fF
C618 a_505_n140# a_149_n140# 0.06fF
C619 a_1275_n194# a_1631_n194# 0.03fF
C620 a_n1275_n140# a_n2699_n140# 0.01fF
C621 a_2343_n194# a_3233_n194# 0.01fF
C622 a_n3411_n140# a_n3589_n140# 0.13fF
C623 a_n3175_n194# a_n1929_n194# 0.01fF
C624 a_n2877_n140# a_n2699_n140# 0.13fF
C625 a_n1039_n194# a_n2463_n194# 0.01fF
C626 a_n2521_n140# a_n3589_n140# 0.02fF
C627 a_2641_n140# a_1395_n140# 0.02fF
C628 a_n207_n140# a_1039_n140# 0.02fF
C629 a_n563_n140# a_n1275_n140# 0.03fF
C630 a_1275_n194# a_1097_n194# 0.10fF
C631 a_n1453_n140# a_n1987_n140# 0.04fF
C632 a_2285_n140# a_2997_n140# 0.03fF
C633 a_n861_n194# a_n1751_n194# 0.01fF
C634 a_n2641_n194# a_n1395_n194# 0.01fF
C635 a_n741_n140# a_n563_n140# 0.13fF
C636 a_n2285_n194# a_n1217_n194# 0.01fF
C637 a_1929_n140# a_2285_n140# 0.06fF
C638 a_207_n194# a_n1217_n194# 0.01fF
C639 a_3531_n140# VSUBS 0.02fF
C640 a_3353_n140# VSUBS 0.02fF
C641 a_3175_n140# VSUBS 0.02fF
C642 a_2997_n140# VSUBS 0.02fF
C643 a_2819_n140# VSUBS 0.02fF
C644 a_2641_n140# VSUBS 0.02fF
C645 a_2463_n140# VSUBS 0.02fF
C646 a_2285_n140# VSUBS 0.02fF
C647 a_2107_n140# VSUBS 0.02fF
C648 a_1929_n140# VSUBS 0.02fF
C649 a_1751_n140# VSUBS 0.02fF
C650 a_1573_n140# VSUBS 0.02fF
C651 a_1395_n140# VSUBS 0.02fF
C652 a_1217_n140# VSUBS 0.02fF
C653 a_1039_n140# VSUBS 0.02fF
C654 a_861_n140# VSUBS 0.02fF
C655 a_683_n140# VSUBS 0.02fF
C656 a_505_n140# VSUBS 0.02fF
C657 a_327_n140# VSUBS 0.02fF
C658 a_149_n140# VSUBS 0.02fF
C659 a_n29_n140# VSUBS 0.02fF
C660 a_n207_n140# VSUBS 0.02fF
C661 a_n385_n140# VSUBS 0.02fF
C662 a_n563_n140# VSUBS 0.02fF
C663 a_n741_n140# VSUBS 0.02fF
C664 a_n919_n140# VSUBS 0.02fF
C665 a_n1097_n140# VSUBS 0.02fF
C666 a_n1275_n140# VSUBS 0.02fF
C667 a_n1453_n140# VSUBS 0.02fF
C668 a_n1631_n140# VSUBS 0.02fF
C669 a_n1809_n140# VSUBS 0.02fF
C670 a_n1987_n140# VSUBS 0.02fF
C671 a_n2165_n140# VSUBS 0.02fF
C672 a_n2343_n140# VSUBS 0.02fF
C673 a_n2521_n140# VSUBS 0.02fF
C674 a_n2699_n140# VSUBS 0.02fF
C675 a_n2877_n140# VSUBS 0.02fF
C676 a_n3055_n140# VSUBS 0.02fF
C677 a_n3233_n140# VSUBS 0.02fF
C678 a_n3411_n140# VSUBS 0.02fF
C679 a_n3589_n140# VSUBS 0.02fF
C680 a_3411_n194# VSUBS 0.29fF
C681 a_3233_n194# VSUBS 0.23fF
C682 a_3055_n194# VSUBS 0.24fF
C683 a_2877_n194# VSUBS 0.25fF
C684 a_2699_n194# VSUBS 0.26fF
C685 a_2521_n194# VSUBS 0.27fF
C686 a_2343_n194# VSUBS 0.28fF
C687 a_2165_n194# VSUBS 0.28fF
C688 a_1987_n194# VSUBS 0.29fF
C689 a_1809_n194# VSUBS 0.29fF
C690 a_1631_n194# VSUBS 0.29fF
C691 a_1453_n194# VSUBS 0.29fF
C692 a_1275_n194# VSUBS 0.29fF
C693 a_1097_n194# VSUBS 0.29fF
C694 a_919_n194# VSUBS 0.29fF
C695 a_741_n194# VSUBS 0.29fF
C696 a_563_n194# VSUBS 0.29fF
C697 a_385_n194# VSUBS 0.29fF
C698 a_207_n194# VSUBS 0.29fF
C699 a_29_n194# VSUBS 0.29fF
C700 a_n149_n194# VSUBS 0.29fF
C701 a_n327_n194# VSUBS 0.29fF
C702 a_n505_n194# VSUBS 0.29fF
C703 a_n683_n194# VSUBS 0.29fF
C704 a_n861_n194# VSUBS 0.29fF
C705 a_n1039_n194# VSUBS 0.29fF
C706 a_n1217_n194# VSUBS 0.29fF
C707 a_n1395_n194# VSUBS 0.29fF
C708 a_n1573_n194# VSUBS 0.29fF
C709 a_n1751_n194# VSUBS 0.29fF
C710 a_n1929_n194# VSUBS 0.29fF
C711 a_n2107_n194# VSUBS 0.29fF
C712 a_n2285_n194# VSUBS 0.29fF
C713 a_n2463_n194# VSUBS 0.29fF
C714 a_n2641_n194# VSUBS 0.29fF
C715 a_n2819_n194# VSUBS 0.29fF
C716 a_n2997_n194# VSUBS 0.29fF
C717 a_n3175_n194# VSUBS 0.29fF
C718 a_n3353_n194# VSUBS 0.29fF
C719 a_n3531_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_7P4E2J a_n149_n194# a_n207_n140# a_207_n194# a_n1217_n194#
+ a_327_n140# a_n1275_n140# a_n861_n194# a_n29_n140# a_n1039_n194# a_149_n140# a_n1097_n140#
+ a_1275_n194# a_29_n194# a_n683_n194# a_1395_n140# a_n741_n140# a_741_n194# a_861_n140#
+ a_1097_n194# a_n505_n194# a_n563_n140# a_563_n194# a_1217_n140# a_683_n140# a_n919_n140#
+ a_919_n194# a_n327_n194# a_1039_n140# a_n385_n140# a_385_n194# a_n1395_n194# a_505_n140#
+ a_n1453_n140# VSUBS
X0 a_n29_n140# a_n149_n194# a_n207_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n563_n140# a_n683_n194# a_n741_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n919_n140# a_n1039_n194# a_n1097_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_505_n140# a_385_n194# a_327_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n385_n140# a_n505_n194# a_n563_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X5 a_1395_n140# a_1275_n194# a_1217_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_327_n140# a_207_n194# a_149_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_149_n140# a_29_n194# a_n29_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_861_n140# a_741_n194# a_683_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n207_n140# a_n327_n194# a_n385_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X10 a_1217_n140# a_1097_n194# a_1039_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n1275_n140# a_n1395_n194# a_n1453_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X12 a_n741_n140# a_n861_n194# a_n919_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n1097_n140# a_n1217_n194# a_n1275_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_683_n140# a_563_n194# a_505_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_1039_n140# a_919_n194# a_861_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n505_n194# a_n1039_n194# 0.02fF
C1 a_n1097_n140# a_505_n140# 0.01fF
C2 a_861_n140# a_1039_n140# 0.13fF
C3 a_563_n194# a_n1039_n194# 0.01fF
C4 a_n741_n140# a_n29_n140# 0.03fF
C5 a_n741_n140# a_n1453_n140# 0.03fF
C6 a_385_n194# a_n327_n194# 0.01fF
C7 a_n683_n194# a_n1395_n194# 0.01fF
C8 a_1275_n194# a_207_n194# 0.01fF
C9 a_n741_n140# a_n563_n140# 0.13fF
C10 a_207_n194# a_741_n194# 0.02fF
C11 a_505_n140# a_327_n140# 0.13fF
C12 a_683_n140# a_n919_n140# 0.01fF
C13 a_149_n140# a_n1275_n140# 0.01fF
C14 a_683_n140# a_1217_n140# 0.04fF
C15 a_n861_n194# a_n1395_n194# 0.02fF
C16 a_29_n194# a_n1217_n194# 0.01fF
C17 a_n505_n194# a_741_n194# 0.01fF
C18 a_n207_n140# a_n1275_n140# 0.02fF
C19 a_1275_n194# a_563_n194# 0.01fF
C20 a_563_n194# a_741_n194# 0.10fF
C21 a_n683_n194# a_919_n194# 0.01fF
C22 a_683_n140# a_1395_n140# 0.03fF
C23 a_29_n194# a_n1039_n194# 0.01fF
C24 a_207_n194# a_n149_n194# 0.03fF
C25 a_n29_n140# a_1039_n140# 0.02fF
C26 a_n1217_n194# a_385_n194# 0.01fF
C27 a_n919_n140# a_149_n140# 0.02fF
C28 a_1217_n140# a_149_n140# 0.02fF
C29 a_n563_n140# a_1039_n140# 0.01fF
C30 a_n385_n140# a_n1275_n140# 0.02fF
C31 a_n505_n194# a_n149_n194# 0.03fF
C32 a_n1217_n194# a_n327_n194# 0.01fF
C33 a_385_n194# a_n1039_n194# 0.01fF
C34 a_n919_n140# a_n207_n140# 0.03fF
C35 a_1217_n140# a_n207_n140# 0.01fF
C36 a_861_n140# a_327_n140# 0.04fF
C37 a_563_n194# a_n149_n194# 0.01fF
C38 a_1395_n140# a_149_n140# 0.02fF
C39 a_29_n194# a_1275_n194# 0.01fF
C40 a_n1039_n194# a_n327_n194# 0.01fF
C41 a_29_n194# a_741_n194# 0.01fF
C42 a_n385_n140# a_n919_n140# 0.04fF
C43 a_1395_n140# a_n207_n140# 0.01fF
C44 a_n385_n140# a_1217_n140# 0.01fF
C45 a_n1097_n140# a_n29_n140# 0.02fF
C46 a_1275_n194# a_385_n194# 0.01fF
C47 a_n1097_n140# a_n1453_n140# 0.06fF
C48 a_741_n194# a_385_n194# 0.03fF
C49 a_n1097_n140# a_n563_n140# 0.04fF
C50 a_29_n194# a_n149_n194# 0.10fF
C51 a_1275_n194# a_n327_n194# 0.01fF
C52 a_n29_n140# a_327_n140# 0.06fF
C53 a_741_n194# a_n327_n194# 0.01fF
C54 a_n1217_n194# a_n1039_n194# 0.10fF
C55 a_683_n140# a_149_n140# 0.04fF
C56 a_n563_n140# a_327_n140# 0.02fF
C57 a_n683_n194# a_207_n194# 0.01fF
C58 a_385_n194# a_n149_n194# 0.02fF
C59 a_683_n140# a_n207_n140# 0.02fF
C60 a_n683_n194# a_n505_n194# 0.10fF
C61 a_n861_n194# a_207_n194# 0.01fF
C62 a_n327_n194# a_n149_n194# 0.10fF
C63 a_505_n140# a_n919_n140# 0.01fF
C64 a_n683_n194# a_563_n194# 0.01fF
C65 a_505_n140# a_1217_n140# 0.03fF
C66 a_n861_n194# a_n505_n194# 0.03fF
C67 a_683_n140# a_n385_n140# 0.02fF
C68 a_149_n140# a_n207_n140# 0.06fF
C69 a_n861_n194# a_563_n194# 0.01fF
C70 a_505_n140# a_1395_n140# 0.02fF
C71 a_n1217_n194# a_n149_n194# 0.01fF
C72 a_n385_n140# a_149_n140# 0.04fF
C73 a_29_n194# a_n683_n194# 0.01fF
C74 a_n741_n140# a_n1097_n140# 0.06fF
C75 a_n385_n140# a_n207_n140# 0.13fF
C76 a_n1039_n194# a_n149_n194# 0.01fF
C77 a_861_n140# a_1217_n140# 0.06fF
C78 a_1275_n194# a_741_n194# 0.02fF
C79 a_n861_n194# a_29_n194# 0.01fF
C80 a_n683_n194# a_385_n194# 0.01fF
C81 a_n741_n140# a_327_n140# 0.02fF
C82 a_683_n140# a_505_n140# 0.13fF
C83 a_n29_n140# a_n1275_n140# 0.02fF
C84 a_n1453_n140# a_n1275_n140# 0.13fF
C85 a_n683_n194# a_n327_n194# 0.03fF
C86 a_1395_n140# a_861_n140# 0.04fF
C87 a_n861_n194# a_385_n194# 0.01fF
C88 a_n563_n140# a_n1275_n140# 0.03fF
C89 a_1275_n194# a_n149_n194# 0.01fF
C90 a_741_n194# a_n149_n194# 0.01fF
C91 a_n861_n194# a_n327_n194# 0.02fF
C92 a_505_n140# a_149_n140# 0.06fF
C93 a_n919_n140# a_n29_n140# 0.02fF
C94 a_1217_n140# a_n29_n140# 0.02fF
C95 a_n919_n140# a_n1453_n140# 0.04fF
C96 a_327_n140# a_1039_n140# 0.03fF
C97 a_n919_n140# a_n563_n140# 0.06fF
C98 a_505_n140# a_n207_n140# 0.03fF
C99 a_n683_n194# a_n1217_n194# 0.02fF
C100 a_683_n140# a_861_n140# 0.13fF
C101 a_1395_n140# a_n29_n140# 0.01fF
C102 a_n861_n194# a_n1217_n194# 0.03fF
C103 a_n683_n194# a_n1039_n194# 0.03fF
C104 a_n385_n140# a_505_n140# 0.02fF
C105 a_n861_n194# a_n1039_n194# 0.10fF
C106 a_861_n140# a_149_n140# 0.03fF
C107 a_n1097_n140# a_327_n140# 0.01fF
C108 a_861_n140# a_n207_n140# 0.02fF
C109 a_n741_n140# a_n1275_n140# 0.04fF
C110 a_683_n140# a_n29_n140# 0.03fF
C111 a_1097_n194# a_919_n194# 0.10fF
C112 a_n683_n194# a_741_n194# 0.01fF
C113 a_683_n140# a_n563_n140# 0.02fF
C114 a_n861_n194# a_741_n194# 0.01fF
C115 a_n385_n140# a_861_n140# 0.02fF
C116 a_n741_n140# a_n919_n140# 0.13fF
C117 a_n683_n194# a_n149_n194# 0.02fF
C118 a_n1395_n194# a_207_n194# 0.01fF
C119 a_149_n140# a_n29_n140# 0.13fF
C120 a_149_n140# a_n1453_n140# 0.01fF
C121 a_n563_n140# a_149_n140# 0.03fF
C122 a_n861_n194# a_n149_n194# 0.01fF
C123 a_n505_n194# a_n1395_n194# 0.01fF
C124 a_n29_n140# a_n207_n140# 0.13fF
C125 a_n207_n140# a_n1453_n140# 0.02fF
C126 a_n563_n140# a_n207_n140# 0.06fF
C127 a_207_n194# a_919_n194# 0.01fF
C128 a_n385_n140# a_n29_n140# 0.06fF
C129 a_n385_n140# a_n1453_n140# 0.02fF
C130 a_1217_n140# a_1039_n140# 0.13fF
C131 a_n385_n140# a_n563_n140# 0.13fF
C132 a_n505_n194# a_919_n194# 0.01fF
C133 a_1097_n194# a_207_n194# 0.01fF
C134 a_505_n140# a_861_n140# 0.06fF
C135 a_563_n194# a_919_n194# 0.03fF
C136 a_n1097_n140# a_n1275_n140# 0.13fF
C137 a_1395_n140# a_1039_n140# 0.06fF
C138 a_29_n194# a_n1395_n194# 0.01fF
C139 a_1097_n194# a_n505_n194# 0.01fF
C140 a_n741_n140# a_683_n140# 0.01fF
C141 a_1097_n194# a_563_n194# 0.02fF
C142 a_327_n140# a_n1275_n140# 0.01fF
C143 a_n1097_n140# a_n919_n140# 0.13fF
C144 a_n861_n194# a_n683_n194# 0.10fF
C145 a_n741_n140# a_149_n140# 0.02fF
C146 a_29_n194# a_919_n194# 0.01fF
C147 a_505_n140# a_n29_n140# 0.04fF
C148 a_n1395_n194# a_n327_n194# 0.01fF
C149 a_505_n140# a_n563_n140# 0.02fF
C150 a_683_n140# a_1039_n140# 0.06fF
C151 a_n919_n140# a_327_n140# 0.02fF
C152 a_n741_n140# a_n207_n140# 0.04fF
C153 a_1217_n140# a_327_n140# 0.02fF
C154 a_1097_n194# a_29_n194# 0.01fF
C155 a_385_n194# a_919_n194# 0.02fF
C156 a_n505_n194# a_207_n194# 0.01fF
C157 a_919_n194# a_n327_n194# 0.01fF
C158 a_n741_n140# a_n385_n140# 0.06fF
C159 a_1395_n140# a_327_n140# 0.02fF
C160 a_1097_n194# a_385_n194# 0.01fF
C161 a_149_n140# a_1039_n140# 0.02fF
C162 a_n1395_n194# a_n1217_n194# 0.10fF
C163 a_207_n194# a_563_n194# 0.03fF
C164 a_861_n140# a_n29_n140# 0.02fF
C165 a_1097_n194# a_n327_n194# 0.01fF
C166 a_n207_n140# a_1039_n140# 0.02fF
C167 a_n505_n194# a_563_n194# 0.01fF
C168 a_n1395_n194# a_n1039_n194# 0.03fF
C169 a_861_n140# a_n563_n140# 0.01fF
C170 a_n385_n140# a_1039_n140# 0.01fF
C171 a_29_n194# a_207_n194# 0.10fF
C172 a_683_n140# a_327_n140# 0.06fF
C173 a_n1097_n140# a_149_n140# 0.02fF
C174 a_29_n194# a_n505_n194# 0.02fF
C175 a_n741_n140# a_505_n140# 0.02fF
C176 a_207_n194# a_385_n194# 0.10fF
C177 a_n29_n140# a_n1453_n140# 0.01fF
C178 a_n1097_n140# a_n207_n140# 0.02fF
C179 a_29_n194# a_563_n194# 0.02fF
C180 a_n563_n140# a_n29_n140# 0.04fF
C181 a_n563_n140# a_n1453_n140# 0.02fF
C182 a_149_n140# a_327_n140# 0.13fF
C183 a_n919_n140# a_n1275_n140# 0.06fF
C184 a_n505_n194# a_385_n194# 0.01fF
C185 a_207_n194# a_n327_n194# 0.02fF
C186 a_n1395_n194# a_n149_n194# 0.01fF
C187 a_1275_n194# a_919_n194# 0.03fF
C188 a_n207_n140# a_327_n140# 0.04fF
C189 a_563_n194# a_385_n194# 0.10fF
C190 a_n1097_n140# a_n385_n140# 0.03fF
C191 a_741_n194# a_919_n194# 0.10fF
C192 a_n505_n194# a_n327_n194# 0.10fF
C193 a_505_n140# a_1039_n140# 0.04fF
C194 a_1097_n194# a_1275_n194# 0.10fF
C195 a_563_n194# a_n327_n194# 0.01fF
C196 a_1097_n194# a_741_n194# 0.03fF
C197 a_n385_n140# a_327_n140# 0.03fF
C198 a_n741_n140# a_861_n140# 0.01fF
C199 a_919_n194# a_n149_n194# 0.01fF
C200 a_207_n194# a_n1217_n194# 0.01fF
C201 a_29_n194# a_385_n194# 0.03fF
C202 a_1395_n140# a_1217_n140# 0.13fF
C203 a_n505_n194# a_n1217_n194# 0.01fF
C204 a_207_n194# a_n1039_n194# 0.01fF
C205 a_1097_n194# a_n149_n194# 0.01fF
C206 a_29_n194# a_n327_n194# 0.03fF
C207 a_1395_n140# VSUBS 0.02fF
C208 a_1217_n140# VSUBS 0.02fF
C209 a_1039_n140# VSUBS 0.02fF
C210 a_861_n140# VSUBS 0.02fF
C211 a_683_n140# VSUBS 0.02fF
C212 a_505_n140# VSUBS 0.02fF
C213 a_327_n140# VSUBS 0.02fF
C214 a_149_n140# VSUBS 0.02fF
C215 a_n29_n140# VSUBS 0.02fF
C216 a_n207_n140# VSUBS 0.02fF
C217 a_n385_n140# VSUBS 0.02fF
C218 a_n563_n140# VSUBS 0.02fF
C219 a_n741_n140# VSUBS 0.02fF
C220 a_n919_n140# VSUBS 0.02fF
C221 a_n1097_n140# VSUBS 0.02fF
C222 a_n1275_n140# VSUBS 0.02fF
C223 a_n1453_n140# VSUBS 0.02fF
C224 a_1275_n194# VSUBS 0.29fF
C225 a_1097_n194# VSUBS 0.23fF
C226 a_919_n194# VSUBS 0.24fF
C227 a_741_n194# VSUBS 0.25fF
C228 a_563_n194# VSUBS 0.26fF
C229 a_385_n194# VSUBS 0.27fF
C230 a_207_n194# VSUBS 0.28fF
C231 a_29_n194# VSUBS 0.28fF
C232 a_n149_n194# VSUBS 0.29fF
C233 a_n327_n194# VSUBS 0.29fF
C234 a_n505_n194# VSUBS 0.29fF
C235 a_n683_n194# VSUBS 0.29fF
C236 a_n861_n194# VSUBS 0.29fF
C237 a_n1039_n194# VSUBS 0.29fF
C238 a_n1217_n194# VSUBS 0.29fF
C239 a_n1395_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_KEEN2X a_n1008_n140# a_2374_n140# a_1306_n140# a_n652_n140#
+ a_652_n194# a_n1662_n194# a_772_n140# a_n2730_n194# a_n1720_n140# a_n60_n194# a_2076_n194#
+ a_1008_n194# a_2196_n140# a_n474_n140# a_n416_n194# a_1128_n140# a_474_n194# a_n1484_n194#
+ a_n2552_n194# a_594_n140# a_n1542_n140# a_n2610_n140# a_1720_n194# a_1840_n140#
+ a_n238_n194# a_n2908_n194# a_3086_n140# a_n296_n140# a_n1898_n140# a_n2966_n140#
+ a_296_n194# a_2018_n140# a_60_n140# a_n1306_n194# a_n2374_n194# a_n1364_n140# a_1542_n194#
+ a_416_n140# a_n2432_n140# a_2610_n194# a_n950_n194# a_1662_n140# a_2730_n140# a_2966_n194#
+ a_1898_n194# a_n2788_n140# a_n118_n140# a_118_n194# a_n2196_n194# a_n1128_n194#
+ a_238_n140# a_n1186_n140# a_n2254_n140# a_2432_n194# a_1364_n194# a_n772_n194# a_2552_n140#
+ a_1484_n140# a_n830_n140# a_2788_n194# a_830_n194# a_n1840_n194# a_950_n140# a_n3086_n194#
+ a_2908_n140# a_1186_n194# a_n2018_n194# a_n2076_n140# a_n3144_n140# a_2254_n194#
+ a_n594_n194# VSUBS
X0 a_2374_n140# a_2254_n194# a_2196_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n2788_n140# a_n2908_n194# a_n2966_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n2432_n140# a_n2552_n194# a_n2610_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1128_n140# a_1008_n194# a_950_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1186_n140# a_n1306_n194# a_n1364_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_772_n140# a_652_n194# a_594_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_1662_n140# a_1542_n194# a_1484_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n2966_n140# a_n3086_n194# a_n3144_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_2730_n140# a_2610_n194# a_2552_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n118_n140# a_n238_n194# a_n296_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_2196_n140# a_2076_n194# a_2018_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X11 a_n2610_n140# a_n2730_n194# a_n2788_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_n2254_n140# a_n2374_n194# a_n2432_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_n652_n140# a_n772_n194# a_n830_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_2018_n140# a_1898_n194# a_1840_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n1008_n140# a_n1128_n194# a_n1186_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_594_n140# a_474_n194# a_416_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X17 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X18 a_3086_n140# a_2966_n194# a_2908_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X19 a_1484_n140# a_1364_n194# a_1306_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X20 a_n1542_n140# a_n1662_n194# a_n1720_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X21 a_2552_n140# a_2432_n194# a_2374_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_950_n140# a_830_n194# a_772_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X23 a_n2076_n140# a_n2196_n194# a_n2254_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X24 a_n830_n140# a_n950_n194# a_n1008_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X25 a_n474_n140# a_n594_n194# a_n652_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X26 a_1840_n140# a_1720_n194# a_1662_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X27 a_416_n140# a_296_n194# a_238_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X28 a_2908_n140# a_2788_n194# a_2730_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X29 a_n1898_n140# a_n2018_n194# a_n2076_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X30 a_n296_n140# a_n416_n194# a_n474_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X31 a_1306_n140# a_1186_n194# a_1128_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X32 a_n1720_n140# a_n1840_n194# a_n1898_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X33 a_n1364_n140# a_n1484_n194# a_n1542_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X34 a_238_n140# a_118_n194# a_60_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_n1542_n140# a_n1008_n140# 0.04fF
C1 a_n772_n194# a_n594_n194# 0.10fF
C2 a_2374_n140# a_772_n140# 0.01fF
C3 a_n1720_n140# a_n3144_n140# 0.01fF
C4 a_2432_n194# a_1364_n194# 0.01fF
C5 a_n1720_n140# a_n652_n140# 0.02fF
C6 a_1008_n194# a_n594_n194# 0.01fF
C7 a_1364_n194# a_652_n194# 0.01fF
C8 a_n2788_n140# a_n2610_n140# 0.13fF
C9 a_830_n194# a_474_n194# 0.03fF
C10 a_1008_n194# a_2254_n194# 0.01fF
C11 a_2432_n194# a_1898_n194# 0.02fF
C12 a_118_n194# a_n416_n194# 0.02fF
C13 a_1128_n140# a_238_n140# 0.02fF
C14 a_1898_n194# a_652_n194# 0.01fF
C15 a_1186_n194# a_n416_n194# 0.01fF
C16 a_1662_n140# a_950_n140# 0.03fF
C17 a_n1186_n140# a_238_n140# 0.01fF
C18 a_n2254_n140# a_n1898_n140# 0.06fF
C19 a_n2552_n194# a_n1840_n194# 0.01fF
C20 a_n1364_n140# a_n1898_n140# 0.04fF
C21 a_n652_n140# a_n1186_n140# 0.04fF
C22 a_n1898_n140# a_n830_n140# 0.02fF
C23 a_1542_n194# a_2254_n194# 0.01fF
C24 a_n2196_n194# a_n1306_n194# 0.01fF
C25 a_n2432_n140# a_n2254_n140# 0.13fF
C26 a_n60_n194# a_652_n194# 0.01fF
C27 a_n1364_n140# a_n296_n140# 0.02fF
C28 a_n296_n140# a_n830_n140# 0.04fF
C29 a_n2432_n140# a_n1364_n140# 0.02fF
C30 a_n474_n140# a_n1008_n140# 0.04fF
C31 a_950_n140# a_60_n140# 0.02fF
C32 a_n2432_n140# a_n830_n140# 0.01fF
C33 a_296_n194# a_n772_n194# 0.01fF
C34 a_n772_n194# a_n950_n194# 0.10fF
C35 a_1364_n194# a_1898_n194# 0.02fF
C36 a_1008_n194# a_296_n194# 0.01fF
C37 a_2552_n140# a_1662_n140# 0.02fF
C38 a_n2610_n140# a_n1008_n140# 0.01fF
C39 a_n2374_n194# a_n2730_n194# 0.03fF
C40 a_1484_n140# a_n118_n140# 0.01fF
C41 a_594_n140# a_416_n140# 0.13fF
C42 a_n2018_n194# a_n1840_n194# 0.10fF
C43 a_474_n194# a_n416_n194# 0.01fF
C44 a_n416_n194# a_n1662_n194# 0.01fF
C45 a_n652_n140# a_238_n140# 0.02fF
C46 a_594_n140# a_1840_n140# 0.02fF
C47 a_2552_n140# a_3086_n140# 0.04fF
C48 a_1364_n194# a_n60_n194# 0.01fF
C49 a_n238_n194# a_652_n194# 0.01fF
C50 a_2374_n140# a_950_n140# 0.01fF
C51 a_n2374_n194# a_n772_n194# 0.01fF
C52 a_n2788_n140# a_n2254_n140# 0.04fF
C53 a_n2788_n140# a_n1364_n140# 0.01fF
C54 a_2196_n140# a_594_n140# 0.01fF
C55 a_1542_n194# a_296_n194# 0.01fF
C56 a_n2966_n140# a_n2076_n140# 0.02fF
C57 a_1364_n194# a_n238_n194# 0.01fF
C58 a_2552_n140# a_2374_n140# 0.13fF
C59 a_n3086_n194# a_n2196_n194# 0.01fF
C60 a_2730_n140# a_1840_n140# 0.02fF
C61 a_2076_n194# a_1720_n194# 0.03fF
C62 a_n296_n140# a_60_n140# 0.06fF
C63 a_2908_n140# a_2552_n140# 0.06fF
C64 a_n60_n194# a_n1484_n194# 0.01fF
C65 a_n2196_n194# a_n1662_n194# 0.02fF
C66 a_2730_n140# a_2196_n140# 0.04fF
C67 a_n2196_n194# a_n2908_n194# 0.01fF
C68 a_2432_n194# a_2610_n194# 0.10fF
C69 a_n2254_n140# a_n1008_n140# 0.02fF
C70 a_1128_n140# a_594_n140# 0.04fF
C71 a_n1364_n140# a_n1008_n140# 0.06fF
C72 a_n1008_n140# a_n830_n140# 0.13fF
C73 a_n238_n194# a_n60_n194# 0.10fF
C74 a_772_n140# a_416_n140# 0.06fF
C75 a_n2552_n194# a_n1128_n194# 0.01fF
C76 a_2788_n194# a_1542_n194# 0.01fF
C77 a_n238_n194# a_n1484_n194# 0.01fF
C78 a_772_n140# a_1840_n140# 0.02fF
C79 a_2432_n194# a_1186_n194# 0.01fF
C80 a_2196_n140# a_772_n140# 0.01fF
C81 a_1364_n194# a_2610_n194# 0.01fF
C82 a_830_n194# a_2076_n194# 0.01fF
C83 a_652_n194# a_118_n194# 0.02fF
C84 a_n2018_n194# a_n1128_n194# 0.01fF
C85 a_2076_n194# a_2966_n194# 0.01fF
C86 a_594_n140# a_238_n140# 0.06fF
C87 a_n2966_n140# a_n1720_n140# 0.02fF
C88 a_2730_n140# a_1128_n140# 0.01fF
C89 a_1186_n194# a_652_n194# 0.02fF
C90 a_594_n140# a_n652_n140# 0.02fF
C91 a_n2018_n194# a_n594_n194# 0.01fF
C92 a_1898_n194# a_2610_n194# 0.01fF
C93 a_n1542_n140# a_n118_n140# 0.01fF
C94 a_n60_n194# a_n1306_n194# 0.01fF
C95 a_1364_n194# a_118_n194# 0.01fF
C96 a_n1840_n194# a_n416_n194# 0.01fF
C97 a_1186_n194# a_1364_n194# 0.10fF
C98 a_n1484_n194# a_n1306_n194# 0.10fF
C99 a_474_n194# a_652_n194# 0.10fF
C100 a_60_n140# a_n1008_n140# 0.02fF
C101 a_1128_n140# a_772_n140# 0.06fF
C102 a_n2552_n194# a_n950_n194# 0.01fF
C103 a_n238_n194# a_n1306_n194# 0.01fF
C104 a_950_n140# a_416_n140# 0.04fF
C105 a_1186_n194# a_1898_n194# 0.01fF
C106 a_2254_n194# a_1720_n194# 0.02fF
C107 a_2018_n140# a_1662_n140# 0.06fF
C108 a_950_n140# a_1840_n140# 0.02fF
C109 a_n60_n194# a_118_n194# 0.10fF
C110 a_1364_n194# a_474_n194# 0.01fF
C111 a_1186_n194# a_n60_n194# 0.01fF
C112 a_n2966_n140# a_n3144_n140# 0.13fF
C113 a_2018_n140# a_3086_n140# 0.02fF
C114 a_n2018_n194# a_n950_n194# 0.01fF
C115 a_2196_n140# a_950_n140# 0.02fF
C116 a_118_n194# a_n1484_n194# 0.01fF
C117 a_n2374_n194# a_n2552_n194# 0.10fF
C118 a_772_n140# a_238_n140# 0.04fF
C119 a_n474_n140# a_n118_n140# 0.06fF
C120 a_n1898_n140# a_n2076_n140# 0.13fF
C121 a_772_n140# a_n652_n140# 0.01fF
C122 a_1898_n194# a_474_n194# 0.01fF
C123 a_n2196_n194# a_n1840_n194# 0.03fF
C124 a_n2432_n140# a_n2076_n140# 0.06fF
C125 a_2552_n140# a_1840_n140# 0.03fF
C126 a_1306_n140# a_1662_n140# 0.06fF
C127 a_n238_n194# a_118_n194# 0.03fF
C128 a_830_n194# a_n594_n194# 0.01fF
C129 a_1186_n194# a_n238_n194# 0.01fF
C130 a_n3086_n194# a_n1484_n194# 0.01fF
C131 a_n2374_n194# a_n2018_n194# 0.03fF
C132 a_296_n194# a_1720_n194# 0.01fF
C133 a_n60_n194# a_474_n194# 0.02fF
C134 a_n60_n194# a_n1662_n194# 0.01fF
C135 a_2018_n140# a_2374_n140# 0.06fF
C136 a_2196_n140# a_2552_n140# 0.06fF
C137 a_1306_n140# a_60_n140# 0.02fF
C138 a_2254_n194# a_830_n194# 0.01fF
C139 a_2254_n194# a_2966_n194# 0.01fF
C140 a_n1662_n194# a_n1484_n194# 0.10fF
C141 a_n1484_n194# a_n2908_n194# 0.01fF
C142 a_2908_n140# a_2018_n140# 0.02fF
C143 a_n296_n140# a_416_n140# 0.03fF
C144 a_n2788_n140# a_n2076_n140# 0.03fF
C145 a_1128_n140# a_950_n140# 0.13fF
C146 a_1306_n140# a_2374_n140# 0.02fF
C147 a_n238_n194# a_474_n194# 0.01fF
C148 a_n238_n194# a_n1662_n194# 0.01fF
C149 a_n416_n194# a_n1128_n194# 0.01fF
C150 a_118_n194# a_n1306_n194# 0.01fF
C151 a_2908_n140# a_1306_n140# 0.01fF
C152 a_n416_n194# a_n594_n194# 0.10fF
C153 a_1008_n194# a_1542_n194# 0.02fF
C154 a_2552_n140# a_1128_n140# 0.01fF
C155 a_830_n194# a_296_n194# 0.02fF
C156 a_n1720_n140# a_n1898_n140# 0.13fF
C157 a_950_n140# a_238_n140# 0.03fF
C158 a_n1720_n140# a_n296_n140# 0.01fF
C159 a_n2432_n140# a_n1720_n140# 0.03fF
C160 a_1186_n194# a_2610_n194# 0.01fF
C161 a_2788_n194# a_1720_n194# 0.01fF
C162 a_950_n140# a_n652_n140# 0.01fF
C163 a_n1364_n140# a_n118_n140# 0.02fF
C164 a_n118_n140# a_n830_n140# 0.03fF
C165 a_n1008_n140# a_n2076_n140# 0.02fF
C166 a_2432_n194# a_2076_n194# 0.03fF
C167 a_n1662_n194# a_n1306_n194# 0.03fF
C168 a_772_n140# a_594_n140# 0.13fF
C169 a_n1542_n140# a_n474_n140# 0.02fF
C170 a_n1306_n194# a_n2908_n194# 0.01fF
C171 a_1128_n140# a_n296_n140# 0.01fF
C172 a_652_n194# a_2076_n194# 0.01fF
C173 a_1186_n194# a_118_n194# 0.01fF
C174 a_n2196_n194# a_n1128_n194# 0.01fF
C175 a_n1720_n140# a_n2788_n140# 0.02fF
C176 a_n1186_n140# a_n1898_n140# 0.03fF
C177 a_n2610_n140# a_n1542_n140# 0.02fF
C178 a_n1186_n140# a_n296_n140# 0.02fF
C179 a_1484_n140# a_1662_n140# 0.13fF
C180 a_296_n194# a_n416_n194# 0.01fF
C181 a_n2432_n140# a_n1186_n140# 0.02fF
C182 a_n2196_n194# a_n594_n194# 0.01fF
C183 a_n416_n194# a_n950_n194# 0.02fF
C184 a_1484_n140# a_3086_n140# 0.01fF
C185 a_n1008_n140# a_416_n140# 0.01fF
C186 a_1484_n140# a_60_n140# 0.01fF
C187 a_1364_n194# a_2076_n194# 0.01fF
C188 a_2788_n194# a_2966_n194# 0.10fF
C189 a_474_n194# a_118_n194# 0.03fF
C190 a_n3144_n140# a_n1898_n140# 0.02fF
C191 a_n296_n140# a_238_n140# 0.04fF
C192 a_n652_n140# a_n1898_n140# 0.02fF
C193 a_1186_n194# a_474_n194# 0.01fF
C194 a_n2432_n140# a_n3144_n140# 0.03fF
C195 a_n652_n140# a_n296_n140# 0.06fF
C196 a_1898_n194# a_2076_n194# 0.10fF
C197 a_n2788_n140# a_n1186_n140# 0.01fF
C198 a_n118_n140# a_60_n140# 0.13fF
C199 a_1484_n140# a_2374_n140# 0.02fF
C200 a_n1840_n194# a_n1484_n194# 0.03fF
C201 a_n3086_n194# a_n1662_n194# 0.01fF
C202 a_2018_n140# a_416_n140# 0.01fF
C203 a_n1720_n140# a_n1008_n140# 0.03fF
C204 a_n3086_n194# a_n2908_n194# 0.10fF
C205 a_n2552_n194# a_n2730_n194# 0.10fF
C206 a_2908_n140# a_1484_n140# 0.01fF
C207 a_2018_n140# a_1840_n140# 0.13fF
C208 a_n238_n194# a_n1840_n194# 0.01fF
C209 a_950_n140# a_594_n140# 0.06fF
C210 a_n1662_n194# a_n2908_n194# 0.01fF
C211 a_n2196_n194# a_n950_n194# 0.01fF
C212 a_n2788_n140# a_n3144_n140# 0.06fF
C213 a_n1542_n140# a_n2254_n140# 0.03fF
C214 a_2018_n140# a_2196_n140# 0.13fF
C215 a_n1542_n140# a_n1364_n140# 0.13fF
C216 a_1306_n140# a_416_n140# 0.02fF
C217 a_n1542_n140# a_n830_n140# 0.03fF
C218 a_n2018_n194# a_n2730_n194# 0.01fF
C219 a_1306_n140# a_1840_n140# 0.04fF
C220 a_652_n194# a_n594_n194# 0.01fF
C221 a_n1186_n140# a_n1008_n140# 0.13fF
C222 a_n2374_n194# a_n2196_n194# 0.10fF
C223 a_2432_n194# a_2254_n194# 0.10fF
C224 a_n2018_n194# a_n772_n194# 0.01fF
C225 a_1306_n140# a_2196_n140# 0.02fF
C226 a_2254_n194# a_652_n194# 0.01fF
C227 a_n1008_n140# a_238_n140# 0.02fF
C228 a_n1840_n194# a_n1306_n194# 0.02fF
C229 a_2018_n140# a_1128_n140# 0.02fF
C230 a_n652_n140# a_n1008_n140# 0.06fF
C231 a_2730_n140# a_2552_n140# 0.13fF
C232 a_n1364_n140# a_n474_n140# 0.02fF
C233 a_1364_n194# a_2254_n194# 0.01fF
C234 a_n474_n140# a_n830_n140# 0.06fF
C235 a_594_n140# a_n296_n140# 0.02fF
C236 a_1008_n194# a_1720_n194# 0.01fF
C237 a_n60_n194# a_n1128_n194# 0.01fF
C238 a_n2610_n140# a_n2254_n140# 0.06fF
C239 a_n2610_n140# a_n1364_n140# 0.02fF
C240 a_n1542_n140# a_60_n140# 0.01fF
C241 a_652_n194# a_296_n194# 0.03fF
C242 a_950_n140# a_772_n140# 0.13fF
C243 a_1306_n140# a_1128_n140# 0.13fF
C244 a_2076_n194# a_2610_n194# 0.02fF
C245 a_652_n194# a_n950_n194# 0.01fF
C246 a_2254_n194# a_1898_n194# 0.03fF
C247 a_n1484_n194# a_n1128_n194# 0.03fF
C248 a_n60_n194# a_n594_n194# 0.02fF
C249 a_1542_n194# a_1720_n194# 0.10fF
C250 a_n594_n194# a_n1484_n194# 0.01fF
C251 a_n238_n194# a_n1128_n194# 0.01fF
C252 a_1364_n194# a_296_n194# 0.01fF
C253 a_830_n194# a_n772_n194# 0.01fF
C254 a_n3086_n194# a_n1840_n194# 0.01fF
C255 a_1306_n140# a_238_n140# 0.02fF
C256 a_n238_n194# a_n594_n194# 0.03fF
C257 a_1008_n194# a_830_n194# 0.10fF
C258 a_1186_n194# a_2076_n194# 0.01fF
C259 a_1484_n140# a_416_n140# 0.02fF
C260 a_1898_n194# a_296_n194# 0.01fF
C261 a_1484_n140# a_1840_n140# 0.06fF
C262 a_n1840_n194# a_n1662_n194# 0.10fF
C263 a_n1840_n194# a_n2908_n194# 0.01fF
C264 a_2432_n194# a_2788_n194# 0.03fF
C265 a_n2966_n140# a_n1898_n140# 0.02fF
C266 a_n474_n140# a_60_n140# 0.04fF
C267 a_n2432_n140# a_n2966_n140# 0.04fF
C268 a_n60_n194# a_296_n194# 0.03fF
C269 a_1484_n140# a_2196_n140# 0.03fF
C270 a_1542_n194# a_830_n194# 0.01fF
C271 a_n118_n140# a_416_n140# 0.04fF
C272 a_772_n140# a_n296_n140# 0.02fF
C273 a_n60_n194# a_n950_n194# 0.01fF
C274 a_1542_n194# a_2966_n194# 0.01fF
C275 a_n2254_n140# a_n830_n140# 0.01fF
C276 a_n2254_n140# a_n1364_n140# 0.02fF
C277 a_474_n194# a_2076_n194# 0.01fF
C278 a_n1364_n140# a_n830_n140# 0.04fF
C279 a_n1306_n194# a_n1128_n194# 0.10fF
C280 a_594_n140# a_n1008_n140# 0.01fF
C281 a_n1484_n194# a_n950_n194# 0.02fF
C282 a_n772_n194# a_n416_n194# 0.03fF
C283 a_2788_n194# a_1364_n194# 0.01fF
C284 a_n594_n194# a_n1306_n194# 0.01fF
C285 a_1008_n194# a_n416_n194# 0.01fF
C286 a_n238_n194# a_296_n194# 0.02fF
C287 a_n2966_n140# a_n2788_n140# 0.13fF
C288 a_n238_n194# a_n950_n194# 0.01fF
C289 a_n1720_n140# a_n118_n140# 0.01fF
C290 a_2552_n140# a_950_n140# 0.01fF
C291 a_n2374_n194# a_n1484_n194# 0.01fF
C292 a_2788_n194# a_1898_n194# 0.01fF
C293 a_n2552_n194# a_n2018_n194# 0.02fF
C294 a_1484_n140# a_1128_n140# 0.06fF
C295 a_2254_n194# a_2610_n194# 0.03fF
C296 a_2018_n140# a_594_n140# 0.01fF
C297 a_118_n194# a_n1128_n194# 0.01fF
C298 a_n2196_n194# a_n2730_n194# 0.02fF
C299 a_118_n194# a_n594_n194# 0.01fF
C300 a_n1542_n140# a_n2076_n140# 0.04fF
C301 a_1128_n140# a_n118_n140# 0.02fF
C302 a_n2196_n194# a_n772_n194# 0.01fF
C303 a_1306_n140# a_594_n140# 0.03fF
C304 a_n1364_n140# a_60_n140# 0.01fF
C305 a_60_n140# a_n830_n140# 0.02fF
C306 a_950_n140# a_n296_n140# 0.02fF
C307 a_n1186_n140# a_n118_n140# 0.02fF
C308 a_1484_n140# a_238_n140# 0.02fF
C309 a_296_n194# a_n1306_n194# 0.01fF
C310 a_1186_n194# a_2254_n194# 0.01fF
C311 a_n1306_n194# a_n950_n194# 0.03fF
C312 a_2730_n140# a_2018_n140# 0.03fF
C313 a_474_n194# a_n1128_n194# 0.01fF
C314 a_n1662_n194# a_n1128_n194# 0.02fF
C315 a_474_n194# a_n594_n194# 0.01fF
C316 a_n594_n194# a_n1662_n194# 0.01fF
C317 a_n118_n140# a_238_n140# 0.06fF
C318 a_n652_n140# a_n118_n140# 0.04fF
C319 a_n2374_n194# a_n1306_n194# 0.01fF
C320 a_2730_n140# a_1306_n140# 0.01fF
C321 a_296_n194# a_118_n194# 0.10fF
C322 a_118_n194# a_n950_n194# 0.01fF
C323 a_1186_n194# a_296_n194# 0.01fF
C324 a_n474_n140# a_n2076_n140# 0.01fF
C325 a_1662_n140# a_3086_n140# 0.01fF
C326 a_2018_n140# a_772_n140# 0.02fF
C327 a_1662_n140# a_60_n140# 0.01fF
C328 a_n2610_n140# a_n2076_n140# 0.04fF
C329 a_n1898_n140# a_n296_n140# 0.01fF
C330 a_n1720_n140# a_n1542_n140# 0.13fF
C331 a_n2432_n140# a_n1898_n140# 0.04fF
C332 a_2788_n194# a_2610_n194# 0.10fF
C333 a_1008_n194# a_2432_n194# 0.01fF
C334 a_1306_n140# a_772_n140# 0.04fF
C335 a_652_n194# a_n772_n194# 0.01fF
C336 a_474_n194# a_296_n194# 0.10fF
C337 a_2374_n140# a_1662_n140# 0.03fF
C338 a_n474_n140# a_416_n140# 0.02fF
C339 a_474_n194# a_n950_n194# 0.01fF
C340 a_n1662_n194# a_n950_n194# 0.01fF
C341 a_1008_n194# a_652_n194# 0.03fF
C342 a_2374_n140# a_3086_n140# 0.03fF
C343 a_n2374_n194# a_n3086_n194# 0.01fF
C344 a_2908_n140# a_1662_n140# 0.02fF
C345 a_n2788_n140# a_n1898_n140# 0.02fF
C346 a_830_n194# a_1720_n194# 0.01fF
C347 a_2432_n194# a_1542_n194# 0.01fF
C348 a_n1542_n140# a_n1186_n140# 0.06fF
C349 a_2908_n140# a_3086_n140# 0.13fF
C350 a_1484_n140# a_594_n140# 0.02fF
C351 a_n2432_n140# a_n2788_n140# 0.06fF
C352 a_1720_n194# a_2966_n194# 0.01fF
C353 a_1186_n194# a_2788_n194# 0.01fF
C354 a_n2374_n194# a_n1662_n194# 0.01fF
C355 a_n2374_n194# a_n2908_n194# 0.02fF
C356 a_1008_n194# a_1364_n194# 0.03fF
C357 a_1542_n194# a_652_n194# 0.01fF
C358 a_n1720_n140# a_n474_n140# 0.02fF
C359 a_n2018_n194# a_n416_n194# 0.01fF
C360 a_2018_n140# a_950_n140# 0.02fF
C361 a_n1542_n140# a_n3144_n140# 0.01fF
C362 a_n2254_n140# a_n2076_n140# 0.13fF
C363 a_594_n140# a_n118_n140# 0.03fF
C364 a_1008_n194# a_1898_n194# 0.01fF
C365 a_n1720_n140# a_n2610_n140# 0.02fF
C366 a_n1364_n140# a_n2076_n140# 0.03fF
C367 a_n830_n140# a_n2076_n140# 0.02fF
C368 a_n1542_n140# a_n652_n140# 0.02fF
C369 a_n1484_n194# a_n2730_n194# 0.01fF
C370 a_2908_n140# a_2374_n140# 0.04fF
C371 a_n1840_n194# a_n1128_n194# 0.01fF
C372 a_n60_n194# a_n772_n194# 0.01fF
C373 a_1542_n194# a_1364_n194# 0.10fF
C374 a_2730_n140# a_1484_n140# 0.02fF
C375 a_1008_n194# a_n60_n194# 0.01fF
C376 a_1128_n140# a_n474_n140# 0.01fF
C377 a_n1898_n140# a_n1008_n140# 0.02fF
C378 a_1306_n140# a_950_n140# 0.06fF
C379 a_n772_n194# a_n1484_n194# 0.01fF
C380 a_2018_n140# a_2552_n140# 0.04fF
C381 a_n1840_n194# a_n594_n194# 0.01fF
C382 a_n296_n140# a_n1008_n140# 0.03fF
C383 a_n2552_n194# a_n2196_n194# 0.03fF
C384 a_n2432_n140# a_n1008_n140# 0.01fF
C385 a_1542_n194# a_1898_n194# 0.03fF
C386 a_n1186_n140# a_n474_n140# 0.03fF
C387 a_n238_n194# a_n772_n194# 0.02fF
C388 a_n830_n140# a_416_n140# 0.02fF
C389 a_n2610_n140# a_n1186_n140# 0.01fF
C390 a_1542_n194# a_n60_n194# 0.01fF
C391 a_1008_n194# a_n238_n194# 0.01fF
C392 a_1306_n140# a_2552_n140# 0.02fF
C393 a_n2018_n194# a_n2196_n194# 0.10fF
C394 a_1484_n140# a_772_n140# 0.03fF
C395 a_n474_n140# a_238_n140# 0.03fF
C396 a_2254_n194# a_2076_n194# 0.10fF
C397 a_n652_n140# a_n474_n140# 0.13fF
C398 a_n2610_n140# a_n3144_n140# 0.04fF
C399 a_n1720_n140# a_n2254_n140# 0.04fF
C400 a_830_n194# a_n416_n194# 0.01fF
C401 a_n1720_n140# a_n1364_n140# 0.06fF
C402 a_n1306_n194# a_n2730_n194# 0.01fF
C403 a_n1720_n140# a_n830_n140# 0.02fF
C404 a_772_n140# a_n118_n140# 0.02fF
C405 a_n1840_n194# a_n950_n194# 0.01fF
C406 a_1306_n140# a_n296_n140# 0.01fF
C407 a_n772_n194# a_n1306_n194# 0.02fF
C408 a_1662_n140# a_416_n140# 0.02fF
C409 a_1662_n140# a_1840_n140# 0.13fF
C410 a_60_n140# a_416_n140# 0.06fF
C411 a_n2374_n194# a_n1840_n194# 0.02fF
C412 a_3086_n140# a_1840_n140# 0.02fF
C413 a_1008_n194# a_2610_n194# 0.01fF
C414 a_2196_n140# a_1662_n140# 0.04fF
C415 a_n2254_n140# a_n1186_n140# 0.02fF
C416 a_n1364_n140# a_n1186_n140# 0.13fF
C417 a_n1186_n140# a_n830_n140# 0.06fF
C418 a_2196_n140# a_3086_n140# 0.02fF
C419 a_n594_n194# a_n1128_n194# 0.02fF
C420 a_118_n194# a_n772_n194# 0.01fF
C421 a_1484_n140# a_950_n140# 0.04fF
C422 a_n3086_n194# a_n2730_n194# 0.03fF
C423 a_1542_n194# a_2610_n194# 0.01fF
C424 a_1008_n194# a_118_n194# 0.01fF
C425 a_n2254_n140# a_n3144_n140# 0.02fF
C426 a_n1364_n140# a_238_n140# 0.01fF
C427 a_2374_n140# a_1840_n140# 0.04fF
C428 a_n830_n140# a_238_n140# 0.02fF
C429 a_n2254_n140# a_n652_n140# 0.01fF
C430 a_1008_n194# a_1186_n194# 0.10fF
C431 a_n1364_n140# a_n652_n140# 0.03fF
C432 a_n652_n140# a_n830_n140# 0.13fF
C433 a_n1662_n194# a_n2730_n194# 0.01fF
C434 a_2432_n194# a_1720_n194# 0.01fF
C435 a_n2908_n194# a_n2730_n194# 0.10fF
C436 a_2196_n140# a_2374_n140# 0.13fF
C437 a_950_n140# a_n118_n140# 0.02fF
C438 a_2908_n140# a_1840_n140# 0.02fF
C439 a_1484_n140# a_2552_n140# 0.02fF
C440 a_594_n140# a_n474_n140# 0.02fF
C441 a_2788_n194# a_2076_n194# 0.01fF
C442 a_1662_n140# a_1128_n140# 0.04fF
C443 a_652_n194# a_1720_n194# 0.01fF
C444 a_1542_n194# a_118_n194# 0.01fF
C445 a_474_n194# a_n772_n194# 0.01fF
C446 a_n772_n194# a_n1662_n194# 0.01fF
C447 a_2908_n140# a_2196_n140# 0.03fF
C448 a_n2966_n140# a_n1542_n140# 0.01fF
C449 a_1186_n194# a_1542_n194# 0.03fF
C450 a_1128_n140# a_60_n140# 0.02fF
C451 a_1008_n194# a_474_n194# 0.02fF
C452 a_296_n194# a_n1128_n194# 0.01fF
C453 a_n2552_n194# a_n1484_n194# 0.01fF
C454 a_n1128_n194# a_n950_n194# 0.10fF
C455 a_n1186_n140# a_60_n140# 0.02fF
C456 a_1364_n194# a_1720_n194# 0.03fF
C457 a_1662_n140# a_238_n140# 0.01fF
C458 a_296_n194# a_n594_n194# 0.01fF
C459 a_n594_n194# a_n950_n194# 0.03fF
C460 a_2432_n194# a_830_n194# 0.01fF
C461 a_2374_n140# a_1128_n140# 0.02fF
C462 a_1542_n194# a_474_n194# 0.01fF
C463 a_2432_n194# a_2966_n194# 0.02fF
C464 a_n2018_n194# a_n1484_n194# 0.02fF
C465 a_1898_n194# a_1720_n194# 0.10fF
C466 a_60_n140# a_238_n140# 0.13fF
C467 a_n2374_n194# a_n1128_n194# 0.01fF
C468 a_830_n194# a_652_n194# 0.10fF
C469 a_1306_n140# a_2018_n140# 0.03fF
C470 a_n652_n140# a_60_n140# 0.03fF
C471 a_n296_n140# a_n118_n140# 0.13fF
C472 a_772_n140# a_n474_n140# 0.02fF
C473 a_1364_n194# a_830_n194# 0.02fF
C474 a_n2966_n140# a_n2610_n140# 0.06fF
C475 a_1364_n194# a_2966_n194# 0.01fF
C476 a_594_n140# a_n830_n140# 0.01fF
C477 a_n2552_n194# a_n1306_n194# 0.01fF
C478 a_296_n194# a_n950_n194# 0.01fF
C479 a_1898_n194# a_830_n194# 0.01fF
C480 a_1898_n194# a_2966_n194# 0.01fF
C481 a_652_n194# a_n416_n194# 0.01fF
C482 a_2788_n194# a_2254_n194# 0.02fF
C483 a_n60_n194# a_830_n194# 0.01fF
C484 a_n2018_n194# a_n1306_n194# 0.01fF
C485 a_n1720_n140# a_n2076_n140# 0.06fF
C486 a_n1840_n194# a_n2730_n194# 0.01fF
C487 a_416_n140# a_1840_n140# 0.01fF
C488 a_n2374_n194# a_n950_n194# 0.01fF
C489 a_n1840_n194# a_n772_n194# 0.01fF
C490 a_1662_n140# a_594_n140# 0.02fF
C491 a_n238_n194# a_830_n194# 0.01fF
C492 a_2196_n140# a_1840_n140# 0.06fF
C493 a_n2966_n140# a_n2254_n140# 0.03fF
C494 a_n118_n140# a_n1008_n140# 0.02fF
C495 a_n2966_n140# a_n1364_n140# 0.01fF
C496 a_n3086_n194# a_n2552_n194# 0.02fF
C497 a_594_n140# a_60_n140# 0.04fF
C498 a_950_n140# a_n474_n140# 0.01fF
C499 a_1720_n194# a_2610_n194# 0.01fF
C500 a_n1186_n140# a_n2076_n140# 0.02fF
C501 a_n1542_n140# a_n1898_n140# 0.06fF
C502 a_772_n140# a_n830_n140# 0.01fF
C503 a_1484_n140# a_2018_n140# 0.04fF
C504 a_n1542_n140# a_n296_n140# 0.02fF
C505 a_1008_n194# a_2076_n194# 0.01fF
C506 a_n60_n194# a_n416_n194# 0.03fF
C507 a_n2432_n140# a_n1542_n140# 0.02fF
C508 a_n2552_n194# a_n1662_n194# 0.01fF
C509 a_n2552_n194# a_n2908_n194# 0.03fF
C510 a_2730_n140# a_1662_n140# 0.02fF
C511 a_n3086_n194# a_n2018_n194# 0.01fF
C512 a_n416_n194# a_n1484_n194# 0.01fF
C513 a_1128_n140# a_416_n140# 0.03fF
C514 a_118_n194# a_1720_n194# 0.01fF
C515 a_n3144_n140# a_n2076_n140# 0.02fF
C516 a_2730_n140# a_3086_n140# 0.06fF
C517 a_n652_n140# a_n2076_n140# 0.01fF
C518 a_1306_n140# a_1484_n140# 0.13fF
C519 a_1186_n194# a_1720_n194# 0.02fF
C520 a_1128_n140# a_1840_n140# 0.03fF
C521 a_n2018_n194# a_n1662_n194# 0.03fF
C522 a_1542_n194# a_2076_n194# 0.02fF
C523 a_n1186_n140# a_416_n140# 0.01fF
C524 a_n238_n194# a_n416_n194# 0.10fF
C525 a_n2018_n194# a_n2908_n194# 0.01fF
C526 a_n2788_n140# a_n1542_n140# 0.02fF
C527 a_2196_n140# a_1128_n140# 0.02fF
C528 a_2610_n194# a_2966_n194# 0.03fF
C529 a_1306_n140# a_n118_n140# 0.01fF
C530 a_2730_n140# a_2374_n140# 0.06fF
C531 a_n1898_n140# a_n474_n140# 0.01fF
C532 a_1662_n140# a_772_n140# 0.02fF
C533 a_238_n140# a_416_n140# 0.13fF
C534 a_n296_n140# a_n474_n140# 0.13fF
C535 a_n652_n140# a_416_n140# 0.02fF
C536 a_474_n194# a_1720_n194# 0.01fF
C537 a_n1128_n194# a_n2730_n194# 0.01fF
C538 a_238_n140# a_1840_n140# 0.01fF
C539 a_n2610_n140# a_n1898_n140# 0.03fF
C540 a_2730_n140# a_2908_n140# 0.13fF
C541 a_772_n140# a_60_n140# 0.03fF
C542 a_n1720_n140# a_n1186_n140# 0.04fF
C543 a_830_n194# a_118_n194# 0.01fF
C544 a_n2196_n194# a_n1484_n194# 0.01fF
C545 a_n2432_n140# a_n2610_n140# 0.13fF
C546 a_1186_n194# a_830_n194# 0.03fF
C547 a_n772_n194# a_n1128_n194# 0.03fF
C548 a_n416_n194# a_n1306_n194# 0.01fF
C549 a_3086_n140# VSUBS 0.02fF
C550 a_2908_n140# VSUBS 0.02fF
C551 a_2730_n140# VSUBS 0.02fF
C552 a_2552_n140# VSUBS 0.02fF
C553 a_2374_n140# VSUBS 0.02fF
C554 a_2196_n140# VSUBS 0.02fF
C555 a_2018_n140# VSUBS 0.02fF
C556 a_1840_n140# VSUBS 0.02fF
C557 a_1662_n140# VSUBS 0.02fF
C558 a_1484_n140# VSUBS 0.02fF
C559 a_1306_n140# VSUBS 0.02fF
C560 a_1128_n140# VSUBS 0.02fF
C561 a_950_n140# VSUBS 0.02fF
C562 a_772_n140# VSUBS 0.02fF
C563 a_594_n140# VSUBS 0.02fF
C564 a_416_n140# VSUBS 0.02fF
C565 a_238_n140# VSUBS 0.02fF
C566 a_60_n140# VSUBS 0.02fF
C567 a_n118_n140# VSUBS 0.02fF
C568 a_n296_n140# VSUBS 0.02fF
C569 a_n474_n140# VSUBS 0.02fF
C570 a_n652_n140# VSUBS 0.02fF
C571 a_n830_n140# VSUBS 0.02fF
C572 a_n1008_n140# VSUBS 0.02fF
C573 a_n1186_n140# VSUBS 0.02fF
C574 a_n1364_n140# VSUBS 0.02fF
C575 a_n1542_n140# VSUBS 0.02fF
C576 a_n1720_n140# VSUBS 0.02fF
C577 a_n1898_n140# VSUBS 0.02fF
C578 a_n2076_n140# VSUBS 0.02fF
C579 a_n2254_n140# VSUBS 0.02fF
C580 a_n2432_n140# VSUBS 0.02fF
C581 a_n2610_n140# VSUBS 0.02fF
C582 a_n2788_n140# VSUBS 0.02fF
C583 a_n2966_n140# VSUBS 0.02fF
C584 a_n3144_n140# VSUBS 0.02fF
C585 a_2966_n194# VSUBS 0.29fF
C586 a_2788_n194# VSUBS 0.23fF
C587 a_2610_n194# VSUBS 0.24fF
C588 a_2432_n194# VSUBS 0.25fF
C589 a_2254_n194# VSUBS 0.26fF
C590 a_2076_n194# VSUBS 0.27fF
C591 a_1898_n194# VSUBS 0.28fF
C592 a_1720_n194# VSUBS 0.28fF
C593 a_1542_n194# VSUBS 0.29fF
C594 a_1364_n194# VSUBS 0.29fF
C595 a_1186_n194# VSUBS 0.29fF
C596 a_1008_n194# VSUBS 0.29fF
C597 a_830_n194# VSUBS 0.29fF
C598 a_652_n194# VSUBS 0.29fF
C599 a_474_n194# VSUBS 0.29fF
C600 a_296_n194# VSUBS 0.29fF
C601 a_118_n194# VSUBS 0.29fF
C602 a_n60_n194# VSUBS 0.29fF
C603 a_n238_n194# VSUBS 0.29fF
C604 a_n416_n194# VSUBS 0.29fF
C605 a_n594_n194# VSUBS 0.29fF
C606 a_n772_n194# VSUBS 0.29fF
C607 a_n950_n194# VSUBS 0.29fF
C608 a_n1128_n194# VSUBS 0.29fF
C609 a_n1306_n194# VSUBS 0.29fF
C610 a_n1484_n194# VSUBS 0.29fF
C611 a_n1662_n194# VSUBS 0.29fF
C612 a_n1840_n194# VSUBS 0.29fF
C613 a_n2018_n194# VSUBS 0.29fF
C614 a_n2196_n194# VSUBS 0.29fF
C615 a_n2374_n194# VSUBS 0.29fF
C616 a_n2552_n194# VSUBS 0.29fF
C617 a_n2730_n194# VSUBS 0.29fF
C618 a_n2908_n194# VSUBS 0.29fF
C619 a_n3086_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__nfet_01v8_VJ4JGY a_n352_n194# a_n60_n194# a_n644_n194# a_n936_n194#
+ a_n410_n140# a_n994_n140# a_n702_n140# a_n232_n140# a_n524_n140# a_524_n194# a_232_n194#
+ a_n816_n140# a_816_n194# a_644_n140# a_352_n140# a_936_n140# a_60_n140# a_174_n140#
+ a_466_n140# a_758_n140# a_n118_n140# VSUBS
X0 a_n232_n140# a_n352_n194# a_n410_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n524_n140# a_n644_n194# a_n702_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n816_n140# a_n936_n194# a_n994_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_60_n140# a_n60_n194# a_n118_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_352_n140# a_232_n194# a_174_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_644_n140# a_524_n194# a_466_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_936_n140# a_816_n194# a_758_n140# VSUBS sky130_fd_pr__nfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
C0 a_524_n194# a_n936_n194# 0.01fF
C1 a_816_n194# a_524_n194# 0.04fF
C2 a_174_n140# a_n994_n140# 0.02fF
C3 a_644_n140# a_936_n140# 0.07fF
C4 a_n352_n194# a_n936_n194# 0.02fF
C5 a_816_n194# a_n352_n194# 0.01fF
C6 a_60_n140# a_n118_n140# 0.13fF
C7 a_n524_n140# a_n702_n140# 0.13fF
C8 a_466_n140# a_n410_n140# 0.02fF
C9 a_n60_n194# a_n936_n194# 0.01fF
C10 a_816_n194# a_n60_n194# 0.01fF
C11 a_644_n140# a_60_n140# 0.03fF
C12 a_n994_n140# a_n524_n140# 0.04fF
C13 a_936_n140# a_n232_n140# 0.02fF
C14 a_n816_n140# a_466_n140# 0.01fF
C15 a_644_n140# a_n118_n140# 0.03fF
C16 a_524_n194# a_n644_n194# 0.01fF
C17 a_n410_n140# a_n702_n140# 0.07fF
C18 a_n352_n194# a_n644_n194# 0.04fF
C19 a_352_n140# a_466_n140# 0.25fF
C20 a_174_n140# a_936_n140# 0.03fF
C21 a_936_n140# a_758_n140# 0.13fF
C22 a_n994_n140# a_n410_n140# 0.03fF
C23 a_60_n140# a_n232_n140# 0.07fF
C24 a_n60_n194# a_n644_n194# 0.02fF
C25 a_n816_n140# a_n702_n140# 0.25fF
C26 a_n118_n140# a_n232_n140# 0.25fF
C27 a_174_n140# a_60_n140# 0.25fF
C28 a_352_n140# a_n702_n140# 0.02fF
C29 a_60_n140# a_758_n140# 0.03fF
C30 a_936_n140# a_n524_n140# 0.01fF
C31 a_n816_n140# a_n994_n140# 0.13fF
C32 a_174_n140# a_n118_n140# 0.07fF
C33 a_n118_n140# a_758_n140# 0.02fF
C34 a_352_n140# a_n994_n140# 0.01fF
C35 a_644_n140# a_n232_n140# 0.02fF
C36 a_60_n140# a_n524_n140# 0.03fF
C37 a_936_n140# a_n410_n140# 0.01fF
C38 a_644_n140# a_174_n140# 0.04fF
C39 a_644_n140# a_758_n140# 0.25fF
C40 a_n118_n140# a_n524_n140# 0.05fF
C41 a_n936_n194# a_n644_n194# 0.04fF
C42 a_816_n194# a_n644_n194# 0.01fF
C43 a_466_n140# a_n702_n140# 0.02fF
C44 a_60_n140# a_n410_n140# 0.04fF
C45 a_644_n140# a_n524_n140# 0.02fF
C46 a_232_n194# a_524_n194# 0.04fF
C47 a_936_n140# a_352_n140# 0.03fF
C48 a_232_n194# a_n352_n194# 0.02fF
C49 a_174_n140# a_n232_n140# 0.05fF
C50 a_n118_n140# a_n410_n140# 0.07fF
C51 a_n232_n140# a_758_n140# 0.02fF
C52 a_466_n140# a_n994_n140# 0.01fF
C53 a_n816_n140# a_60_n140# 0.02fF
C54 a_174_n140# a_758_n140# 0.03fF
C55 a_n60_n194# a_232_n194# 0.04fF
C56 a_n816_n140# a_n118_n140# 0.03fF
C57 a_60_n140# a_352_n140# 0.07fF
C58 a_644_n140# a_n410_n140# 0.02fF
C59 a_n232_n140# a_n524_n140# 0.07fF
C60 a_n994_n140# a_n702_n140# 0.07fF
C61 a_352_n140# a_n118_n140# 0.04fF
C62 a_174_n140# a_n524_n140# 0.03fF
C63 a_644_n140# a_n816_n140# 0.01fF
C64 a_758_n140# a_n524_n140# 0.01fF
C65 a_936_n140# a_466_n140# 0.04fF
C66 a_644_n140# a_352_n140# 0.07fF
C67 a_n232_n140# a_n410_n140# 0.13fF
C68 a_174_n140# a_n410_n140# 0.03fF
C69 a_758_n140# a_n410_n140# 0.02fF
C70 a_232_n194# a_n936_n194# 0.01fF
C71 a_816_n194# a_232_n194# 0.02fF
C72 a_n816_n140# a_n232_n140# 0.03fF
C73 a_60_n140# a_466_n140# 0.05fF
C74 a_936_n140# a_n702_n140# 0.01fF
C75 a_466_n140# a_n118_n140# 0.03fF
C76 a_352_n140# a_n232_n140# 0.03fF
C77 a_174_n140# a_n816_n140# 0.02fF
C78 a_n816_n140# a_758_n140# 0.01fF
C79 a_n410_n140# a_n524_n140# 0.25fF
C80 a_60_n140# a_n702_n140# 0.03fF
C81 a_174_n140# a_352_n140# 0.13fF
C82 a_352_n140# a_758_n140# 0.05fF
C83 a_644_n140# a_466_n140# 0.13fF
C84 a_n118_n140# a_n702_n140# 0.03fF
C85 a_232_n194# a_n644_n194# 0.01fF
C86 a_n816_n140# a_n524_n140# 0.07fF
C87 a_60_n140# a_n994_n140# 0.02fF
C88 a_n352_n194# a_524_n194# 0.01fF
C89 a_n994_n140# a_n118_n140# 0.02fF
C90 a_352_n140# a_n524_n140# 0.02fF
C91 a_644_n140# a_n702_n140# 0.01fF
C92 a_n60_n194# a_524_n194# 0.02fF
C93 a_466_n140# a_n232_n140# 0.03fF
C94 a_n60_n194# a_n352_n194# 0.04fF
C95 a_n816_n140# a_n410_n140# 0.05fF
C96 a_644_n140# a_n994_n140# 0.01fF
C97 a_174_n140# a_466_n140# 0.07fF
C98 a_466_n140# a_758_n140# 0.07fF
C99 a_352_n140# a_n410_n140# 0.03fF
C100 a_936_n140# a_60_n140# 0.02fF
C101 a_n232_n140# a_n702_n140# 0.04fF
C102 a_936_n140# a_n118_n140# 0.02fF
C103 a_n816_n140# a_352_n140# 0.02fF
C104 a_n994_n140# a_n232_n140# 0.03fF
C105 a_466_n140# a_n524_n140# 0.02fF
C106 a_174_n140# a_n702_n140# 0.02fF
C107 a_758_n140# a_n702_n140# 0.01fF
C108 a_936_n140# VSUBS 0.02fF
C109 a_758_n140# VSUBS 0.02fF
C110 a_644_n140# VSUBS 0.02fF
C111 a_466_n140# VSUBS 0.02fF
C112 a_352_n140# VSUBS 0.02fF
C113 a_174_n140# VSUBS 0.02fF
C114 a_60_n140# VSUBS 0.02fF
C115 a_n118_n140# VSUBS 0.02fF
C116 a_n232_n140# VSUBS 0.02fF
C117 a_n410_n140# VSUBS 0.02fF
C118 a_n524_n140# VSUBS 0.02fF
C119 a_n702_n140# VSUBS 0.02fF
C120 a_n816_n140# VSUBS 0.02fF
C121 a_n994_n140# VSUBS 0.02fF
C122 a_816_n194# VSUBS 0.29fF
C123 a_524_n194# VSUBS 0.24fF
C124 a_232_n194# VSUBS 0.26fF
C125 a_n60_n194# VSUBS 0.27fF
C126 a_n352_n194# VSUBS 0.29fF
C127 a_n644_n194# VSUBS 0.29fF
C128 a_n936_n194# VSUBS 0.35fF
.ends

.subckt sky130_fd_pr__pfet_01v8_E4DCBA a_n1008_n140# a_n416_n205# a_1306_n140# a_n652_n140#
+ a_474_n205# a_n1484_n205# a_772_n140# a_n1720_n140# a_1720_n205# a_n238_n205# a_n474_n140#
+ a_296_n205# a_1128_n140# a_594_n140# a_1542_n205# a_n1306_n205# w_n2112_n240# a_n1542_n140#
+ a_n950_n205# a_1840_n140# a_1898_n205# a_n296_n140# a_n1898_n140# a_2018_n140# a_60_n140#
+ a_118_n205# a_n1128_n205# a_n1364_n140# a_1364_n205# a_416_n140# a_n772_n205# a_1662_n140#
+ a_830_n205# a_n1840_n205# a_n118_n140# a_1186_n205# a_n2018_n205# a_238_n140# a_n1186_n140#
+ a_n594_n205# a_1484_n140# a_n830_n140# a_652_n205# a_n1662_n205# a_950_n140# a_n60_n205#
+ a_n2076_n140# a_1008_n205# VSUBS
X0 a_1662_n140# a_1542_n205# a_1484_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_n118_n140# a_n238_n205# a_n296_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n652_n140# a_n772_n205# a_n830_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_2018_n140# a_1898_n205# a_1840_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_n1008_n140# a_n1128_n205# a_n1186_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_594_n140# a_474_n205# a_416_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_60_n140# a_n60_n205# a_n118_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X7 a_1484_n140# a_1364_n205# a_1306_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X8 a_n1542_n140# a_n1662_n205# a_n1720_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_950_n140# a_830_n205# a_772_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n830_n140# a_n950_n205# a_n1008_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n474_n140# a_n594_n205# a_n652_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_1840_n140# a_1720_n205# a_1662_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_416_n140# a_296_n205# a_238_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X14 a_n1898_n140# a_n2018_n205# a_n2076_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X15 a_n296_n140# a_n416_n205# a_n474_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X16 a_n1720_n140# a_n1840_n205# a_n1898_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X17 a_1306_n140# a_1186_n205# a_1128_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X18 a_n1364_n140# a_n1484_n205# a_n1542_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X19 a_238_n140# a_118_n205# a_60_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X20 a_1128_n140# a_1008_n205# a_950_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X21 a_n1186_n140# a_n1306_n205# a_n1364_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X22 a_772_n140# a_652_n205# a_594_n140# w_n2112_n240# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_830_n205# a_1542_n205# 0.01fF
C1 w_n2112_n240# a_1840_n140# 0.02fF
C2 a_n1008_n140# a_n474_n140# 0.04fF
C3 w_n2112_n240# a_416_n140# 0.02fF
C4 a_830_n205# a_n772_n205# 0.01fF
C5 a_n652_n140# a_238_n140# 0.02fF
C6 a_n1128_n205# a_n1306_n205# 0.11fF
C7 a_60_n140# a_238_n140# 0.13fF
C8 a_n2076_n140# a_n474_n140# 0.01fF
C9 a_474_n205# a_n238_n205# 0.01fF
C10 a_474_n205# a_1186_n205# 0.01fF
C11 a_n1898_n140# a_n1186_n140# 0.03fF
C12 a_n830_n140# a_n118_n140# 0.03fF
C13 a_474_n205# a_296_n205# 0.11fF
C14 a_1128_n140# w_n2112_n240# 0.02fF
C15 a_n772_n205# a_n594_n205# 0.11fF
C16 a_n950_n205# a_652_n205# 0.01fF
C17 a_1306_n140# a_n296_n140# 0.01fF
C18 a_n416_n205# a_1008_n205# 0.01fF
C19 a_n950_n205# a_n1484_n205# 0.02fF
C20 a_594_n140# w_n2112_n240# 0.02fF
C21 a_n772_n205# a_n1840_n205# 0.01fF
C22 a_1484_n140# a_238_n140# 0.02fF
C23 a_n652_n140# a_n118_n140# 0.04fF
C24 a_950_n140# a_1840_n140# 0.02fF
C25 a_n1542_n140# a_n296_n140# 0.02fF
C26 a_n118_n140# a_60_n140# 0.13fF
C27 a_950_n140# a_416_n140# 0.04fF
C28 a_n60_n205# a_1008_n205# 0.01fF
C29 a_n1128_n205# w_n2112_n240# 0.24fF
C30 a_n950_n205# a_n1662_n205# 0.01fF
C31 a_n1542_n140# a_n474_n140# 0.02fF
C32 w_n2112_n240# a_n1720_n140# 0.02fF
C33 a_n1720_n140# a_n1364_n140# 0.06fF
C34 a_n2018_n205# a_n1306_n205# 0.01fF
C35 a_n238_n205# a_n1306_n205# 0.01fF
C36 a_950_n140# a_1128_n140# 0.13fF
C37 a_n296_n140# a_n1898_n140# 0.01fF
C38 a_652_n205# a_n416_n205# 0.01fF
C39 a_1484_n140# a_n118_n140# 0.01fF
C40 a_772_n140# a_1662_n140# 0.02fF
C41 a_n1484_n205# a_n416_n205# 0.01fF
C42 a_1364_n205# a_n238_n205# 0.01fF
C43 a_296_n205# a_n1306_n205# 0.01fF
C44 a_594_n140# a_950_n140# 0.06fF
C45 a_1364_n205# a_1186_n205# 0.11fF
C46 a_n1008_n140# w_n2112_n240# 0.02fF
C47 a_118_n205# a_1008_n205# 0.01fF
C48 a_772_n140# a_1306_n140# 0.04fF
C49 a_n1008_n140# a_n1364_n140# 0.06fF
C50 a_1898_n205# a_1186_n205# 0.01fF
C51 a_296_n205# a_1364_n205# 0.01fF
C52 a_n296_n140# a_n1186_n140# 0.02fF
C53 a_n1898_n140# a_n474_n140# 0.01fF
C54 a_652_n205# a_n60_n205# 0.01fF
C55 a_n1484_n205# a_n60_n205# 0.01fF
C56 a_296_n205# a_1898_n205# 0.01fF
C57 w_n2112_n240# a_n2076_n140# 0.02fF
C58 a_n1128_n205# a_n594_n205# 0.02fF
C59 a_n2076_n140# a_n1364_n140# 0.03fF
C60 a_n1662_n205# a_n416_n205# 0.01fF
C61 a_n1840_n205# a_n1128_n205# 0.01fF
C62 a_n830_n140# a_416_n140# 0.02fF
C63 a_n474_n140# a_n1186_n140# 0.03fF
C64 w_n2112_n240# a_n238_n205# 0.24fF
C65 a_n2018_n205# w_n2112_n240# 0.31fF
C66 a_118_n205# a_652_n205# 0.02fF
C67 a_n1662_n205# a_n60_n205# 0.01fF
C68 a_118_n205# a_n1484_n205# 0.01fF
C69 w_n2112_n240# a_1186_n205# 0.21fF
C70 a_296_n205# w_n2112_n240# 0.24fF
C71 a_n652_n140# a_416_n140# 0.02fF
C72 w_n2112_n240# a_1662_n140# 0.02fF
C73 a_1720_n205# a_1008_n205# 0.01fF
C74 a_830_n205# a_n238_n205# 0.01fF
C75 a_60_n140# a_416_n140# 0.06fF
C76 a_830_n205# a_1186_n205# 0.03fF
C77 a_1306_n140# w_n2112_n240# 0.02fF
C78 a_594_n140# a_n830_n140# 0.01fF
C79 a_830_n205# a_296_n205# 0.02fF
C80 a_n1542_n140# w_n2112_n240# 0.02fF
C81 a_n1542_n140# a_n1364_n140# 0.13fF
C82 a_1484_n140# a_1840_n140# 0.06fF
C83 a_1542_n205# a_1008_n205# 0.02fF
C84 a_1128_n140# a_60_n140# 0.02fF
C85 a_n238_n205# a_n594_n205# 0.03fF
C86 a_n2018_n205# a_n594_n205# 0.01fF
C87 a_n950_n205# a_n416_n205# 0.02fF
C88 a_n296_n140# a_n474_n140# 0.13fF
C89 a_1484_n140# a_416_n140# 0.02fF
C90 a_594_n140# a_n652_n140# 0.02fF
C91 a_n1840_n205# a_n238_n205# 0.01fF
C92 a_n1840_n205# a_n2018_n205# 0.11fF
C93 a_594_n140# a_60_n140# 0.04fF
C94 a_n830_n140# a_n1720_n140# 0.02fF
C95 a_652_n205# a_1720_n205# 0.01fF
C96 a_296_n205# a_n594_n205# 0.01fF
C97 a_950_n140# a_1662_n140# 0.03fF
C98 w_n2112_n240# a_n1898_n140# 0.02fF
C99 a_n1898_n140# a_n1364_n140# 0.04fF
C100 a_n950_n205# a_n60_n205# 0.01fF
C101 a_1306_n140# a_950_n140# 0.06fF
C102 a_1484_n140# a_1128_n140# 0.06fF
C103 a_772_n140# a_n296_n140# 0.02fF
C104 a_n830_n140# a_n1008_n140# 0.13fF
C105 a_n652_n140# a_n1720_n140# 0.02fF
C106 a_594_n140# a_1484_n140# 0.02fF
C107 a_1542_n205# a_652_n205# 0.01fF
C108 w_n2112_n240# a_n1186_n140# 0.02fF
C109 a_n1186_n140# a_n1364_n140# 0.13fF
C110 a_n772_n205# a_652_n205# 0.01fF
C111 a_n830_n140# a_n2076_n140# 0.02fF
C112 a_474_n205# a_1364_n205# 0.01fF
C113 a_n772_n205# a_n1484_n205# 0.01fF
C114 a_n652_n140# a_n1008_n140# 0.06fF
C115 a_n950_n205# a_118_n205# 0.01fF
C116 a_772_n140# a_n474_n140# 0.02fF
C117 a_474_n205# a_1898_n205# 0.01fF
C118 a_n1008_n140# a_60_n140# 0.02fF
C119 a_n416_n205# a_n60_n205# 0.03fF
C120 a_n652_n140# a_n2076_n140# 0.01fF
C121 a_n772_n205# a_n1662_n205# 0.01fF
C122 w_n2112_n240# a_n296_n140# 0.02fF
C123 a_474_n205# w_n2112_n240# 0.24fF
C124 a_n296_n140# a_n1364_n140# 0.02fF
C125 a_118_n205# a_n416_n205# 0.02fF
C126 a_2018_n140# a_1840_n140# 0.13fF
C127 a_n1542_n140# a_n830_n140# 0.03fF
C128 a_2018_n140# a_416_n140# 0.01fF
C129 a_474_n205# a_830_n205# 0.03fF
C130 a_60_n140# a_1662_n140# 0.01fF
C131 w_n2112_n240# a_n474_n140# 0.02fF
C132 a_n474_n140# a_n1364_n140# 0.02fF
C133 a_118_n205# a_n60_n205# 0.11fF
C134 a_1306_n140# a_60_n140# 0.02fF
C135 a_n1128_n205# a_n1484_n205# 0.03fF
C136 a_1364_n205# a_1898_n205# 0.02fF
C137 a_n652_n140# a_n1542_n140# 0.02fF
C138 a_n118_n140# a_238_n140# 0.06fF
C139 a_2018_n140# a_1128_n140# 0.02fF
C140 a_n1542_n140# a_60_n140# 0.01fF
C141 a_n830_n140# a_n1898_n140# 0.02fF
C142 a_474_n205# a_n594_n205# 0.01fF
C143 a_594_n140# a_2018_n140# 0.01fF
C144 a_1484_n140# a_1662_n140# 0.13fF
C145 a_950_n140# a_n296_n140# 0.02fF
C146 a_n950_n205# a_n772_n205# 0.11fF
C147 a_n238_n205# a_1008_n205# 0.01fF
C148 a_772_n140# w_n2112_n240# 0.02fF
C149 a_1186_n205# a_1008_n205# 0.11fF
C150 a_1484_n140# a_1306_n140# 0.13fF
C151 w_n2112_n240# a_n1306_n205# 0.24fF
C152 a_n1662_n205# a_n1128_n205# 0.02fF
C153 a_n830_n140# a_n1186_n140# 0.06fF
C154 a_n652_n140# a_n1898_n140# 0.02fF
C155 a_296_n205# a_1008_n205# 0.01fF
C156 w_n2112_n240# a_1364_n205# 0.20fF
C157 a_950_n140# a_n474_n140# 0.01fF
C158 w_n2112_n240# a_1898_n205# 0.24fF
C159 a_n652_n140# a_n1186_n140# 0.04fF
C160 a_830_n205# a_1364_n205# 0.02fF
C161 a_60_n140# a_n1186_n140# 0.02fF
C162 a_652_n205# a_n238_n205# 0.01fF
C163 a_n772_n205# a_n416_n205# 0.03fF
C164 a_830_n205# a_1898_n205# 0.01fF
C165 a_n1484_n205# a_n238_n205# 0.01fF
C166 a_n2018_n205# a_n1484_n205# 0.02fF
C167 a_652_n205# a_1186_n205# 0.02fF
C168 a_772_n140# a_950_n140# 0.13fF
C169 a_652_n205# a_296_n205# 0.03fF
C170 a_n594_n205# a_n1306_n205# 0.01fF
C171 a_1542_n205# a_n60_n205# 0.01fF
C172 a_118_n205# a_1720_n205# 0.01fF
C173 a_n1840_n205# a_n1306_n205# 0.02fF
C174 a_n772_n205# a_n60_n205# 0.01fF
C175 a_n830_n140# a_n296_n140# 0.04fF
C176 w_n2112_n240# a_n1364_n140# 0.02fF
C177 a_1840_n140# a_238_n140# 0.01fF
C178 a_n950_n205# a_n1128_n205# 0.11fF
C179 a_n1662_n205# a_n238_n205# 0.01fF
C180 a_n1662_n205# a_n2018_n205# 0.03fF
C181 a_416_n140# a_238_n140# 0.13fF
C182 a_830_n205# w_n2112_n240# 0.23fF
C183 a_118_n205# a_1542_n205# 0.01fF
C184 a_n652_n140# a_n296_n140# 0.06fF
C185 a_n830_n140# a_n474_n140# 0.06fF
C186 a_n296_n140# a_60_n140# 0.06fF
C187 a_118_n205# a_n772_n205# 0.01fF
C188 a_2018_n140# a_1662_n140# 0.06fF
C189 a_1128_n140# a_238_n140# 0.02fF
C190 w_n2112_n240# a_n594_n205# 0.24fF
C191 a_2018_n140# a_1306_n140# 0.03fF
C192 a_n652_n140# a_n474_n140# 0.13fF
C193 a_950_n140# w_n2112_n240# 0.02fF
C194 a_n1128_n205# a_n416_n205# 0.01fF
C195 a_594_n140# a_238_n140# 0.06fF
C196 a_n118_n140# a_416_n140# 0.04fF
C197 a_60_n140# a_n474_n140# 0.04fF
C198 a_n1840_n205# w_n2112_n240# 0.24fF
C199 a_772_n140# a_n830_n140# 0.01fF
C200 a_830_n205# a_n594_n205# 0.01fF
C201 a_n1128_n205# a_n60_n205# 0.01fF
C202 a_474_n205# a_1008_n205# 0.02fF
C203 a_1128_n140# a_n118_n140# 0.02fF
C204 a_n950_n205# a_n238_n205# 0.01fF
C205 a_n950_n205# a_n2018_n205# 0.01fF
C206 a_772_n140# a_n652_n140# 0.01fF
C207 a_1542_n205# a_1720_n205# 0.11fF
C208 a_772_n140# a_60_n140# 0.03fF
C209 a_n950_n205# a_296_n205# 0.01fF
C210 a_594_n140# a_n118_n140# 0.03fF
C211 a_n1840_n205# a_n594_n205# 0.01fF
C212 a_n1008_n140# a_238_n140# 0.02fF
C213 a_118_n205# a_n1128_n205# 0.01fF
C214 a_772_n140# a_1484_n140# 0.03fF
C215 a_n830_n140# w_n2112_n240# 0.02fF
C216 a_474_n205# a_652_n205# 0.11fF
C217 a_n830_n140# a_n1364_n140# 0.04fF
C218 a_n416_n205# a_n238_n205# 0.11fF
C219 a_n2018_n205# a_n416_n205# 0.01fF
C220 a_n118_n140# a_n1720_n140# 0.01fF
C221 a_n416_n205# a_1186_n205# 0.01fF
C222 a_296_n205# a_n416_n205# 0.01fF
C223 a_n652_n140# w_n2112_n240# 0.02fF
C224 a_n1008_n140# a_n118_n140# 0.02fF
C225 a_n652_n140# a_n1364_n140# 0.03fF
C226 a_n238_n205# a_n60_n205# 0.11fF
C227 a_1840_n140# a_416_n140# 0.01fF
C228 w_n2112_n240# a_60_n140# 0.02fF
C229 a_n60_n205# a_1186_n205# 0.01fF
C230 a_1364_n205# a_1008_n205# 0.03fF
C231 a_60_n140# a_n1364_n140# 0.01fF
C232 a_296_n205# a_n60_n205# 0.03fF
C233 a_1898_n205# a_1008_n205# 0.01fF
C234 a_1662_n140# a_238_n140# 0.01fF
C235 a_1306_n140# a_238_n140# 0.02fF
C236 a_1128_n140# a_1840_n140# 0.03fF
C237 a_118_n205# a_n238_n205# 0.03fF
C238 a_1128_n140# a_416_n140# 0.03fF
C239 a_1484_n140# w_n2112_n240# 0.02fF
C240 a_118_n205# a_1186_n205# 0.01fF
C241 a_594_n140# a_1840_n140# 0.02fF
C242 a_n1484_n205# a_n1306_n205# 0.11fF
C243 a_118_n205# a_296_n205# 0.11fF
C244 a_594_n140# a_416_n140# 0.13fF
C245 a_n652_n140# a_950_n140# 0.01fF
C246 a_652_n205# a_1364_n205# 0.01fF
C247 w_n2112_n240# a_1008_n205# 0.22fF
C248 a_950_n140# a_60_n140# 0.02fF
C249 a_n772_n205# a_n1128_n205# 0.03fF
C250 a_652_n205# a_1898_n205# 0.01fF
C251 a_1306_n140# a_n118_n140# 0.01fF
C252 a_830_n205# a_1008_n205# 0.11fF
C253 a_594_n140# a_1128_n140# 0.04fF
C254 a_n1662_n205# a_n1306_n205# 0.03fF
C255 a_n1542_n140# a_n118_n140# 0.01fF
C256 a_474_n205# a_n950_n205# 0.01fF
C257 a_772_n140# a_2018_n140# 0.02fF
C258 a_1484_n140# a_950_n140# 0.04fF
C259 a_n1186_n140# a_238_n140# 0.01fF
C260 a_1720_n205# a_1186_n205# 0.02fF
C261 a_652_n205# w_n2112_n240# 0.24fF
C262 a_n1484_n205# w_n2112_n240# 0.24fF
C263 a_n594_n205# a_1008_n205# 0.01fF
C264 a_n1008_n140# a_416_n140# 0.01fF
C265 a_296_n205# a_1720_n205# 0.01fF
C266 a_830_n205# a_652_n205# 0.11fF
C267 a_n652_n140# a_n830_n140# 0.13fF
C268 a_1542_n205# a_1186_n205# 0.03fF
C269 a_474_n205# a_n416_n205# 0.01fF
C270 a_n772_n205# a_n238_n205# 0.02fF
C271 a_n830_n140# a_60_n140# 0.02fF
C272 a_n772_n205# a_n2018_n205# 0.01fF
C273 a_n118_n140# a_n1186_n140# 0.02fF
C274 a_1542_n205# a_296_n205# 0.01fF
C275 a_n1662_n205# w_n2112_n240# 0.24fF
C276 a_n772_n205# a_296_n205# 0.01fF
C277 a_594_n140# a_n1008_n140# 0.01fF
C278 a_n950_n205# a_n1306_n205# 0.03fF
C279 a_2018_n140# w_n2112_n240# 0.02fF
C280 a_652_n205# a_n594_n205# 0.01fF
C281 a_474_n205# a_n60_n205# 0.02fF
C282 a_n296_n140# a_238_n140# 0.04fF
C283 a_n1484_n205# a_n594_n205# 0.01fF
C284 a_1840_n140# a_1662_n140# 0.13fF
C285 a_n652_n140# a_60_n140# 0.03fF
C286 a_n1840_n205# a_n1484_n205# 0.03fF
C287 a_416_n140# a_1662_n140# 0.02fF
C288 a_1306_n140# a_1840_n140# 0.04fF
C289 a_1306_n140# a_416_n140# 0.02fF
C290 a_n1008_n140# a_n1720_n140# 0.03fF
C291 a_n474_n140# a_238_n140# 0.03fF
C292 a_474_n205# a_118_n205# 0.03fF
C293 a_n1662_n205# a_n594_n205# 0.01fF
C294 a_1128_n140# a_1662_n140# 0.04fF
C295 a_1484_n140# a_60_n140# 0.01fF
C296 a_n118_n140# a_n296_n140# 0.13fF
C297 a_n416_n205# a_n1306_n205# 0.01fF
C298 a_n1840_n205# a_n1662_n205# 0.11fF
C299 a_n1720_n140# a_n2076_n140# 0.06fF
C300 a_1306_n140# a_1128_n140# 0.13fF
C301 a_594_n140# a_1662_n140# 0.02fF
C302 a_2018_n140# a_950_n140# 0.02fF
C303 a_n950_n205# w_n2112_n240# 0.24fF
C304 a_772_n140# a_238_n140# 0.04fF
C305 a_594_n140# a_1306_n140# 0.03fF
C306 a_n1128_n205# a_n238_n205# 0.01fF
C307 a_n2018_n205# a_n1128_n205# 0.01fF
C308 a_n60_n205# a_n1306_n205# 0.01fF
C309 a_n118_n140# a_n474_n140# 0.06fF
C310 a_n1008_n140# a_n2076_n140# 0.02fF
C311 a_n1128_n205# a_296_n205# 0.01fF
C312 a_1364_n205# a_n60_n205# 0.01fF
C313 a_n1186_n140# a_416_n140# 0.01fF
C314 a_474_n205# a_1720_n205# 0.01fF
C315 a_118_n205# a_n1306_n205# 0.01fF
C316 a_772_n140# a_n118_n140# 0.02fF
C317 a_n416_n205# w_n2112_n240# 0.24fF
C318 a_n950_n205# a_n594_n205# 0.03fF
C319 a_n1542_n140# a_n1720_n140# 0.13fF
C320 a_118_n205# a_1364_n205# 0.01fF
C321 a_n950_n205# a_n1840_n205# 0.01fF
C322 a_830_n205# a_n416_n205# 0.01fF
C323 a_474_n205# a_1542_n205# 0.01fF
C324 w_n2112_n240# a_n60_n205# 0.24fF
C325 a_n1542_n140# a_n1008_n140# 0.04fF
C326 w_n2112_n240# a_238_n140# 0.02fF
C327 a_n1364_n140# a_238_n140# 0.01fF
C328 a_474_n205# a_n772_n205# 0.01fF
C329 a_n1720_n140# a_n1898_n140# 0.13fF
C330 a_n238_n205# a_1186_n205# 0.01fF
C331 a_830_n205# a_n60_n205# 0.01fF
C332 a_n1542_n140# a_n2076_n140# 0.04fF
C333 a_296_n205# a_n238_n205# 0.02fF
C334 a_n296_n140# a_416_n140# 0.03fF
C335 a_296_n205# a_1186_n205# 0.01fF
C336 a_n416_n205# a_n594_n205# 0.11fF
C337 a_652_n205# a_1008_n205# 0.03fF
C338 a_n1840_n205# a_n416_n205# 0.01fF
C339 a_n1008_n140# a_n1898_n140# 0.02fF
C340 a_118_n205# w_n2112_n240# 0.24fF
C341 a_n1720_n140# a_n1186_n140# 0.04fF
C342 w_n2112_n240# a_n118_n140# 0.02fF
C343 a_n118_n140# a_n1364_n140# 0.02fF
C344 a_1364_n205# a_1720_n205# 0.03fF
C345 a_1306_n140# a_1662_n140# 0.06fF
C346 a_n474_n140# a_416_n140# 0.02fF
C347 a_1128_n140# a_n296_n140# 0.01fF
C348 a_n60_n205# a_n594_n205# 0.02fF
C349 a_n2076_n140# a_n1898_n140# 0.13fF
C350 a_830_n205# a_118_n205# 0.01fF
C351 a_1898_n205# a_1720_n205# 0.11fF
C352 a_950_n140# a_238_n140# 0.03fF
C353 a_n1008_n140# a_n1186_n140# 0.13fF
C354 a_594_n140# a_n296_n140# 0.02fF
C355 a_2018_n140# a_1484_n140# 0.04fF
C356 a_n772_n205# a_n1306_n205# 0.02fF
C357 a_1542_n205# a_1364_n205# 0.11fF
C358 a_1128_n140# a_n474_n140# 0.01fF
C359 a_772_n140# a_1840_n140# 0.02fF
C360 a_n2076_n140# a_n1186_n140# 0.02fF
C361 a_772_n140# a_416_n140# 0.06fF
C362 a_1542_n205# a_1898_n205# 0.03fF
C363 a_118_n205# a_n594_n205# 0.01fF
C364 a_594_n140# a_n474_n140# 0.02fF
C365 a_474_n205# a_n1128_n205# 0.01fF
C366 w_n2112_n240# a_1720_n205# 0.18fF
C367 a_950_n140# a_n118_n140# 0.02fF
C368 a_n1720_n140# a_n296_n140# 0.01fF
C369 a_772_n140# a_1128_n140# 0.06fF
C370 a_n1542_n140# a_n1898_n140# 0.06fF
C371 a_830_n205# a_1720_n205# 0.01fF
C372 a_n1662_n205# a_n1484_n205# 0.11fF
C373 a_n1008_n140# a_n296_n140# 0.03fF
C374 a_772_n140# a_594_n140# 0.13fF
C375 a_n1720_n140# a_n474_n140# 0.02fF
C376 a_1542_n205# w_n2112_n240# 0.19fF
C377 a_n830_n140# a_238_n140# 0.02fF
C378 a_n772_n205# w_n2112_n240# 0.24fF
C379 a_n1542_n140# a_n1186_n140# 0.06fF
C380 w_n2112_n240# VSUBS 6.08fF
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6QKDBA a_n207_n140# a_n1039_n205# a_1275_n205#
+ a_29_n205# a_327_n140# a_n1275_n140# a_n683_n205# a_741_n205# a_n29_n140# a_149_n140#
+ a_n1097_n140# a_1097_n205# a_1395_n140# a_n505_n205# a_n741_n140# a_563_n205# a_861_n140#
+ a_919_n205# a_n327_n205# a_n563_n140# a_385_n205# a_1217_n140# a_n1395_n205# a_683_n140#
+ a_n919_n140# w_n1489_n240# a_n149_n205# a_1039_n140# a_n385_n140# a_207_n205# a_n1217_n205#
+ a_505_n140# a_n1453_n140# a_n861_n205# VSUBS
X0 a_n919_n140# a_n1039_n205# a_n1097_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X1 a_505_n140# a_385_n205# a_327_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X2 a_n385_n140# a_n505_n205# a_n563_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X3 a_1395_n140# a_1275_n205# a_1217_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X4 a_327_n140# a_207_n205# a_149_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X5 a_149_n140# a_29_n205# a_n29_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X6 a_861_n140# a_741_n205# a_683_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X7 a_n207_n140# a_n327_n205# a_n385_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X8 a_1217_n140# a_1097_n205# a_1039_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X9 a_n1275_n140# a_n1395_n205# a_n1453_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=4.06e+11p ps=3.38e+06u w=1.4e+06u l=600000u
X10 a_n741_n140# a_n861_n205# a_n919_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=4.06e+11p pd=3.38e+06u as=0p ps=0u w=1.4e+06u l=600000u
X11 a_n1097_n140# a_n1217_n205# a_n1275_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X12 a_683_n140# a_563_n205# a_505_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X13 a_1039_n140# a_919_n205# a_861_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X14 a_n29_n140# a_n149_n205# a_n207_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
X15 a_n563_n140# a_n683_n205# a_n741_n140# w_n1489_n240# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.4e+06u l=600000u
C0 a_919_n205# a_385_n205# 0.02fF
C1 a_327_n140# a_1395_n140# 0.02fF
C2 a_1097_n205# a_29_n205# 0.01fF
C3 a_n741_n140# a_n919_n140# 0.13fF
C4 a_n29_n140# a_n385_n140# 0.06fF
C5 a_327_n140# a_861_n140# 0.04fF
C6 a_n919_n140# a_n207_n140# 0.03fF
C7 a_563_n205# a_n861_n205# 0.01fF
C8 a_29_n205# a_563_n205# 0.02fF
C9 a_741_n205# a_1275_n205# 0.02fF
C10 a_1217_n140# a_505_n140# 0.03fF
C11 a_1275_n205# a_207_n205# 0.01fF
C12 a_n1097_n140# a_n1275_n140# 0.13fF
C13 a_741_n205# a_n327_n205# 0.01fF
C14 a_n327_n205# a_207_n205# 0.02fF
C15 a_n149_n205# a_385_n205# 0.02fF
C16 w_n1489_n240# a_n683_n205# 0.24fF
C17 w_n1489_n240# a_683_n140# 0.02fF
C18 a_1395_n140# a_861_n140# 0.04fF
C19 a_n1217_n205# a_n1039_n205# 0.11fF
C20 a_29_n205# a_n861_n205# 0.01fF
C21 a_n563_n140# a_505_n140# 0.02fF
C22 a_n741_n140# a_n1275_n140# 0.04fF
C23 a_n1275_n140# a_n207_n140# 0.02fF
C24 a_n563_n140# a_n1453_n140# 0.02fF
C25 a_683_n140# a_1039_n140# 0.06fF
C26 a_n327_n205# a_n683_n205# 0.03fF
C27 a_327_n140# a_149_n140# 0.13fF
C28 a_741_n205# a_385_n205# 0.03fF
C29 a_385_n205# a_207_n205# 0.11fF
C30 a_n1395_n205# a_n1039_n205# 0.03fF
C31 a_n29_n140# a_1217_n140# 0.02fF
C32 a_n741_n140# a_683_n140# 0.01fF
C33 a_1395_n140# a_149_n140# 0.02fF
C34 a_505_n140# w_n1489_n240# 0.02fF
C35 a_n1217_n205# a_n861_n205# 0.03fF
C36 a_683_n140# a_n207_n140# 0.02fF
C37 a_n1217_n205# a_29_n205# 0.01fF
C38 a_n29_n140# a_n563_n140# 0.04fF
C39 a_861_n140# a_149_n140# 0.03fF
C40 w_n1489_n240# a_n1453_n140# 0.02fF
C41 a_919_n205# a_n505_n205# 0.01fF
C42 a_327_n140# a_n919_n140# 0.02fF
C43 a_1217_n140# a_n385_n140# 0.01fF
C44 a_n683_n205# a_385_n205# 0.01fF
C45 w_n1489_n240# a_n1039_n205# 0.24fF
C46 a_505_n140# a_1039_n140# 0.04fF
C47 a_n1097_n140# a_505_n140# 0.01fF
C48 a_n563_n140# a_n385_n140# 0.13fF
C49 a_n1395_n205# a_n861_n205# 0.02fF
C50 a_n149_n205# a_n505_n205# 0.03fF
C51 a_n1395_n205# a_29_n205# 0.01fF
C52 a_n1097_n140# a_n1453_n140# 0.06fF
C53 a_1097_n205# w_n1489_n240# 0.18fF
C54 a_327_n140# a_n1275_n140# 0.01fF
C55 a_505_n140# a_n741_n140# 0.02fF
C56 a_n29_n140# w_n1489_n240# 0.02fF
C57 a_505_n140# a_n207_n140# 0.03fF
C58 a_n327_n205# a_n1039_n205# 0.01fF
C59 a_n741_n140# a_n1453_n140# 0.03fF
C60 a_n1453_n140# a_n207_n140# 0.02fF
C61 w_n1489_n240# a_563_n205# 0.21fF
C62 a_1097_n205# a_1275_n205# 0.11fF
C63 w_n1489_n240# a_n861_n205# 0.24fF
C64 a_1097_n205# a_n327_n205# 0.01fF
C65 w_n1489_n240# a_n385_n140# 0.02fF
C66 a_n29_n140# a_1039_n140# 0.02fF
C67 w_n1489_n240# a_29_n205# 0.24fF
C68 a_741_n205# a_n505_n205# 0.01fF
C69 a_n505_n205# a_207_n205# 0.01fF
C70 a_n1097_n140# a_n29_n140# 0.02fF
C71 a_327_n140# a_683_n140# 0.06fF
C72 a_n1395_n205# a_n1217_n205# 0.11fF
C73 a_919_n205# a_n149_n205# 0.01fF
C74 a_n919_n140# a_149_n140# 0.02fF
C75 a_563_n205# a_1275_n205# 0.01fF
C76 a_563_n205# a_n327_n205# 0.01fF
C77 a_n29_n140# a_n741_n140# 0.03fF
C78 a_385_n205# a_n1039_n205# 0.01fF
C79 a_1395_n140# a_683_n140# 0.03fF
C80 a_n29_n140# a_n207_n140# 0.13fF
C81 a_n385_n140# a_1039_n140# 0.01fF
C82 a_n327_n205# a_n861_n205# 0.02fF
C83 a_29_n205# a_1275_n205# 0.01fF
C84 a_29_n205# a_n327_n205# 0.03fF
C85 a_n1097_n140# a_n385_n140# 0.03fF
C86 a_861_n140# a_683_n140# 0.13fF
C87 a_n505_n205# a_n683_n205# 0.11fF
C88 a_1097_n205# a_385_n205# 0.01fF
C89 a_n741_n140# a_n385_n140# 0.06fF
C90 w_n1489_n240# a_n1217_n205# 0.24fF
C91 a_n1275_n140# a_149_n140# 0.01fF
C92 a_919_n205# a_741_n205# 0.11fF
C93 a_n385_n140# a_n207_n140# 0.13fF
C94 a_919_n205# a_207_n205# 0.01fF
C95 a_327_n140# a_505_n140# 0.13fF
C96 a_563_n205# a_385_n205# 0.11fF
C97 a_1217_n140# w_n1489_n240# 0.02fF
C98 a_385_n205# a_n861_n205# 0.01fF
C99 a_29_n205# a_385_n205# 0.03fF
C100 a_1395_n140# a_505_n140# 0.02fF
C101 a_741_n205# a_n149_n205# 0.01fF
C102 a_n1217_n205# a_n327_n205# 0.01fF
C103 a_n149_n205# a_207_n205# 0.03fF
C104 a_n563_n140# w_n1489_n240# 0.02fF
C105 a_n919_n140# a_n1275_n140# 0.06fF
C106 a_919_n205# a_n683_n205# 0.01fF
C107 w_n1489_n240# a_n1395_n205# 0.31fF
C108 a_683_n140# a_149_n140# 0.04fF
C109 a_505_n140# a_861_n140# 0.06fF
C110 a_1217_n140# a_1039_n140# 0.13fF
C111 a_n563_n140# a_1039_n140# 0.01fF
C112 a_327_n140# a_n29_n140# 0.06fF
C113 a_n149_n205# a_n683_n205# 0.02fF
C114 a_n1097_n140# a_n563_n140# 0.04fF
C115 a_n505_n205# a_n1039_n205# 0.02fF
C116 a_n1395_n205# a_n327_n205# 0.01fF
C117 a_1217_n140# a_n207_n140# 0.01fF
C118 a_741_n205# a_207_n205# 0.02fF
C119 a_n919_n140# a_683_n140# 0.01fF
C120 a_n1217_n205# a_385_n205# 0.01fF
C121 a_n29_n140# a_1395_n140# 0.01fF
C122 a_n563_n140# a_n741_n140# 0.13fF
C123 a_n563_n140# a_n207_n140# 0.06fF
C124 a_1097_n205# a_n505_n205# 0.01fF
C125 a_327_n140# a_n385_n140# 0.03fF
C126 a_n29_n140# a_861_n140# 0.02fF
C127 a_505_n140# a_149_n140# 0.06fF
C128 a_149_n140# a_n1453_n140# 0.01fF
C129 w_n1489_n240# a_1039_n140# 0.02fF
C130 w_n1489_n240# a_1275_n205# 0.24fF
C131 a_741_n205# a_n683_n205# 0.01fF
C132 a_n683_n205# a_207_n205# 0.01fF
C133 w_n1489_n240# a_n327_n205# 0.24fF
C134 a_563_n205# a_n505_n205# 0.01fF
C135 a_n1097_n140# w_n1489_n240# 0.02fF
C136 a_861_n140# a_n385_n140# 0.02fF
C137 a_n505_n205# a_n861_n205# 0.03fF
C138 a_29_n205# a_n505_n205# 0.02fF
C139 a_n741_n140# w_n1489_n240# 0.02fF
C140 a_505_n140# a_n919_n140# 0.01fF
C141 w_n1489_n240# a_n207_n140# 0.02fF
C142 a_n919_n140# a_n1453_n140# 0.04fF
C143 a_1275_n205# a_n327_n205# 0.01fF
C144 a_1097_n205# a_919_n205# 0.11fF
C145 a_n29_n140# a_149_n140# 0.13fF
C146 a_n149_n205# a_n1039_n205# 0.01fF
C147 w_n1489_n240# a_385_n205# 0.22fF
C148 a_327_n140# a_1217_n140# 0.02fF
C149 a_919_n205# a_563_n205# 0.03fF
C150 a_n1097_n140# a_n741_n140# 0.06fF
C151 a_1039_n140# a_n207_n140# 0.02fF
C152 a_n1097_n140# a_n207_n140# 0.02fF
C153 a_1097_n205# a_n149_n205# 0.01fF
C154 a_n385_n140# a_149_n140# 0.04fF
C155 a_n1275_n140# a_n1453_n140# 0.13fF
C156 a_n1217_n205# a_n505_n205# 0.01fF
C157 a_327_n140# a_n563_n140# 0.02fF
C158 a_919_n205# a_29_n205# 0.01fF
C159 a_1217_n140# a_1395_n140# 0.13fF
C160 a_n29_n140# a_n919_n140# 0.02fF
C161 a_n741_n140# a_n207_n140# 0.04fF
C162 a_1275_n205# a_385_n205# 0.01fF
C163 a_n327_n205# a_385_n205# 0.01fF
C164 a_1217_n140# a_861_n140# 0.06fF
C165 a_563_n205# a_n149_n205# 0.01fF
C166 a_207_n205# a_n1039_n205# 0.01fF
C167 a_n149_n205# a_n861_n205# 0.01fF
C168 a_505_n140# a_683_n140# 0.13fF
C169 a_29_n205# a_n149_n205# 0.11fF
C170 a_n563_n140# a_861_n140# 0.01fF
C171 a_n919_n140# a_n385_n140# 0.04fF
C172 a_1097_n205# a_741_n205# 0.03fF
C173 a_1097_n205# a_207_n205# 0.01fF
C174 a_n1395_n205# a_n505_n205# 0.01fF
C175 a_n29_n140# a_n1275_n140# 0.02fF
C176 a_327_n140# w_n1489_n240# 0.02fF
C177 a_n683_n205# a_n1039_n205# 0.03fF
C178 a_741_n205# a_563_n205# 0.11fF
C179 a_563_n205# a_207_n205# 0.03fF
C180 a_1395_n140# w_n1489_n240# 0.02fF
C181 a_1217_n140# a_149_n140# 0.02fF
C182 a_n1275_n140# a_n385_n140# 0.02fF
C183 a_741_n205# a_n861_n205# 0.01fF
C184 a_207_n205# a_n861_n205# 0.01fF
C185 a_741_n205# a_29_n205# 0.01fF
C186 a_29_n205# a_207_n205# 0.11fF
C187 a_861_n140# w_n1489_n240# 0.02fF
C188 a_327_n140# a_1039_n140# 0.03fF
C189 w_n1489_n240# a_n505_n205# 0.24fF
C190 a_n1217_n205# a_n149_n205# 0.01fF
C191 a_n1097_n140# a_327_n140# 0.01fF
C192 a_n29_n140# a_683_n140# 0.03fF
C193 a_n563_n140# a_149_n140# 0.03fF
C194 a_563_n205# a_n683_n205# 0.01fF
C195 a_1395_n140# a_1039_n140# 0.06fF
C196 a_327_n140# a_n741_n140# 0.02fF
C197 a_327_n140# a_n207_n140# 0.04fF
C198 a_861_n140# a_1039_n140# 0.13fF
C199 a_n683_n205# a_n861_n205# 0.11fF
C200 a_29_n205# a_n683_n205# 0.01fF
C201 a_683_n140# a_n385_n140# 0.02fF
C202 a_n327_n205# a_n505_n205# 0.11fF
C203 a_n1395_n205# a_n149_n205# 0.01fF
C204 a_n563_n140# a_n919_n140# 0.06fF
C205 a_1395_n140# a_n207_n140# 0.01fF
C206 a_n1217_n205# a_207_n205# 0.01fF
C207 a_861_n140# a_n741_n140# 0.01fF
C208 w_n1489_n240# a_149_n140# 0.02fF
C209 a_919_n205# w_n1489_n240# 0.19fF
C210 a_861_n140# a_n207_n140# 0.02fF
C211 a_n29_n140# a_505_n140# 0.04fF
C212 a_n29_n140# a_n1453_n140# 0.01fF
C213 a_n563_n140# a_n1275_n140# 0.03fF
C214 a_n505_n205# a_385_n205# 0.01fF
C215 a_n1217_n205# a_n683_n205# 0.02fF
C216 w_n1489_n240# a_n149_n205# 0.24fF
C217 a_1039_n140# a_149_n140# 0.02fF
C218 a_919_n205# a_1275_n205# 0.03fF
C219 a_n1395_n205# a_207_n205# 0.01fF
C220 a_919_n205# a_n327_n205# 0.01fF
C221 a_505_n140# a_n385_n140# 0.02fF
C222 a_n1097_n140# a_149_n140# 0.02fF
C223 a_n919_n140# w_n1489_n240# 0.02fF
C224 a_n385_n140# a_n1453_n140# 0.02fF
C225 a_563_n205# a_n1039_n205# 0.01fF
C226 a_1217_n140# a_683_n140# 0.04fF
C227 a_n741_n140# a_149_n140# 0.02fF
C228 a_149_n140# a_n207_n140# 0.06fF
C229 a_1275_n205# a_n149_n205# 0.01fF
C230 a_n861_n205# a_n1039_n205# 0.11fF
C231 a_n327_n205# a_n149_n205# 0.11fF
C232 a_29_n205# a_n1039_n205# 0.01fF
C233 a_n563_n140# a_683_n140# 0.02fF
C234 a_n1395_n205# a_n683_n205# 0.01fF
C235 a_1097_n205# a_563_n205# 0.02fF
C236 a_n1097_n140# a_n919_n140# 0.13fF
C237 w_n1489_n240# a_n1275_n140# 0.02fF
C238 w_n1489_n240# a_741_n205# 0.20fF
C239 w_n1489_n240# a_207_n205# 0.23fF
C240 w_n1489_n240# VSUBS 4.29fF
.ends

.subckt ota sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480#
+ m1_11825_n9711# sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# m1_12118_n9704# sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# m1_12410_n9718# m1_n6302_n3889# sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# sc_cmfb_0/transmission_gate_9/in m1_2463_n5585#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# m1_n947_n12836# sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480#
+ m1_11534_n9706# m1_11242_n9716# m1_n2176_n12171# sc_cmfb_0/transmission_gate_8/in
+ sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# p2_b
+ sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# sc_cmfb_0/transmission_gate_6/in ip
+ sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# m1_2462_n3318# cm m1_n208_n2883# in
+ sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS m1_6690_n8907# p1_b i_bias m1_n5574_n13620#
+ sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ sc_cmfb_0/transmission_gate_7/in bias_a sc_cmfb_0/transmission_gate_3/out bias_b
+ bias_d op p2 m1_1038_n2886# VDD sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# cmc
+ bias_c p1 on m1_n1659_n11581#
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_0 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_1 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_2 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_3 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_4 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_0 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_1 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_5 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_2 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_BASQVB_0 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias
+ i_bias i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_6 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_3 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_0 m1_n1659_n11581# bias_d VSS bias_d bias_a m1_n947_n12836#
+ m1_n1659_n11581# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# on op bias_d
+ bias_d op op on op bias_d VSS on m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n947_n12836#
+ bias_d bias_d bias_d VSS m1_n1659_n11581# m1_n1659_n11581# on VSS m1_n1659_n11581#
+ on m1_n947_n12836# m1_n947_n12836# bias_d bias_d op bias_d op bias_d m1_n947_n12836#
+ bias_d bias_d op VSS on VSS VSS on op bias_d bias_d m1_n1659_n11581# on on bias_d
+ bias_d bias_d VSS bias_d VSS m1_n947_n12836# m1_n1659_n11581# m1_n2176_n12171# VSS
+ m1_n947_n12836# bias_d bias_d op VSS m1_n947_n12836# bias_d m1_n1659_n11581# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_1 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias
+ bias_c i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_VU7MNH_7 bias_b bias_c bias_c bias_b bias_c bias_b bias_b
+ bias_c bias_b bias_b bias_b bias_b bias_b bias_c bias_b bias_c bias_b bias_b bias_b
+ VSS sky130_fd_pr__nfet_01v8_lvt_VU7MNH
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_4 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_1 m1_n947_n12836# bias_d bias_d bias_d op m1_n947_n12836#
+ m1_n2176_n12171# bias_d VSS bias_d VSS bias_d m1_n1659_n11581# on VSS bias_d bias_d
+ on bias_a bias_a bias_a bias_d bias_d bias_a m1_n1659_n11581# VSS bias_d on op VSS
+ VSS bias_d bias_d bias_d m1_n947_n12836# m1_n2176_n12171# bias_a bias_d m1_n947_n12836#
+ bias_a m1_n2176_n12171# m1_n1659_n11581# bias_d bias_d bias_a bias_d op VSS m1_n2176_n12171#
+ bias_d VSS bias_a bias_d VSS op bias_d bias_a on bias_d bias_d m1_n1659_n11581#
+ op on VSS bias_d bias_d on bias_d bias_d m1_n2176_n12171# VSS m1_n1659_n11581# bias_d
+ m1_n947_n12836# bias_d VSS bias_a op m1_n947_n12836# bias_d m1_n2176_n12171# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_2 bias_c VSS i_bias VSS i_bias i_bias i_bias i_bias
+ bias_c i_bias VSS i_bias VSS VSS bias_c bias_c i_bias i_bias i_bias bias_c VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_5 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_UFQYRB_2 m1_n947_n12836# bias_d VSS bias_d bias_a m1_n1659_n11581#
+ m1_n947_n12836# bias_d bias_d bias_d bias_d bias_d m1_n2176_n12171# op on bias_d
+ bias_d on on op on bias_d VSS op m1_n2176_n12171# bias_d bias_d VSS bias_a m1_n1659_n11581#
+ bias_d bias_d bias_d VSS m1_n947_n12836# m1_n947_n12836# op VSS m1_n947_n12836#
+ op m1_n1659_n11581# m1_n1659_n11581# bias_d bias_d on bias_d on bias_d m1_n1659_n11581#
+ bias_d bias_d on VSS op VSS VSS op on bias_d bias_d m1_n947_n12836# op op bias_d
+ bias_d bias_d VSS bias_d VSS m1_n1659_n11581# m1_n947_n12836# m1_n2176_n12171# VSS
+ m1_n1659_n11581# bias_d bias_d on VSS m1_n1659_n11581# bias_d m1_n947_n12836# VSS
+ sky130_fd_pr__nfet_01v8_UFQYRB
Xsky130_fd_pr__nfet_01v8_BASQVB_3 i_bias VSS i_bias VSS i_bias bias_c i_bias i_bias
+ i_bias i_bias VSS i_bias VSS VSS i_bias i_bias i_bias bias_c i_bias i_bias VSS VSS
+ i_bias VSS sky130_fd_pr__nfet_01v8_BASQVB
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_10 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_11 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_6 m1_n5574_n13620# m1_n208_n2883# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_12 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_7 m1_1038_n2886# m1_n5574_n13620# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_7P4E2J_0 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_KEEN2X_10 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS cmc cmc bias_a VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS cmc bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_13 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_8 m1_1038_n2886# m1_1038_n2886# m1_1038_n2886#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_KEEN2X_11 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS bias_a bias_a cmc VSS m1_n5574_n13620# cmc VSS bias_a bias_a
+ cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS bias_a cmc VSS VSS
+ m1_n5574_n13620# m1_n5574_n13620# bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc
+ VSS VSS bias_a cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620#
+ bias_a bias_a cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# bias_a cmc
+ cmc VSS VSS m1_n5574_n13620# bias_a cmc bias_a m1_n5574_n13620# m1_n5574_n13620#
+ VSS cmc bias_a VSS m1_n5574_n13620# bias_a cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_7P4E2J_1 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ bias_d bias_a m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_d
+ m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_a m1_6690_n8907# bias_a VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_9 m1_n5574_n13620# m1_1038_n2886# ip VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_14 m1_n208_n2883# m1_n5574_n13620# in VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_7P4E2J_2 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d bias_a
+ m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_a bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_7P4E2J_3 m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ bias_d bias_d m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d m1_6690_n8907# m1_6690_n8907#
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d
+ m1_6690_n8907# m1_6690_n8907# m1_6690_n8907# bias_d bias_d m1_6690_n8907# bias_d
+ m1_6690_n8907# bias_d VSS sky130_fd_pr__nfet_01v8_7P4E2J
Xsky130_fd_pr__nfet_01v8_lvt_TRAZV8_15 m1_n208_n2883# m1_n208_n2883# m1_n208_n2883#
+ VSS sky130_fd_pr__nfet_01v8_lvt_TRAZV8
Xsky130_fd_pr__nfet_01v8_KEEN2X_12 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS bias_a bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# bias_a VSS bias_a bias_a VSS
+ VSS m1_n5574_n13620# m1_n5574_n13620# cmc m1_n5574_n13620# VSS cmc bias_a VSS bias_a
+ VSS VSS cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS m1_n5574_n13620#
+ bias_a bias_a cmc m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc bias_a
+ bias_a VSS VSS m1_n5574_n13620# cmc cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS
+ cmc bias_a VSS m1_n5574_n13620# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_VJ4JGY_0 cm cm cm cm cm cm cm m1_11534_n9706# m1_11242_n9716#
+ cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711# cm cm cm cm VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_1 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490#
+ m1_11534_n9706# m1_11242_n9716# cm cm cm cm m1_12410_n9718# m1_12118_n9704# cm m1_11825_n9711#
+ m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_2 cm cm cm cm m1_11356_n10481# cm m1_11063_n10490#
+ m1_11534_n11258# m1_11244_n11260# cm cm cm cm m1_12410_n11263# m1_12118_n11263#
+ cm m1_11826_n11260# m1_11940_n10482# m1_12232_n10488# cm m1_11648_n10486# VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__nfet_01v8_VJ4JGY_3 cm cm cm cm VSS cm VSS m1_11534_n11258# m1_11244_n11260#
+ cm cm cm cm m1_12410_n11263# m1_12118_n11263# cm m1_11826_n11260# VSS VSS cm VSS
+ VSS sky130_fd_pr__nfet_01v8_VJ4JGY
Xsky130_fd_pr__pfet_01v8_E4DCBA_0 VDD bias_c m1_6690_n8907# op bias_c bias_c m1_1038_n2886#
+ bias_b bias_c VDD m1_n208_n2883# bias_c VDD on bias_c VDD VDD m1_2463_n5585# VDD
+ m1_2462_n3318# m1_2462_n3318# op m1_2463_n5585# m1_2462_n3318# VDD VDD VDD bias_b
+ bias_c m1_1038_n2886# bias_c m1_6690_n8907# VDD bias_c VDD VDD m1_2463_n5585# on
+ VDD bias_c m1_2462_n3318# m1_n208_n2883# bias_c bias_c VDD VDD m1_2463_n5585# VDD
+ VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_2 on VDD op on VDD bias_c m1_n208_n2883# on bias_c
+ bias_c VDD VDD m1_n208_n2883# op bias_c bias_c VDD m1_1038_n2886# bias_c m1_n208_n2883#
+ m1_n208_n2883# m1_n6302_n3889# m1_1038_n2886# m1_n208_n2883# m1_n6302_n3889# bias_c
+ bias_c on bias_c VDD bias_c op bias_c bias_c cm bias_c m1_1038_n2886# cm m1_1038_n2886#
+ VDD m1_n208_n2883# m1_1038_n2886# bias_c bias_c op bias_c m1_1038_n2886# bias_c
+ VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_1 op VDD on op VDD bias_c m1_1038_n2886# op bias_c
+ bias_c VDD VDD m1_1038_n2886# on bias_c bias_c VDD m1_n208_n2883# bias_c m1_1038_n2886#
+ m1_1038_n2886# m1_n6302_n3889# m1_n208_n2883# m1_1038_n2886# m1_n6302_n3889# bias_c
+ bias_c op bias_c VDD bias_c on bias_c bias_c cm bias_c m1_n208_n2883# cm m1_n208_n2883#
+ VDD m1_1038_n2886# m1_n208_n2883# bias_c bias_c on bias_c m1_n208_n2883# bias_c
+ VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsky130_fd_pr__pfet_01v8_E4DCBA_3 VDD bias_c bias_b on bias_c bias_c m1_n208_n2883#
+ m1_6690_n8907# bias_c VDD m1_1038_n2886# bias_c VDD op bias_c VDD VDD m1_2462_n3318#
+ VDD m1_2463_n5585# m1_2463_n5585# on m1_2462_n3318# m1_2463_n5585# VDD VDD VDD m1_6690_n8907#
+ bias_c m1_n208_n2883# bias_c bias_b VDD bias_c VDD VDD m1_2462_n3318# op VDD bias_c
+ m1_2463_n5585# m1_1038_n2886# bias_c bias_c VDD VDD m1_2462_n3318# VDD VSS sky130_fd_pr__pfet_01v8_E4DCBA
Xsc_cmfb_0 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_4/out sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580#
+ sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480#
+ bias_a sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# p2_b sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480#
+ p1 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480#
+ p2 VDD sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# sc_cmfb_0/transmission_gate_3/out sc_cmfb_0/transmission_gate_6/in
+ cmc sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# on sc_cmfb_0/transmission_gate_8/in
+ sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580#
+ sc_cmfb_0/transmission_gate_7/in cm sc_cmfb_0/transmission_gate_9/in sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480#
+ sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# p1_b VSS op sc_cmfb
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_0 m1_n208_n2883# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_1038_n2886# VDD VDD VDD bias_b VDD bias_b m1_1038_n2886# bias_b bias_b
+ m1_1038_n2886# bias_b VDD VDD VDD m1_n208_n2883# VDD bias_b VDD VDD bias_b VDD m1_n208_n2883#
+ VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_4 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS cmc cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS cmc cmc VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# bias_a m1_n5574_n13620# VSS bias_a cmc VSS cmc VSS VSS bias_a bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS m1_n5574_n13620# cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ bias_a bias_a m1_n5574_n13620# m1_n5574_n13620# VSS bias_a cmc VSS m1_n5574_n13620#
+ cmc cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_1 m1_2463_n5585# bias_b m1_2462_n3318# bias_b
+ VDD m1_2463_n5585# bias_b bias_b VDD m1_2462_n3318# VDD bias_b m1_2462_n3318# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2462_n3318# m1_2463_n5585#
+ VDD m1_1038_n2886# VDD bias_b VDD VDD bias_b bias_b m1_n208_n2883# m1_2463_n5585#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_5 VSS m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc
+ VSS bias_a VSS VSS bias_a cmc VSS m1_n5574_n13620# bias_a VSS cmc cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a VSS VSS bias_a VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# cmc m1_n5574_n13620# VSS bias_a cmc VSS bias_a VSS VSS cmc bias_a
+ m1_n5574_n13620# m1_n5574_n13620# VSS bias_a VSS VSS VSS cmc bias_a m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# cmc bias_a bias_a VSS VSS m1_n5574_n13620# cmc
+ cmc cmc m1_n5574_n13620# m1_n5574_n13620# VSS cmc cmc VSS m1_n5574_n13620# bias_a
+ bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_3 m1_2462_n3318# bias_b m1_2463_n5585# bias_b
+ VDD m1_2462_n3318# bias_b bias_b VDD m1_2463_n5585# VDD bias_b m1_2463_n5585# bias_b
+ VDD bias_b m1_1038_n2886# bias_b bias_b m1_n208_n2883# bias_b m1_2463_n5585# m1_2462_n3318#
+ VDD m1_1038_n2886# VDD bias_b VDD VDD bias_b bias_b m1_n208_n2883# m1_2462_n3318#
+ bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_2 m1_n6302_n3889# bias_b m1_n6302_n3889# bias_b
+ VDD m1_n6302_n3889# bias_b bias_b VDD m1_n6302_n3889# VDD bias_b m1_n6302_n3889#
+ bias_b VDD bias_b m1_n208_n2883# bias_b bias_b m1_1038_n2886# bias_b m1_n6302_n3889#
+ m1_n6302_n3889# VDD m1_n208_n2883# VDD bias_b VDD VDD bias_b bias_b m1_1038_n2886#
+ m1_n6302_n3889# bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_6 VSS VSS VSS VSS bias_a bias_a m1_n947_n12836# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n1659_n11581# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n947_n12836# bias_a m1_n1659_n11581# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n1659_n11581# m1_n947_n12836# bias_a bias_a bias_a
+ m1_n1659_n11581# m1_n2176_n12171# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__pfet_01v8_lvt_6QKDBA_4 m1_1038_n2886# bias_b VDD bias_b VDD VDD bias_b
+ bias_b VDD m1_n208_n2883# VDD VDD VDD bias_b VDD bias_b m1_n208_n2883# bias_b bias_b
+ m1_n208_n2883# bias_b VDD VDD VDD m1_1038_n2886# VDD bias_b VDD VDD bias_b VDD m1_1038_n2886#
+ VDD bias_b VSS sky130_fd_pr__pfet_01v8_lvt_6QKDBA
Xsky130_fd_pr__nfet_01v8_KEEN2X_7 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n1659_n11581# m1_n947_n12836# bias_a m1_n947_n12836# bias_a
+ bias_a bias_a VSS m1_n1659_n11581# m1_n2176_n12171# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n947_n12836# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n947_n12836# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n2176_n12171# m1_n1659_n11581# m1_n1659_n11581# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_KEEN2X_9 VSS m1_n5574_n13620# m1_n5574_n13620# VSS bias_a
+ bias_a VSS cmc VSS VSS cmc bias_a VSS m1_n5574_n13620# cmc VSS bias_a bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# m1_n5574_n13620# cmc VSS VSS cmc VSS VSS m1_n5574_n13620#
+ m1_n5574_n13620# bias_a m1_n5574_n13620# VSS cmc bias_a VSS cmc VSS VSS bias_a cmc
+ m1_n5574_n13620# m1_n5574_n13620# VSS cmc VSS VSS VSS bias_a cmc m1_n5574_n13620#
+ m1_n5574_n13620# m1_n5574_n13620# bias_a cmc cmc VSS VSS m1_n5574_n13620# bias_a
+ bias_a bias_a m1_n5574_n13620# m1_n5574_n13620# VSS bias_a bias_a VSS m1_n5574_n13620#
+ cmc cmc VSS sky130_fd_pr__nfet_01v8_KEEN2X
Xsky130_fd_pr__nfet_01v8_KEEN2X_8 VSS VSS VSS VSS bias_a bias_a m1_n1659_n11581# bias_a
+ VSS VSS bias_a bias_a m1_n947_n12836# m1_n947_n12836# bias_a m1_n1659_n11581# bias_a
+ bias_a bias_a VSS m1_n2176_n12171# m1_n1659_n11581# bias_a m1_n947_n12836# VSS bias_a
+ m1_n2176_n12171# VSS m1_n1659_n11581# m1_n2176_n12171# bias_a VSS VSS bias_a bias_a
+ VSS bias_a m1_n1659_n11581# VSS bias_a bias_a VSS VSS m1_n2176_n12171# bias_a VSS
+ VSS VSS bias_a bias_a VSS m1_n947_n12836# m1_n1659_n11581# bias_a bias_a bias_a
+ m1_n947_n12836# m1_n2176_n12171# m1_n947_n12836# bias_a bias_a bias_a VSS m1_n2176_n12171#
+ m1_n2176_n12171# bias_a bias_a VSS m1_n2176_n12171# bias_a bias_a VSS sky130_fd_pr__nfet_01v8_KEEN2X
C0 bias_b m1_1038_n2886# 10.79fF
C1 cm bias_a 0.62fF
C2 m1_12410_n9718# m1_11242_n9716# 0.02fF
C3 ip m1_n5574_n13620# 1.01fF
C4 m1_11826_n11260# m1_11244_n11260# 0.03fF
C5 VDD op 5.61fF
C6 m1_2463_n5585# m1_n208_n2883# 3.39fF
C7 on m1_n208_n2883# 0.40fF
C8 p1 op 0.00fF
C9 m1_2463_n5585# bias_c 2.57fF
C10 m1_11534_n11258# m1_12118_n11263# 0.03fF
C11 m1_11940_n10482# m1_11356_n10481# 0.03fF
C12 on bias_c 4.92fF
C13 m1_11940_n10482# m1_11648_n10486# 0.07fF
C14 VDD bias_a 0.11fF
C15 VDD sc_cmfb_0/transmission_gate_4/out 0.01fF
C16 p1 bias_a 0.04fF
C17 VDD cm 3.69fF
C18 p1 sc_cmfb_0/transmission_gate_4/out -0.00fF
C19 sc_cmfb_0/transmission_gate_8/in bias_a 0.02fF
C20 m1_12410_n9718# m1_11825_n9711# 0.03fF
C21 p1 cm 0.17fF
C22 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# bias_a 0.05fF
C23 cm m1_11534_n9706# 0.65fF
C24 bias_b in 0.09fF
C25 sc_cmfb_0/transmission_gate_8/in cm 0.04fF
C26 m1_11940_n10482# m1_11063_n10490# 0.02fF
C27 m1_2463_n5585# m1_1038_n2886# 3.88fF
C28 bias_b op 0.14fF
C29 on m1_1038_n2886# 3.37fF
C30 m1_n5574_n13620# m1_n208_n2883# 2.49fF
C31 m1_2462_n3318# m1_n208_n2883# 3.03fF
C32 on cmc 1.17fF
C33 m1_n5574_n13620# bias_c 0.50fF
C34 m1_2462_n3318# bias_c 4.04fF
C35 m1_6690_n8907# bias_d 35.87fF
C36 bias_b cm 0.36fF
C37 m1_11826_n11260# m1_12118_n11263# 0.07fF
C38 p1 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.00fF
C39 sc_cmfb_0/transmission_gate_8/in sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.08fF
C40 m1_n5574_n13620# m1_1038_n2886# 2.45fF
C41 m1_2462_n3318# m1_1038_n2886# 4.36fF
C42 m1_12118_n9704# m1_11242_n9716# 0.02fF
C43 cmc m1_n5574_n13620# 54.64fF
C44 m1_12118_n9704# m1_12118_n11263# 0.01fF
C45 sc_cmfb_0/transmission_gate_7/in cm 0.04fF
C46 m1_12410_n9718# m1_12410_n11263# 0.01fF
C47 on m1_n2176_n12171# 8.63fF
C48 m1_n1659_n11581# m1_n947_n12836# 9.35fF
C49 bias_b VDD 41.24fF
C50 m1_2463_n5585# op 0.25fF
C51 cm m1_11244_n11260# 0.55fF
C52 m1_n947_n12836# bias_d 16.58fF
C53 op on 7.65fF
C54 m1_11534_n11258# m1_12410_n11263# 0.02fF
C55 m1_11825_n9711# m1_11826_n11260# 0.01fF
C56 m1_12232_n10488# cm 0.57fF
C57 on bias_a 4.51fF
C58 m1_11825_n9711# m1_12118_n9704# 0.07fF
C59 m1_6690_n8907# m1_n208_n2883# 0.10fF
C60 m1_2463_n5585# cm 0.52fF
C61 m1_6690_n8907# bias_c 1.61fF
C62 cm on 1.01fF
C63 m1_n5574_n13620# m1_n2176_n12171# 0.57fF
C64 in m1_n5574_n13620# 2.04fF
C65 m1_n1659_n11581# bias_d 12.63fF
C66 i_bias ip 0.17fF
C67 op m1_n5574_n13620# 0.17fF
C68 m1_2462_n3318# op 0.28fF
C69 m1_n6302_n3889# m1_n208_n2883# 3.54fF
C70 m1_n6302_n3889# bias_c 3.58fF
C71 m1_2463_n5585# VDD 7.63fF
C72 m1_2462_n3318# bias_a 0.11fF
C73 m1_n5574_n13620# bias_a 21.14fF
C74 m1_6690_n8907# m1_1038_n2886# 0.28fF
C75 VDD on 5.69fF
C76 m1_6690_n8907# cmc 0.56fF
C77 p2_b p2 0.00fF
C78 p1 on 0.01fF
C79 cm m1_11242_n9716# 0.68fF
C80 cm m1_2462_n3318# 1.44fF
C81 cm m1_n5574_n13620# 0.02fF
C82 m1_11826_n11260# m1_12410_n11263# 0.03fF
C83 cm m1_12118_n11263# 0.57fF
C84 m1_n6302_n3889# m1_1038_n2886# 2.81fF
C85 i_bias m1_n208_n2883# 0.24fF
C86 i_bias bias_c 12.15fF
C87 m1_2463_n5585# bias_b 6.62fF
C88 VDD m1_2462_n3318# 7.01fF
C89 cm m1_11356_n10481# 0.58fF
C90 VDD m1_n5574_n13620# 0.03fF
C91 bias_b on 0.07fF
C92 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# cm 0.01fF
C93 m1_11534_n9706# m1_11242_n9716# 0.07fF
C94 cm m1_11648_n10486# 0.59fF
C95 cm m1_11825_n9711# 0.65fF
C96 m1_6690_n8907# m1_n2176_n12171# 0.00fF
C97 m1_n947_n12836# cmc 0.37fF
C98 cmc p2_b 0.01fF
C99 m1_6690_n8907# op 2.49fF
C100 i_bias m1_1038_n2886# 0.27fF
C101 cm m1_11063_n10490# 0.61fF
C102 m1_6690_n8907# bias_a 2.54fF
C103 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# p1 0.00fF
C104 m1_n6302_n3889# op 0.17fF
C105 bias_b m1_2462_n3318# 3.43fF
C106 bias_b m1_n5574_n13620# 0.11fF
C107 ip m1_n208_n2883# 1.08fF
C108 m1_6690_n8907# sc_cmfb_0/transmission_gate_4/out 0.01fF
C109 m1_11825_n9711# m1_11534_n9706# 0.07fF
C110 cm m1_6690_n8907# 4.14fF
C111 ip bias_c 0.11fF
C112 m1_n1659_n11581# cmc 0.44fF
C113 sc_cmfb_0/transmission_gate_9/in on 0.00fF
C114 cmc bias_d 0.03fF
C115 m1_2463_n5585# on 0.09fF
C116 m1_n947_n12836# m1_n2176_n12171# 10.60fF
C117 m1_n6302_n3889# cm 2.61fF
C118 m1_11534_n11258# m1_11826_n11260# 0.07fF
C119 m1_12410_n9718# m1_12118_n9704# 0.07fF
C120 cm m1_12410_n11263# 0.58fF
C121 op m1_n947_n12836# 1.19fF
C122 m1_11244_n11260# m1_11242_n9716# 0.01fF
C123 i_bias in 0.29fF
C124 VDD m1_6690_n8907# 3.64fF
C125 ip m1_1038_n2886# 1.68fF
C126 m1_11244_n11260# m1_12118_n11263# 0.02fF
C127 m1_n947_n12836# bias_a 21.86fF
C128 bias_c m1_n208_n2883# 8.21fF
C129 m1_n1659_n11581# m1_n2176_n12171# 10.31fF
C130 m1_n6302_n3889# VDD 3.85fF
C131 m1_2463_n5585# m1_2462_n3318# 4.55fF
C132 sc_cmfb_0/transmission_gate_7/in sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.02fF
C133 on m1_n5574_n13620# 0.06fF
C134 m1_2462_n3318# on 0.27fF
C135 bias_d m1_n2176_n12171# 8.59fF
C136 m1_n1659_n11581# op 8.09fF
C137 op bias_d 12.45fF
C138 cmc p2 0.00fF
C139 bias_b m1_6690_n8907# 0.39fF
C140 m1_n1659_n11581# bias_a 20.90fF
C141 m1_12232_n10488# m1_11356_n10481# 0.02fF
C142 m1_n208_n2883# m1_1038_n2886# 17.20fF
C143 cmc m1_n208_n2883# 0.14fF
C144 m1_12232_n10488# m1_11648_n10486# 0.03fF
C145 bias_c m1_1038_n2886# 7.06fF
C146 VDD p2_b 0.00fF
C147 ip in 3.13fF
C148 bias_d bias_a 8.20fF
C149 cmc bias_c 0.07fF
C150 m1_n6302_n3889# bias_b 2.49fF
C151 cm bias_d 0.08fF
C152 m1_11940_n10482# cm 0.59fF
C153 m1_12232_n10488# m1_11063_n10490# 0.02fF
C154 m1_12410_n9718# cm 0.64fF
C155 cmc m1_1038_n2886# 0.17fF
C156 m1_11534_n11258# cm 0.58fF
C157 m1_2463_n5585# m1_6690_n8907# 0.36fF
C158 m1_n2176_n12171# m1_n208_n2883# 0.09fF
C159 in m1_n208_n2883# 3.17fF
C160 cmc p1_b 0.03fF
C161 m1_11244_n11260# m1_12410_n11263# 0.02fF
C162 m1_6690_n8907# on 1.68fF
C163 m1_11825_n9711# m1_11242_n9716# 0.03fF
C164 bias_c m1_n2176_n12171# 0.02fF
C165 in bias_c 0.44fF
C166 op m1_n208_n2883# 3.85fF
C167 op bias_c 5.30fF
C168 m1_12410_n9718# m1_11534_n9706# 0.02fF
C169 m1_2463_n5585# m1_n6302_n3889# 0.56fF
C170 m1_n6302_n3889# on 0.08fF
C171 bias_a m1_n208_n2883# 0.04fF
C172 m1_11534_n11258# m1_11534_n9706# 0.01fF
C173 bias_a bias_c 0.00fF
C174 m1_11356_n10481# m1_11648_n10486# 0.07fF
C175 cm m1_n208_n2883# 0.17fF
C176 m1_n2176_n12171# m1_1038_n2886# 0.11fF
C177 in m1_1038_n2886# 1.58fF
C178 cm bias_c 3.39fF
C179 cmc m1_n2176_n12171# 1.14fF
C180 cmc in 0.04fF
C181 m1_6690_n8907# m1_n5574_n13620# 0.08fF
C182 m1_6690_n8907# m1_2462_n3318# 2.72fF
C183 op m1_1038_n2886# 0.78fF
C184 op cmc 1.53fF
C185 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# op 0.00fF
C186 m1_n947_n12836# on 8.70fF
C187 cm m1_11826_n11260# 0.58fF
C188 m1_11063_n10490# m1_11356_n10481# 0.07fF
C189 bias_b ip 0.07fF
C190 m1_n6302_n3889# m1_2462_n3318# 0.57fF
C191 m1_11063_n10490# m1_11648_n10486# 0.03fF
C192 bias_a m1_1038_n2886# 0.07fF
C193 VDD m1_n208_n2883# 15.19fF
C194 cmc bias_a 12.12fF
C195 VDD bias_c 10.55fF
C196 cm m1_1038_n2886# 1.34fF
C197 cm m1_12118_n9704# 0.64fF
C198 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# sc_cmfb_0/transmission_gate_4/out 0.00fF
C199 cm cmc 0.79fF
C200 m1_12118_n11263# m1_12410_n11263# 0.07fF
C201 bias_a p1_b 0.01fF
C202 cm p1_b 0.09fF
C203 m1_n1659_n11581# on 1.52fF
C204 op sc_cmfb_0/transmission_gate_3/out 0.00fF
C205 m1_12232_n10488# m1_11940_n10482# 0.07fF
C206 m1_n947_n12836# m1_n5574_n13620# 0.12fF
C207 on bias_d 13.96fF
C208 op m1_n2176_n12171# 1.95fF
C209 m1_11534_n11258# m1_11244_n11260# 0.07fF
C210 VDD m1_1038_n2886# 15.36fF
C211 i_bias m1_n5574_n13620# 0.12fF
C212 bias_b m1_n208_n2883# 9.15fF
C213 VDD cmc 0.08fF
C214 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VDD 0.02fF
C215 m1_11534_n9706# m1_12118_n9704# 0.03fF
C216 bias_b bias_c 25.24fF
C217 p1 cmc 0.00fF
C218 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# p1 -0.00fF
C219 bias_a m1_n2176_n12171# 23.78fF
C220 VDD p1_b -0.01fF
C221 p1 p1_b -0.00fF
C222 op bias_a 2.42fF
C223 m1_n1659_n11581# m1_n5574_n13620# 0.14fF
C224 cm op 0.76fF
C225 m1_1038_n2886# VSS -75.81fF
C226 m1_n208_n2883# VSS -83.40fF
C227 m1_n6302_n3889# VSS 10.46fF
C228 m1_2463_n5585# VSS 0.31fF
C229 sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VSS 1.37fF
C230 sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VSS 1.37fF
C231 sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VSS 1.37fF
C232 sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VSS 1.37fF
C233 sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# VSS 1.37fF
C234 sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VSS 1.37fF
C235 sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# VSS 1.37fF
C236 sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VSS 1.37fF
C237 sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VSS 1.37fF
C238 sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VSS 1.37fF
C239 sc_cmfb_0/transmission_gate_9/in VSS -27.99fF
C240 sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VSS 1.37fF
C241 sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VSS 1.37fF
C242 sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VSS 1.37fF
C243 sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VSS 1.37fF
C244 sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VSS 1.37fF
C245 p2 VSS 9.44fF
C246 p2_b VSS 3.15fF
C247 sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# VSS 1.37fF
C248 sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VSS 1.37fF
C249 sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# VSS 1.37fF
C250 sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VSS 1.37fF
C251 sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VSS 1.35fF
C252 sc_cmfb_0/transmission_gate_8/in VSS -0.37fF
C253 sc_cmfb_0/transmission_gate_6/in VSS 2.41fF
C254 sc_cmfb_0/transmission_gate_7/in VSS 1.93fF
C255 cm VSS -12.64fF
C256 p1 VSS 9.90fF
C257 op VSS -11.38fF
C258 sc_cmfb_0/transmission_gate_4/out VSS 0.87fF
C259 p1_b VSS 1.49fF
C260 VDD VSS 364.29fF
C261 on VSS -76.62fF
C262 sc_cmfb_0/transmission_gate_3/out VSS -4.68fF
C263 m1_2462_n3318# VSS -13.18fF
C264 m1_12410_n11263# VSS 0.18fF
C265 m1_12118_n11263# VSS 0.31fF
C266 m1_11826_n11260# VSS 0.32fF
C267 m1_11534_n11258# VSS 0.23fF
C268 m1_11244_n11260# VSS 0.24fF
C269 m1_12232_n10488# VSS 0.24fF
C270 m1_11940_n10482# VSS 0.35fF
C271 m1_11648_n10486# VSS 0.25fF
C272 m1_11356_n10481# VSS 0.27fF
C273 m1_11063_n10490# VSS 0.27fF
C274 m1_12410_n9718# VSS 0.17fF
C275 m1_12118_n9704# VSS 0.28fF
C276 m1_11825_n9711# VSS 0.29fF
C277 m1_11534_n9706# VSS 0.22fF
C278 m1_11242_n9716# VSS 0.23fF
C279 cmc VSS 33.96fF
C280 bias_a VSS -227.80fF
C281 m1_n5574_n13620# VSS 202.89fF
C282 m1_6690_n8907# VSS -73.62fF
C283 bias_c VSS 46.67fF
C284 i_bias VSS 34.74fF
C285 m1_n1659_n11581# VSS 8.89fF
C286 m1_n947_n12836# VSS 15.59fF
C287 in VSS 2.39fF
C288 m1_n2176_n12171# VSS 17.22fF
C289 bias_d VSS 120.47fF
C290 bias_b VSS 12.98fF
C291 ip VSS 2.32fF
.ends

.subckt sky130_fd_pr__nfet_01v8_E56BNL a_n33_32# a_15_n90# a_n73_n90# VSUBS
X0 a_15_n90# a_n33_32# a_n73_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
C0 a_n73_n90# a_15_n90# 0.14fF
C1 a_15_n90# a_n33_32# 0.01fF
C2 a_n73_n90# a_n33_32# 0.01fF
C3 a_15_n90# VSUBS 0.02fF
C4 a_n73_n90# VSUBS 0.02fF
C5 a_n33_32# VSUBS 0.15fF
.ends

.subckt switch_5t out en_b transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD in en VSS transmission_gate_1/in
Xtransmission_gate_0 en VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in transmission_gate_1/in VSS en_b transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_1/in out VSS en_b transmission_gate
Xsky130_fd_pr__nfet_01v8_E56BNL_0 en_b transmission_gate_1/in VSS VSS sky130_fd_pr__nfet_01v8_E56BNL
C0 out en_b 0.02fF
C1 en in 0.13fF
C2 transmission_gate_1/in en_b 0.23fF
C3 out VDD 0.16fF
C4 VDD transmission_gate_1/in 0.42fF
C5 en en_b 0.06fF
C6 out transmission_gate_1/in 0.72fF
C7 en_b in 0.12fF
C8 VDD in 0.10fF
C9 en transmission_gate_1/in 0.09fF
C10 out in 0.43fF
C11 transmission_gate_1/in in 0.68fF
C12 VDD en_b 0.57fF
C13 en VSS 3.45fF
C14 out VSS 0.90fF
C15 en_b VSS 0.55fF
C16 VDD VSS 10.85fF
C17 transmission_gate_1/in VSS 2.10fF
C18 in VSS 1.01fF
.ends

.subckt sky130_fd_sc_hd__inv_1 Y A VGND VPWR VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
C0 A VGND 0.05fF
C1 VPWR VGND 0.05fF
C2 VPB A 0.08fF
C3 VPB VPWR 0.21fF
C4 Y A 0.05fF
C5 Y VPWR 0.22fF
C6 Y VGND 0.17fF
C7 Y VPB 0.06fF
C8 A VPWR 0.05fF
C9 VGND VNB 0.25fF
C10 Y VNB 0.06fF
C11 VPWR VNB 0.06fF
C12 A VNB 0.13fF
C13 VPB VNB 0.34fF
.ends

.subckt a_mux2_en transmission_gate_1/en_b switch_5t_0/in switch_5t_1/transmission_gate_1/in
+ VDD switch_5t_0/transmission_gate_1/in in0 s0 out en switch_5t_1/in VSS in1 switch_5t_1/en
Xswitch_5t_0 out switch_5t_1/en switch_5t_0/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD switch_5t_0/in s0 VSS switch_5t_0/transmission_gate_1/in switch_5t
Xswitch_5t_1 out s0 switch_5t_1/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD switch_5t_1/in switch_5t_1/en VSS switch_5t_1/transmission_gate_1/in switch_5t
Xtransmission_gate_0 en VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in0 switch_5t_1/in VSS transmission_gate_1/en_b transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in1 switch_5t_0/in VSS transmission_gate_1/en_b transmission_gate
Xsky130_fd_sc_hd__inv_1_1 switch_5t_1/en s0 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 transmission_gate_1/en_b en VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
C0 switch_5t_0/transmission_gate_1/in VDD 0.06fF
C1 switch_5t_0/transmission_gate_1/in s0 0.07fF
C2 switch_5t_0/in in1 0.03fF
C3 transmission_gate_1/en_b switch_5t_1/in 0.09fF
C4 switch_5t_1/transmission_gate_1/in switch_5t_1/in 0.02fF
C5 in1 in0 0.51fF
C6 en switch_5t_1/in 0.07fF
C7 switch_5t_0/transmission_gate_1/in transmission_gate_1/en_b 0.01fF
C8 switch_5t_1/transmission_gate_1/in out 0.21fF
C9 switch_5t_1/en switch_5t_1/in 0.21fF
C10 out switch_5t_1/en 0.03fF
C11 switch_5t_0/transmission_gate_1/in switch_5t_1/transmission_gate_1/in 0.33fF
C12 switch_5t_0/in switch_5t_1/in 0.36fF
C13 s0 VDD 0.21fF
C14 switch_5t_0/transmission_gate_1/in switch_5t_1/en 0.03fF
C15 in0 switch_5t_1/in 0.02fF
C16 switch_5t_0/transmission_gate_1/in switch_5t_0/in 0.06fF
C17 transmission_gate_1/en_b VDD 0.28fF
C18 switch_5t_1/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# en 0.00fF
C19 s0 transmission_gate_1/en_b 0.04fF
C20 switch_5t_0/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# switch_5t_0/in 0.00fF
C21 switch_5t_1/transmission_gate_1/in VDD 0.25fF
C22 switch_5t_1/transmission_gate_1/in s0 0.12fF
C23 en VDD 0.04fF
C24 s0 en 0.18fF
C25 switch_5t_1/en VDD 0.09fF
C26 switch_5t_1/en s0 0.78fF
C27 switch_5t_0/in VDD 0.17fF
C28 in1 switch_5t_1/in 0.08fF
C29 switch_5t_0/in s0 0.02fF
C30 transmission_gate_1/en_b en 0.44fF
C31 in0 VDD 0.07fF
C32 switch_5t_1/en transmission_gate_1/en_b 0.05fF
C33 s0 in0 0.02fF
C34 switch_5t_0/in transmission_gate_1/en_b 0.14fF
C35 switch_5t_1/transmission_gate_1/in switch_5t_1/en 0.10fF
C36 switch_5t_1/en en 0.24fF
C37 switch_5t_1/transmission_gate_1/in switch_5t_0/in 0.06fF
C38 in0 transmission_gate_1/en_b 0.12fF
C39 switch_5t_0/in en 0.13fF
C40 switch_5t_1/en switch_5t_0/in 0.06fF
C41 switch_5t_0/transmission_gate_1/in switch_5t_1/in 0.07fF
C42 switch_5t_0/transmission_gate_1/in out 0.15fF
C43 in1 VDD -0.15fF
C44 in0 en 0.05fF
C45 in1 s0 0.00fF
C46 switch_5t_1/en in0 0.03fF
C47 switch_5t_0/in in0 0.08fF
C48 switch_5t_1/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# switch_5t_1/in 0.00fF
C49 in1 transmission_gate_1/en_b 0.10fF
C50 switch_5t_1/in VDD 0.35fF
C51 s0 switch_5t_1/in 0.14fF
C52 out VDD 0.35fF
C53 out s0 0.14fF
C54 in1 en 0.05fF
C55 VDD VSS 29.38fF
C56 en VSS 5.89fF
C57 switch_5t_0/in VSS 1.76fF
C58 in1 VSS 0.51fF
C59 transmission_gate_1/en_b VSS 0.96fF
C60 switch_5t_1/in VSS 1.12fF
C61 in0 VSS 0.58fF
C62 switch_5t_1/en VSS 7.48fF
C63 out VSS 0.88fF
C64 s0 VSS 5.14fF
C65 switch_5t_1/transmission_gate_1/in VSS 1.97fF
C66 switch_5t_0/transmission_gate_1/in VSS 1.72fF
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VPWR X a_1290_413# a_757_363#
+ a_1478_413# a_277_47# VNB VPB a_750_97# a_27_413# a_923_363# a_193_47# a_834_97#
+ a_247_21# a_668_97# a_193_413# a_27_47#
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=2.226e+11p pd=2.74e+06u as=2.184e+11p ps=2.72e+06u w=420000u l=150000u
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=6.142e+11p pd=7.3e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=2.1715e+11p pd=2.72e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=7.039e+11p ps=8e+06u w=420000u l=150000u
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.822e+11p pd=3.5e+06u as=2.171e+11p ps=2.72e+06u w=420000u l=150000u
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=2.184e+11p pd=2.72e+06u as=2.7965e+11p ps=3.21e+06u w=420000u l=150000u
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.083e+11p ps=1.36e+06u w=420000u l=150000u
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.84175e+11p ps=1.98e+06u w=420000u l=150000u
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.8025e+11p pd=1.99e+06u as=0p ps=0u w=420000u l=150000u
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0205e+11p ps=2.57e+06u w=420000u l=150000u
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.171e+11p pd=2.72e+06u as=0p ps=0u w=420000u l=150000u
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 A0 A3 0.01fF
C1 a_750_97# a_27_47# 0.01fF
C2 a_27_413# S0 0.00fF
C3 a_193_413# a_27_47# 0.02fF
C4 a_750_97# S1 0.06fF
C5 a_750_97# A2 0.03fF
C6 A1 A3 0.01fF
C7 A0 VGND 0.04fF
C8 a_1290_413# A3 0.02fF
C9 a_750_97# a_277_47# 0.44fF
C10 VPB X 0.05fF
C11 a_193_413# a_277_47# 0.12fF
C12 a_247_21# a_668_97# 0.04fF
C13 A1 VGND 0.03fF
C14 a_750_97# S0 0.16fF
C15 a_750_97# a_923_363# 0.00fF
C16 a_1290_413# VGND 0.17fF
C17 a_193_413# S0 0.02fF
C18 a_750_97# a_27_413# 0.01fF
C19 a_668_97# a_1478_413# 0.01fF
C20 a_193_413# a_27_413# 0.12fF
C21 a_247_21# VPWR 0.21fF
C22 a_247_21# a_757_363# 0.06fF
C23 a_1290_413# X 0.03fF
C24 a_1478_413# VPWR 0.34fF
C25 a_1478_413# a_757_363# 0.01fF
C26 a_193_413# a_750_97# 0.01fF
C27 a_834_97# a_1290_413# 0.02fF
C28 a_247_21# a_27_47# 0.07fF
C29 a_247_21# S1 0.04fF
C30 a_247_21# A2 0.04fF
C31 A3 VGND 0.02fF
C32 a_1478_413# a_27_47# 0.01fF
C33 a_247_21# a_277_47# 0.60fF
C34 a_1478_413# S1 0.02fF
C35 a_1478_413# A2 0.01fF
C36 A3 X 0.00fF
C37 a_277_47# a_1478_413# 0.18fF
C38 a_247_21# S0 0.45fF
C39 a_247_21# a_27_413# 0.02fF
C40 VPB VPWR 0.82fF
C41 a_1478_413# S0 0.01fF
C42 a_193_47# a_27_47# 0.02fF
C43 A0 VPWR 0.04fF
C44 X VGND 0.08fF
C45 VPB a_757_363# 0.04fF
C46 a_27_413# a_1478_413# 0.00fF
C47 a_834_97# A3 0.05fF
C48 a_1290_413# a_668_97# 0.01fF
C49 a_247_21# a_750_97# 0.24fF
C50 A1 VPWR 0.04fF
C51 a_247_21# a_193_413# 0.17fF
C52 a_1290_413# VPWR 0.17fF
C53 a_834_97# VGND 0.18fF
C54 a_750_97# a_1478_413# 0.24fF
C55 a_1290_413# a_757_363# 0.03fF
C56 VPB S1 0.17fF
C57 A0 a_27_47# 0.07fF
C58 a_193_413# a_1478_413# 0.00fF
C59 VPB A2 0.07fF
C60 a_834_97# X 0.01fF
C61 A0 S1 0.01fF
C62 A0 A2 0.01fF
C63 a_277_47# VPB 0.05fF
C64 A0 a_277_47# 0.11fF
C65 A1 a_27_47# 0.06fF
C66 VPB S0 0.30fF
C67 A1 S1 0.01fF
C68 a_1290_413# a_27_47# 0.01fF
C69 A1 A2 0.01fF
C70 a_668_97# A3 0.02fF
C71 a_27_413# VPB 0.04fF
C72 A0 S0 0.03fF
C73 a_1290_413# S1 0.22fF
C74 a_1290_413# A2 0.03fF
C75 A1 a_277_47# 0.02fF
C76 a_27_413# A0 0.08fF
C77 a_1290_413# a_277_47# 0.60fF
C78 A3 VPWR 0.02fF
C79 a_668_97# VGND 0.37fF
C80 A1 S0 0.02fF
C81 A3 a_757_363# 0.04fF
C82 a_27_413# A1 0.06fF
C83 a_1290_413# S0 0.02fF
C84 a_750_97# VPB 0.08fF
C85 a_1290_413# a_27_413# 0.00fF
C86 a_193_413# VPB 0.05fF
C87 a_668_97# X 0.00fF
C88 VPWR VGND 0.27fF
C89 a_750_97# A0 0.01fF
C90 a_193_413# A0 0.01fF
C91 a_757_363# VGND 0.03fF
C92 a_247_21# a_1478_413# 0.02fF
C93 VPWR X 0.09fF
C94 a_750_97# A1 0.01fF
C95 A3 S1 0.05fF
C96 A3 A2 0.20fF
C97 X a_757_363# 0.01fF
C98 a_834_97# a_668_97# 0.11fF
C99 a_750_97# a_1290_413# 0.23fF
C100 a_277_47# A3 0.02fF
C101 a_193_413# a_1290_413# 0.01fF
C102 a_27_47# VGND 0.39fF
C103 a_834_97# VPWR 0.03fF
C104 S1 VGND 0.04fF
C105 A2 VGND 0.02fF
C106 A3 S0 0.04fF
C107 a_277_47# VGND 0.54fF
C108 a_834_97# a_757_363# 0.04fF
C109 X a_27_47# 0.00fF
C110 X S1 0.01fF
C111 A2 X 0.00fF
C112 a_277_47# X 0.04fF
C113 S0 VGND 0.06fF
C114 a_247_21# VPB 0.23fF
C115 a_27_413# VGND 0.03fF
C116 a_834_97# a_27_47# 0.01fF
C117 a_247_21# A0 0.12fF
C118 a_750_97# A3 0.05fF
C119 X S0 0.00fF
C120 a_834_97# A2 0.07fF
C121 VPB a_1478_413# 0.11fF
C122 a_27_413# X 0.00fF
C123 A0 a_1478_413# 0.00fF
C124 a_834_97# a_277_47# 0.05fF
C125 a_247_21# A1 0.05fF
C126 a_668_97# VPWR 0.02fF
C127 a_750_97# VGND 0.22fF
C128 a_247_21# a_1290_413# 0.04fF
C129 a_193_413# VGND 0.02fF
C130 a_668_97# a_757_363# 0.02fF
C131 a_1290_413# a_1478_413# 0.15fF
C132 a_750_97# X 0.04fF
C133 a_193_413# X 0.00fF
C134 VPWR a_757_363# 0.40fF
C135 a_668_97# a_27_47# 0.02fF
C136 a_750_97# a_834_97# 0.08fF
C137 a_277_47# a_668_97# 0.01fF
C138 VPWR a_27_47# 0.03fF
C139 A0 VPB 0.10fF
C140 VPWR S1 0.05fF
C141 VPWR A2 0.04fF
C142 a_247_21# A3 0.09fF
C143 a_277_47# VPWR 0.26fF
C144 a_668_97# S0 0.03fF
C145 A2 a_757_363# 0.05fF
C146 A3 a_1478_413# 0.01fF
C147 A1 VPB 0.14fF
C148 a_277_47# a_757_363# 0.03fF
C149 a_247_21# VGND 0.23fF
C150 a_1290_413# VPB 0.13fF
C151 A0 A1 0.17fF
C152 VPWR S0 0.07fF
C153 a_923_363# VPWR 0.01fF
C154 a_1290_413# A0 0.01fF
C155 a_27_413# VPWR 0.15fF
C156 S0 a_757_363# 0.04fF
C157 a_1478_413# VGND 0.31fF
C158 a_923_363# a_757_363# 0.02fF
C159 a_247_21# X 0.01fF
C160 a_27_413# a_757_363# 0.01fF
C161 A2 S1 0.09fF
C162 a_750_97# a_668_97# 0.11fF
C163 a_277_47# a_27_47# 0.14fF
C164 a_1290_413# A1 0.01fF
C165 a_1478_413# X 0.22fF
C166 a_277_47# S1 0.06fF
C167 a_277_47# A2 0.02fF
C168 a_750_97# VPWR 0.32fF
C169 S0 a_27_47# 0.02fF
C170 a_247_21# a_834_97# 0.05fF
C171 a_193_413# VPWR 0.31fF
C172 a_27_413# a_27_47# 0.04fF
C173 S0 S1 0.03fF
C174 a_750_97# a_757_363# 0.21fF
C175 A2 S0 0.03fF
C176 a_193_47# VGND 0.00fF
C177 a_193_413# a_757_363# 0.03fF
C178 a_277_47# S0 0.07fF
C179 a_834_97# a_1478_413# 0.01fF
C180 VPB A3 0.07fF
C181 a_27_413# a_277_47# 0.11fF
C182 VGND VNB 1.06fF
C183 X VNB 0.05fF
C184 S1 VNB 0.21fF
C185 A2 VNB 0.08fF
C186 A3 VNB 0.09fF
C187 S0 VNB 0.34fF
C188 VPWR VNB 0.41fF
C189 A0 VNB 0.10fF
C190 A1 VNB 0.15fF
C191 VPB VNB 1.93fF
C192 a_834_97# VNB 0.02fF
C193 a_668_97# VNB 0.03fF
C194 a_27_47# VNB 0.03fF
C195 a_1478_413# VNB 0.11fF
C196 a_1290_413# VNB 0.15fF
C197 a_750_97# VNB 0.03fF
C198 a_277_47# VNB 0.07fF
C199 a_247_21# VNB 0.27fF
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_XAYTAL a_n129_n203# a_n173_n100# w_n311_n319#
+ VSUBS
X0 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=1.28e+12p pd=1.056e+07u as=0p ps=0u w=1e+06u l=150000u
X1 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n173_n100# a_n129_n203# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 w_n311_n319# a_n173_n100# 0.42fF
C1 w_n311_n319# a_n129_n203# 0.51fF
C2 a_n173_n100# a_n129_n203# 0.30fF
C3 w_n311_n319# VSUBS 1.19fF
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X a_110_47# VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.045e+12p pd=2.809e+07u as=5.6e+11p ps=5.12e+06u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.24e+12p ps=2.048e+07u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.8e+06u as=1.2789e+12p ps=1.533e+07u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.408e+11p ps=1.12e+07u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_110_47# VGND 0.78fF
C1 X VPWR 2.96fF
C2 VPWR VPB 0.78fF
C3 X VPB 0.03fF
C4 VPWR A 0.07fF
C5 VPWR a_110_47# 0.98fF
C6 X A 0.00fF
C7 VPWR VGND 0.28fF
C8 X a_110_47# 2.36fF
C9 VPB A 0.23fF
C10 X VGND 1.95fF
C11 a_110_47# VPB 0.81fF
C12 a_110_47# A 0.51fF
C13 VGND A 0.10fF
C14 VGND VNB 1.05fF
C15 X VNB 0.10fF
C16 VPWR VNB 0.39fF
C17 A VNB 0.43fF
C18 VPB VNB 1.85fF
C19 a_110_47# VNB 1.28fF
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=1.05e+06u
C0 VPWR VPB 0.27fF
C1 VPWR VGND 0.82fF
C2 VGND VPB 0.25fF
C3 VPWR VNB 0.41fF
C4 VGND VNB 0.37fF
C5 VPB VNB 0.43fF
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=2.89e+06u
C0 VPB VPWR 0.37fF
C1 VGND VPWR 1.92fF
C2 VGND VPB 0.55fF
C3 VPWR VNB 0.86fF
C4 VGND VNB 0.56fF
C5 VPB VNB 0.78fF
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=4.73e+06u
C0 VGND VPB 0.87fF
C1 VPWR VGND 3.03fF
C2 VPWR VPB 0.47fF
C3 VPWR VNB 1.33fF
C4 VGND VNB 0.77fF
C5 VPB VNB 1.14fF
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VPWR X VNB VPB a_283_47# a_390_47#
+ a_27_47#
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.173e+11p pd=2.17e+06u as=6.517e+11p ps=5.37e+06u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.173e+11p ps=2.17e+06u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=4.027e+11p pd=3.97e+06u as=1.7225e+11p ps=1.83e+06u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=3.55e+11p pd=2.71e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.491e+11p pd=1.55e+06u as=0p ps=0u w=420000u l=150000u
C0 VPWR A 0.02fF
C1 X A 0.00fF
C2 VGND a_283_47# 0.14fF
C3 a_27_47# a_390_47# 0.05fF
C4 a_27_47# VPB 0.16fF
C5 VPB a_390_47# 0.06fF
C6 a_283_47# VPWR 0.17fF
C7 a_283_47# X 0.04fF
C8 a_27_47# A 0.29fF
C9 A a_390_47# 0.01fF
C10 VGND VPWR 0.11fF
C11 VGND X 0.14fF
C12 A VPB 0.06fF
C13 VPWR X 0.19fF
C14 a_283_47# a_27_47# 0.18fF
C15 a_283_47# a_390_47# 0.44fF
C16 VGND a_27_47# 0.24fF
C17 VGND a_390_47# 0.14fF
C18 a_283_47# VPB 0.12fF
C19 a_283_47# A 0.02fF
C20 VPWR a_27_47# 0.31fF
C21 VPWR a_390_47# 0.16fF
C22 VGND A 0.02fF
C23 X a_27_47# 0.02fF
C24 X a_390_47# 0.12fF
C25 VPWR VPB 0.32fF
C26 X VPB 0.05fF
C27 VGND VNB 0.43fF
C28 X VNB 0.05fF
C29 VPWR VNB 0.16fF
C30 A VNB 0.13fF
C31 VPB VNB 0.78fF
C32 a_390_47# VNB 0.10fF
C33 a_283_47# VNB 0.18fF
C34 a_27_47# VNB 0.18fF
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB a_27_47#
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.08e+12p pd=1.016e+07u as=1.33e+12p ps=1.266e+07u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 Y VPB 0.02fF
C1 VPB A 0.18fF
C2 VPWR VPB 0.43fF
C3 B VPB 0.21fF
C4 Y a_27_47# 0.41fF
C5 Y VGND 0.13fF
C6 Y A 0.35fF
C7 a_27_47# VGND 0.77fF
C8 Y VPWR 1.44fF
C9 a_27_47# A 0.10fF
C10 a_27_47# VPWR 0.07fF
C11 Y B 0.30fF
C12 A VGND 0.08fF
C13 VPWR VGND 0.12fF
C14 B a_27_47# 0.33fF
C15 VPWR A 0.09fF
C16 B VGND 0.10fF
C17 B A 0.16fF
C18 B VPWR 0.12fF
C19 VGND VNB 0.48fF
C20 Y VNB 0.01fF
C21 VPWR VNB 0.18fF
C22 A VNB 0.26fF
C23 B VNB 0.30fF
C24 VPB VNB 0.87fF
C25 a_27_47# VNB 0.06fF
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=4.524e+11p pd=4.52e+06u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=2.86e+11p pd=3.24e+06u as=0p ps=0u w=550000u l=590000u
C0 VPWR VPB 0.24fF
C1 VGND VPB 0.16fF
C2 VPWR VGND 0.54fF
C3 VPWR VNB 0.28fF
C4 VGND VNB 0.31fF
C5 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__dfxbp_1 CLK D VGND VPWR Q Q_N a_975_413# a_891_413# VNB VPB
+ a_466_413# a_592_47# a_1059_315# a_193_47# a_561_413# a_634_159# a_381_47# a_1017_47#
+ a_1490_369# a_27_47#
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=9.432e+11p ps=1.006e+07u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=1.368e+11p pd=1.48e+06u as=1.978e+11p ps=1.99e+06u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.32905e+12p pd=1.228e+07u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X4 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=0p ps=0u w=420000u l=150000u
X5 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.392e+11p ps=1.53e+06u w=420000u l=150000u
X6 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1059_315# a_1490_369# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.19e+11p pd=2.15e+06u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.68e+06u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.32e+11p ps=1.49e+06u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.242e+11p ps=1.41e+06u w=360000u l=150000u
X17 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.626e+11p ps=1.66e+06u w=360000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X22 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X23 Q_N a_1490_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q_N a_1490_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X27 VPWR a_1059_315# a_1490_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
C0 D a_1059_315# 0.02fF
C1 D VPWR 0.03fF
C2 D a_1490_369# 0.01fF
C3 Q_N D 0.00fF
C4 a_891_413# a_1059_315# 0.44fF
C5 VPWR a_891_413# 0.20fF
C6 a_466_413# Q 0.02fF
C7 CLK a_466_413# 0.01fF
C8 a_975_413# a_891_413# 0.02fF
C9 VPB a_1059_315# 0.24fF
C10 Q_N a_891_413# 0.02fF
C11 a_1490_369# a_891_413# 0.04fF
C12 VPB VPWR 0.73fF
C13 a_1490_369# VPB 0.06fF
C14 Q_N VPB 0.05fF
C15 D a_466_413# 0.03fF
C16 CLK Q 0.00fF
C17 a_592_47# a_466_413# 0.01fF
C18 a_193_47# VGND 0.24fF
C19 a_466_413# a_891_413# 0.04fF
C20 a_193_47# a_381_47# 0.22fF
C21 a_381_47# VGND 0.09fF
C22 VPB a_466_413# 0.08fF
C23 a_634_159# a_193_47# 0.21fF
C24 D Q 0.00fF
C25 a_193_47# a_27_47# 1.69fF
C26 D CLK 0.04fF
C27 a_634_159# VGND 0.18fF
C28 a_27_47# VGND 0.30fF
C29 a_634_159# a_381_47# 0.03fF
C30 a_27_47# a_381_47# 0.16fF
C31 a_1017_47# VGND 0.00fF
C32 Q a_891_413# 0.04fF
C33 CLK a_891_413# 0.01fF
C34 a_634_159# a_27_47# 0.29fF
C35 VPB Q 0.02fF
C36 VPB CLK 0.14fF
C37 a_193_47# a_1059_315# 0.13fF
C38 a_193_47# VPWR 0.37fF
C39 VPWR a_561_413# 0.01fF
C40 VGND a_1059_315# 0.22fF
C41 VPWR VGND 0.26fF
C42 a_381_47# a_1059_315# 0.01fF
C43 VPWR a_381_47# 0.13fF
C44 D a_891_413# 0.01fF
C45 a_193_47# a_1490_369# 0.03fF
C46 Q_N a_193_47# 0.02fF
C47 a_1490_369# VGND 0.12fF
C48 Q_N VGND 0.11fF
C49 a_1490_369# a_381_47# 0.01fF
C50 Q_N a_381_47# 0.01fF
C51 D VPB 0.13fF
C52 a_634_159# a_1059_315# 0.06fF
C53 a_634_159# VPWR 0.21fF
C54 a_27_47# a_1059_315# 0.14fF
C55 VPWR a_27_47# 0.60fF
C56 a_634_159# a_1490_369# 0.02fF
C57 Q_N a_634_159# 0.01fF
C58 a_1490_369# a_27_47# 0.03fF
C59 Q_N a_27_47# 0.02fF
C60 VPB a_891_413# 0.08fF
C61 a_193_47# a_466_413# 0.20fF
C62 a_466_413# a_561_413# 0.01fF
C63 a_466_413# VGND 0.15fF
C64 a_381_47# a_466_413# 0.09fF
C65 VPWR a_1059_315# 0.37fF
C66 a_975_413# VPWR 0.01fF
C67 a_1490_369# a_1059_315# 0.18fF
C68 a_634_159# a_466_413# 0.36fF
C69 Q_N a_1059_315# 0.03fF
C70 a_1490_369# VPWR 0.29fF
C71 Q_N VPWR 0.25fF
C72 a_27_47# a_466_413# 0.51fF
C73 a_193_47# Q 0.03fF
C74 a_193_47# CLK 0.06fF
C75 Q_N a_1490_369# 0.14fF
C76 Q VGND 0.14fF
C77 CLK VGND 0.04fF
C78 a_381_47# Q 0.01fF
C79 CLK a_381_47# 0.01fF
C80 a_466_413# a_1059_315# 0.05fF
C81 VPWR a_466_413# 0.31fF
C82 a_634_159# Q 0.02fF
C83 a_634_159# CLK 0.01fF
C84 a_27_47# Q 0.03fF
C85 CLK a_27_47# 0.33fF
C86 D a_193_47# 0.30fF
C87 D VGND 0.05fF
C88 a_1490_369# a_466_413# 0.02fF
C89 Q_N a_466_413# 0.01fF
C90 D a_381_47# 0.21fF
C91 a_193_47# a_891_413# 0.38fF
C92 a_592_47# VGND 0.00fF
C93 a_891_413# VGND 0.18fF
C94 a_381_47# a_891_413# 0.02fF
C95 D a_634_159# 0.04fF
C96 D a_27_47# 0.17fF
C97 a_193_47# VPB 0.21fF
C98 Q a_1059_315# 0.19fF
C99 CLK a_1059_315# 0.01fF
C100 VPWR Q 0.24fF
C101 CLK VPWR 0.03fF
C102 VPB a_381_47# 0.03fF
C103 a_634_159# a_891_413# 0.10fF
C104 a_27_47# a_891_413# 0.09fF
C105 a_1490_369# Q 0.31fF
C106 Q_N Q 0.05fF
C107 Q_N CLK 0.00fF
C108 a_1490_369# CLK 0.00fF
C109 a_1017_47# a_891_413# 0.01fF
C110 a_634_159# VPB 0.08fF
C111 VPB a_27_47# 0.30fF
C112 Q_N VNB 0.05fF
C113 Q VNB 0.01fF
C114 VGND VNB 0.95fF
C115 VPWR VNB 0.37fF
C116 D VNB 0.12fF
C117 CLK VNB 0.18fF
C118 VPB VNB 1.76fF
C119 a_381_47# VNB 0.03fF
C120 a_1490_369# VNB 0.09fF
C121 a_891_413# VNB 0.12fF
C122 a_1059_315# VNB 0.24fF
C123 a_466_413# VNB 0.11fF
C124 a_634_159# VNB 0.12fF
C125 a_193_47# VNB 0.21fF
C126 a_27_47# VNB 0.31fF
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=5.2e+11p pd=5.04e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 VPWR VPB 0.24fF
C1 Y A 0.11fF
C2 A B 0.07fF
C3 Y VPB 0.02fF
C4 VGND a_113_47# 0.01fF
C5 VPWR VGND 0.05fF
C6 VPB B 0.06fF
C7 Y a_113_47# 0.01fF
C8 Y VPWR 0.40fF
C9 Y VGND 0.21fF
C10 VPWR B 0.06fF
C11 VPB A 0.06fF
C12 VGND B 0.06fF
C13 VPWR A 0.05fF
C14 Y B 0.05fF
C15 VGND A 0.02fF
C16 VGND VNB 0.23fF
C17 Y VNB 0.05fF
C18 VPWR VNB 0.06fF
C19 A VNB 0.10fF
C20 B VNB 0.10fF
C21 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=2.268e+11p pd=2.22e+06u as=4.536e+11p ps=4.44e+06u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=1.197e+11p pd=1.41e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 VGND VPWR 0.04fF
C1 Y A 0.26fF
C2 Y VPB 0.00fF
C3 Y VPWR 0.35fF
C4 A VPB 0.14fF
C5 VGND Y 0.17fF
C6 A VPWR 0.04fF
C7 VGND A 0.05fF
C8 VPB VPWR 0.23fF
C9 VGND VNB 0.23fF
C10 Y VNB 0.04fF
C11 VPWR VNB 0.06fF
C12 A VNB 0.24fF
C13 VPB VNB 0.34fF
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB a_505_21# a_439_47# a_218_47#
+ a_76_199# a_218_374#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=4.553e+11p pd=4.29e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=1.533e+11p pd=1.57e+06u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=5.155e+11p pd=4.31e+06u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=3.864e+11p pd=2.68e+06u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.995e+11p ps=1.79e+06u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
C0 A1 S 0.25fF
C1 A1 A0 0.41fF
C2 A1 VPB 0.06fF
C3 a_76_199# VPWR 0.15fF
C4 S A0 0.09fF
C5 VGND VPWR 0.12fF
C6 VPWR a_505_21# 0.12fF
C7 S VPB 0.24fF
C8 A1 X 0.04fF
C9 a_218_374# S 0.01fF
C10 A0 VPB 0.08fF
C11 VGND a_439_47# 0.01fF
C12 X S 0.08fF
C13 a_76_199# VGND 0.24fF
C14 a_76_199# a_505_21# 0.04fF
C15 a_76_199# a_218_47# 0.01fF
C16 X A0 0.02fF
C17 X VPB 0.06fF
C18 VGND a_505_21# 0.16fF
C19 VGND a_218_47# 0.01fF
C20 A1 VPWR 0.04fF
C21 a_535_374# S 0.01fF
C22 A1 a_439_47# 0.00fF
C23 S VPWR 0.64fF
C24 VPWR A0 0.01fF
C25 a_76_199# A1 0.41fF
C26 VPWR VPB 0.44fF
C27 VGND A1 0.12fF
C28 A1 a_505_21# 0.16fF
C29 a_439_47# A0 0.01fF
C30 a_76_199# S 0.54fF
C31 a_76_199# A0 0.14fF
C32 X VPWR 0.23fF
C33 VGND S 0.07fF
C34 S a_505_21# 0.26fF
C35 a_76_199# VPB 0.08fF
C36 a_76_199# a_218_374# 0.00fF
C37 VGND A0 0.08fF
C38 A0 a_505_21# 0.08fF
C39 a_505_21# VPB 0.09fF
C40 a_76_199# X 0.18fF
C41 VGND X 0.09fF
C42 X a_505_21# 0.02fF
C43 VGND VNB 0.48fF
C44 A1 VNB 0.09fF
C45 A0 VNB 0.08fF
C46 S VNB 0.17fF
C47 VPWR VNB 0.18fF
C48 X VNB 0.06fF
C49 VPB VNB 0.87fF
C50 a_505_21# VNB 0.15fF
C51 a_76_199# VNB 0.11fF
.ends

.subckt clock_v2 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A sky130_fd_sc_hd__mux2_1_0/a_439_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__dfxbp_1_1/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__clkinv_1_2/Y
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__dfxbp_1_1/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__mux2_1_0/a_76_199#
+ p2_b sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47#
+ sky130_fd_sc_hd__clkbuf_16_14/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47#
+ sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47#
+ Ad_b sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47#
+ A_b sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47#
+ sky130_fd_sc_hd__clkbuf_16_15/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__nand2_4_0/B
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47#
+ sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47#
+ sky130_fd_sc_hd__clkinv_4_7/Y sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Bd p1d_b sky130_fd_sc_hd__clkdlybuf4s50_1_125/X
+ sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47#
+ sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__nand2_1_1/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47#
+ sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47#
+ sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__dfxbp_1_0/a_891_413#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_4_1/B
+ sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# p2d sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__mux2_1_0/S Ad sky130_fd_sc_hd__dfxbp_1_1/a_592_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__nand2_4_3/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_975_413# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47#
+ sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47#
+ sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413#
+ sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__nand2_4_1/Y
+ sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X
+ sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__dfxbp_1_1/a_193_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47#
+ p1 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# p1_b sky130_fd_sc_hd__clkdlybuf4s50_1_154/X
+ sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47#
+ sky130_fd_sc_hd__clkbuf_16_2/a_110_47# sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__dfxbp_1_0/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_4/Y sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47#
+ B p1d sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47#
+ sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47#
+ sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47#
+ sky130_fd_sc_hd__nand2_1_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/X sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/A clk sky130_fd_sc_hd__clkdlybuf4s50_1_56/X
+ sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A
+ sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47#
+ Bd_b sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/X p2d_b sky130_fd_sc_hd__clkdlybuf4s50_1_127/X
+ B_b sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__dfxbp_1_0/a_634_159#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47#
+ sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_136/A p2 sky130_fd_sc_hd__clkinv_4_5/Y
+ sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
+ sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkbuf_16_7/a_110_47#
+ VSUBS sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VDD VSS sky130_fd_sc_hd__clkdlybuf4s50_1_93/A
+ sky130_fd_sc_hd__nand2_4_2/Y
Xsky130_fd_sc_hd__clkbuf_16_11 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD p1d_b sky130_fd_sc_hd__clkbuf_16_11/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_248 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_237 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_226 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_215 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_204 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_90 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_170 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_12 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD p2d_b sky130_fd_sc_hd__clkbuf_16_12/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_249 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_238 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_227 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_216 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_205 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_80 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_91 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_160 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_13 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD p2d sky130_fd_sc_hd__clkbuf_16_13/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_239 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_228 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_217 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_206 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_0 sky130_fd_sc_hd__clkinv_1_0/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_70 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_81 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_92 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_150 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_161 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_14 sky130_fd_sc_hd__clkinv_4_10/Y VSS VDD p2_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_10 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_4_10/Y
+ sky130_fd_sc_hd__clkinv_4_10/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_229 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_218 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_207 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_1 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_60 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_71 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_82 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_93 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_140 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_151 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_162 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_15 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD p2 sky130_fd_sc_hd__clkbuf_16_15/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_4_11 sky130_fd_sc_hd__nand2_4_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/A
+ sky130_fd_sc_hd__clkinv_4_11/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_219 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_208 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_2 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_130 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_72 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_61 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_50 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_83 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_94 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_152 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_141 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_163 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_4_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/Y VSUBS VDD sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_209 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_3 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS VDD sky130_fd_sc_hd__nand2_4_0/B
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_62 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_120 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_40 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_73 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_84 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_95 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_131 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_142 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_153 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_164 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/Y VSUBS VDD sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkinv_4_0 sky130_fd_sc_hd__nand2_4_0/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/A
+ sky130_fd_sc_hd__clkinv_4_0/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_52 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_110 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_63 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_74 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_85 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_121 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_96 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_132 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_154 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_143 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_165 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__nand2_4_2 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__nand2_4_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/Y VSUBS VDD sky130_fd_sc_hd__nand2_4_2/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__decap_4_190 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_5 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__clkinv_4_1/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_53 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_42 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_64 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_75 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_86 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_111 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_97 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_122 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_100 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_133 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_166 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_155 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_144 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_191 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_180 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_4_3 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_4_3/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_3/Y VSUBS VDD sky130_fd_sc_hd__nand2_4_3/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_6 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__clkinv_4_2/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_54 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_65 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_123 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_76 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_87 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_98 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_112 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_101 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_167 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_156 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_134 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_145 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_4_170 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_192 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_181 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__clkinv_4_3/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_55 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_66 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_113 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_77 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_124 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_88 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_102 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_99 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_168 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_157 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_146 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_135 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_193 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_160 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_171 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_182 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_8 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/X
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__clkinv_4_4/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_125 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_45 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_67 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_78 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_114 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_89 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_103 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_169 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_147 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_158 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_136 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_150 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_161 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_172 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_183 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_194 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_5 sky130_fd_sc_hd__nand2_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_4_5/Y
+ sky130_fd_sc_hd__clkinv_4_5/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_4_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_57 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_126 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_46 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_115 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_68 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_104 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_79 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_159 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_137 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_148 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_195 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_140 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_151 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_162 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_173 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_184 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_4_6 sky130_fd_sc_hd__nand2_4_2/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/A
+ sky130_fd_sc_hd__clkinv_4_6/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_190 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_127 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_36 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_58 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_69 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_116 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_105 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_149 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_138 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_196 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_141 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_130 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_152 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_163 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_174 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_185 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_90 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_7 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_4_7/Y
+ sky130_fd_sc_hd__clkinv_4_7/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_90 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_59 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_37 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_191 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_180 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_117 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_128 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_106 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_139 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_120 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_142 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_131 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_153 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_164 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_175 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_186 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_197 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_80 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_8 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD sky130_fd_sc_hd__clkinv_4_8/Y
+ sky130_fd_sc_hd__clkinv_4_8/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_91 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_80 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_129 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_107 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_38 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_118 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_49 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_121 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_110 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_143 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_132 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_154 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_165 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_176 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_198 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_187 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_92 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkinv_4_9 sky130_fd_sc_hd__nand2_4_3/Y VSS VDD sky130_fd_sc_hd__clkinv_4_9/Y
+ sky130_fd_sc_hd__clkinv_4_9/w_82_21# VSUBS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__decap_8_92 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_70 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_193 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_182 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_81 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_119 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_108 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_39 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_100 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_122 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_111 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_144 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_133 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_155 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_166 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_177 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_199 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_188 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_71 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_82 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_93 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_0 p2 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__mux2_1_0/S
+ sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__dfxbp_1_0/a_975_413# sky130_fd_sc_hd__dfxbp_1_0/a_891_413#
+ VSUBS VDD sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_592_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__dfxbp_1_0/a_1017_47#
+ sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_93 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_71 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_60 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_172 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_82 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_150 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_109 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_101 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_123 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_112 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_145 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_134 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_156 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_167 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_178 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_189 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_50 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_61 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__dfxbp_1_1 clk sky130_fd_sc_hd__dfxbp_1_1/D VSS VDD sky130_fd_sc_hd__nand2_1_1/A
+ sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__dfxbp_1_1/a_975_413# sky130_fd_sc_hd__dfxbp_1_1/a_891_413#
+ VSUBS VDD sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_592_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_561_413#
+ sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# sky130_fd_sc_hd__dfxbp_1_1/a_1017_47#
+ sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__decap_8_94 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_72 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_61 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_50 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_195 sky130_fd_sc_hd__clkinv_4_9/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/X
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_184 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_173 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_140 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_83 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_162 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_102 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_124 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_113 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_146 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_135 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_157 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_168 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_179 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_73 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_84 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_95 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_95 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_73 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_62 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_51 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_40 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_84 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_141 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_196 sky130_fd_sc_hd__clkinv_1_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_174 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_152 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_163 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_103 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_125 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_114 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_136 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_147 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_158 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_169 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_52 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_63 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_96 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_74 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_63 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_52 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_41 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_96 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_197 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_186 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_164 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_131 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_85 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_142 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD B sky130_fd_sc_hd__clkbuf_16_0/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_104 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_115 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_137 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_126 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_148 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_159 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_42 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_20 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_31 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_75 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_86 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_97 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_1/B VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_97 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_75 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_64 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_53 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_198 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_42 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_187 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_121 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_86 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_132 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_154 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_1 sky130_fd_sc_hd__nand2_4_0/Y VSS VDD Bd sky130_fd_sc_hd__clkbuf_16_1/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_116 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_105 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_138 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_127 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_149 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_10 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_54 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_32 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_65 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_87 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_10 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_98 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_21 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_65 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_76 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_54 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_43 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_199 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_3/B VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_177 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_100 sky130_fd_sc_hd__clkinv_1_2/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_87 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_122 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS VDD
+ sky130_fd_sc_hd__nand2_1_4/B VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_32 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_2 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD B_b sky130_fd_sc_hd__clkbuf_16_2/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_117 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_106 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_139 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_128 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_22 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_44 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_11 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_77 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_99 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/X
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_11 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_99 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_77 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_66 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_55 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_44 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_178 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_167 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_112 sky130_fd_sc_hd__clkinv_4_8/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_101 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_22 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_88 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_123 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_134 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_33 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkbuf_16_3 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD Bd_b sky130_fd_sc_hd__clkbuf_16_3/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_107 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_118 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_129 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_56 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_34 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_67 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_78 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_89 sky130_fd_sc_hd__clkinv_1_1/Y VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A
+ VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_67 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_12 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_56 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_45 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_78 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_34 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_157 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_102 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_23 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_89 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_113 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_146 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_168 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_12_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_4 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD Ad_b sky130_fd_sc_hd__clkbuf_16_4/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_4_119 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_108 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_24 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_13 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_68 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_0/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_46 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_68 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_57 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_79 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_24 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_35 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_169 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_2/B VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_103 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS VDD
+ sky130_fd_sc_hd__nand2_4_2/B VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_125 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_136 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_147 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_158 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_5 sky130_fd_sc_hd__nand2_4_1/Y VSS VDD Ad sky130_fd_sc_hd__clkbuf_16_5/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_12_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_4_109 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkdlybuf4s50_1_25 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_47 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_58 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_36 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_69 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_69 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_14 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_58 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_47 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_104 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_25 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_36 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_159 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_6 sky130_fd_sc_hd__clkinv_4_4/Y VSS VDD A_b sky130_fd_sc_hd__clkbuf_16_6/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_15 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_48 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_59 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_15 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_59 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_48 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_26 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_116 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_127 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_138 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_37 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_149 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkbuf_16_7 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD A sky130_fd_sc_hd__clkbuf_16_7/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_49 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS VDD
+ sky130_fd_sc_hd__nand2_1_1/B VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_27 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_38 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_250 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_16 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_49 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_38 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_117 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_27 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_0 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_0/A VSUBS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_8 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD p1 sky130_fd_sc_hd__clkbuf_16_8/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__decap_8_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_17 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_39 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_251 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_240 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_17 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_39 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_107 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_118 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_129 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_8_28 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nand2_1_1 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_1/A VSUBS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkbuf_16_9 sky130_fd_sc_hd__clkinv_4_7/Y VSS VDD p1_b sky130_fd_sc_hd__clkbuf_16_9/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_0 sky130_fd_sc_hd__clkinv_4_1/A VSS VDD sky130_fd_sc_hd__clkinv_1_0/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_18 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__clkdlybuf4s50_1_29 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_252 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_241 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_230 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_18 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_29 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_108 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_2 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_1_2/B
+ VSS VDD sky130_fd_sc_hd__nand2_4_2/A VSUBS VDD sky130_fd_sc_hd__nand2_1_2/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_1 sky130_fd_sc_hd__clkinv_4_5/Y VSS VDD sky130_fd_sc_hd__clkinv_1_1/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_253 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_242 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_231 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_220 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_8_19 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__clkdlybuf4s50_1_109 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS VDD
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSUBS VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47#
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__nand2_1_3/A clk VSS VDD sky130_fd_sc_hd__nand2_4_3/A
+ VSUBS VDD sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_2 sky130_fd_sc_hd__clkinv_4_7/A VSS VDD sky130_fd_sc_hd__clkinv_1_2/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_254 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_243 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_232 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_221 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_210 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__nand2_1_4 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/B
+ VSS VDD sky130_fd_sc_hd__nand2_1_4/Y VSUBS VDD sky130_fd_sc_hd__nand2_1_4/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__clkinv_1_3 sky130_fd_sc_hd__clkinv_1_3/A VSS VDD sky130_fd_sc_hd__clkinv_1_3/Y
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_255 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_244 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_233 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_222 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_211 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_200 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux2_1_0 Ad_b Bd_b sky130_fd_sc_hd__mux2_1_0/S VSS VDD sky130_fd_sc_hd__mux2_1_0/X
+ VSUBS VDD sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/a_439_47#
+ sky130_fd_sc_hd__mux2_1_0/a_218_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374#
+ sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkinv_1_4 sky130_fd_sc_hd__nand2_1_4/Y VSS VDD sky130_fd_sc_hd__nand2_1_3/A
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_245 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_234 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_223 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_212 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_201 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkinv_1_5 sky130_fd_sc_hd__nand2_1_1/A VSS VDD sky130_fd_sc_hd__nand2_1_0/B
+ VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_246 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_235 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_224 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_213 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_202 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_30 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_16_10 sky130_fd_sc_hd__nand2_4_2/Y VSS VDD p1d sky130_fd_sc_hd__clkbuf_16_10/a_110_47#
+ VSUBS VDD sky130_fd_sc_hd__clkbuf_16
Xsky130_fd_sc_hd__clkinv_1_6 clk VSS VDD sky130_fd_sc_hd__nand2_1_2/A VSUBS VDD sky130_fd_sc_hd__clkinv_1
Xsky130_fd_sc_hd__decap_4_247 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_236 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_225 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_214 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_203 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_12_31 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_12_20 VSS VDD VSUBS VDD sky130_fd_sc_hd__decap_12
C0 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.15fF
C1 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C2 sky130_fd_sc_hd__clkinv_4_9/Y Ad_b 0.03fF
C3 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.08fF
C4 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.34fF
C5 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.01fF
C6 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C7 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C8 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.07fF
C9 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C10 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.02fF
C11 sky130_fd_sc_hd__mux2_1_0/S Bd_b 0.12fF
C12 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C13 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C14 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C15 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C16 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C17 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C18 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C19 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_8/Y 0.68fF
C20 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C21 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.02fF
C22 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C23 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C24 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.03fF
C25 VDD sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.46fF
C26 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__nand2_4_2/A 0.13fF
C27 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C28 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.00fF
C29 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.00fF
C30 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C31 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.10fF
C32 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# Ad_b 0.06fF
C33 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C34 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C35 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C36 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# -0.00fF
C37 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C38 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.09fF
C39 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 1.13fF
C40 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C41 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.00fF
C42 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.15fF
C43 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.31fF
C44 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C45 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C46 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C47 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.19fF
C48 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.16fF
C49 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.05fF
C50 sky130_fd_sc_hd__clkinv_4_5/Y VSUBS 0.27fF
C51 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.04fF
C52 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.04fF
C53 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.08fF
C54 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.01fF
C55 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C56 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.01fF
C57 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.05fF
C58 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C59 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C60 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C61 sky130_fd_sc_hd__dfxbp_1_1/D clk 0.04fF
C62 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.01fF
C63 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.09fF
C64 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C65 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C66 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C67 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C68 p1 p1d 0.20fF
C69 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# -0.00fF
C70 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.06fF
C71 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.07fF
C72 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__nand2_1_1/B 0.03fF
C73 VDD sky130_fd_sc_hd__nand2_4_3/Y 6.10fF
C74 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkinv_1_2/Y 0.03fF
C75 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Bd_b 0.10fF
C76 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.10fF
C77 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C78 Ad_b sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C79 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.00fF
C80 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.02fF
C81 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.02fF
C82 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.16fF
C83 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_561_413# 0.01fF
C84 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.04fF
C85 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.08fF
C86 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C87 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.19fF
C88 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.03fF
C89 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_3/A 0.49fF
C90 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C91 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C92 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.15fF
C93 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.00fF
C94 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.05fF
C95 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.02fF
C96 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.00fF
C97 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C98 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C99 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 1.48fF
C100 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C101 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C102 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C103 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.04fF
C104 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C105 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C106 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.05fF
C107 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C108 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_2/B 0.23fF
C109 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C110 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C111 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.05fF
C112 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Ad_b 0.12fF
C113 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__mux2_1_0/S 0.03fF
C114 sky130_fd_sc_hd__nand2_4_1/B Ad_b 0.06fF
C115 p1d_b sky130_fd_sc_hd__clkinv_4_8/Y 0.03fF
C116 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.42fF
C117 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.04fF
C118 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C119 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C120 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C121 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__nand2_4_0/A 2.21fF
C122 sky130_fd_sc_hd__clkinv_4_2/Y Bd_b 0.10fF
C123 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.15fF
C124 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C125 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C126 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C127 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C128 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C129 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C130 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C131 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.05fF
C132 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C133 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_7/Y 0.02fF
C134 sky130_fd_sc_hd__clkinv_4_10/Y VSUBS 0.01fF
C135 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.08fF
C136 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.14fF
C137 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.02fF
C138 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.02fF
C139 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C140 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C141 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C142 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C143 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.02fF
C144 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C145 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkinv_4_9/w_82_21# 0.05fF
C146 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C147 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 2.24fF
C148 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.03fF
C149 VDD Bd 1.53fF
C150 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C151 VDD B 1.54fF
C152 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C153 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.00fF
C154 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C155 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.27fF
C156 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C157 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C158 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C159 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C160 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C161 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C162 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C163 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C164 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C165 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C166 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C167 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.01fF
C168 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C169 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.01fF
C170 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C171 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C172 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C173 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C174 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C175 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C176 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.13fF
C177 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C178 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.04fF
C179 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.15fF
C180 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C181 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/D 0.02fF
C182 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 1.14fF
C183 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C184 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 2.25fF
C185 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C186 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C187 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C188 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.12fF
C189 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C190 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C191 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 2.26fF
C192 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.10fF
C193 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.10fF
C194 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/A -0.58fF
C195 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C196 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C197 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.14fF
C198 VSUBS sky130_fd_sc_hd__nand2_4_0/A -0.18fF
C199 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.00fF
C200 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C201 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkinv_1_2/Y 0.69fF
C202 p1d_b sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.06fF
C203 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.08fF
C204 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C205 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C206 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C207 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.18fF
C208 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C209 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C210 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C211 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C212 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.09fF
C213 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.03fF
C214 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C215 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C216 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C217 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# -0.00fF
C218 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C219 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.33fF
C220 sky130_fd_sc_hd__nand2_4_3/B Bd_b 0.03fF
C221 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.04fF
C222 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.04fF
C223 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C224 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.01fF
C225 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.15fF
C226 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.34fF
C227 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.03fF
C228 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C229 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C230 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# 0.00fF
C231 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C232 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C233 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.13fF
C234 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.15fF
C235 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C236 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C237 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C238 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.07fF
C239 sky130_fd_sc_hd__clkinv_4_4/w_82_21# sky130_fd_sc_hd__clkinv_4_4/Y -0.00fF
C240 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__nand2_4_1/B 0.02fF
C241 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C242 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C243 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.23fF
C244 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C245 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0.04fF
C246 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.04fF
C247 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.31fF
C248 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C249 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C250 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C251 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C252 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C253 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C254 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C255 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C256 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C257 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.05fF
C258 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C259 sky130_fd_sc_hd__nand2_4_0/Y Bd_b 0.00fF
C260 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.08fF
C261 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.00fF
C262 sky130_fd_sc_hd__nand2_4_3/A Bd_b 0.27fF
C263 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0.03fF
C264 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C265 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.07fF
C266 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C267 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.01fF
C268 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.00fF
C269 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C270 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C271 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C272 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C273 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.05fF
C274 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C275 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C276 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.02fF
C277 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C278 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C279 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C280 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.04fF
C281 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.04fF
C282 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.19fF
C283 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.13fF
C284 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.02fF
C285 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0.02fF
C286 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.02fF
C287 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.02fF
C288 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.19fF
C289 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# Bd_b 0.06fF
C290 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.10fF
C291 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.03fF
C292 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.05fF
C293 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.10fF
C294 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.16fF
C295 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.74fF
C296 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_1_0/B 0.00fF
C297 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C298 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.08fF
C299 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.01fF
C300 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C301 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD 1.07fF
C302 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.08fF
C303 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C304 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C305 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C306 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C307 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.15fF
C308 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.04fF
C309 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C310 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.03fF
C311 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C312 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.20fF
C313 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.04fF
C314 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.04fF
C315 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C316 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.03fF
C317 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C318 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C319 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.02fF
C320 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C321 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__nand2_1_1/B 0.03fF
C322 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 1.16fF
C323 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_1/Y 0.33fF
C324 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A -0.00fF
C325 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C326 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C327 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C328 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.04fF
C329 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VDD 0.16fF
C330 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_1_3/Y 0.37fF
C331 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VDD 0.35fF
C332 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.08fF
C333 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C334 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.08fF
C335 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.19fF
C336 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C337 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C338 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C339 p2d_b sky130_fd_sc_hd__clkinv_4_9/Y 0.03fF
C340 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A sky130_fd_sc_hd__nand2_1_1/B 0.07fF
C341 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C342 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C343 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C344 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.01fF
C345 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C346 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C347 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C348 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C349 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C350 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C351 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C352 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C353 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.01fF
C354 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.02fF
C355 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.15fF
C356 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/A -0.81fF
C357 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.16fF
C358 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C359 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C360 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C361 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.07fF
C362 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VDD 0.13fF
C363 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.34fF
C364 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C365 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C366 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.08fF
C367 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C368 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C369 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.01fF
C370 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.00fF
C371 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A -0.00fF
C372 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 1.35fF
C373 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C374 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C375 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C376 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C377 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C378 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C379 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C380 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C381 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C382 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C383 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.03fF
C384 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.13fF
C385 VDD sky130_fd_sc_hd__dfxbp_1_1/a_27_47# 0.35fF
C386 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C387 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.14fF
C388 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X -0.00fF
C389 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.11fF
C390 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.03fF
C391 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.15fF
C392 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C393 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C394 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C395 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C396 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C397 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.09fF
C398 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C399 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# -0.00fF
C400 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C401 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.03fF
C402 B_b sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.06fF
C403 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C404 VDD Ad 1.64fF
C405 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C406 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C407 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.25fF
C408 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C409 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C410 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C411 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C412 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C413 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C414 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C415 sky130_fd_sc_hd__clkinv_4_10/w_82_21# sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C416 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C417 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_0/B 0.12fF
C418 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.19fF
C419 sky130_fd_sc_hd__mux2_1_0/a_505_21# Bd_b 0.04fF
C420 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.02fF
C421 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C422 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C423 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C424 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C425 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.03fF
C426 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.00fF
C427 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.15fF
C428 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.05fF
C429 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C430 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C431 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.02fF
C432 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C433 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C434 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C435 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C436 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C437 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C438 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.16fF
C439 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A -0.00fF
C440 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.15fF
C441 p1_b p1d 0.52fF
C442 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C443 sky130_fd_sc_hd__clkinv_4_9/Y Bd_b 0.00fF
C444 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_1_1/Y 0.12fF
C445 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.21fF
C446 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.03fF
C447 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C448 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C449 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C450 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C451 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C452 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.08fF
C453 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.73fF
C454 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C455 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C456 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.05fF
C457 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.03fF
C458 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C459 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C460 Ad_b Bd_b 4.81fF
C461 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A -0.00fF
C462 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VDD 0.33fF
C463 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C464 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C465 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C466 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.08fF
C467 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.00fF
C468 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 1.22fF
C469 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C470 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.03fF
C471 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.08fF
C472 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C473 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C474 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C475 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C476 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C477 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C478 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C479 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.02fF
C480 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C481 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C482 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C483 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C484 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C485 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# Ad_b 0.07fF
C486 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# Bd_b 0.05fF
C487 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C488 sky130_fd_sc_hd__nand2_1_1/B clk 0.00fF
C489 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A -0.00fF
C490 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.02fF
C491 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C492 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.08fF
C493 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.04fF
C494 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C495 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C496 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C497 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C498 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C499 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.02fF
C500 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.18fF
C501 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__mux2_1_0/X 0.05fF
C502 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.15fF
C503 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.32fF
C504 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.03fF
C505 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.06fF
C506 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.07fF
C507 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C508 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C509 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C510 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.05fF
C511 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.02fF
C512 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C513 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.02fF
C514 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C515 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C516 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C517 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C518 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C519 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C520 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.06fF
C521 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C522 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C523 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C524 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VDD 0.23fF
C525 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.08fF
C526 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.04fF
C527 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.22fF
C528 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/A 0.73fF
C529 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.01fF
C530 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C531 VDD sky130_fd_sc_hd__clkinv_4_4/Y 0.57fF
C532 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C533 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C534 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# A 0.06fF
C535 Ad sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.06fF
C536 Bd_b sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C537 p2 sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C538 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.02fF
C539 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.00fF
C540 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C541 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.02fF
C542 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.15fF
C543 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.05fF
C544 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.05fF
C545 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C546 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.05fF
C547 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C548 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C549 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C550 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C551 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C552 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C553 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C554 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C555 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.09fF
C556 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C557 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C558 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X -0.00fF
C559 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C560 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_2/A 0.05fF
C561 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C562 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C563 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C564 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Bd_b 0.14fF
C565 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C566 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C567 sky130_fd_sc_hd__clkinv_4_5/Y Ad_b 0.31fF
C568 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__mux2_1_0/X 0.05fF
C569 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C570 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.08fF
C571 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.31fF
C572 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C573 sky130_fd_sc_hd__nand2_4_1/B Bd_b 0.07fF
C574 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.01fF
C575 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.02fF
C576 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C577 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.00fF
C578 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.08fF
C579 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C580 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.89fF
C581 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C582 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/Y 0.73fF
C583 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C584 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.00fF
C585 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C586 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C587 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.04fF
C588 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C589 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C590 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C591 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.14fF
C592 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C593 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.02fF
C594 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C595 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C596 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C597 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C598 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.01fF
C599 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.13fF
C600 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.07fF
C601 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.04fF
C602 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.02fF
C603 VDD sky130_fd_sc_hd__clkinv_4_3/Y 1.73fF
C604 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.03fF
C605 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.02fF
C606 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_1_2/A 0.00fF
C607 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C608 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.15fF
C609 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C610 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.18fF
C611 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C612 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C613 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_592_47# 0.00fF
C614 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X -0.00fF
C615 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C616 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C617 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C618 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.04fF
C619 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C620 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C621 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.08fF
C622 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A -0.00fF
C623 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C624 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C625 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A -0.00fF
C626 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.11fF
C627 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 1.22fF
C628 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C629 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.01fF
C630 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkinv_4_7/Y 0.14fF
C631 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C632 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.02fF
C633 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.33fF
C634 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# Ad_b 0.16fF
C635 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.09fF
C636 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C637 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X -0.00fF
C638 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VDD 0.77fF
C639 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Ad_b 0.12fF
C640 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.14fF
C641 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C642 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C643 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C644 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C645 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C646 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_4_9/Y 0.14fF
C647 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 1.33fF
C648 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.22fF
C649 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.11fF
C650 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/D 0.10fF
C651 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.03fF
C652 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C653 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.02fF
C654 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C655 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.03fF
C656 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.03fF
C657 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C658 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C659 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C660 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.06fF
C661 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C662 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C663 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# 0.01fF
C664 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C665 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C666 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.32fF
C667 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C668 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_1_3/A 0.12fF
C669 VDD B_b 0.77fF
C670 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.00fF
C671 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.05fF
C672 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/A -0.69fF
C673 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X -0.00fF
C674 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.04fF
C675 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.01fF
C676 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.03fF
C677 sky130_fd_sc_hd__nand2_1_4/a_113_47# sky130_fd_sc_hd__nand2_1_4/Y -0.01fF
C678 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__nand2_1_1/A 0.03fF
C679 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__nand2_4_0/A 0.77fF
C680 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C681 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.15fF
C682 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.15fF
C683 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.02fF
C684 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/X -0.10fF
C685 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.02fF
C686 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C687 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C688 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C689 VSUBS sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C690 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C691 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C692 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C693 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C694 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# -0.00fF
C695 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.15fF
C696 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_4_1/B 0.11fF
C697 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.01fF
C698 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C699 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C700 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.07fF
C701 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.30fF
C702 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C703 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C704 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.05fF
C705 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.05fF
C706 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C707 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C708 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C709 VDD sky130_fd_sc_hd__nand2_1_1/A 13.45fF
C710 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.07fF
C711 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C712 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C713 p2_b VDD 0.77fF
C714 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C715 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_1_1/B 0.95fF
C716 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C717 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C718 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C719 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.08fF
C720 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.08fF
C721 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C722 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C723 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.17fF
C724 sky130_fd_sc_hd__clkinv_4_6/w_82_21# sky130_fd_sc_hd__nand2_4_2/A -0.30fF
C725 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.00fF
C726 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# 0.05fF
C727 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.01fF
C728 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.01fF
C729 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0.01fF
C730 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.01fF
C731 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C732 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.18fF
C733 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C734 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C735 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.07fF
C736 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C737 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.03fF
C738 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C739 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C740 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C741 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.30fF
C742 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C743 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C744 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C745 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C746 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.02fF
C747 Ad A_b 0.53fF
C748 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C749 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C750 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.14fF
C751 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.03fF
C752 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C753 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C754 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C755 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.02fF
C756 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.10fF
C757 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.07fF
C758 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C759 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.00fF
C760 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 1.14fF
C761 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/A 0.45fF
C762 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C763 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C764 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.09fF
C765 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C766 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A -0.00fF
C767 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C768 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C769 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C770 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C771 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C772 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C773 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.04fF
C774 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C775 p2 sky130_fd_sc_hd__nand2_4_3/B 0.06fF
C776 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_4/B 0.40fF
C777 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C778 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X -0.00fF
C779 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C780 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.05fF
C781 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.05fF
C782 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C783 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C784 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C785 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C786 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.02fF
C787 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.10fF
C788 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# 0.00fF
C789 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 6.53fF
C790 sky130_fd_sc_hd__clkinv_4_1/A B 0.00fF
C791 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.01fF
C792 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.03fF
C793 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.13fF
C794 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C795 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.16fF
C796 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C797 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.23fF
C798 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C799 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.01fF
C800 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C801 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.10fF
C802 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C803 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C804 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VDD -0.21fF
C805 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.18fF
C806 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C807 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.04fF
C808 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.09fF
C809 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C810 sky130_fd_sc_hd__nand2_4_1/Y Ad 0.00fF
C811 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.01fF
C812 p2 sky130_fd_sc_hd__nand2_4_3/A 0.34fF
C813 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C814 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.02fF
C815 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# 0.15fF
C816 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.02fF
C817 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.01fF
C818 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.01fF
C819 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.01fF
C820 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C821 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C822 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 1.13fF
C823 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.03fF
C824 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C825 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.07fF
C826 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C827 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C828 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.01fF
C829 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C830 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C831 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C832 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkinv_4_9/Y 0.08fF
C833 sky130_fd_sc_hd__clkinv_4_4/Y A_b 0.03fF
C834 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.05fF
C835 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VDD 0.16fF
C836 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C837 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.04fF
C838 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.04fF
C839 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.02fF
C840 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C841 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C842 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VDD 0.18fF
C843 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_1_4/B 0.07fF
C844 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# -0.08fF
C845 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.30fF
C846 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.05fF
C847 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.09fF
C848 p1d_b sky130_fd_sc_hd__clkbuf_16_11/a_110_47# 0.10fF
C849 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C850 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.02fF
C851 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C852 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VDD 1.14fF
C853 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.05fF
C854 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.05fF
C855 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C856 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.00fF
C857 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C858 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.02fF
C859 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.03fF
C860 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.09fF
C861 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.13fF
C862 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.16fF
C863 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VDD 0.10fF
C864 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__nand2_1_1/A 0.07fF
C865 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.17fF
C866 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C867 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C868 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.04fF
C869 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 2.24fF
C870 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C871 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.03fF
C872 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.02fF
C873 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C874 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C875 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C876 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C877 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C878 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.47fF
C879 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.01fF
C880 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C881 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.05fF
C882 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.01fF
C883 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1 -0.03fF
C884 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.05fF
C885 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.05fF
C886 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C887 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_47# -0.00fF
C888 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C889 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C890 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C891 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C892 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/A -0.21fF
C893 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.02fF
C894 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C895 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C896 VDD sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.21fF
C897 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.08fF
C898 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C899 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# -0.00fF
C900 p2d p2d_b 0.52fF
C901 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C902 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C903 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 3.21fF
C904 VDD sky130_fd_sc_hd__nand2_4_2/B 0.51fF
C905 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_1/A 0.47fF
C906 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.08fF
C907 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C908 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.05fF
C909 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C910 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.02fF
C911 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.10fF
C912 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C913 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.10fF
C914 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.04fF
C915 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.04fF
C916 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A -0.00fF
C917 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.03fF
C918 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.12fF
C919 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.18fF
C920 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.03fF
C921 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C922 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C923 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.13fF
C924 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C925 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.19fF
C926 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C927 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.00fF
C928 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.01fF
C929 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X -0.00fF
C930 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.30fF
C931 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C932 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C933 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.02fF
C934 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.03fF
C935 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.01fF
C936 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_4_1/A 1.35fF
C937 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C938 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C939 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C940 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C941 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.00fF
C942 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C943 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C944 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.16fF
C945 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C946 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C947 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C948 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C949 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C950 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.03fF
C951 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0.12fF
C952 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.01fF
C953 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.03fF
C954 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.15fF
C955 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C956 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C957 VDD sky130_fd_sc_hd__clkinv_1_1/Y 0.41fF
C958 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C959 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.01fF
C960 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.02fF
C961 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C962 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C963 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C964 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C965 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clk 0.05fF
C966 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C967 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.31fF
C968 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.21fF
C969 VDD sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.42fF
C970 sky130_fd_sc_hd__nand2_4_0/a_27_47# VDD 0.04fF
C971 sky130_fd_sc_hd__clkinv_4_8/w_82_21# sky130_fd_sc_hd__clkinv_4_8/Y -0.00fF
C972 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C973 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C974 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C975 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C976 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.01fF
C977 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.02fF
C978 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.01fF
C979 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C980 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C981 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 1.12fF
C982 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.06fF
C983 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.02fF
C984 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C985 A Ad_b 0.26fF
C986 p2_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.12fF
C987 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C988 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C989 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C990 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 1.27fF
C991 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C992 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.08fF
C993 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.08fF
C994 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.02fF
C995 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.00fF
C996 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.00fF
C997 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C998 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C999 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C1000 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C1001 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C1002 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C1003 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# Bd_b 0.06fF
C1004 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_1/A 0.08fF
C1005 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.03fF
C1006 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C1007 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C1008 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1009 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.95fF
C1010 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.05fF
C1011 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C1012 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.01fF
C1013 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C1014 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/B 0.11fF
C1015 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C1016 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.15fF
C1017 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C1018 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C1019 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.04fF
C1020 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.04fF
C1021 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_1/A 0.10fF
C1022 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.17fF
C1023 VDD sky130_fd_sc_hd__mux2_1_0/X 0.62fF
C1024 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.67fF
C1025 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.02fF
C1026 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.01fF
C1027 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C1028 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.02fF
C1029 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C1030 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.03fF
C1031 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.06fF
C1032 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__nand2_4_0/A 0.49fF
C1033 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.33fF
C1034 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C1035 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C1036 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C1037 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C1038 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C1039 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C1040 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C1041 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C1042 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C1043 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C1044 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C1045 p2 sky130_fd_sc_hd__clkinv_4_9/Y 0.04fF
C1046 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.05fF
C1047 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C1048 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.01fF
C1049 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.01fF
C1050 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C1051 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.09fF
C1052 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.05fF
C1053 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.31fF
C1054 p2 Ad_b 1.13fF
C1055 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# 0.84fF
C1056 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.30fF
C1057 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C1058 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.02fF
C1059 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.18fF
C1060 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.15fF
C1061 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__dfxbp_1_0/a_592_47# -0.00fF
C1062 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.33fF
C1063 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.04fF
C1064 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C1065 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_3/A 0.25fF
C1066 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.12fF
C1067 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C1068 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C1069 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD -0.70fF
C1070 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.02fF
C1071 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C1072 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.01fF
C1073 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkinv_4_3/Y -0.00fF
C1074 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C1075 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C1076 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C1077 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# p2 0.02fF
C1078 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C1079 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C1080 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C1081 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C1082 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C1083 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C1084 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C1085 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.04fF
C1086 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C1087 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Ad_b 0.07fF
C1088 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C1089 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C1090 sky130_fd_sc_hd__clkinv_4_5/Y Bd_b 0.46fF
C1091 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# A 0.02fF
C1092 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.05fF
C1093 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C1094 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.06fF
C1095 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C1096 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.01fF
C1097 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C1098 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C1099 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C1100 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C1101 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# 0.46fF
C1102 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.02fF
C1103 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.44fF
C1104 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.02fF
C1105 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.01fF
C1106 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X Bd_b 0.00fF
C1107 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C1108 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C1109 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C1110 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VDD 0.36fF
C1111 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C1112 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1113 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A -0.00fF
C1114 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C1115 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.01fF
C1116 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C1117 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C1118 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C1119 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.04fF
C1120 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C1121 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C1122 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C1123 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C1124 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.08fF
C1125 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.07fF
C1126 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C1127 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C1128 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C1129 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkinv_4_1/A 0.12fF
C1130 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/a_975_413# 0.00fF
C1131 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C1132 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.09fF
C1133 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.19fF
C1134 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C1135 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C1136 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C1137 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.07fF
C1138 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C1139 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C1140 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C1141 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C1142 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C1143 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.01fF
C1144 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.02fF
C1145 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.01fF
C1146 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.04fF
C1147 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C1148 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.13fF
C1149 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C1150 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C1151 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C1152 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.11fF
C1153 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.17fF
C1154 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# Bd_b 0.10fF
C1155 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C1156 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.35fF
C1157 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C1158 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C1159 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.00fF
C1160 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.22fF
C1161 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C1162 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# 0.09fF
C1163 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A Bd_b 0.14fF
C1164 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.01fF
C1165 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C1166 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C1167 VDD sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.11fF
C1168 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C1169 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C1170 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.09fF
C1171 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C1172 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/D 0.08fF
C1173 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C1174 p2 sky130_fd_sc_hd__nand2_4_1/B 0.04fF
C1175 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A -0.00fF
C1176 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.19fF
C1177 sky130_fd_sc_hd__clkinv_4_5/w_82_21# sky130_fd_sc_hd__nand2_4_1/A -0.30fF
C1178 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C1179 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C1180 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C1181 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.05fF
C1182 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C1183 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.03fF
C1184 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C1185 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.04fF
C1186 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.04fF
C1187 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.02fF
C1188 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C1189 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C1190 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C1191 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 1.21fF
C1192 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__clkinv_1_1/Y 0.73fF
C1193 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C1194 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.17fF
C1195 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.04fF
C1196 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.04fF
C1197 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C1198 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.11fF
C1199 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C1200 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.23fF
C1201 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.02fF
C1202 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C1203 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# 0.01fF
C1204 VSUBS sky130_fd_sc_hd__nand2_1_0/B 0.00fF
C1205 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.03fF
C1206 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C1207 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.02fF
C1208 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 1.18fF
C1209 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VDD 0.10fF
C1210 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.01fF
C1211 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.15fF
C1212 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.02fF
C1213 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.01fF
C1214 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.05fF
C1215 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C1216 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C1217 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C1218 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.00fF
C1219 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.15fF
C1220 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C1221 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.02fF
C1222 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.02fF
C1223 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.08fF
C1224 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C1225 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.03fF
C1226 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.17fF
C1227 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C1228 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.02fF
C1229 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C1230 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C1231 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C1232 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.03fF
C1233 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C1234 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.00fF
C1235 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C1236 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C1237 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C1238 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C1239 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C1240 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.33fF
C1241 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C1242 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C1243 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C1244 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C1245 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C1246 VSUBS sky130_fd_sc_hd__clkinv_4_1/Y 0.01fF
C1247 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.05fF
C1248 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C1249 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C1250 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.05fF
C1251 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.01fF
C1252 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C1253 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C1254 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0.02fF
C1255 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.02fF
C1256 p2d_b sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.14fF
C1257 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.15fF
C1258 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C1259 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C1260 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.03fF
C1261 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C1262 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C1263 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.11fF
C1264 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C1265 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C1266 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C1267 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.04fF
C1268 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C1269 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C1270 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 1.22fF
C1271 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C1272 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C1273 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C1274 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C1275 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C1276 sky130_fd_sc_hd__nand2_1_1/A clk 0.06fF
C1277 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.45fF
C1278 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C1279 sky130_fd_sc_hd__nand2_1_4/B Ad_b 0.02fF
C1280 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.14fF
C1281 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C1282 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C1283 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.18fF
C1284 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C1285 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C1286 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2d_b 0.12fF
C1287 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.03fF
C1288 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C1289 sky130_fd_sc_hd__nand2_4_2/Y p1d 0.00fF
C1290 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C1291 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.01fF
C1292 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C1293 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C1294 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_1/A 0.18fF
C1295 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C1296 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C1297 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C1298 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.01fF
C1299 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C1300 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C1301 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C1302 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C1303 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.32fF
C1304 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.14fF
C1305 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C1306 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# -0.00fF
C1307 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C1308 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.04fF
C1309 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C1310 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.03fF
C1311 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C1312 sky130_fd_sc_hd__clkinv_4_7/A VDD 4.01fF
C1313 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.04fF
C1314 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.04fF
C1315 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.11fF
C1316 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C1317 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C1318 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C1319 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.19fF
C1320 p1 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.12fF
C1321 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1_b 0.12fF
C1322 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.08fF
C1323 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.02fF
C1324 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.35fF
C1325 VDD sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.30fF
C1326 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C1327 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.02fF
C1328 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.02fF
C1329 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.11fF
C1330 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C1331 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_1_4/Y -0.43fF
C1332 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C1333 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C1334 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.15fF
C1335 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C1336 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.04fF
C1337 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.04fF
C1338 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C1339 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C1340 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.07fF
C1341 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C1342 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C1343 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C1344 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.00fF
C1345 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.03fF
C1346 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.45fF
C1347 p2d sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.02fF
C1348 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.09fF
C1349 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.00fF
C1350 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.00fF
C1351 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C1352 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C1353 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C1354 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C1355 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C1356 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C1357 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VDD 0.16fF
C1358 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.10fF
C1359 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.16fF
C1360 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.01fF
C1361 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# 0.09fF
C1362 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.03fF
C1363 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.10fF
C1364 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.23fF
C1365 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C1366 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.01fF
C1367 p1d_b sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.12fF
C1368 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C1369 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.02fF
C1370 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C1371 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.02fF
C1372 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C1373 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C1374 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C1375 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C1376 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.11fF
C1377 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C1378 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C1379 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VDD 0.06fF
C1380 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.15fF
C1381 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.03fF
C1382 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C1383 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C1384 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.31fF
C1385 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.02fF
C1386 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C1387 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.08fF
C1388 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C1389 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C1390 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.02fF
C1391 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# -0.00fF
C1392 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.01fF
C1393 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.05fF
C1394 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2d 0.12fF
C1395 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C1396 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C1397 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C1398 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C1399 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.11fF
C1400 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C1401 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.07fF
C1402 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C1403 VDD sky130_fd_sc_hd__dfxbp_1_1/a_634_159# -0.06fF
C1404 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C1405 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C1406 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C1407 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_0/w_82_21# 0.05fF
C1408 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.05fF
C1409 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.05fF
C1410 sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.05fF
C1411 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C1412 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C1413 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C1414 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.08fF
C1415 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C1416 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C1417 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C1418 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C1419 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.05fF
C1420 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.02fF
C1421 VSUBS sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C1422 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C1423 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C1424 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.13fF
C1425 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.02fF
C1426 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C1427 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.01fF
C1428 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C1429 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.02fF
C1430 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.14fF
C1431 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0.06fF
C1432 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C1433 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.14fF
C1434 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.12fF
C1435 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.01fF
C1436 p1d_b VDD 0.80fF
C1437 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C1438 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C1439 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C1440 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C1441 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C1442 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.16fF
C1443 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C1444 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C1445 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C1446 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.05fF
C1447 VDD sky130_fd_sc_hd__nand2_4_1/A 11.01fF
C1448 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C1449 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C1450 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C1451 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C1452 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C1453 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C1454 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C1455 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C1456 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C1457 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C1458 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.00fF
C1459 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.02fF
C1460 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.04fF
C1461 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.04fF
C1462 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.06fF
C1463 p2 p2d_b 0.09fF
C1464 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.04fF
C1465 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.04fF
C1466 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C1467 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C1468 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C1469 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clk 0.01fF
C1470 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C1471 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C1472 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.18fF
C1473 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.14fF
C1474 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C1475 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C1476 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.02fF
C1477 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C1478 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C1479 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C1480 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C1481 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C1482 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.02fF
C1483 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C1484 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C1485 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VDD 0.22fF
C1486 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.04fF
C1487 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.03fF
C1488 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C1489 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.03fF
C1490 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.09fF
C1491 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0.00fF
C1492 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.02fF
C1493 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.31fF
C1494 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.04fF
C1495 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1496 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C1497 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# -0.08fF
C1498 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.01fF
C1499 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.02fF
C1500 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0.08fF
C1501 VSUBS sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C1502 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C1503 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C1504 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C1505 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C1506 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.11fF
C1507 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C1508 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.02fF
C1509 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C1510 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C1511 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD -0.63fF
C1512 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.04fF
C1513 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.09fF
C1514 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C1515 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1516 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_0/A 0.21fF
C1517 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.00fF
C1518 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C1519 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.02fF
C1520 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C1521 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.04fF
C1522 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.04fF
C1523 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 1.21fF
C1524 p2_b sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.12fF
C1525 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C1526 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C1527 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C1528 sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C1529 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# Bd 0.02fF
C1530 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C1531 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.01fF
C1532 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C1533 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.01fF
C1534 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# Bd 0.06fF
C1535 B sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.06fF
C1536 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.14fF
C1537 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/B 0.02fF
C1538 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# B 0.02fF
C1539 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.03fF
C1540 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0.01fF
C1541 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.05fF
C1542 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C1543 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.17fF
C1544 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C1545 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C1546 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C1547 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C1548 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C1549 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C1550 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C1551 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C1552 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C1553 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.10fF
C1554 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 3.20fF
C1555 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C1556 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.04fF
C1557 VDD A_b 0.82fF
C1558 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VDD 0.35fF
C1559 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.01fF
C1560 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.15fF
C1561 p2 Bd_b 0.56fF
C1562 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.00fF
C1563 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# 0.15fF
C1564 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.18fF
C1565 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C1566 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.25fF
C1567 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.01fF
C1568 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.34fF
C1569 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C1570 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__dfxbp_1_0/a_975_413# 0.01fF
C1571 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.19fF
C1572 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.04fF
C1573 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.04fF
C1574 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C1575 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.31fF
C1576 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C1577 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C1578 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.16fF
C1579 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.04fF
C1580 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1581 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.07fF
C1582 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.35fF
C1583 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C1584 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.12fF
C1585 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.05fF
C1586 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.11fF
C1587 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.12fF
C1588 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.01fF
C1589 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C1590 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# p2 0.02fF
C1591 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C1592 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C1593 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C1594 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C1595 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.04fF
C1596 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_1_4/B 0.11fF
C1597 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C1598 p2d p2 0.20fF
C1599 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.26fF
C1600 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C1601 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_1/Y 0.20fF
C1602 VSUBS sky130_fd_sc_hd__nand2_4_3/Y -0.26fF
C1603 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C1604 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C1605 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C1606 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C1607 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C1608 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.04fF
C1609 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.04fF
C1610 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.04fF
C1611 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X Bd_b 0.07fF
C1612 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.03fF
C1613 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C1614 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C1615 sky130_fd_sc_hd__clkinv_4_5/Y A 0.00fF
C1616 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.03fF
C1617 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.15fF
C1618 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.63fF
C1619 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C1620 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C1621 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.05fF
C1622 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0.18fF
C1623 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C1624 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C1625 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C1626 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C1627 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.19fF
C1628 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VDD 0.20fF
C1629 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.23fF
C1630 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.01fF
C1631 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C1632 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C1633 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C1634 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# sky130_fd_sc_hd__nand2_1_4/B 0.02fF
C1635 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.41fF
C1636 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_3/A 0.21fF
C1637 sky130_fd_sc_hd__nand2_4_1/Y VDD 6.27fF
C1638 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.04fF
C1639 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C1640 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.04fF
C1641 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.04fF
C1642 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.04fF
C1643 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C1644 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C1645 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C1646 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.04fF
C1647 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C1648 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# sky130_fd_sc_hd__clkinv_4_1/Y 0.08fF
C1649 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.03fF
C1650 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C1651 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.00fF
C1652 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C1653 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 2.24fF
C1654 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.09fF
C1655 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/X -0.16fF
C1656 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C1657 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C1658 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C1659 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C1660 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C1661 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.03fF
C1662 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C1663 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C1664 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.07fF
C1665 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C1666 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C1667 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.84fF
C1668 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.02fF
C1669 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C1670 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C1671 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.14fF
C1672 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.04fF
C1673 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# A 0.12fF
C1674 A_b sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.12fF
C1675 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.09fF
C1676 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.02fF
C1677 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.30fF
C1678 p2 sky130_fd_sc_hd__clkinv_4_5/Y 0.16fF
C1679 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.04fF
C1680 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C1681 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C1682 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C1683 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C1684 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C1685 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.10fF
C1686 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# sky130_fd_sc_hd__dfxbp_1_1/D 0.07fF
C1687 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C1688 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.01fF
C1689 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.06fF
C1690 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.04fF
C1691 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# 0.12fF
C1692 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C1693 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/A -0.24fF
C1694 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.34fF
C1695 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C1696 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C1697 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C1698 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C1699 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.08fF
C1700 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C1701 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.14fF
C1702 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C1703 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X -0.00fF
C1704 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_4_3/A 0.73fF
C1705 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_3/A 0.02fF
C1706 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C1707 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C1708 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C1709 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.08fF
C1710 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.12fF
C1711 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C1712 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0.01fF
C1713 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C1714 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.02fF
C1715 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 2.25fF
C1716 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.00fF
C1717 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C1718 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.01fF
C1719 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.10fF
C1720 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C1721 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C1722 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.01fF
C1723 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.03fF
C1724 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.03fF
C1725 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.15fF
C1726 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C1727 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.02fF
C1728 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.02fF
C1729 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C1730 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C1731 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C1732 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.15fF
C1733 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C1734 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C1735 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.09fF
C1736 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.03fF
C1737 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C1738 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.55fF
C1739 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.31fF
C1740 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.31fF
C1741 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C1742 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.03fF
C1743 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.11fF
C1744 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# p1_b 0.10fF
C1745 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VDD 0.35fF
C1746 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.14fF
C1747 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C1748 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.10fF
C1749 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C1750 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/A -0.75fF
C1751 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C1752 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.02fF
C1753 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C1754 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C1755 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C1756 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C1757 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.02fF
C1758 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C1759 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.09fF
C1760 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.02fF
C1761 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C1762 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.11fF
C1763 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C1764 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.07fF
C1765 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C1766 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.05fF
C1767 VDD clk 1.78fF
C1768 sky130_fd_sc_hd__nand2_1_4/B Bd_b 0.02fF
C1769 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C1770 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C1771 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.12fF
C1772 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C1773 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.03fF
C1774 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X -0.00fF
C1775 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_1_0/A 0.06fF
C1776 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.02fF
C1777 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.02fF
C1778 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.01fF
C1779 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.01fF
C1780 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.33fF
C1781 sky130_fd_sc_hd__clkinv_1_3/A VDD 4.68fF
C1782 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C1783 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C1784 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C1785 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C1786 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C1787 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C1788 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C1789 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C1790 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C1791 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C1792 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.08fF
C1793 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.14fF
C1794 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.08fF
C1795 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C1796 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.30fF
C1797 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.05fF
C1798 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C1799 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C1800 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C1801 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C1802 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.08fF
C1803 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C1804 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C1805 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# -0.00fF
C1806 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.01fF
C1807 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C1808 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C1809 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C1810 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.44fF
C1811 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.05fF
C1812 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.00fF
C1813 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C1814 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.15fF
C1815 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C1816 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.02fF
C1817 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.01fF
C1818 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C1819 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 1.17fF
C1820 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C1821 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C1822 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/A 0.62fF
C1823 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C1824 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.00fF
C1825 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C1826 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C1827 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C1828 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_1_3/A 0.04fF
C1829 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.05fF
C1830 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/X -0.15fF
C1831 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C1832 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C1833 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.02fF
C1834 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.00fF
C1835 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C1836 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.02fF
C1837 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C1838 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.05fF
C1839 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C1840 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C1841 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C1842 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C1843 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.12fF
C1844 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.02fF
C1845 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.04fF
C1846 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.04fF
C1847 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.00fF
C1848 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.05fF
C1849 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.12fF
C1850 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.15fF
C1851 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.03fF
C1852 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C1853 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C1854 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C1855 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.02fF
C1856 sky130_fd_sc_hd__clkinv_4_1/A VDD 4.66fF
C1857 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.05fF
C1858 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C1859 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C1860 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C1861 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# 0.32fF
C1862 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.03fF
C1863 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.02fF
C1864 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__nand2_1_2/B 0.00fF
C1865 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C1866 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/B 0.16fF
C1867 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_4/B 0.14fF
C1868 sky130_fd_sc_hd__dfxbp_1_0/a_561_413# VDD 0.00fF
C1869 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.09fF
C1870 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C1871 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.18fF
C1872 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C1873 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C1874 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C1875 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C1876 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# 0.31fF
C1877 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C1878 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.02fF
C1879 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.30fF
C1880 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.62fF
C1881 p2 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.06fF
C1882 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C1883 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C1884 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C1885 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C1886 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C1887 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C1888 VDD sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.08fF
C1889 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# 0.06fF
C1890 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C1891 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C1892 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C1893 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C1894 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.03fF
C1895 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.03fF
C1896 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C1897 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.01fF
C1898 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.01fF
C1899 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C1900 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C1901 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C1902 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.03fF
C1903 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.00fF
C1904 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.08fF
C1905 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C1906 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 1.12fF
C1907 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C1908 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C1909 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C1910 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.15fF
C1911 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.02fF
C1912 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.02fF
C1913 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.02fF
C1914 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.02fF
C1915 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0.06fF
C1916 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C1917 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.00fF
C1918 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C1919 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_3/A 0.62fF
C1920 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.03fF
C1921 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C1922 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1923 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.00fF
C1924 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.10fF
C1925 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C1926 sky130_fd_sc_hd__mux2_1_0/a_439_47# Ad_b 0.02fF
C1927 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.15fF
C1928 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.01fF
C1929 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C1930 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C1931 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.15fF
C1932 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2 0.02fF
C1933 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VDD 0.15fF
C1934 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C1935 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C1936 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C1937 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C1938 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C1939 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C1940 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.07fF
C1941 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C1942 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C1943 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C1944 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C1945 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C1946 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C1947 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.04fF
C1948 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C1949 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C1950 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C1951 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.07fF
C1952 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.06fF
C1953 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C1954 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C1955 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.02fF
C1956 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.05fF
C1957 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C1958 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C1959 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A -0.00fF
C1960 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.11fF
C1961 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.15fF
C1962 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# -0.00fF
C1963 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C1964 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C1965 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C1966 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.07fF
C1967 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C1968 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C1969 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.03fF
C1970 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.08fF
C1971 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.00fF
C1972 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C1973 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C1974 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.02fF
C1975 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C1976 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.01fF
C1977 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C1978 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.08fF
C1979 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.05fF
C1980 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.05fF
C1981 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.08fF
C1982 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.18fF
C1983 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.06fF
C1984 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.02fF
C1985 VDD sky130_fd_sc_hd__clkinv_4_7/Y 0.55fF
C1986 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.10fF
C1987 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C1988 sky130_fd_sc_hd__clkinv_4_1/w_82_21# sky130_fd_sc_hd__clkinv_4_1/Y 0.04fF
C1989 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C1990 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C1991 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1 0.02fF
C1992 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.01fF
C1993 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C1994 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# Ad_b 0.01fF
C1995 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C1996 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# -0.00fF
C1997 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 1.35fF
C1998 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.19fF
C1999 VDD sky130_fd_sc_hd__nand2_1_0/A 1.27fF
C2000 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 1.12fF
C2001 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C2002 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VDD 0.54fF
C2003 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.00fF
C2004 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.08fF
C2005 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C2006 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.01fF
C2007 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.01fF
C2008 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C2009 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C2010 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C2011 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C2012 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.55fF
C2013 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.02fF
C2014 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.02fF
C2015 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C2016 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C2017 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.03fF
C2018 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C2019 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.06fF
C2020 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.01fF
C2021 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.01fF
C2022 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.18fF
C2023 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.04fF
C2024 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VDD 0.39fF
C2025 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.15fF
C2026 sky130_fd_sc_hd__nand2_4_0/Y Bd 0.00fF
C2027 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 1.29fF
C2028 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.03fF
C2029 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C2030 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2031 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C2032 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C2033 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C2034 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C2035 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VDD 0.49fF
C2036 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C2037 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C2038 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.19fF
C2039 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.07fF
C2040 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C2041 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.04fF
C2042 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VDD 0.17fF
C2043 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VDD 0.11fF
C2044 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.15fF
C2045 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.03fF
C2046 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C2047 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C2048 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.12fF
C2049 p2 A 0.02fF
C2050 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C2051 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C2052 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.15fF
C2053 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.13fF
C2054 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.17fF
C2055 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C2056 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/B 0.07fF
C2057 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.15fF
C2058 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.02fF
C2059 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.37fF
C2060 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.14fF
C2061 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.03fF
C2062 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.25fF
C2063 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.62fF
C2064 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C2065 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C2066 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C2067 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.08fF
C2068 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C2069 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 6.27fF
C2070 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.17fF
C2071 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C2072 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C2073 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.02fF
C2074 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C2075 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C2076 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.04fF
C2077 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.04fF
C2078 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.30fF
C2079 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.07fF
C2080 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.01fF
C2081 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C2082 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C2083 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# B_b 0.15fF
C2084 Bd sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.15fF
C2085 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.02fF
C2086 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C2087 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# B_b 0.12fF
C2088 B sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.12fF
C2089 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C2090 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C2091 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/Y 0.32fF
C2092 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C2093 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C2094 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.03fF
C2095 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C2096 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.03fF
C2097 VSUBS sky130_fd_sc_hd__clkinv_4_4/Y 0.00fF
C2098 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.02fF
C2099 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C2100 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.06fF
C2101 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C2102 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C2103 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C2104 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C2105 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0.08fF
C2106 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.02fF
C2107 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C2108 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C2109 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C2110 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C2111 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C2112 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C2113 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.01fF
C2114 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.02fF
C2115 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.12fF
C2116 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# 0.13fF
C2117 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C2118 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.09fF
C2119 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VDD 0.15fF
C2120 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.12fF
C2121 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C2122 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.02fF
C2123 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Ad 0.05fF
C2124 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.97fF
C2125 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.40fF
C2126 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.00fF
C2127 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.00fF
C2128 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__nand2_1_4/B 0.10fF
C2129 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C2130 VDD sky130_fd_sc_hd__nand2_1_3/A 4.52fF
C2131 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C2132 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C2133 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C2134 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.02fF
C2135 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.00fF
C2136 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.00fF
C2137 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C2138 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__nand2_4_3/Y 0.66fF
C2139 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# 0.01fF
C2140 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.07fF
C2141 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.11fF
C2142 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.50fF
C2143 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.02fF
C2144 VDD sky130_fd_sc_hd__nand2_1_2/B 1.61fF
C2145 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.04fF
C2146 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.04fF
C2147 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C2148 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C2149 sky130_fd_sc_hd__nand2_4_3/Y Ad_b 0.00fF
C2150 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.10fF
C2151 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.45fF
C2152 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# 0.05fF
C2153 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.02fF
C2154 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.10fF
C2155 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.15fF
C2156 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.03fF
C2157 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C2158 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C2159 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.30fF
C2160 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.03fF
C2161 VSUBS sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C2162 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.03fF
C2163 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.07fF
C2164 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C2165 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C2166 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C2167 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.10fF
C2168 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_3/Y 0.01fF
C2169 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0.06fF
C2170 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.04fF
C2171 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.04fF
C2172 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.17fF
C2173 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C2174 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C2175 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.04fF
C2176 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.30fF
C2177 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C2178 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C2179 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C2180 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C2181 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.02fF
C2182 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C2183 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.02fF
C2184 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.10fF
C2185 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.07fF
C2186 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C2187 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/X -0.28fF
C2188 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/B 0.07fF
C2189 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C2190 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C2191 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.01fF
C2192 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.00fF
C2193 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.07fF
C2194 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C2195 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.10fF
C2196 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C2197 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C2198 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C2199 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.08fF
C2200 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C2201 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A -0.00fF
C2202 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C2203 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.16fF
C2204 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.05fF
C2205 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C2206 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.08fF
C2207 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C2208 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C2209 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C2210 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.18fF
C2211 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.05fF
C2212 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C2213 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 1.09fF
C2214 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.33fF
C2215 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_1_2/B 0.00fF
C2216 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0.01fF
C2217 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/A 0.46fF
C2218 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.03fF
C2219 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C2220 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C2221 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.01fF
C2222 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.07fF
C2223 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C2224 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C2225 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.00fF
C2226 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C2227 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C2228 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C2229 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.31fF
C2230 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.03fF
C2231 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C2232 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C2233 VSUBS sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C2234 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C2235 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C2236 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C2237 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.01fF
C2238 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C2239 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C2240 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_4_1/B 0.00fF
C2241 sky130_fd_sc_hd__nand2_4_3/a_27_47# VDD 0.05fF
C2242 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/X -0.72fF
C2243 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.06fF
C2244 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C2245 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.34fF
C2246 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C2247 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.18fF
C2248 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.04fF
C2249 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C2250 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C2251 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C2252 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.03fF
C2253 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.17fF
C2254 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.07fF
C2255 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.18fF
C2256 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C2257 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C2258 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C2259 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.04fF
C2260 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C2261 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C2262 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C2263 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.15fF
C2264 sky130_fd_sc_hd__clkinv_4_8/Y sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2265 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.04fF
C2266 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.04fF
C2267 sky130_fd_sc_hd__nand2_4_0/B VDD 0.55fF
C2268 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.17fF
C2269 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C2270 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.08fF
C2271 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C2272 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.33fF
C2273 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C2274 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C2275 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.08fF
C2276 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X -0.00fF
C2277 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.02fF
C2278 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.02fF
C2279 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.00fF
C2280 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.06fF
C2281 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A -0.00fF
C2282 sky130_fd_sc_hd__clkinv_4_9/w_82_21# sky130_fd_sc_hd__nand2_4_3/Y 0.03fF
C2283 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C2284 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C2285 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C2286 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.04fF
C2287 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.01fF
C2288 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.03fF
C2289 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C2290 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C2291 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C2292 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C2293 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C2294 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.00fF
C2295 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C2296 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A -0.00fF
C2297 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C2298 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C2299 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C2300 sky130_fd_sc_hd__clkinv_1_3/A clk 0.00fF
C2301 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_3/A 0.13fF
C2302 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.31fF
C2303 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C2304 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C2305 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.01fF
C2306 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.00fF
C2307 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C2308 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/A -0.61fF
C2309 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.01fF
C2310 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.01fF
C2311 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.02fF
C2312 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.05fF
C2313 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.04fF
C2314 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.04fF
C2315 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# 0.09fF
C2316 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C2317 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C2318 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.07fF
C2319 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.03fF
C2320 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.10fF
C2321 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C2322 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.09fF
C2323 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.07fF
C2324 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.06fF
C2325 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.05fF
C2326 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C2327 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 2.24fF
C2328 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.00fF
C2329 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.00fF
C2330 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C2331 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0.05fF
C2332 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.10fF
C2333 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.10fF
C2334 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C2335 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.10fF
C2336 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C2337 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.08fF
C2338 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.02fF
C2339 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# 0.17fF
C2340 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C2341 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_1_2/B 0.03fF
C2342 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.11fF
C2343 sky130_fd_sc_hd__dfxbp_1_0/a_975_413# VDD 0.00fF
C2344 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.08fF
C2345 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C2346 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C2347 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.15fF
C2348 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.01fF
C2349 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C2350 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C2351 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.04fF
C2352 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.04fF
C2353 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.08fF
C2354 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.02fF
C2355 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.19fF
C2356 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A -0.00fF
C2357 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.14fF
C2358 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.01fF
C2359 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C2360 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.00fF
C2361 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C2362 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C2363 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__mux2_1_0/S 0.08fF
C2364 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C2365 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C2366 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.05fF
C2367 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.09fF
C2368 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C2369 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C2370 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.02fF
C2371 VDD sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# 0.19fF
C2372 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.07fF
C2373 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C2374 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C2375 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.02fF
C2376 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.02fF
C2377 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1_b 0.06fF
C2378 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.01fF
C2379 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.03fF
C2380 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.98fF
C2381 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C2382 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.08fF
C2383 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0.12fF
C2384 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C2385 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.10fF
C2386 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.00fF
C2387 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C2388 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Ad_b 0.05fF
C2389 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.05fF
C2390 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.04fF
C2391 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.04fF
C2392 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C2393 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__nand2_4_0/A 0.16fF
C2394 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C2395 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.01fF
C2396 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C2397 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.03fF
C2398 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C2399 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C2400 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C2401 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C2402 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/A -0.61fF
C2403 sky130_fd_sc_hd__mux2_1_0/a_439_47# Bd_b 0.00fF
C2404 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.00fF
C2405 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C2406 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C2407 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.04fF
C2408 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C2409 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.02fF
C2410 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.04fF
C2411 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.04fF
C2412 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C2413 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C2414 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C2415 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C2416 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 1.11fF
C2417 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C2418 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C2419 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C2420 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.00fF
C2421 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C2422 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C2423 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.03fF
C2424 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Ad_b 0.05fF
C2425 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.07fF
C2426 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.02fF
C2427 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.02fF
C2428 VSUBS sky130_fd_sc_hd__nand2_4_2/B -0.05fF
C2429 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C2430 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.01fF
C2431 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C2432 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C2433 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.12fF
C2434 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.01fF
C2435 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.00fF
C2436 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VDD 0.51fF
C2437 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C2438 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.01fF
C2439 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C2440 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C2441 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C2442 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.02fF
C2443 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C2444 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C2445 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.01fF
C2446 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# 0.07fF
C2447 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C2448 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.65fF
C2449 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.15fF
C2450 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.14fF
C2451 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C2452 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0.04fF
C2453 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.04fF
C2454 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# 0.33fF
C2455 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.10fF
C2456 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.07fF
C2457 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.04fF
C2458 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.04fF
C2459 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# Ad_b 0.00fF
C2460 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/S 0.06fF
C2461 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# Bd_b 0.01fF
C2462 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.36fF
C2463 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C2464 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.09fF
C2465 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.01fF
C2466 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# p1d 0.06fF
C2467 p1 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.06fF
C2468 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0.05fF
C2469 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.04fF
C2470 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSUBS -0.05fF
C2471 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 1.12fF
C2472 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C2473 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C2474 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.07fF
C2475 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C2476 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.02fF
C2477 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.10fF
C2478 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C2479 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C2480 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C2481 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.03fF
C2482 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.05fF
C2483 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.05fF
C2484 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C2485 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.05fF
C2486 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 1.38fF
C2487 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C2488 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C2489 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0.06fF
C2490 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.12fF
C2491 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.01fF
C2492 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.03fF
C2493 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.05fF
C2494 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.05fF
C2495 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.10fF
C2496 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C2497 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.03fF
C2498 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.01fF
C2499 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.04fF
C2500 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C2501 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C2502 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.01fF
C2503 sky130_fd_sc_hd__nand2_4_2/a_27_47# VDD 0.04fF
C2504 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C2505 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.05fF
C2506 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.02fF
C2507 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# 0.08fF
C2508 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.08fF
C2509 Ad Ad_b 0.60fF
C2510 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VDD 0.16fF
C2511 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C2512 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C2513 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C2514 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.31fF
C2515 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_0/B 0.03fF
C2516 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C2517 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.12fF
C2518 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.08fF
C2519 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C2520 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.15fF
C2521 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# sky130_fd_sc_hd__dfxbp_1_0/a_1017_47# -0.00fF
C2522 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C2523 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.00fF
C2524 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2525 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.22fF
C2526 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.13fF
C2527 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C2528 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C2529 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/X 0.01fF
C2530 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C2531 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C2532 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C2533 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.00fF
C2534 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.15fF
C2535 VSUBS sky130_fd_sc_hd__mux2_1_0/X -0.01fF
C2536 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.19fF
C2537 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C2538 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.05fF
C2539 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C2540 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.01fF
C2541 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.01fF
C2542 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.01fF
C2543 VDD p1 1.45fF
C2544 sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C2545 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.11fF
C2546 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.00fF
C2547 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.00fF
C2548 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.08fF
C2549 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.08fF
C2550 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C2551 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.01fF
C2552 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# p2 0.00fF
C2553 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C2554 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# sky130_fd_sc_hd__clkinv_1_3/A 0.02fF
C2555 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.01fF
C2556 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.04fF
C2557 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.00fF
C2558 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.01fF
C2559 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C2560 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.01fF
C2561 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C2562 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.04fF
C2563 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.02fF
C2564 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.02fF
C2565 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C2566 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C2567 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C2568 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C2569 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C2570 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.14fF
C2571 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.04fF
C2572 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.04fF
C2573 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.03fF
C2574 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C2575 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.01fF
C2576 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.01fF
C2577 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.01fF
C2578 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C2579 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C2580 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C2581 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C2582 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C2583 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.00fF
C2584 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 3.21fF
C2585 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C2586 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.03fF
C2587 VDD sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.37fF
C2588 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C2589 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C2590 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C2591 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C2592 VDD sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0.54fF
C2593 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.03fF
C2594 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.10fF
C2595 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C2596 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C2597 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C2598 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.24fF
C2599 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C2600 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# sky130_fd_sc_hd__nand2_1_4/B 0.13fF
C2601 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C2602 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A -0.00fF
C2603 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.30fF
C2604 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.02fF
C2605 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C2606 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_4_3/A 0.30fF
C2607 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.04fF
C2608 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C2609 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C2610 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C2611 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.02fF
C2612 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.02fF
C2613 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.01fF
C2614 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.00fF
C2615 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.01fF
C2616 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C2617 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C2618 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C2619 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# B_b 0.12fF
C2620 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C2621 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C2622 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.08fF
C2623 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.05fF
C2624 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_3/Y 0.03fF
C2625 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.02fF
C2626 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.01fF
C2627 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.03fF
C2628 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C2629 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.01fF
C2630 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C2631 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C2632 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.01fF
C2633 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.08fF
C2634 VDD sky130_fd_sc_hd__nand2_1_2/A -0.72fF
C2635 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C2636 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.01fF
C2637 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C2638 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C2639 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C2640 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C2641 sky130_fd_sc_hd__nand2_4_3/Y Bd_b 0.00fF
C2642 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C2643 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C2644 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C2645 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C2646 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.00fF
C2647 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.09fF
C2648 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C2649 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# Ad 0.12fF
C2650 sky130_fd_sc_hd__clkinv_4_7/A p1 0.00fF
C2651 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.07fF
C2652 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.15fF
C2653 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C2654 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkinv_1_1/Y 0.12fF
C2655 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.04fF
C2656 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_1_0/A 0.01fF
C2657 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C2658 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.15fF
C2659 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.04fF
C2660 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C2661 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C2662 sky130_fd_sc_hd__nand2_1_3/A clk 0.02fF
C2663 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.08fF
C2664 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C2665 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C2666 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C2667 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/a_27_47# 0.00fF
C2668 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C2669 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_3/Y 0.01fF
C2670 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__mux2_1_0/S 0.02fF
C2671 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C2672 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0.05fF
C2673 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.01fF
C2674 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.01fF
C2675 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.01fF
C2676 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C2677 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.15fF
C2678 p2d sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C2679 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VDD 6.44fF
C2680 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.02fF
C2681 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_4_10/w_82_21# 0.04fF
C2682 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.16fF
C2683 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C2684 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C2685 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_3/A 0.16fF
C2686 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.31fF
C2687 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_4_3/A 2.16fF
C2688 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C2689 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 1.12fF
C2690 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.08fF
C2691 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C2692 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C2693 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C2694 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.04fF
C2695 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.04fF
C2696 sky130_fd_sc_hd__nand2_1_2/B clk 0.04fF
C2697 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C2698 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.00fF
C2699 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C2700 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C2701 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C2702 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C2703 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C2704 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.01fF
C2705 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0.06fF
C2706 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C2707 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C2708 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.03fF
C2709 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.08fF
C2710 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C2711 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.02fF
C2712 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C2713 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkinv_4_2/Y 0.08fF
C2714 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C2715 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C2716 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.00fF
C2717 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C2718 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C2719 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C2720 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C2721 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C2722 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C2723 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C2724 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C2725 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C2726 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.02fF
C2727 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.02fF
C2728 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C2729 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C2730 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.14fF
C2731 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.05fF
C2732 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C2733 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C2734 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.16fF
C2735 sky130_fd_sc_hd__clkinv_4_3/Y Ad_b 0.07fF
C2736 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.14fF
C2737 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C2738 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_1_2/A 0.01fF
C2739 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C2740 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X -0.00fF
C2741 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.07fF
C2742 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C2743 Bd Bd_b 0.47fF
C2744 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.04fF
C2745 B Bd_b 0.08fF
C2746 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.02fF
C2747 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.51fF
C2748 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.04fF
C2749 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C2750 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.00fF
C2751 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C2752 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C2753 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.03fF
C2754 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.10fF
C2755 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.04fF
C2756 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.02fF
C2757 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VDD 0.21fF
C2758 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.01fF
C2759 VDD sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.20fF
C2760 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.98fF
C2761 VSUBS VDD -5.81fF
C2762 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.18fF
C2763 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C2764 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.00fF
C2765 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C2766 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.26fF
C2767 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.03fF
C2768 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C2769 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 1.33fF
C2770 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.09fF
C2771 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.03fF
C2772 p1d_b p1 0.08fF
C2773 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C2774 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.19fF
C2775 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.01fF
C2776 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.17fF
C2777 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C2778 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C2779 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C2780 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.09fF
C2781 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C2782 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C2783 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.02fF
C2784 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VDD 0.40fF
C2785 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.14fF
C2786 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C2787 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C2788 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C2789 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_3/A 0.04fF
C2790 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.04fF
C2791 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.02fF
C2792 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C2793 VDD sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.16fF
C2794 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C2795 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C2796 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Ad_b 0.04fF
C2797 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__nand2_4_2/A 0.42fF
C2798 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.32fF
C2799 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.09fF
C2800 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# -0.00fF
C2801 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.08fF
C2802 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.01fF
C2803 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.01fF
C2804 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C2805 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.08fF
C2806 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.14fF
C2807 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.19fF
C2808 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.16fF
C2809 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.02fF
C2810 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.03fF
C2811 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C2812 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C2813 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.00fF
C2814 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C2815 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.01fF
C2816 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A -0.00fF
C2817 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.07fF
C2818 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.00fF
C2819 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.08fF
C2820 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C2821 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C2822 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# sky130_fd_sc_hd__nand2_1_0/A 0.10fF
C2823 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C2824 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C2825 sky130_fd_sc_hd__nand2_1_1/A Ad_b 0.55fF
C2826 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C2827 VDD sky130_fd_sc_hd__mux2_1_0/S -0.29fF
C2828 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.08fF
C2829 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A -0.00fF
C2830 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C2831 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C2832 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.02fF
C2833 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.11fF
C2834 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A -0.00fF
C2835 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.00fF
C2836 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X -0.00fF
C2837 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C2838 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.78fF
C2839 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C2840 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.01fF
C2841 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.01fF
C2842 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.01fF
C2843 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.07fF
C2844 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C2845 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C2846 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.01fF
C2847 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C2848 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__nand2_4_3/Y 0.19fF
C2849 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C2850 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.03fF
C2851 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C2852 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.06fF
C2853 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.04fF
C2854 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_1_1/A 0.06fF
C2855 sky130_fd_sc_hd__clkinv_1_1/Y sky130_fd_sc_hd__nand2_4_3/A 0.03fF
C2856 sky130_fd_sc_hd__clkinv_4_7/A VSUBS 0.25fF
C2857 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C2858 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C2859 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.01fF
C2860 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.01fF
C2861 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.04fF
C2862 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 2.25fF
C2863 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.01fF
C2864 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.01fF
C2865 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C2866 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C2867 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.11fF
C2868 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.19fF
C2869 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C2870 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C2871 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C2872 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.01fF
C2873 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.00fF
C2874 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.00fF
C2875 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C2876 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C2877 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C2878 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 2.82fF
C2879 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C2880 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C2881 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.04fF
C2882 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C2883 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.04fF
C2884 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# 0.14fF
C2885 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.01fF
C2886 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_4/B 0.00fF
C2887 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.05fF
C2888 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.02fF
C2889 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.08fF
C2890 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.01fF
C2891 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C2892 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C2893 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.12fF
C2894 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.04fF
C2895 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C2896 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C2897 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.00fF
C2898 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C2899 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.01fF
C2900 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C2901 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.01fF
C2902 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C2903 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C2904 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C2905 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.14fF
C2906 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.01fF
C2907 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.07fF
C2908 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C2909 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Ad_b 0.09fF
C2910 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.01fF
C2911 VDD sky130_fd_sc_hd__clkbuf_16_5/a_110_47# -0.06fF
C2912 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# -0.01fF
C2913 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_4/Y 0.06fF
C2914 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__nand2_4_0/A 0.06fF
C2915 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C2916 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C2917 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.00fF
C2918 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.03fF
C2919 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C2920 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.04fF
C2921 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.04fF
C2922 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C2923 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.05fF
C2924 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C2925 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.02fF
C2926 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.00fF
C2927 VDD sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.10fF
C2928 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.19fF
C2929 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.11fF
C2930 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__mux2_1_0/X 0.07fF
C2931 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C2932 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C2933 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.00fF
C2934 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 1.48fF
C2935 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__nand2_1_0/A 0.02fF
C2936 p1_b sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.15fF
C2937 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# p1d 0.15fF
C2938 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.27fF
C2939 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C2940 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C2941 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C2942 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X Bd_b 0.05fF
C2943 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C2944 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C2945 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C2946 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C2947 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C2948 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.19fF
C2949 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.00fF
C2950 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C2951 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C2952 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C2953 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.03fF
C2954 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.04fF
C2955 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.04fF
C2956 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.01fF
C2957 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.02fF
C2958 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C2959 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.41fF
C2960 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.11fF
C2961 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A -0.00fF
C2962 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X Bd_b 0.05fF
C2963 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C2964 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C2965 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.03fF
C2966 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.01fF
C2967 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.03fF
C2968 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.05fF
C2969 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.03fF
C2970 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSUBS -0.01fF
C2971 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_4_3/A 0.13fF
C2972 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.01fF
C2973 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.09fF
C2974 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C2975 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C2976 VDD sky130_fd_sc_hd__clkinv_4_2/Y 1.52fF
C2977 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.02fF
C2978 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# 0.34fF
C2979 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.03fF
C2980 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/X -0.16fF
C2981 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C2982 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/B 0.11fF
C2983 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_4/Y 0.04fF
C2984 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.03fF
C2985 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.02fF
C2986 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C2987 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C2988 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.03fF
C2989 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.05fF
C2990 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C2991 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.03fF
C2992 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.02fF
C2993 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.02fF
C2994 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.00fF
C2995 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.00fF
C2996 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.03fF
C2997 VDD p1_b 1.24fF
C2998 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.04fF
C2999 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.04fF
C3000 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C3001 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C3002 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C3003 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.05fF
C3004 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.05fF
C3005 VSUBS sky130_fd_sc_hd__nand2_4_1/A -0.20fF
C3006 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.30fF
C3007 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0.15fF
C3008 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C3009 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C3010 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C3011 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.23fF
C3012 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# Bd_b 0.01fF
C3013 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# Ad_b 0.01fF
C3014 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.24fF
C3015 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__nand2_4_3/Y 0.02fF
C3016 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0.34fF
C3017 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.00fF
C3018 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.00fF
C3019 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C3020 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.07fF
C3021 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C3022 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C3023 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C3024 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.01fF
C3025 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C3026 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.02fF
C3027 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.04fF
C3028 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C3029 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.15fF
C3030 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C3031 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X -0.00fF
C3032 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C3033 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C3034 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C3035 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.01fF
C3036 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C3037 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.05fF
C3038 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C3039 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.01fF
C3040 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C3041 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 1.05fF
C3042 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.01fF
C3043 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C3044 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C3045 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C3046 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.15fF
C3047 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# 0.08fF
C3048 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__nand2_4_3/Y 0.04fF
C3049 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C3050 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C3051 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.14fF
C3052 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C3053 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.02fF
C3054 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.01fF
C3055 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C3056 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.17fF
C3057 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__mux2_1_0/S 0.05fF
C3058 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.12fF
C3059 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.49fF
C3060 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.10fF
C3061 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.01fF
C3062 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.02fF
C3063 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.02fF
C3064 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.07fF
C3065 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.04fF
C3066 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.04fF
C3067 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.04fF
C3068 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.15fF
C3069 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C3070 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/X -0.60fF
C3071 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# p2 -0.00fF
C3072 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C3073 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C3074 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0.09fF
C3075 VDD sky130_fd_sc_hd__nand2_4_3/B 0.58fF
C3076 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# Ad_b 0.02fF
C3077 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.00fF
C3078 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.00fF
C3079 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.05fF
C3080 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.05fF
C3081 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C3082 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C3083 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.32fF
C3084 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.11fF
C3085 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3086 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.09fF
C3087 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C3088 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.05fF
C3089 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C3090 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0.02fF
C3091 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C3092 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.01fF
C3093 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C3094 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C3095 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.13fF
C3096 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C3097 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.00fF
C3098 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.00fF
C3099 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.02fF
C3100 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C3101 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C3102 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.02fF
C3103 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.02fF
C3104 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.07fF
C3105 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.08fF
C3106 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C3107 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.02fF
C3108 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C3109 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.08fF
C3110 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.31fF
C3111 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C3112 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.01fF
C3113 sky130_fd_sc_hd__nand2_4_0/Y VDD 6.10fF
C3114 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.18fF
C3115 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3116 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C3117 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C3118 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.17fF
C3119 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.01fF
C3120 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.03fF
C3121 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3122 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C3123 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C3124 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C3125 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.04fF
C3126 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.04fF
C3127 VDD sky130_fd_sc_hd__nand2_4_3/A 10.99fF
C3128 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.02fF
C3129 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/B 0.02fF
C3130 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.00fF
C3131 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/A -0.59fF
C3132 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C3133 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.00fF
C3134 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C3135 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C3136 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C3137 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.00fF
C3138 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 2.24fF
C3139 sky130_fd_sc_hd__mux2_1_0/X Ad_b 0.00fF
C3140 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# 0.01fF
C3141 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__nand2_4_0/B 0.02fF
C3142 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.12fF
C3143 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.04fF
C3144 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.04fF
C3145 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.05fF
C3146 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C3147 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C3148 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.30fF
C3149 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.01fF
C3150 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C3151 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C3152 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C3153 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.05fF
C3154 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C3155 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.02fF
C3156 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.01fF
C3157 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.00fF
C3158 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.00fF
C3159 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C3160 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.01fF
C3161 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.00fF
C3162 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C3163 sky130_fd_sc_hd__clkinv_4_4/Y Bd_b 0.08fF
C3164 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.03fF
C3165 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C3166 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.01fF
C3167 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C3168 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.07fF
C3169 VDD sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.22fF
C3170 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C3171 sky130_fd_sc_hd__nand2_4_1/Y VSUBS -0.31fF
C3172 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.12fF
C3173 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.15fF
C3174 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C3175 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.08fF
C3176 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C3177 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C3178 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Ad_b 0.02fF
C3179 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.02fF
C3180 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.02fF
C3181 p2d_b sky130_fd_sc_hd__clkbuf_16_11/a_110_47# 0.02fF
C3182 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VDD 0.17fF
C3183 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3184 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C3185 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.15fF
C3186 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.15fF
C3187 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.04fF
C3188 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C3189 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C3190 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C3191 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C3192 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C3193 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C3194 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C3195 sky130_fd_sc_hd__nand2_1_2/A clk 0.05fF
C3196 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0.00fF
C3197 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.08fF
C3198 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.01fF
C3199 p1d_b p1_b 0.19fF
C3200 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C3201 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C3202 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C3203 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C3204 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C3205 sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C3206 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C3207 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.00fF
C3208 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.00fF
C3209 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C3210 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C3211 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C3212 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C3213 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.02fF
C3214 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C3215 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C3216 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C3217 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C3218 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C3219 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# A_b 0.15fF
C3220 Ad sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.15fF
C3221 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.02fF
C3222 p2 sky130_fd_sc_hd__nand2_4_3/Y 0.09fF
C3223 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.01fF
C3224 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.09fF
C3225 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C3226 sky130_fd_sc_hd__clkinv_4_3/Y Bd_b 0.18fF
C3227 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C3228 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.15fF
C3229 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0.10fF
C3230 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.01fF
C3231 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C3232 VDD sky130_fd_sc_hd__clkinv_1_2/Y 0.21fF
C3233 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C3234 p2_b p2d_b 0.22fF
C3235 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkbuf_16_11/a_110_47# 0.04fF
C3236 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.08fF
C3237 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C3238 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C3239 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C3240 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C3241 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C3242 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.18fF
C3243 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.04fF
C3244 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C3245 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C3246 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0.02fF
C3247 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.31fF
C3248 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C3249 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C3250 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C3251 sky130_fd_sc_hd__clkinv_1_0/Y VDD 0.26fF
C3252 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.15fF
C3253 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkinv_4_4/Y 0.02fF
C3254 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.02fF
C3255 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C3256 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VDD 0.31fF
C3257 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.55fF
C3258 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C3259 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.06fF
C3260 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkinv_4_8/Y 0.03fF
C3261 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C3262 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C3263 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C3264 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.00fF
C3265 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Ad_b 0.07fF
C3266 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 1.21fF
C3267 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_1/A 0.02fF
C3268 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.03fF
C3269 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C3270 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C3271 VDD sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.34fF
C3272 B_b Bd_b 0.20fF
C3273 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C3274 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.14fF
C3275 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A Bd_b 0.05fF
C3276 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.04fF
C3277 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.04fF
C3278 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.16fF
C3279 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C3280 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.02fF
C3281 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.03fF
C3282 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C3283 VSUBS clk 0.00fF
C3284 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.15fF
C3285 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.01fF
C3286 sky130_fd_sc_hd__clkinv_4_9/Y VDD 1.49fF
C3287 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.08fF
C3288 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.01fF
C3289 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C3290 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3291 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.05fF
C3292 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.19fF
C3293 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__clkinv_4_4/Y 0.07fF
C3294 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.03fF
C3295 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.02fF
C3296 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C3297 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.02fF
C3298 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.00fF
C3299 sky130_fd_sc_hd__nand2_1_1/A Bd_b 1.60fF
C3300 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C3301 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C3302 VDD Ad_b 5.95fF
C3303 sky130_fd_sc_hd__clkinv_1_3/A VSUBS 0.38fF
C3304 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C3305 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C3306 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.00fF
C3307 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C3308 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_1_2/Y 0.36fF
C3309 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.34fF
C3310 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.45fF
C3311 sky130_fd_sc_hd__nand2_4_2/B sky130_fd_sc_hd__nand2_4_2/A 0.80fF
C3312 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C3313 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.01fF
C3314 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_4_3/A 0.32fF
C3315 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C3316 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C3317 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.04fF
C3318 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.64fF
C3319 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.05fF
C3320 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.05fF
C3321 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C3322 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C3323 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_1_1/A 0.10fF
C3324 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C3325 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VDD 0.53fF
C3326 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A -0.00fF
C3327 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.02fF
C3328 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C3329 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# 0.05fF
C3330 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C3331 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C3332 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.05fF
C3333 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C3334 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C3335 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkinv_4_3/Y 0.04fF
C3336 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.07fF
C3337 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.01fF
C3338 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.03fF
C3339 p2d p2_b 0.53fF
C3340 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C3341 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X -0.00fF
C3342 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.00fF
C3343 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.01fF
C3344 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.01fF
C3345 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.03fF
C3346 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C3347 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C3348 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C3349 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.03fF
C3350 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.11fF
C3351 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C3352 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C3353 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.00fF
C3354 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.01fF
C3355 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C3356 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.04fF
C3357 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C3358 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.00fF
C3359 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C3360 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C3361 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.01fF
C3362 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.04fF
C3363 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.04fF
C3364 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C3365 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C3366 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C3367 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.10fF
C3368 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.04fF
C3369 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.01fF
C3370 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C3371 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.02fF
C3372 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.02fF
C3373 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C3374 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C3375 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.02fF
C3376 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.02fF
C3377 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.01fF
C3378 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.03fF
C3379 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A -0.00fF
C3380 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C3381 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.00fF
C3382 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C3383 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.08fF
C3384 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C3385 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.10fF
C3386 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__mux2_1_0/S 0.04fF
C3387 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.97fF
C3388 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A Bd_b 0.07fF
C3389 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.08fF
C3390 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.19fF
C3391 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A -0.00fF
C3392 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C3393 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C3394 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C3395 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.03fF
C3396 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkinv_4_3/Y 0.01fF
C3397 VDD sky130_fd_sc_hd__nand2_1_4/Y 0.45fF
C3398 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.22fF
C3399 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.19fF
C3400 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.01fF
C3401 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.01fF
C3402 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C3403 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.01fF
C3404 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.11fF
C3405 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.08fF
C3406 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.06fF
C3407 VDD sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.12fF
C3408 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.05fF
C3409 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C3410 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C3411 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# -0.00fF
C3412 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.01fF
C3413 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C3414 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__nand2_4_1/B 0.07fF
C3415 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.08fF
C3416 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkinv_4_1/A 0.01fF
C3417 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C3418 sky130_fd_sc_hd__clkinv_4_1/A VSUBS 0.38fF
C3419 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.03fF
C3420 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.02fF
C3421 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C3422 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C3423 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.04fF
C3424 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.01fF
C3425 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.08fF
C3426 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.07fF
C3427 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.05fF
C3428 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C3429 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C3430 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C3431 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.01fF
C3432 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.02fF
C3433 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.02fF
C3434 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C3435 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C3436 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C3437 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C3438 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# Ad_b 0.12fF
C3439 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C3440 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.03fF
C3441 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C3442 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.01fF
C3443 VDD sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.67fF
C3444 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.01fF
C3445 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.01fF
C3446 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.01fF
C3447 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_1/A 0.37fF
C3448 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.02fF
C3449 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.02fF
C3450 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.03fF
C3451 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.01fF
C3452 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.01fF
C3453 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0.01fF
C3454 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0.02fF
C3455 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C3456 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.04fF
C3457 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.04fF
C3458 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C3459 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.02fF
C3460 VDD sky130_fd_sc_hd__nand2_4_1/B 0.69fF
C3461 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.01fF
C3462 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C3463 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C3464 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C3465 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C3466 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.03fF
C3467 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.04fF
C3468 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.00fF
C3469 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C3470 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.04fF
C3471 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.04fF
C3472 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.18fF
C3473 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# 0.17fF
C3474 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C3475 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 1.36fF
C3476 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C3477 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C3478 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.31fF
C3479 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C3480 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C3481 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C3482 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.00fF
C3483 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.02fF
C3484 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.01fF
C3485 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C3486 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.04fF
C3487 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.04fF
C3488 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.04fF
C3489 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkinv_4_8/Y 0.04fF
C3490 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.01fF
C3491 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C3492 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C3493 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# 0.10fF
C3494 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.27fF
C3495 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C3496 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.01fF
C3497 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C3498 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.01fF
C3499 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.15fF
C3500 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.04fF
C3501 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C3502 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# 0.15fF
C3503 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.15fF
C3504 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 1.20fF
C3505 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.02fF
C3506 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C3507 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.17fF
C3508 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# Bd_b 0.01fF
C3509 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.05fF
C3510 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C3511 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3512 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C3513 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.14fF
C3514 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.01fF
C3515 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.02fF
C3516 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.04fF
C3517 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C3518 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C3519 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.01fF
C3520 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C3521 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C3522 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.04fF
C3523 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.04fF
C3524 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.17fF
C3525 sky130_fd_sc_hd__nand2_1_0/a_113_47# sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C3526 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_1/Y 0.03fF
C3527 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C3528 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.29fF
C3529 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.01fF
C3530 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.02fF
C3531 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/B 0.14fF
C3532 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.02fF
C3533 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C3534 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.37fF
C3535 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.00fF
C3536 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.02fF
C3537 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.02fF
C3538 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.00fF
C3539 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.02fF
C3540 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# sky130_fd_sc_hd__nand2_4_2/A 0.34fF
C3541 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C3542 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C3543 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.03fF
C3544 VSUBS sky130_fd_sc_hd__clkinv_4_7/Y 0.00fF
C3545 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.02fF
C3546 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.02fF
C3547 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.07fF
C3548 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C3549 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C3550 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.31fF
C3551 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C3552 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C3553 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.03fF
C3554 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C3555 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.07fF
C3556 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.32fF
C3557 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.15fF
C3558 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.08fF
C3559 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# 0.04fF
C3560 p2_b sky130_fd_sc_hd__clkinv_4_10/Y 0.03fF
C3561 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C3562 Ad A 0.19fF
C3563 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.09fF
C3564 VSUBS sky130_fd_sc_hd__nand2_1_0/A 0.01fF
C3565 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C3566 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C3567 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C3568 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.14fF
C3569 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.14fF
C3570 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.02fF
C3571 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.00fF
C3572 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C3573 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C3574 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.09fF
C3575 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C3576 sky130_fd_sc_hd__nand2_4_1/A Ad_b 0.48fF
C3577 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.01fF
C3578 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.04fF
C3579 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.20fF
C3580 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.09fF
C3581 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C3582 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C3583 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.31fF
C3584 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_1_2/A 0.26fF
C3585 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.01fF
C3586 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.01fF
C3587 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.01fF
C3588 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C3589 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C3590 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.04fF
C3591 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 2.82fF
C3592 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C3593 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# Bd_b 0.46fF
C3594 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C3595 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0.00fF
C3596 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C3597 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.14fF
C3598 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.01fF
C3599 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.01fF
C3600 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C3601 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C3602 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.03fF
C3603 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.08fF
C3604 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C3605 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.01fF
C3606 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.00fF
C3607 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.05fF
C3608 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C3609 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.07fF
C3610 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3611 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.08fF
C3612 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C3613 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.13fF
C3614 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.03fF
C3615 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C3616 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C3617 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.02fF
C3618 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.01fF
C3619 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.10fF
C3620 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# p1d 0.12fF
C3621 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VDD -0.76fF
C3622 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.06fF
C3623 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C3624 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C3625 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.02fF
C3626 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.01fF
C3627 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C3628 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C3629 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Ad_b 0.02fF
C3630 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.14fF
C3631 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.05fF
C3632 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.11fF
C3633 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3634 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C3635 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 1.48fF
C3636 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C3637 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C3638 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C3639 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.01fF
C3640 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C3641 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C3642 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C3643 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.08fF
C3644 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C3645 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.02fF
C3646 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C3647 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.05fF
C3648 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.03fF
C3649 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_2/Y 0.68fF
C3650 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C3651 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C3652 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C3653 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C3654 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.00fF
C3655 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C3656 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.01fF
C3657 sky130_fd_sc_hd__nand2_4_1/A sky130_fd_sc_hd__nand2_1_4/Y 0.04fF
C3658 sky130_fd_sc_hd__mux2_1_0/X Bd_b 0.01fF
C3659 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.07fF
C3660 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.04fF
C3661 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.88fF
C3662 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C3663 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.01fF
C3664 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.01fF
C3665 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.01fF
C3666 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C3667 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C3668 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/B 0.11fF
C3669 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.04fF
C3670 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.04fF
C3671 sky130_fd_sc_hd__clkinv_4_4/w_82_21# sky130_fd_sc_hd__clkinv_4_5/Y 0.03fF
C3672 sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C3673 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.06fF
C3674 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C3675 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.01fF
C3676 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.10fF
C3677 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C3678 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C3679 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.06fF
C3680 VDD sky130_fd_sc_hd__nand2_4_2/A 5.81fF
C3681 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C3682 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 1.32fF
C3683 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A sky130_fd_sc_hd__nand2_4_3/A 0.47fF
C3684 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.00fF
C3685 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.00fF
C3686 A_b Ad_b 0.33fF
C3687 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.07fF
C3688 sky130_fd_sc_hd__clkinv_4_0/w_82_21# sky130_fd_sc_hd__nand2_4_0/A -0.29fF
C3689 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.09fF
C3690 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.05fF
C3691 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.04fF
C3692 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.04fF
C3693 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C3694 VSUBS sky130_fd_sc_hd__nand2_1_3/A -0.00fF
C3695 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C3696 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.04fF
C3697 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.02fF
C3698 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C3699 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C3700 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.16fF
C3701 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3702 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_11/a_110_47# 0.04fF
C3703 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# 0.25fF
C3704 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.05fF
C3705 sky130_fd_sc_hd__nand2_4_3/A clk 0.03fF
C3706 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C3707 sky130_fd_sc_hd__clkinv_4_5/w_82_21# sky130_fd_sc_hd__clkinv_4_5/Y -0.00fF
C3708 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C3709 sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C3710 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X Bd_b 0.02fF
C3711 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# 0.71fF
C3712 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.04fF
C3713 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.04fF
C3714 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C3715 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C3716 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_4/Y 0.01fF
C3717 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_1/A 0.87fF
C3718 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0.02fF
C3719 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C3720 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C3721 sky130_fd_sc_hd__clkinv_4_11/w_82_21# sky130_fd_sc_hd__clkinv_1_3/A 0.05fF
C3722 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkinv_1_1/Y 0.37fF
C3723 VSUBS sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C3724 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_4_3/A 1.25fF
C3725 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.15fF
C3726 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.18fF
C3727 sky130_fd_sc_hd__clkinv_4_3/w_82_21# sky130_fd_sc_hd__clkinv_4_3/Y -0.00fF
C3728 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C3729 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.08fF
C3730 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C3731 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C3732 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C3733 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C3734 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C3735 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.00fF
C3736 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C3737 p2_b sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.15fF
C3738 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C3739 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C3740 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.02fF
C3741 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.02fF
C3742 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C3743 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.01fF
C3744 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C3745 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C3746 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C3747 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C3748 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.00fF
C3749 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C3750 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C3751 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.04fF
C3752 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.03fF
C3753 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C3754 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.01fF
C3755 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C3756 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.19fF
C3757 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C3758 sky130_fd_sc_hd__nand2_4_1/Y Ad_b 0.00fF
C3759 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C3760 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C3761 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.01fF
C3762 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C3763 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C3764 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C3765 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p2_b 0.06fF
C3766 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_1_1/A 0.05fF
C3767 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__nand2_4_2/A 1.13fF
C3768 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.10fF
C3769 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X -0.00fF
C3770 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C3771 p2d_b VDD 0.79fF
C3772 sky130_fd_sc_hd__clkinv_4_7/Y p1_b 0.03fF
C3773 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.03fF
C3774 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C3775 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.09fF
C3776 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.03fF
C3777 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C3778 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C3779 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C3780 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_2/B 0.07fF
C3781 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# A_b 0.06fF
C3782 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.01fF
C3783 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.03fF
C3784 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.51fF
C3785 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.19fF
C3786 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/Y 0.73fF
C3787 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.04fF
C3788 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.04fF
C3789 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0.09fF
C3790 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.05fF
C3791 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C3792 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C3793 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C3794 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C3795 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.03fF
C3796 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VDD 0.18fF
C3797 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0.08fF
C3798 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.05fF
C3799 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# sky130_fd_sc_hd__nand2_4_1/A 0.08fF
C3800 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.31fF
C3801 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C3802 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C3803 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C3804 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.01fF
C3805 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.31fF
C3806 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X Bd_b 0.07fF
C3807 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C3808 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.01fF
C3809 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.12fF
C3810 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.04fF
C3811 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.06fF
C3812 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C3813 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C3814 p2 sky130_fd_sc_hd__clkinv_4_3/Y 0.03fF
C3815 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.19fF
C3816 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VDD 1.07fF
C3817 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.00fF
C3818 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C3819 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0.01fF
C3820 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.01fF
C3821 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.14fF
C3822 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.02fF
C3823 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.01fF
C3824 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.03fF
C3825 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.08fF
C3826 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__mux2_1_0/X 0.03fF
C3827 sky130_fd_sc_hd__nand2_4_2/Y VDD 5.75fF
C3828 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.04fF
C3829 sky130_fd_sc_hd__nand2_4_3/a_27_47# VSUBS -0.05fF
C3830 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C3831 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C3832 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.02fF
C3833 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X sky130_fd_sc_hd__nand2_1_3/A 0.01fF
C3834 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C3835 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.02fF
C3836 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C3837 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C3838 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C3839 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C3840 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C3841 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C3842 VDD Bd_b 8.01fF
C3843 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.08fF
C3844 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C3845 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C3846 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C3847 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C3848 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C3849 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.17fF
C3850 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C3851 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C3852 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.04fF
C3853 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.31fF
C3854 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C3855 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.01fF
C3856 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C3857 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VDD 0.34fF
C3858 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.01fF
C3859 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.01fF
C3860 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.03fF
C3861 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.10fF
C3862 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__nand2_1_0/B 0.06fF
C3863 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.01fF
C3864 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C3865 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.01fF
C3866 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.02fF
C3867 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.01fF
C3868 sky130_fd_sc_hd__nand2_4_0/B VSUBS -0.02fF
C3869 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C3870 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__nand2_4_1/B 0.16fF
C3871 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.05fF
C3872 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C3873 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C3874 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C3875 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.00fF
C3876 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VDD 0.36fF
C3877 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C3878 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.04fF
C3879 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.04fF
C3880 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C3881 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C3882 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C3883 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.04fF
C3884 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 2.83fF
C3885 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.02fF
C3886 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0.08fF
C3887 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Ad_b 0.03fF
C3888 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C3889 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.24fF
C3890 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.02fF
C3891 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X -0.00fF
C3892 p2d VDD 1.53fF
C3893 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.11fF
C3894 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.07fF
C3895 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 2.83fF
C3896 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.00fF
C3897 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.01fF
C3898 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.01fF
C3899 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X sky130_fd_sc_hd__nand2_1_2/B 0.03fF
C3900 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_150/X -0.28fF
C3901 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C3902 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.01fF
C3903 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.07fF
C3904 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.04fF
C3905 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.00fF
C3906 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C3907 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.01fF
C3908 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.02fF
C3909 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.02fF
C3910 sky130_fd_sc_hd__clkinv_4_6/w_82_21# sky130_fd_sc_hd__clkinv_4_7/A -0.00fF
C3911 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C3912 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C3913 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.08fF
C3914 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.19fF
C3915 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C3916 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C3917 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C3918 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_9/Y 0.68fF
C3919 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C3920 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.02fF
C3921 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C3922 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.01fF
C3923 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.01fF
C3924 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.07fF
C3925 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.01fF
C3926 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C3927 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C3928 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.02fF
C3929 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C3930 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.00fF
C3931 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.00fF
C3932 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C3933 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.01fF
C3934 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C3935 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.00fF
C3936 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.02fF
C3937 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C3938 sky130_fd_sc_hd__clkinv_1_3/A Ad_b 0.25fF
C3939 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.10fF
C3940 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.03fF
C3941 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# -0.07fF
C3942 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.10fF
C3943 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.03fF
C3944 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.00fF
C3945 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C3946 p2 sky130_fd_sc_hd__nand2_1_1/A 0.01fF
C3947 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.04fF
C3948 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.04fF
C3949 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C3950 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C3951 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C3952 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.10fF
C3953 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.09fF
C3954 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.02fF
C3955 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.02fF
C3956 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.00fF
C3957 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 3.22fF
C3958 p2_b p2 0.47fF
C3959 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C3960 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_7/A 0.72fF
C3961 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C3962 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.07fF
C3963 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.08fF
C3964 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.33fF
C3965 VDD sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.06fF
C3966 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.08fF
C3967 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.00fF
C3968 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.00fF
C3969 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.07fF
C3970 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.01fF
C3971 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.01fF
C3972 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.03fF
C3973 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C3974 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.05fF
C3975 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.53fF
C3976 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkinv_1_3/A 0.04fF
C3977 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.11fF
C3978 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.14fF
C3979 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C3980 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C3981 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C3982 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0.00fF
C3983 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.01fF
C3984 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__nand2_4_0/Y 0.16fF
C3985 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C3986 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C3987 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_1_0/Y 0.37fF
C3988 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/X -0.30fF
C3989 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C3990 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C3991 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C3992 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C3993 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C3994 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.00fF
C3995 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C3996 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.03fF
C3997 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# Bd_b 0.10fF
C3998 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__nand2_1_1/A 0.05fF
C3999 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C4000 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C4001 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C4002 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C4003 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.08fF
C4004 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0.02fF
C4005 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.02fF
C4006 sky130_fd_sc_hd__clkinv_4_5/Y VDD 4.38fF
C4007 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.30fF
C4008 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.11fF
C4009 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C4010 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C4011 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.01fF
C4012 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C4013 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.00fF
C4014 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C4015 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C4016 p1d_b p2d_b 0.11fF
C4017 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# -0.00fF
C4018 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.04fF
C4019 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4020 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.32fF
C4021 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.02fF
C4022 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.02fF
C4023 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.01fF
C4024 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C4025 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# 0.15fF
C4026 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C4027 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.03fF
C4028 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.03fF
C4029 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.18fF
C4030 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.09fF
C4031 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.03fF
C4032 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C4033 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C4034 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C4035 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.29fF
C4036 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C4037 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.34fF
C4038 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.00fF
C4039 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C4040 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.01fF
C4041 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.01fF
C4042 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.01fF
C4043 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C4044 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.08fF
C4045 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.07fF
C4046 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.02fF
C4047 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.02fF
C4048 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C4049 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.02fF
C4050 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C4051 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.15fF
C4052 p2d_b sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.07fF
C4053 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C4054 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.03fF
C4055 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4056 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C4057 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C4058 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C4059 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C4060 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.00fF
C4061 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.11fF
C4062 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.04fF
C4063 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.04fF
C4064 VDD sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.45fF
C4065 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.01fF
C4066 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.01fF
C4067 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.01fF
C4068 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.15fF
C4069 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.11fF
C4070 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C4071 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# 0.00fF
C4072 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.01fF
C4073 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C4074 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C4075 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.25fF
C4076 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_4_3/A 0.69fF
C4077 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C4078 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 6.89fF
C4079 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C4080 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C4081 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.01fF
C4082 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.05fF
C4083 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.00fF
C4084 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C4085 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C4086 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.01fF
C4087 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.00fF
C4088 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkinv_1_2/Y 0.05fF
C4089 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.14fF
C4090 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C4091 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.14fF
C4092 sky130_fd_sc_hd__clkinv_4_10/Y VDD 0.49fF
C4093 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C4094 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C4095 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# 0.04fF
C4096 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C4097 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.00fF
C4098 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.00fF
C4099 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.00fF
C4100 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.02fF
C4101 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__nand2_4_2/B 0.00fF
C4102 sky130_fd_sc_hd__nand2_4_1/A Bd_b 0.66fF
C4103 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.14fF
C4104 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C4105 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.01fF
C4106 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C4107 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C4108 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.14fF
C4109 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.04fF
C4110 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C4111 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C4112 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.00fF
C4113 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C4114 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.19fF
C4115 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0.02fF
C4116 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4117 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.02fF
C4118 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.25fF
C4119 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.01fF
C4120 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.05fF
C4121 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.02fF
C4122 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.02fF
C4123 sky130_fd_sc_hd__nand2_4_2/a_27_47# VSUBS -0.05fF
C4124 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0.00fF
C4125 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.00fF
C4126 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.15fF
C4127 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.19fF
C4128 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkinv_1_2/Y 0.00fF
C4129 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.00fF
C4130 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C4131 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C4132 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.08fF
C4133 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__nand2_4_1/A 0.03fF
C4134 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.01fF
C4135 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C4136 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C4137 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C4138 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.08fF
C4139 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.03fF
C4140 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.08fF
C4141 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C4142 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.01fF
C4143 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.03fF
C4144 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.04fF
C4145 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.04fF
C4146 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.01fF
C4147 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C4148 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# p1d 0.05fF
C4149 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.09fF
C4150 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C4151 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.05fF
C4152 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A -0.00fF
C4153 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4154 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X Bd_b 0.02fF
C4155 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.14fF
C4156 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C4157 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.05fF
C4158 p2d sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.15fF
C4159 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C4160 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C4161 VDD sky130_fd_sc_hd__nand2_4_0/A 16.63fF
C4162 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C4163 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C4164 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.00fF
C4165 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.00fF
C4166 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C4167 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.03fF
C4168 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.02fF
C4169 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.02fF
C4170 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.31fF
C4171 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.03fF
C4172 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.06fF
C4173 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__clkinv_1_2/Y 0.01fF
C4174 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C4175 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C4176 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Ad_b 0.04fF
C4177 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/B 0.07fF
C4178 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C4179 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C4180 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.08fF
C4181 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_4/B 0.92fF
C4182 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.00fF
C4183 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C4184 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.07fF
C4185 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0.02fF
C4186 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.02fF
C4187 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C4188 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C4189 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.22fF
C4190 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C4191 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C4192 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.01fF
C4193 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.01fF
C4194 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.01fF
C4195 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C4196 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4197 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.02fF
C4198 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C4199 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.00fF
C4200 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4201 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.04fF
C4202 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.04fF
C4203 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C4204 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.01fF
C4205 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.01fF
C4206 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A -0.00fF
C4207 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.01fF
C4208 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C4209 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.01fF
C4210 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkinv_4_7/w_82_21# 0.03fF
C4211 VDD p1d 1.51fF
C4212 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.00fF
C4213 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C4214 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C4215 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0.16fF
C4216 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.06fF
C4217 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkinv_4_8/Y 0.02fF
C4218 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_4_1/A 1.26fF
C4219 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C4220 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C4221 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C4222 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.02fF
C4223 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# 0.18fF
C4224 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.02fF
C4225 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkinv_4_1/w_82_21# 0.03fF
C4226 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.01fF
C4227 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C4228 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.00fF
C4229 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.01fF
C4230 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C4231 VSUBS sky130_fd_sc_hd__nand2_1_2/A -0.02fF
C4232 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X sky130_fd_sc_hd__nand2_4_1/A 0.01fF
C4233 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.01fF
C4234 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C4235 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.15fF
C4236 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C4237 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C4238 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0.00fF
C4239 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C4240 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VDD 0.37fF
C4241 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.01fF
C4242 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VDD 0.14fF
C4243 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.01fF
C4244 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.10fF
C4245 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__nand2_4_0/B 0.16fF
C4246 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.00fF
C4247 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A sky130_fd_sc_hd__nand2_1_4/B 0.04fF
C4248 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C4249 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C4250 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C4251 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.04fF
C4252 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C4253 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C4254 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C4255 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.04fF
C4256 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.04fF
C4257 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.00fF
C4258 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/A -0.00fF
C4259 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.01fF
C4260 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C4261 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C4262 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.08fF
C4263 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 2.25fF
C4264 sky130_fd_sc_hd__nand2_4_1/Y Bd_b 0.22fF
C4265 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C4266 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.14fF
C4267 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.03fF
C4268 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C4269 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.00fF
C4270 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C4271 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VDD 0.42fF
C4272 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.08fF
C4273 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VDD -0.18fF
C4274 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/X -0.00fF
C4275 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.02fF
C4276 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_4_1/A 2.16fF
C4277 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A sky130_fd_sc_hd__nand2_4_2/A 0.41fF
C4278 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__nand2_4_1/B 0.02fF
C4279 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 1.23fF
C4280 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.05fF
C4281 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.08fF
C4282 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4283 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.02fF
C4284 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkinv_1_1/Y 0.05fF
C4285 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0.09fF
C4286 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C4287 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C4288 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_1_2/A 0.00fF
C4289 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# 0.11fF
C4290 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C4291 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.01fF
C4292 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.01fF
C4293 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C4294 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.03fF
C4295 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.01fF
C4296 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C4297 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C4298 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.08fF
C4299 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.19fF
C4300 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.08fF
C4301 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.03fF
C4302 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.02fF
C4303 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.01fF
C4304 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C4305 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VDD 0.16fF
C4306 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C4307 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.16fF
C4308 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.08fF
C4309 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C4310 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C4311 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C4312 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C4313 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.33fF
C4314 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C4315 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.18fF
C4316 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.08fF
C4317 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C4318 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C4319 sky130_fd_sc_hd__nand2_1_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.05fF
C4320 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/A -0.00fF
C4321 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.11fF
C4322 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.01fF
C4323 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.00fF
C4324 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C4325 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.02fF
C4326 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0.02fF
C4327 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/A -0.00fF
C4328 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.04fF
C4329 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.08fF
C4330 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.01fF
C4331 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C4332 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C4333 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.04fF
C4334 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.03fF
C4335 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.01fF
C4336 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C4337 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.01fF
C4338 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C4339 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C4340 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.02fF
C4341 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.15fF
C4342 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.05fF
C4343 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.00fF
C4344 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 1.06fF
C4345 p1 p1_b 0.47fF
C4346 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# A_b 0.09fF
C4347 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.00fF
C4348 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.03fF
C4349 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.01fF
C4350 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.01fF
C4351 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VDD 0.17fF
C4352 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.00fF
C4353 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C4354 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.01fF
C4355 VDD A 1.54fF
C4356 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 1.22fF
C4357 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.15fF
C4358 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.01fF
C4359 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.00fF
C4360 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C4361 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C4362 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkinv_4_5/Y 0.73fF
C4363 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.15fF
C4364 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.04fF
C4365 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.04fF
C4366 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VDD 0.17fF
C4367 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.08fF
C4368 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.23fF
C4369 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.04fF
C4370 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C4371 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C4372 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.01fF
C4373 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.01fF
C4374 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.02fF
C4375 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0.02fF
C4376 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.02fF
C4377 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C4378 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VDD 0.08fF
C4379 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.02fF
C4380 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.01fF
C4381 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.01fF
C4382 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.01fF
C4383 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0.00fF
C4384 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C4385 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4386 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.15fF
C4387 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A Bd_b 0.03fF
C4388 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C4389 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.14fF
C4390 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.01fF
C4391 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.08fF
C4392 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C4393 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.03fF
C4394 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C4395 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C4396 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C4397 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.05fF
C4398 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# 0.35fF
C4399 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.05fF
C4400 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__nand2_4_3/a_27_47# 0.01fF
C4401 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.01fF
C4402 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__clkinv_1_1/Y 0.08fF
C4403 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X -0.00fF
C4404 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C4405 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/S 0.05fF
C4406 VSUBS sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4407 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0.01fF
C4408 p1d_b p1d 0.47fF
C4409 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.08fF
C4410 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C4411 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C4412 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.02fF
C4413 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.32fF
C4414 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C4415 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.11fF
C4416 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.02fF
C4417 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.02fF
C4418 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C4419 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C4420 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.07fF
C4421 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.00fF
C4422 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.00fF
C4423 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C4424 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.02fF
C4425 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.11fF
C4426 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.02fF
C4427 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C4428 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C4429 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.02fF
C4430 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.10fF
C4431 sky130_fd_sc_hd__clkinv_1_3/A Bd_b 0.22fF
C4432 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.07fF
C4433 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C4434 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.04fF
C4435 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.00fF
C4436 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.07fF
C4437 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.07fF
C4438 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.01fF
C4439 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.01fF
C4440 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.01fF
C4441 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C4442 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.00fF
C4443 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C4444 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C4445 p2 VDD 4.24fF
C4446 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.10fF
C4447 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C4448 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C4449 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.02fF
C4450 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.04fF
C4451 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.02fF
C4452 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.14fF
C4453 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0.00fF
C4454 VDD sky130_fd_sc_hd__dfxbp_1_1/a_561_413# 0.01fF
C4455 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C4456 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0.31fF
C4457 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.05fF
C4458 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.05fF
C4459 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C4460 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.18fF
C4461 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.14fF
C4462 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkinv_1_3/A 0.03fF
C4463 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.01fF
C4464 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.04fF
C4465 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C4466 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C4467 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C4468 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.02fF
C4469 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.03fF
C4470 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 1.33fF
C4471 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__mux2_1_0/X 0.02fF
C4472 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.00fF
C4473 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C4474 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.00fF
C4475 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C4476 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C4477 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C4478 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C4479 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C4480 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.05fF
C4481 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.34fF
C4482 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 1.11fF
C4483 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C4484 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C4485 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.00fF
C4486 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C4487 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# p1d_b 0.02fF
C4488 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.02fF
C4489 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 1.14fF
C4490 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# A 0.04fF
C4491 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/D 0.91fF
C4492 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C4493 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# -0.08fF
C4494 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.01fF
C4495 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.07fF
C4496 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.09fF
C4497 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.01fF
C4498 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.02fF
C4499 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.02fF
C4500 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.01fF
C4501 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4502 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.01fF
C4503 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.00fF
C4504 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VDD 0.19fF
C4505 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C4506 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C4507 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C4508 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C4509 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4510 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.02fF
C4511 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.02fF
C4512 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0.01fF
C4513 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 2.24fF
C4514 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C4515 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.01fF
C4516 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.01fF
C4517 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.03fF
C4518 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C4519 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.01fF
C4520 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C4521 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C4522 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C4523 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.15fF
C4524 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.02fF
C4525 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C4526 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C4527 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C4528 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C4529 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.16fF
C4530 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.17fF
C4531 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C4532 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.00fF
C4533 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.02fF
C4534 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0.02fF
C4535 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0.02fF
C4536 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.07fF
C4537 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.08fF
C4538 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.33fF
C4539 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A sky130_fd_sc_hd__nand2_4_2/A 2.12fF
C4540 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.04fF
C4541 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.04fF
C4542 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.33fF
C4543 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C4544 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.42fF
C4545 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C4546 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.02fF
C4547 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C4548 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C4549 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4550 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0.00fF
C4551 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.04fF
C4552 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.04fF
C4553 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C4554 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C4555 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C4556 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C4557 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.02fF
C4558 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.11fF
C4559 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0.12fF
C4560 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.09fF
C4561 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C4562 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.01fF
C4563 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.01fF
C4564 VSUBS sky130_fd_sc_hd__clkinv_4_2/Y 0.01fF
C4565 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.02fF
C4566 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.14fF
C4567 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.02fF
C4568 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# sky130_fd_sc_hd__nand2_4_3/A 0.10fF
C4569 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.01fF
C4570 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C4571 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.00fF
C4572 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C4573 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.01fF
C4574 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.13fF
C4575 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkinv_4_5/Y 0.02fF
C4576 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.14fF
C4577 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.00fF
C4578 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.05fF
C4579 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.05fF
C4580 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0.31fF
C4581 B Bd 0.20fF
C4582 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C4583 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.00fF
C4584 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C4585 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C4586 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.01fF
C4587 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# sky130_fd_sc_hd__nand2_4_2/A 0.02fF
C4588 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.00fF
C4589 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 1.17fF
C4590 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.03fF
C4591 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.01fF
C4592 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# p2d_b 0.03fF
C4593 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.14fF
C4594 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 1.09fF
C4595 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C4596 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.01fF
C4597 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.14fF
C4598 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.08fF
C4599 sky130_fd_sc_hd__nand2_4_0/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.00fF
C4600 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.41fF
C4601 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.31fF
C4602 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.07fF
C4603 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C4604 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C4605 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__nand2_1_2/B 0.05fF
C4606 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.07fF
C4607 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.01fF
C4608 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.03fF
C4609 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C4610 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C4611 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C4612 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C4613 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.00fF
C4614 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.00fF
C4615 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C4616 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.16fF
C4617 sky130_fd_sc_hd__nand2_1_2/B sky130_fd_sc_hd__nand2_4_2/A 0.03fF
C4618 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C4619 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C4620 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.00fF
C4621 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.07fF
C4622 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.19fF
C4623 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.16fF
C4624 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.00fF
C4625 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.35fF
C4626 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.07fF
C4627 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.01fF
C4628 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_7/Y 0.19fF
C4629 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.04fF
C4630 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.04fF
C4631 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.04fF
C4632 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0.01fF
C4633 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C4634 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.00fF
C4635 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0.08fF
C4636 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.01fF
C4637 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C4638 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.04fF
C4639 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.04fF
C4640 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.01fF
C4641 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.01fF
C4642 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0.01fF
C4643 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.01fF
C4644 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/B 0.02fF
C4645 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.06fF
C4646 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.04fF
C4647 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C4648 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C4649 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkinv_1_3/A 0.32fF
C4650 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.01fF
C4651 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_4_3/Y 0.13fF
C4652 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.10fF
C4653 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C4654 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.03fF
C4655 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C4656 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.03fF
C4657 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C4658 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.04fF
C4659 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.08fF
C4660 VSUBS sky130_fd_sc_hd__nand2_4_3/B -0.02fF
C4661 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4662 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C4663 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C4664 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C4665 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.02fF
C4666 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.00fF
C4667 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.01fF
C4668 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C4669 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0.02fF
C4670 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.00fF
C4671 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A Bd_b 0.05fF
C4672 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_0/B 0.14fF
C4673 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0.01fF
C4674 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.01fF
C4675 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C4676 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C4677 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.08fF
C4678 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.31fF
C4679 sky130_fd_sc_hd__clkinv_4_1/Y B_b 0.03fF
C4680 p2 sky130_fd_sc_hd__nand2_4_1/A 0.17fF
C4681 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.26fF
C4682 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.14fF
C4683 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C4684 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C4685 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.01fF
C4686 VDD sky130_fd_sc_hd__nand2_1_4/B 2.14fF
C4687 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# sky130_fd_sc_hd__dfxbp_1_1/D 0.41fF
C4688 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C4689 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.10fF
C4690 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C4691 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.02fF
C4692 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C4693 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4694 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.10fF
C4695 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C4696 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C4697 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C4698 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VDD 0.15fF
C4699 p2d sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.06fF
C4700 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A sky130_fd_sc_hd__nand2_4_3/A 0.46fF
C4701 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.05fF
C4702 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C4703 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C4704 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C4705 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C4706 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.01fF
C4707 A_b A 0.47fF
C4708 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.05fF
C4709 sky130_fd_sc_hd__nand2_4_0/Y VSUBS -0.26fF
C4710 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.04fF
C4711 p2 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0.12fF
C4712 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_163/A -0.00fF
C4713 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.02fF
C4714 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.02fF
C4715 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C4716 VSUBS sky130_fd_sc_hd__nand2_4_3/A -0.18fF
C4717 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.01fF
C4718 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.01fF
C4719 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.01fF
C4720 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.12fF
C4721 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C4722 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__nand2_4_1/A 0.13fF
C4723 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.05fF
C4724 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.05fF
C4725 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.01fF
C4726 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C4727 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.03fF
C4728 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.03fF
C4729 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.02fF
C4730 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0.02fF
C4731 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# 0.13fF
C4732 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.00fF
C4733 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.00fF
C4734 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.00fF
C4735 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.00fF
C4736 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__nand2_4_0/Y 0.01fF
C4737 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.01fF
C4738 sky130_fd_sc_hd__clkinv_4_3/w_82_21# sky130_fd_sc_hd__nand2_4_1/Y 0.03fF
C4739 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C4740 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A sky130_fd_sc_hd__nand2_1_2/B 0.02fF
C4741 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.01fF
C4742 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.00fF
C4743 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C4744 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.03fF
C4745 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0.00fF
C4746 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C4747 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.30fF
C4748 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C4749 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.03fF
C4750 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__nand2_4_2/A 0.13fF
C4751 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.09fF
C4752 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C4753 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.01fF
C4754 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.02fF
C4755 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.01fF
C4756 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.01fF
C4757 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.01fF
C4758 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.15fF
C4759 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.01fF
C4760 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C4761 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.02fF
C4762 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__nand2_1_4/Y 0.00fF
C4763 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C4764 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.00fF
C4765 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C4766 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C4767 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__mux2_1_0/S 0.11fF
C4768 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.36fF
C4769 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.01fF
C4770 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C4771 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.02fF
C4772 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.04fF
C4773 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkinv_1_0/Y 0.00fF
C4774 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.03fF
C4775 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.08fF
C4776 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.02fF
C4777 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C4778 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C4779 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C4780 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 1.15fF
C4781 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.07fF
C4782 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A sky130_fd_sc_hd__nand2_4_1/A 0.06fF
C4783 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0.01fF
C4784 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.05fF
C4785 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.01fF
C4786 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0.01fF
C4787 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__nand2_4_1/B 0.03fF
C4788 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 1.27fF
C4789 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__clkinv_1_3/Y 0.04fF
C4790 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4791 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.19fF
C4792 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# 0.07fF
C4793 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.00fF
C4794 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.00fF
C4795 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.23fF
C4796 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.07fF
C4797 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.02fF
C4798 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.02fF
C4799 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C4800 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4801 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.02fF
C4802 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__nand2_4_0/A 1.27fF
C4803 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C4804 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C4805 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.04fF
C4806 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.03fF
C4807 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkinv_1_2/Y 0.12fF
C4808 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.16fF
C4809 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkinv_4_8/Y 0.07fF
C4810 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C4811 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.17fF
C4812 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C4813 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C4814 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0.33fF
C4815 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.02fF
C4816 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C4817 p2 sky130_fd_sc_hd__nand2_4_1/Y 0.00fF
C4818 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.01fF
C4819 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 1.32fF
C4820 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.00fF
C4821 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C4822 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.03fF
C4823 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.01fF
C4824 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.01fF
C4825 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C4826 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.01fF
C4827 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C4828 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C4829 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C4830 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C4831 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.33fF
C4832 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.02fF
C4833 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.08fF
C4834 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.18fF
C4835 sky130_fd_sc_hd__clkinv_4_7/w_82_21# sky130_fd_sc_hd__clkinv_4_7/Y -0.00fF
C4836 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.00fF
C4837 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C4838 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C4839 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.01fF
C4840 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C4841 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VDD 0.24fF
C4842 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.00fF
C4843 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.04fF
C4844 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.03fF
C4845 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X -0.00fF
C4846 sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.02fF
C4847 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C4848 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C4849 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C4850 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.13fF
C4851 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# sky130_fd_sc_hd__nand2_4_0/A 0.09fF
C4852 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C4853 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.00fF
C4854 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C4855 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C4856 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.00fF
C4857 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0.15fF
C4858 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__nand2_1_3/A 0.07fF
C4859 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_149/X -0.30fF
C4860 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0.01fF
C4861 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.01fF
C4862 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C4863 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VDD 0.15fF
C4864 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.11fF
C4865 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.02fF
C4866 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.00fF
C4867 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.04fF
C4868 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.66fF
C4869 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.02fF
C4870 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.02fF
C4871 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C4872 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VDD 0.11fF
C4873 sky130_fd_sc_hd__nand2_1_4/B sky130_fd_sc_hd__nand2_4_1/A 0.31fF
C4874 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C4875 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C4876 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Ad_b 0.03fF
C4877 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.11fF
C4878 sky130_fd_sc_hd__clkinv_4_9/Y VSUBS 0.01fF
C4879 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.04fF
C4880 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.02fF
C4881 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C4882 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.01fF
C4883 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.01fF
C4884 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.01fF
C4885 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# 0.20fF
C4886 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.01fF
C4887 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C4888 sky130_fd_sc_hd__dfxbp_1_0/Q_N Ad_b 0.01fF
C4889 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# sky130_fd_sc_hd__clkinv_1_3/Y 0.01fF
C4890 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0.00fF
C4891 VSUBS Ad_b 0.00fF
C4892 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.01fF
C4893 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.17fF
C4894 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_127/X -0.25fF
C4895 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.01fF
C4896 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.34fF
C4897 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.00fF
C4898 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.07fF
C4899 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.00fF
C4900 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C4901 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.02fF
C4902 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 2.25fF
C4903 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0.08fF
C4904 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0.34fF
C4905 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkinv_4_8/w_82_21# 0.03fF
C4906 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C4907 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.07fF
C4908 sky130_fd_sc_hd__nand2_1_0/A sky130_fd_sc_hd__nand2_4_0/A 0.21fF
C4909 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.05fF
C4910 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.05fF
C4911 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.07fF
C4912 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.02fF
C4913 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.07fF
C4914 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.02fF
C4915 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.02fF
C4916 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C4917 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C4918 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.07fF
C4919 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.18fF
C4920 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/S 0.11fF
C4921 sky130_fd_sc_hd__mux2_1_0/a_76_199# Ad_b 0.02fF
C4922 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__nand2_1_4/B 0.01fF
C4923 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.00fF
C4924 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.00fF
C4925 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.15fF
C4926 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0.03fF
C4927 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0.01fF
C4928 VDD sky130_fd_sc_hd__dfxbp_1_1/a_975_413# 0.01fF
C4929 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_592_47# 0.01fF
C4930 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.31fF
C4931 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C4932 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.04fF
C4933 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.04fF
C4934 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__nand2_1_1/B 0.69fF
C4935 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.11fF
C4936 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.00fF
C4937 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.18fF
C4938 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.13fF
C4939 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0.33fF
C4940 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C4941 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__nand2_4_0/A 0.47fF
C4942 sky130_fd_sc_hd__nand2_4_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.13fF
C4943 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.03fF
C4944 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.01fF
C4945 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.04fF
C4946 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# 0.01fF
C4947 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 1.12fF
C4948 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C4949 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.04fF
C4950 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.01fF
C4951 sky130_fd_sc_hd__mux2_1_0/S Ad_b 0.17fF
C4952 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_8/X -0.70fF
C4953 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.00fF
C4954 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.01fF
C4955 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.00fF
C4956 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.04fF
C4957 VDD sky130_fd_sc_hd__dfxbp_1_1/D 0.61fF
C4958 VSUBS sky130_fd_sc_hd__nand2_1_4/Y -0.62fF
C4959 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C4960 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.10fF
C4961 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C4962 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C4963 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.01fF
C4964 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# -0.00fF
C4965 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C4966 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C4967 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.07fF
C4968 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C4969 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.01fF
C4970 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C4971 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0.01fF
C4972 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.01fF
C4973 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C4974 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C4975 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# sky130_fd_sc_hd__nand2_1_3/A 0.00fF
C4976 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.01fF
C4977 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.08fF
C4978 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.02fF
C4979 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.11fF
C4980 sky130_fd_sc_hd__clkinv_4_2/w_82_21# sky130_fd_sc_hd__clkinv_4_2/Y 0.05fF
C4981 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__nand2_4_3/B 0.01fF
C4982 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.01fF
C4983 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.01fF
C4984 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__mux2_1_0/S 0.00fF
C4985 sky130_fd_sc_hd__nand2_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C4986 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.00fF
C4987 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C4988 sky130_fd_sc_hd__nand2_4_3/B sky130_fd_sc_hd__nand2_4_3/A 0.87fF
C4989 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.07fF
C4990 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# -0.00fF
C4991 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.05fF
C4992 p2 sky130_fd_sc_hd__clkinv_1_3/A 0.24fF
C4993 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C4994 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C4995 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.07fF
C4996 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.07fF
C4997 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.15fF
C4998 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.14fF
C4999 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.03fF
C5000 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C5001 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C5002 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.15fF
C5003 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.03fF
C5004 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.01fF
C5005 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0.01fF
C5006 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.01fF
C5007 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.01fF
C5008 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 1.06fF
C5009 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.35fF
C5010 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.15fF
C5011 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.06fF
C5012 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.09fF
C5013 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C5014 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.04fF
C5015 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.04fF
C5016 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.01fF
C5017 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C5018 sky130_fd_sc_hd__clkinv_1_3/Y sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C5019 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C5020 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C5021 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# 0.00fF
C5022 VSUBS sky130_fd_sc_hd__nand2_4_1/B -0.05fF
C5023 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.14fF
C5024 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.00fF
C5025 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C5026 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0.01fF
C5027 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0.02fF
C5028 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.00fF
C5029 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C5030 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C5031 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C5032 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0.06fF
C5033 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# sky130_fd_sc_hd__nand2_1_1/B 0.00fF
C5034 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C5035 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0.01fF
C5036 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.02fF
C5037 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.02fF
C5038 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.00fF
C5039 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# Ad_b 0.22fF
C5040 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# sky130_fd_sc_hd__nand2_4_3/A 0.06fF
C5041 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VDD 0.24fF
C5042 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.00fF
C5043 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C5044 sky130_fd_sc_hd__clkinv_4_11/w_82_21# sky130_fd_sc_hd__nand2_4_3/A -0.29fF
C5045 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C5046 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.00fF
C5047 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__nand2_1_4/Y 0.02fF
C5048 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.19fF
C5049 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.12fF
C5050 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.01fF
C5051 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.00fF
C5052 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.01fF
C5053 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0.01fF
C5054 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C5055 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.16fF
C5056 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.00fF
C5057 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.00fF
C5058 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.08fF
C5059 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.00fF
C5060 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.34fF
C5061 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.11fF
C5062 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.03fF
C5063 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0.00fF
C5064 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.19fF
C5065 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.31fF
C5066 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0.09fF
C5067 VDD sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.25fF
C5068 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.08fF
C5069 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.00fF
C5070 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.00fF
C5071 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A sky130_fd_sc_hd__nand2_4_0/A 0.01fF
C5072 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.02fF
C5073 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.01fF
C5074 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.00fF
C5075 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.01fF
C5076 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# sky130_fd_sc_hd__clkinv_1_1/Y 0.00fF
C5077 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.02fF
C5078 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.00fF
C5079 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.82fF
C5080 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.03fF
C5081 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.01fF
C5082 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.03fF
C5083 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.03fF
C5084 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.05fF
C5085 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.01fF
C5086 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C5087 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.01fF
C5088 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.01fF
C5089 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C5090 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.01fF
C5091 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.01fF
C5092 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C5093 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.03fF
C5094 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.01fF
C5095 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.01fF
C5096 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0.00fF
C5097 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.00fF
C5098 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.08fF
C5099 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.01fF
C5100 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/A -0.00fF
C5101 sky130_fd_sc_hd__nand2_1_2/A sky130_fd_sc_hd__nand2_4_2/A 0.15fF
C5102 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C5103 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.03fF
C5104 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.12fF
C5105 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0.01fF
C5106 Bd B_b 0.53fF
C5107 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.01fF
C5108 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.01fF
C5109 B B_b 0.47fF
C5110 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C5111 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.17fF
C5112 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.00fF
C5113 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0.00fF
C5114 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.07fF
C5115 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0.02fF
C5116 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# -0.00fF
C5117 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.03fF
C5118 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0.32fF
C5119 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0.01fF
C5120 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.01fF
C5121 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0.01fF
C5122 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C5123 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C5124 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.19fF
C5125 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.02fF
C5126 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.00fF
C5127 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VDD 0.17fF
C5128 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.01fF
C5129 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.02fF
C5130 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.01fF
C5131 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C5132 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A -0.00fF
C5133 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.00fF
C5134 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0.02fF
C5135 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0.02fF
C5136 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_44/X -0.00fF
C5137 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.26fF
C5138 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# sky130_fd_sc_hd__dfxbp_1_1/a_561_413# 0.01fF
C5139 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.02fF
C5140 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.01fF
C5141 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.00fF
C5142 sky130_fd_sc_hd__nand2_4_0/Y sky130_fd_sc_hd__clkinv_4_2/w_82_21# 0.03fF
C5143 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.02fF
C5144 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.01fF
C5145 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.01fF
C5146 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.02fF
C5147 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C5148 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.04fF
C5149 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.04fF
C5150 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# sky130_fd_sc_hd__clkinv_4_7/Y 0.01fF
C5151 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.00fF
C5152 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C5153 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0.01fF
C5154 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0.01fF
C5155 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# sky130_fd_sc_hd__nand2_4_2/B 0.01fF
C5156 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.38fF
C5157 sky130_fd_sc_hd__clkinv_4_7/A sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.01fF
C5158 VDD sky130_fd_sc_hd__nand2_1_0/B 1.07fF
C5159 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__nand2_4_2/a_27_47# 0.02fF
C5160 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C5161 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C5162 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C5163 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.62fF
C5164 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C5165 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.03fF
C5166 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.01fF
C5167 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.08fF
C5168 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.02fF
C5169 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C5170 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# sky130_fd_sc_hd__dfxbp_1_1/D -0.03fF
C5171 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C5172 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.03fF
C5173 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.01fF
C5174 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.00fF
C5175 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.00fF
C5176 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0.02fF
C5177 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.02fF
C5178 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.02fF
C5179 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.05fF
C5180 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.10fF
C5181 VDD sky130_fd_sc_hd__clkinv_4_1/Y 0.49fF
C5182 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.00fF
C5183 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0.00fF
C5184 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C5185 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.00fF
C5186 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.01fF
C5187 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.08fF
C5188 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.00fF
C5189 sky130_fd_sc_hd__nand2_4_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0.01fF
C5190 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.02fF
C5191 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.01fF
C5192 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0.01fF
C5193 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.31fF
C5194 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.04fF
C5195 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0.04fF
C5196 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C5197 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.01fF
C5198 sky130_fd_sc_hd__nand2_4_3/B Ad_b 0.04fF
C5199 sky130_fd_sc_hd__nand2_1_4/B clk 0.07fF
C5200 VSUBS sky130_fd_sc_hd__nand2_4_2/A -0.22fF
C5201 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C5202 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__nand2_4_2/A 0.13fF
C5203 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0.00fF
C5204 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0.00fF
C5205 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.02fF
C5206 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.00fF
C5207 p2 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.02fF
C5208 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0.01fF
C5209 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C5210 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.03fF
C5211 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A sky130_fd_sc_hd__nand2_4_2/A 0.06fF
C5212 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0.03fF
C5213 sky130_fd_sc_hd__clkinv_1_0/Y sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.05fF
C5214 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0.15fF
C5215 p2 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.03fF
C5216 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.00fF
C5217 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C5218 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.00fF
C5219 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__nand2_1_1/B 0.05fF
C5220 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__nand2_1_4/B 0.12fF
C5221 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.03fF
C5222 sky130_fd_sc_hd__nand2_4_0/B sky130_fd_sc_hd__nand2_4_0/A 1.15fF
C5223 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C5224 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.36fF
C5225 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.02fF
C5226 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# 0.09fF
C5227 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# Bd_b 0.12fF
C5228 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# sky130_fd_sc_hd__nand2_1_1/B 0.01fF
C5229 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.05fF
C5230 sky130_fd_sc_hd__clkinv_4_9/Y sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C5231 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.01fF
C5232 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# Bd_b 0.02fF
C5233 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.02fF
C5234 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.02fF
C5235 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C5236 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.04fF
C5237 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.11fF
C5238 sky130_fd_sc_hd__nand2_4_3/Y sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0.01fF
C5239 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X sky130_fd_sc_hd__nand2_1_3/A 0.09fF
C5240 sky130_fd_sc_hd__nand2_4_3/A Ad_b 0.32fF
C5241 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.01fF
C5242 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C5243 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.00fF
C5244 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__nand2_4_1/B 0.01fF
C5245 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0.00fF
C5246 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.00fF
C5247 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C5248 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.08fF
C5249 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.01fF
C5250 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.11fF
C5251 p1d_b sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.02fF
C5252 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0.03fF
C5253 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.08fF
C5254 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.08fF
C5255 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.06fF
C5256 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_3/A 0.11fF
C5257 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C5258 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.00fF
C5259 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.01fF
C5260 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.19fF
C5261 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C5262 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.00fF
C5263 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C5264 VDD sky130_fd_sc_hd__clkinv_1_3/Y 0.29fF
C5265 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.07fF
C5266 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# 0.05fF
C5267 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.00fF
C5268 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.00fF
C5269 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.03fF
C5270 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# -0.00fF
C5271 sky130_fd_sc_hd__clkinv_4_5/Y sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# 0.07fF
C5272 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.01fF
C5273 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.03fF
C5274 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.12fF
C5275 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.01fF
C5276 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.01fF
C5277 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.10fF
C5278 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.31fF
C5279 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.00fF
C5280 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.01fF
C5281 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.01fF
C5282 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0.01fF
C5283 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# sky130_fd_sc_hd__nand2_4_0/B 0.01fF
C5284 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.01fF
C5285 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.01fF
C5286 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__nand2_1_1/A 0.00fF
C5287 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.14fF
C5288 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0.00fF
C5289 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0.00fF
C5290 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C5291 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.08fF
C5292 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C5293 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C5294 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0.00fF
C5295 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0.00fF
C5296 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.17fF
C5297 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.03fF
C5298 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C5299 sky130_fd_sc_hd__nand2_4_3/A sky130_fd_sc_hd__nand2_1_4/Y 0.06fF
C5300 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.49fF
C5301 sky130_fd_sc_hd__clkinv_4_1/A sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.06fF
C5302 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_152/X -0.00fF
C5303 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C5304 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkinv_1_1/Y 0.03fF
C5305 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C5306 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C5307 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.00fF
C5308 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C5309 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.03fF
C5310 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.00fF
C5311 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.00fF
C5312 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.00fF
C5313 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.15fF
C5314 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0.01fF
C5315 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.07fF
C5316 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.02fF
C5317 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VDD 0.30fF
C5318 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.02fF
C5319 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0.02fF
C5320 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.19fF
C5321 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.00fF
C5322 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.08fF
C5323 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5324 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.02fF
C5325 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.01fF
C5326 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.01fF
C5327 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.04fF
C5328 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.04fF
C5329 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.00fF
C5330 Bd sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.12fF
C5331 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C5332 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.02fF
C5333 B sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.02fF
C5334 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.05fF
C5335 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.05fF
C5336 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.10fF
C5337 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0.31fF
C5338 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.01fF
C5339 sky130_fd_sc_hd__nand2_4_1/B sky130_fd_sc_hd__nand2_4_3/A 0.02fF
C5340 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0.02fF
C5341 VDD sky130_fd_sc_hd__clkinv_4_8/Y 1.51fF
C5342 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VDD 0.59fF
C5343 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.08fF
C5344 sky130_fd_sc_hd__nand2_4_2/Y VSUBS -0.31fF
C5345 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.01fF
C5346 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.07fF
C5347 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A Bd_b 0.03fF
C5348 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.10fF
C5349 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0.01fF
C5350 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C5351 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.03fF
C5352 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.14fF
C5353 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.02fF
C5354 sky130_fd_sc_hd__clkinv_4_10/Y sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.01fF
C5355 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 1.48fF
C5356 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# sky130_fd_sc_hd__nand2_4_0/A 0.76fF
C5357 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# 0.16fF
C5358 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0.01fF
C5359 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.08fF
C5360 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.08fF
C5361 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.11fF
C5362 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.01fF
C5363 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.00fF
C5364 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0.09fF
C5365 sky130_fd_sc_hd__dfxbp_1_0/Q_N Bd_b 0.01fF
C5366 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374# 0.01fF
C5367 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.03fF
C5368 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C5369 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C5370 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 1.12fF
C5371 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.03fF
C5372 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.01fF
C5373 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C5374 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.00fF
C5375 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0.01fF
C5376 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.00fF
C5377 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0.00fF
C5378 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.00fF
C5379 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_27_47# 0.08fF
C5380 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0.14fF
C5381 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.17fF
C5382 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.00fF
C5383 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.00fF
C5384 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.34fF
C5385 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.21fF
C5386 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.01fF
C5387 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C5388 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0.00fF
C5389 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.00fF
C5390 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.00fF
C5391 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.21fF
C5392 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.02fF
C5393 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.01fF
C5394 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.01fF
C5395 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.01fF
C5396 sky130_fd_sc_hd__nand2_4_3/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0.05fF
C5397 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0.01fF
C5398 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.01fF
C5399 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.01fF
C5400 sky130_fd_sc_hd__nand2_4_2/Y sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.05fF
C5401 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.08fF
C5402 sky130_fd_sc_hd__mux2_1_0/a_76_199# Bd_b 0.02fF
C5403 sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__mux2_1_0/S 0.01fF
C5404 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.01fF
C5405 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.01fF
C5406 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.01fF
C5407 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__clkinv_4_4/Y 0.14fF
C5408 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.14fF
C5409 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A sky130_fd_sc_hd__nand2_1_2/B 0.02fF
C5410 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# 0.10fF
C5411 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.00fF
C5412 sky130_fd_sc_hd__nand2_1_1/A sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# 0.01fF
C5413 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.01fF
C5414 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.15fF
C5415 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.01fF
C5416 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.02fF
C5417 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0.01fF
C5418 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.01fF
C5419 VDD sky130_fd_sc_hd__nand2_1_1/B 1.42fF
C5420 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C5421 sky130_fd_sc_hd__clkinv_1_3/A sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.06fF
C5422 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.16fF
C5423 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.04fF
C5424 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.04fF
C5425 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0.02fF
C5426 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.01fF
C5427 VDD sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0.30fF
C5428 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.00fF
C5429 clk VSS 17.23fF
C5430 p1d VSS 14.97fF
C5431 sky130_fd_sc_hd__clkbuf_16_10/a_110_47# VSS 1.46fF
C5432 sky130_fd_sc_hd__nand2_1_0/B VSS 20.35fF
C5433 sky130_fd_sc_hd__nand2_1_4/Y VSS 34.81fF
C5434 Bd_b VSS 36.76fF
C5435 Ad_b VSS 11.76fF
C5436 sky130_fd_sc_hd__mux2_1_0/S VSS 10.43fF
C5437 sky130_fd_sc_hd__mux2_1_0/a_439_47# VSS 0.01fF
C5438 sky130_fd_sc_hd__mux2_1_0/a_218_47# VSS 0.01fF
C5439 sky130_fd_sc_hd__mux2_1_0/a_505_21# VSS 0.30fF
C5440 sky130_fd_sc_hd__mux2_1_0/a_76_199# VSS 0.29fF
C5441 sky130_fd_sc_hd__mux2_1_0/X VSS 43.23fF
C5442 sky130_fd_sc_hd__nand2_1_4/a_113_47# VSS 0.01fF
C5443 sky130_fd_sc_hd__clkinv_1_2/Y VSS 25.04fF
C5444 sky130_fd_sc_hd__nand2_4_3/A VSS 26.29fF
C5445 sky130_fd_sc_hd__nand2_1_3/A VSS 19.61fF
C5446 sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS -0.00fF
C5447 sky130_fd_sc_hd__clkdlybuf4s50_1_112/X VSS 9.23fF
C5448 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# VSS 0.21fF
C5449 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# VSS 0.27fF
C5450 sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# VSS 0.37fF
C5451 sky130_fd_sc_hd__clkinv_1_1/Y VSS 32.90fF
C5452 sky130_fd_sc_hd__nand2_4_2/A VSS 17.61fF
C5453 sky130_fd_sc_hd__nand2_1_2/A VSS 10.61fF
C5454 sky130_fd_sc_hd__nand2_1_2/B VSS 11.61fF
C5455 sky130_fd_sc_hd__clkdlybuf4s50_1_109/X VSS 9.33fF
C5456 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# VSS 0.20fF
C5457 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# VSS 0.28fF
C5458 sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# VSS 0.38fF
C5459 sky130_fd_sc_hd__clkdlybuf4s50_1_31/A VSS 25.89fF
C5460 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# VSS 0.20fF
C5461 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# VSS 0.27fF
C5462 sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# VSS 0.42fF
C5463 sky130_fd_sc_hd__clkdlybuf4s50_1_20/A VSS 24.24fF
C5464 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# VSS 0.20fF
C5465 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# VSS 0.27fF
C5466 sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# VSS 0.41fF
C5467 p1_b VSS 15.64fF
C5468 sky130_fd_sc_hd__clkinv_4_7/Y VSS 28.94fF
C5469 sky130_fd_sc_hd__clkbuf_16_9/a_110_47# VSS 1.58fF
C5470 sky130_fd_sc_hd__nand2_4_1/A VSS 26.18fF
C5471 sky130_fd_sc_hd__nand2_1_1/B VSS 13.67fF
C5472 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.01fF
C5473 sky130_fd_sc_hd__clkdlybuf4s50_1_131/X VSS 20.94fF
C5474 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# VSS 0.21fF
C5475 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# VSS 0.28fF
C5476 sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# VSS 0.39fF
C5477 sky130_fd_sc_hd__clkdlybuf4s50_1_121/A VSS 24.15fF
C5478 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# VSS 0.21fF
C5479 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# VSS 0.29fF
C5480 sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# VSS 0.43fF
C5481 sky130_fd_sc_hd__clkdlybuf4s50_1_108/X VSS 12.28fF
C5482 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# VSS 0.20fF
C5483 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# VSS 0.28fF
C5484 sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# VSS 0.37fF
C5485 sky130_fd_sc_hd__clkdlybuf4s50_1_49/A VSS 28.20fF
C5486 sky130_fd_sc_hd__clkdlybuf4s50_1_39/A VSS 44.62fF
C5487 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# VSS 0.22fF
C5488 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# VSS 0.30fF
C5489 sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# VSS 0.40fF
C5490 sky130_fd_sc_hd__clkdlybuf4s50_1_24/X VSS 14.40fF
C5491 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# VSS 0.22fF
C5492 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# VSS 0.27fF
C5493 sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# VSS 0.36fF
C5494 p1 VSS 7.25fF
C5495 sky130_fd_sc_hd__clkbuf_16_8/a_110_47# VSS 1.41fF
C5496 sky130_fd_sc_hd__nand2_4_0/A VSS 22.99fF
C5497 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS -0.00fF
C5498 sky130_fd_sc_hd__clkdlybuf4s50_1_118/A VSS 21.61fF
C5499 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# VSS 0.22fF
C5500 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# VSS 0.29fF
C5501 sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# VSS 0.42fF
C5502 sky130_fd_sc_hd__clkdlybuf4s50_1_38/A VSS 23.36fF
C5503 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# VSS 0.22fF
C5504 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# VSS 0.27fF
C5505 sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# VSS 0.36fF
C5506 sky130_fd_sc_hd__clkdlybuf4s50_1_29/A VSS 21.64fF
C5507 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# VSS 0.21fF
C5508 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# VSS 0.27fF
C5509 sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# VSS 0.41fF
C5510 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# VSS 0.23fF
C5511 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# VSS 0.35fF
C5512 sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# VSS 0.81fF
C5513 A VSS 28.24fF
C5514 sky130_fd_sc_hd__clkbuf_16_7/a_110_47# VSS 1.45fF
C5515 sky130_fd_sc_hd__clkdlybuf4s50_1_152/X VSS 14.41fF
C5516 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# VSS 0.23fF
C5517 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# VSS 0.31fF
C5518 sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# VSS 0.41fF
C5519 sky130_fd_sc_hd__clkdlybuf4s50_1_140/A VSS 25.87fF
C5520 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# VSS 0.21fF
C5521 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# VSS 0.29fF
C5522 sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# VSS 0.43fF
C5523 sky130_fd_sc_hd__clkdlybuf4s50_1_129/X VSS 21.30fF
C5524 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# VSS 0.21fF
C5525 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# VSS 0.29fF
C5526 sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# VSS 0.40fF
C5527 sky130_fd_sc_hd__clkdlybuf4s50_1_117/A VSS 15.49fF
C5528 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# VSS 0.21fF
C5529 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# VSS 0.29fF
C5530 sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# VSS 0.42fF
C5531 sky130_fd_sc_hd__clkdlybuf4s50_1_61/A VSS 21.27fF
C5532 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# VSS 0.21fF
C5533 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# VSS 0.29fF
C5534 sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# VSS 0.41fF
C5535 sky130_fd_sc_hd__clkdlybuf4s50_1_48/A VSS 24.27fF
C5536 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# VSS 0.21fF
C5537 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# VSS 0.30fF
C5538 sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# VSS 0.40fF
C5539 sky130_fd_sc_hd__clkdlybuf4s50_1_17/X VSS 20.79fF
C5540 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# VSS 0.23fF
C5541 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# VSS 0.30fF
C5542 sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# VSS 0.40fF
C5543 A_b VSS 15.73fF
C5544 sky130_fd_sc_hd__clkinv_4_4/Y VSS 28.94fF
C5545 sky130_fd_sc_hd__clkbuf_16_6/a_110_47# VSS 1.58fF
C5546 sky130_fd_sc_hd__clkdlybuf4s50_1_162/A VSS 43.46fF
C5547 sky130_fd_sc_hd__clkdlybuf4s50_1_168/X VSS 23.70fF
C5548 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# VSS 0.21fF
C5549 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# VSS 0.27fF
C5550 sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# VSS 0.41fF
C5551 sky130_fd_sc_hd__clkdlybuf4s50_1_113/A VSS 11.05fF
C5552 sky130_fd_sc_hd__clkdlybuf4s50_1_107/X VSS 5.52fF
C5553 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# VSS 0.21fF
C5554 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# VSS 0.29fF
C5555 sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# VSS 0.38fF
C5556 sky130_fd_sc_hd__clkdlybuf4s50_1_69/X VSS 14.27fF
C5557 sky130_fd_sc_hd__clkdlybuf4s50_1_71/X VSS 25.25fF
C5558 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# VSS 0.20fF
C5559 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# VSS 0.28fF
C5560 sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# VSS 0.39fF
C5561 sky130_fd_sc_hd__clkdlybuf4s50_1_38/X VSS 41.35fF
C5562 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# VSS 0.23fF
C5563 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# VSS 0.30fF
C5564 sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# VSS 0.40fF
C5565 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# VSS 0.21fF
C5566 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# VSS 0.26fF
C5567 sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# VSS 0.35fF
C5568 sky130_fd_sc_hd__clkdlybuf4s50_1_47/X VSS 22.13fF
C5569 sky130_fd_sc_hd__clkdlybuf4s50_1_48/X VSS 14.28fF
C5570 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# VSS 0.21fF
C5571 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# VSS 0.27fF
C5572 sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# VSS 0.41fF
C5573 sky130_fd_sc_hd__clkdlybuf4s50_1_27/A VSS 22.79fF
C5574 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# VSS 0.20fF
C5575 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# VSS 0.27fF
C5576 sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# VSS 0.41fF
C5577 Ad VSS 12.34fF
C5578 sky130_fd_sc_hd__clkbuf_16_5/a_110_47# VSS 1.46fF
C5579 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# VSS 0.21fF
C5580 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# VSS 0.26fF
C5581 sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# VSS 0.35fF
C5582 sky130_fd_sc_hd__clkdlybuf4s50_1_150/X VSS 43.41fF
C5583 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# VSS 0.21fF
C5584 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# VSS 0.28fF
C5585 sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# VSS 0.39fF
C5586 sky130_fd_sc_hd__clkdlybuf4s50_1_138/A VSS 21.62fF
C5587 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# VSS 0.22fF
C5588 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# VSS 0.29fF
C5589 sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# VSS 0.42fF
C5590 sky130_fd_sc_hd__clkdlybuf4s50_1_127/X VSS 11.42fF
C5591 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# VSS 0.21fF
C5592 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# VSS 0.28fF
C5593 sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# VSS 0.39fF
C5594 sky130_fd_sc_hd__nand2_4_2/B VSS 55.18fF
C5595 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# VSS 0.19fF
C5596 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# VSS 0.26fF
C5597 sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# VSS 0.38fF
C5598 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# VSS 0.23fF
C5599 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# VSS 0.35fF
C5600 sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# VSS 0.81fF
C5601 sky130_fd_sc_hd__nand2_1_0/A VSS 15.18fF
C5602 sky130_fd_sc_hd__clkdlybuf4s50_1_68/A VSS 23.05fF
C5603 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# VSS 0.22fF
C5604 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# VSS 0.35fF
C5605 sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# VSS 0.82fF
C5606 sky130_fd_sc_hd__clkdlybuf4s50_1_15/X VSS 21.13fF
C5607 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# VSS 0.23fF
C5608 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# VSS 0.31fF
C5609 sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# VSS 0.41fF
C5610 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# VSS 0.18fF
C5611 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# VSS 0.26fF
C5612 sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# VSS 0.40fF
C5613 sky130_fd_sc_hd__clkbuf_16_4/a_110_47# VSS 1.64fF
C5614 sky130_fd_sc_hd__clkdlybuf4s50_1_172/X VSS 24.27fF
C5615 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# VSS 0.21fF
C5616 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# VSS 0.30fF
C5617 sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# VSS 0.40fF
C5618 sky130_fd_sc_hd__clkdlybuf4s50_1_149/X VSS 26.31fF
C5619 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# VSS 0.22fF
C5620 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# VSS 0.30fF
C5621 sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# VSS 0.40fF
C5622 sky130_fd_sc_hd__clkdlybuf4s50_1_116/A VSS 21.26fF
C5623 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# VSS 0.21fF
C5624 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# VSS 0.29fF
C5625 sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# VSS 0.41fF
C5626 sky130_fd_sc_hd__clkdlybuf4s50_1_103/A VSS 18.11fF
C5627 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# VSS 0.19fF
C5628 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# VSS 0.25fF
C5629 sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# VSS 0.37fF
C5630 sky130_fd_sc_hd__clkdlybuf4s50_1_167/X VSS 19.93fF
C5631 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# VSS 0.22fF
C5632 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# VSS 0.27fF
C5633 sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# VSS 0.36fF
C5634 sky130_fd_sc_hd__clkdlybuf4s50_1_93/A VSS 12.29fF
C5635 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# VSS 0.22fF
C5636 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# VSS 0.35fF
C5637 sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# VSS 0.57fF
C5638 sky130_fd_sc_hd__clkdlybuf4s50_1_80/A VSS 21.27fF
C5639 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# VSS 0.22fF
C5640 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# VSS 0.29fF
C5641 sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# VSS 0.42fF
C5642 sky130_fd_sc_hd__clkdlybuf4s50_1_67/X VSS 14.36fF
C5643 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# VSS 0.19fF
C5644 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# VSS 0.27fF
C5645 sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# VSS 0.41fF
C5646 sky130_fd_sc_hd__clkdlybuf4s50_1_36/X VSS 27.69fF
C5647 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# VSS 0.23fF
C5648 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# VSS 0.31fF
C5649 sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# VSS 0.41fF
C5650 sky130_fd_sc_hd__clkdlybuf4s50_1_58/X VSS 21.39fF
C5651 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# VSS 0.22fF
C5652 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# VSS 0.29fF
C5653 sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# VSS 0.39fF
C5654 sky130_fd_sc_hd__clkinv_4_2/Y VSS 38.86fF
C5655 sky130_fd_sc_hd__clkbuf_16_3/a_110_47# VSS 1.56fF
C5656 sky130_fd_sc_hd__clkdlybuf4s50_1_136/A VSS 22.77fF
C5657 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# VSS 0.21fF
C5658 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# VSS 0.29fF
C5659 sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# VSS 0.42fF
C5660 sky130_fd_sc_hd__clkdlybuf4s50_1_132/A VSS 14.27fF
C5661 sky130_fd_sc_hd__clkdlybuf4s50_1_125/X VSS 25.25fF
C5662 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# VSS 0.20fF
C5663 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# VSS 0.28fF
C5664 sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# VSS 0.39fF
C5665 sky130_fd_sc_hd__clkdlybuf4s50_1_102/A VSS 19.57fF
C5666 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# VSS 0.19fF
C5667 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# VSS 0.26fF
C5668 sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# VSS 0.38fF
C5669 sky130_fd_sc_hd__clkinv_4_8/Y VSS 11.48fF
C5670 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# VSS 0.19fF
C5671 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# VSS 0.24fF
C5672 sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# VSS 0.32fF
C5673 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# VSS 0.18fF
C5674 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# VSS 0.26fF
C5675 sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# VSS 0.40fF
C5676 sky130_fd_sc_hd__clkdlybuf4s50_1_180/A VSS 22.12fF
C5677 sky130_fd_sc_hd__clkdlybuf4s50_1_187/X VSS 20.13fF
C5678 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# VSS 0.21fF
C5679 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# VSS 0.28fF
C5680 sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# VSS 0.41fF
C5681 sky130_fd_sc_hd__clkinv_4_3/Y VSS 43.40fF
C5682 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# VSS 0.20fF
C5683 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# VSS 0.24fF
C5684 sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# VSS 0.33fF
C5685 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# VSS 0.20fF
C5686 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# VSS 0.25fF
C5687 sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# VSS 0.34fF
C5688 sky130_fd_sc_hd__clkdlybuf4s50_1_13/X VSS 11.31fF
C5689 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# VSS 0.22fF
C5690 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# VSS 0.30fF
C5691 sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# VSS 0.40fF
C5692 sky130_fd_sc_hd__clkdlybuf4s50_1_44/X VSS 36.82fF
C5693 sky130_fd_sc_hd__clkdlybuf4s50_1_44/A VSS 20.30fF
C5694 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# VSS 0.21fF
C5695 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# VSS 0.28fF
C5696 sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# VSS 0.41fF
C5697 sky130_fd_sc_hd__clkdlybuf4s50_1_24/A VSS 38.72fF
C5698 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# VSS 0.20fF
C5699 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# VSS 0.27fF
C5700 sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# VSS 0.42fF
C5701 B_b VSS 21.34fF
C5702 sky130_fd_sc_hd__clkinv_4_1/Y VSS 58.18fF
C5703 sky130_fd_sc_hd__clkbuf_16_2/a_110_47# VSS 1.52fF
C5704 sky130_fd_sc_hd__nand2_1_4/B VSS 40.85fF
C5705 sky130_fd_sc_hd__clkdlybuf4s50_1_142/X VSS 23.05fF
C5706 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# VSS 0.22fF
C5707 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# VSS 0.33fF
C5708 sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# VSS 0.80fF
C5709 sky130_fd_sc_hd__clkdlybuf4s50_1_101/A VSS 8.39fF
C5710 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# VSS 0.20fF
C5711 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# VSS 0.27fF
C5712 sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# VSS 0.49fF
C5713 sky130_fd_sc_hd__clkdlybuf4s50_1_186/X VSS 14.39fF
C5714 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# VSS 0.22fF
C5715 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# VSS 0.27fF
C5716 sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# VSS 0.36fF
C5717 sky130_fd_sc_hd__nand2_4_3/B VSS 73.02fF
C5718 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# VSS 0.20fF
C5719 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# VSS 0.27fF
C5720 sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# VSS 0.40fF
C5721 sky130_fd_sc_hd__clkdlybuf4s50_1_87/X VSS 19.82fF
C5722 sky130_fd_sc_hd__clkdlybuf4s50_1_90/X VSS 20.12fF
C5723 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# VSS 0.22fF
C5724 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# VSS 0.30fF
C5725 sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# VSS 0.41fF
C5726 sky130_fd_sc_hd__clkdlybuf4s50_1_67/A VSS 25.87fF
C5727 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# VSS 0.21fF
C5728 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# VSS 0.29fF
C5729 sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# VSS 0.43fF
C5730 sky130_fd_sc_hd__clkdlybuf4s50_1_34/X VSS 50.92fF
C5731 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# VSS 0.22fF
C5732 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# VSS 0.30fF
C5733 sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# VSS 0.40fF
C5734 sky130_fd_sc_hd__clkdlybuf4s50_1_56/X VSS 14.39fF
C5735 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# VSS 0.21fF
C5736 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# VSS 0.29fF
C5737 sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# VSS 0.40fF
C5738 sky130_fd_sc_hd__clkdlybuf4s50_1_8/X VSS 26.56fF
C5739 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# VSS 0.22fF
C5740 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# VSS 0.31fF
C5741 sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# VSS 0.39fF
C5742 Bd VSS 15.05fF
C5743 sky130_fd_sc_hd__clkbuf_16_1/a_110_47# VSS 1.51fF
C5744 sky130_fd_sc_hd__clkdlybuf4s50_1_158/X VSS 35.62fF
C5745 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# VSS 0.22fF
C5746 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# VSS 0.29fF
C5747 sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# VSS 0.39fF
C5748 sky130_fd_sc_hd__clkdlybuf4s50_1_134/A VSS 21.27fF
C5749 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# VSS 0.21fF
C5750 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# VSS 0.29fF
C5751 sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# VSS 0.41fF
C5752 sky130_fd_sc_hd__clkdlybuf4s50_1_131/A VSS 14.44fF
C5753 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# VSS 0.19fF
C5754 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# VSS 0.27fF
C5755 sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# VSS 0.41fF
C5756 sky130_fd_sc_hd__clkdlybuf4s50_1_190/X VSS 14.05fF
C5757 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# VSS 0.23fF
C5758 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# VSS 0.31fF
C5759 sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# VSS 0.42fF
C5760 sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VSS 24.15fF
C5761 sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VSS 25.83fF
C5762 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VSS 0.22fF
C5763 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VSS 0.31fF
C5764 sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VSS 0.45fF
C5765 sky130_fd_sc_hd__nand2_4_1/B VSS 72.99fF
C5766 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# VSS 0.21fF
C5767 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# VSS 0.29fF
C5768 sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# VSS 0.41fF
C5769 sky130_fd_sc_hd__clkdlybuf4s50_1_86/X VSS 14.41fF
C5770 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# VSS 0.19fF
C5771 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# VSS 0.27fF
C5772 sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# VSS 0.41fF
C5773 sky130_fd_sc_hd__clkdlybuf4s50_1_77/X VSS 20.94fF
C5774 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# VSS 0.21fF
C5775 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# VSS 0.28fF
C5776 sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# VSS 0.39fF
C5777 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# VSS 0.18fF
C5778 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# VSS 0.26fF
C5779 sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# VSS 0.40fF
C5780 sky130_fd_sc_hd__clkdlybuf4s50_1_22/A VSS 36.43fF
C5781 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# VSS 0.21fF
C5782 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# VSS 0.27fF
C5783 sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# VSS 0.41fF
C5784 sky130_fd_sc_hd__clkdlybuf4s50_1_42/A VSS 10.02fF
C5785 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# VSS 0.22fF
C5786 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# VSS 0.31fF
C5787 sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# VSS 0.40fF
C5788 B VSS 14.98fF
C5789 sky130_fd_sc_hd__clkbuf_16_0/a_110_47# VSS 1.49fF
C5790 sky130_fd_sc_hd__clkdlybuf4s50_1_147/X VSS 38.89fF
C5791 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# VSS 0.21fF
C5792 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# VSS 0.29fF
C5793 sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# VSS 0.40fF
C5794 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# VSS 0.20fF
C5795 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# VSS 0.25fF
C5796 sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# VSS 0.34fF
C5797 sky130_fd_sc_hd__clkdlybuf4s50_1_167/A VSS 50.91fF
C5798 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# VSS 0.20fF
C5799 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# VSS 0.27fF
C5800 sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# VSS 0.42fF
C5801 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# VSS 0.18fF
C5802 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# VSS 0.26fF
C5803 sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# VSS 0.40fF
C5804 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# VSS 0.20fF
C5805 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# VSS 0.28fF
C5806 sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# VSS 0.40fF
C5807 sky130_fd_sc_hd__clkdlybuf4s50_1_99/X VSS 41.22fF
C5808 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# VSS 0.22fF
C5809 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# VSS 0.29fF
C5810 sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# VSS 0.39fF
C5811 sky130_fd_sc_hd__clkdlybuf4s50_1_65/A VSS 21.62fF
C5812 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# VSS 0.22fF
C5813 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# VSS 0.29fF
C5814 sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# VSS 0.42fF
C5815 sky130_fd_sc_hd__clkdlybuf4s50_1_54/X VSS 26.29fF
C5816 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# VSS 0.21fF
C5817 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# VSS 0.28fF
C5818 sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# VSS 0.39fF
C5819 sky130_fd_sc_hd__clkdlybuf4s50_1_164/A VSS 43.38fF
C5820 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# VSS 0.21fF
C5821 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# VSS 0.27fF
C5822 sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# VSS 0.41fF
C5823 sky130_fd_sc_hd__clkdlybuf4s50_1_157/X VSS 20.96fF
C5824 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# VSS 0.23fF
C5825 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# VSS 0.30fF
C5826 sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# VSS 0.40fF
C5827 sky130_fd_sc_hd__clkdlybuf4s50_1_177/X VSS 20.79fF
C5828 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# VSS 0.23fF
C5829 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# VSS 0.30fF
C5830 sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# VSS 0.40fF
C5831 sky130_fd_sc_hd__clkdlybuf4s50_1_197/A VSS 12.67fF
C5832 sky130_fd_sc_hd__clkinv_1_3/Y VSS 32.97fF
C5833 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# VSS 0.20fF
C5834 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# VSS 0.28fF
C5835 sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# VSS 0.53fF
C5836 sky130_fd_sc_hd__clkdlybuf4s50_1_169/A VSS 22.84fF
C5837 sky130_fd_sc_hd__clkdlybuf4s50_1_146/X VSS 22.22fF
C5838 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# VSS 0.22fF
C5839 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# VSS 0.30fF
C5840 sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# VSS 0.40fF
C5841 sky130_fd_sc_hd__clkdlybuf4s50_1_97/A VSS 24.09fF
C5842 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# VSS 0.23fF
C5843 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# VSS 0.32fF
C5844 sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# VSS 0.45fF
C5845 sky130_fd_sc_hd__clkdlybuf4s50_1_86/A VSS 24.16fF
C5846 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# VSS 0.22fF
C5847 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# VSS 0.30fF
C5848 sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# VSS 0.44fF
C5849 sky130_fd_sc_hd__clkdlybuf4s50_1_75/X VSS 21.30fF
C5850 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# VSS 0.21fF
C5851 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# VSS 0.29fF
C5852 sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# VSS 0.40fF
C5853 sky130_fd_sc_hd__clkdlybuf4s50_1_163/A VSS 44.28fF
C5854 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# VSS 0.20fF
C5855 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# VSS 0.27fF
C5856 sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# VSS 0.41fF
C5857 sky130_fd_sc_hd__clkdlybuf4s50_1_158/A VSS 20.42fF
C5858 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# VSS 0.19fF
C5859 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# VSS 0.27fF
C5860 sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# VSS 0.41fF
C5861 sky130_fd_sc_hd__clkdlybuf4s50_1_174/X VSS 21.13fF
C5862 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# VSS 0.23fF
C5863 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# VSS 0.31fF
C5864 sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# VSS 0.41fF
C5865 sky130_fd_sc_hd__clkdlybuf4s50_1_186/A VSS 24.13fF
C5866 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# VSS 0.21fF
C5867 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# VSS 0.28fF
C5868 sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# VSS 0.42fF
C5869 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# VSS 0.22fF
C5870 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# VSS 0.27fF
C5871 sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# VSS 0.36fF
C5872 sky130_fd_sc_hd__dfxbp_1_1/D VSS 8.30fF
C5873 sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# VSS -0.00fF
C5874 sky130_fd_sc_hd__dfxbp_1_1/a_592_47# VSS -0.00fF
C5875 sky130_fd_sc_hd__dfxbp_1_1/a_381_47# VSS 0.05fF
C5876 sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# VSS 0.16fF
C5877 sky130_fd_sc_hd__dfxbp_1_1/a_891_413# VSS 0.19fF
C5878 sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# VSS 0.36fF
C5879 sky130_fd_sc_hd__dfxbp_1_1/a_466_413# VSS 0.16fF
C5880 sky130_fd_sc_hd__dfxbp_1_1/a_634_159# VSS 0.04fF
C5881 sky130_fd_sc_hd__dfxbp_1_1/a_193_47# VSS 0.33fF
C5882 sky130_fd_sc_hd__dfxbp_1_1/a_27_47# VSS 0.53fF
C5883 sky130_fd_sc_hd__clkdlybuf4s50_1_63/A VSS 22.77fF
C5884 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# VSS 0.21fF
C5885 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# VSS 0.29fF
C5886 sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# VSS 0.42fF
C5887 sky130_fd_sc_hd__clkdlybuf4s50_1_52/X VSS 23.85fF
C5888 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# VSS 0.21fF
C5889 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# VSS 0.29fF
C5890 sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# VSS 0.40fF
C5891 sky130_fd_sc_hd__clkdlybuf4s50_1_154/X VSS 23.27fF
C5892 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# VSS 0.21fF
C5893 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# VSS 0.29fF
C5894 sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# VSS 0.40fF
C5895 sky130_fd_sc_hd__clkdlybuf4s50_1_173/X VSS 11.31fF
C5896 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# VSS 0.22fF
C5897 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# VSS 0.30fF
C5898 sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# VSS 0.40fF
C5899 sky130_fd_sc_hd__dfxbp_1_0/Q_N VSS 0.22fF
C5900 sky130_fd_sc_hd__nand2_1_1/A VSS 49.47fF
C5901 sky130_fd_sc_hd__dfxbp_1_0/a_1017_47# VSS 0.22fF
C5902 sky130_fd_sc_hd__dfxbp_1_0/a_592_47# VSS 0.01fF
C5903 sky130_fd_sc_hd__dfxbp_1_0/a_381_47# VSS 0.08fF
C5904 sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# VSS 0.16fF
C5905 sky130_fd_sc_hd__dfxbp_1_0/a_891_413# VSS 0.21fF
C5906 sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# VSS 0.36fF
C5907 sky130_fd_sc_hd__dfxbp_1_0/a_466_413# VSS 0.19fF
C5908 sky130_fd_sc_hd__dfxbp_1_0/a_634_159# VSS 0.20fF
C5909 sky130_fd_sc_hd__dfxbp_1_0/a_193_47# VSS 0.38fF
C5910 sky130_fd_sc_hd__dfxbp_1_0/a_27_47# VSS 0.57fF
C5911 sky130_fd_sc_hd__clkdlybuf4s50_1_95/A VSS 25.77fF
C5912 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# VSS 0.23fF
C5913 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# VSS 0.33fF
C5914 sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# VSS 0.45fF
C5915 sky130_fd_sc_hd__clkdlybuf4s50_1_84/A VSS 21.62fF
C5916 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# VSS 0.22fF
C5917 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# VSS 0.30fF
C5918 sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# VSS 0.43fF
C5919 sky130_fd_sc_hd__clkdlybuf4s50_1_73/X VSS 11.42fF
C5920 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# VSS 0.21fF
C5921 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# VSS 0.28fF
C5922 sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# VSS 0.39fF
C5923 sky130_fd_sc_hd__clkdlybuf4s50_1_184/A VSS 21.57fF
C5924 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# VSS 0.21fF
C5925 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# VSS 0.28fF
C5926 sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# VSS 0.42fF
C5927 sky130_fd_sc_hd__clkdlybuf4s50_1_195/X VSS 35.17fF
C5928 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# VSS 0.24fF
C5929 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# VSS 0.31fF
C5930 sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# VSS 0.41fF
C5931 sky130_fd_sc_hd__nand2_4_3/Y VSS 112.88fF
C5932 sky130_fd_sc_hd__clkinv_4_9/w_82_21# VSS 0.00fF
C5933 sky130_fd_sc_hd__clkdlybuf4s50_1_96/X VSS 42.03fF
C5934 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# VSS 0.21fF
C5935 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# VSS 0.29fF
C5936 sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# VSS 0.39fF
C5937 sky130_fd_sc_hd__clkinv_4_8/w_82_21# VSS 0.01fF
C5938 VDD VSS -38063.93fF
C5939 VSUBS VSS 14.41fF
C5940 sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VSS 15.50fF
C5941 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VSS 0.22fF
C5942 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VSS 0.29fF
C5943 sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VSS 0.42fF
C5944 sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VSS 15.51fF
C5945 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VSS 0.20fF
C5946 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VSS 0.27fF
C5947 sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VSS 0.41fF
C5948 sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VSS 35.90fF
C5949 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VSS 0.23fF
C5950 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VSS 0.31fF
C5951 sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VSS 0.41fF
C5952 sky130_fd_sc_hd__clkinv_4_7/w_82_21# VSS 0.01fF
C5953 sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VSS 51.45fF
C5954 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VSS 0.21fF
C5955 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VSS 0.29fF
C5956 sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VSS 0.39fF
C5957 sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VSS 43.41fF
C5958 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VSS 0.23fF
C5959 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VSS 0.31fF
C5960 sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VSS 0.41fF
C5961 sky130_fd_sc_hd__clkinv_4_7/A VSS 79.83fF
C5962 sky130_fd_sc_hd__clkinv_4_6/w_82_21# VSS 0.00fF
C5963 sky130_fd_sc_hd__clkinv_4_5/Y VSS 118.80fF
C5964 sky130_fd_sc_hd__clkinv_4_5/w_82_21# VSS 0.01fF
C5965 sky130_fd_sc_hd__clkinv_4_4/w_82_21# VSS 0.01fF
C5966 sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VSS 21.27fF
C5967 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VSS 0.22fF
C5968 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VSS 0.31fF
C5969 sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VSS 0.41fF
C5970 sky130_fd_sc_hd__clkinv_4_3/w_82_21# VSS 0.01fF
C5971 sky130_fd_sc_hd__nand2_4_0/Y VSS 65.47fF
C5972 sky130_fd_sc_hd__clkinv_4_2/w_82_21# VSS 0.00fF
C5973 sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VSS 20.83fF
C5974 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VSS 0.22fF
C5975 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# VSS 0.30fF
C5976 sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VSS 0.39fF
C5977 sky130_fd_sc_hd__nand2_4_3/a_27_47# VSS 0.38fF
C5978 sky130_fd_sc_hd__clkinv_4_1/A VSS 127.69fF
C5979 sky130_fd_sc_hd__clkinv_4_1/w_82_21# VSS -0.03fF
C5980 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VSS 0.21fF
C5981 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VSS 0.27fF
C5982 sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# VSS 0.35fF
C5983 sky130_fd_sc_hd__nand2_4_2/Y VSS 64.92fF
C5984 sky130_fd_sc_hd__nand2_4_2/a_27_47# VSS 0.35fF
C5985 sky130_fd_sc_hd__clkinv_4_0/w_82_21# VSS -0.00fF
C5986 sky130_fd_sc_hd__nand2_4_1/Y VSS 67.41fF
C5987 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.40fF
C5988 sky130_fd_sc_hd__nand2_4_0/B VSS 72.96fF
C5989 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VSS 0.19fF
C5990 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VSS 0.27fF
C5991 sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VSS 0.39fF
C5992 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.35fF
C5993 sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VSS 24.11fF
C5994 sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VSS 25.78fF
C5995 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VSS 0.19fF
C5996 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VSS 0.25fF
C5997 sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VSS 0.38fF
C5998 sky130_fd_sc_hd__clkinv_4_11/w_82_21# VSS -0.00fF
C5999 p2 VSS 59.01fF
C6000 sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VSS 1.52fF
C6001 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VSS 0.19fF
C6002 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VSS 0.27fF
C6003 sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VSS 0.39fF
C6004 sky130_fd_sc_hd__clkinv_1_3/A VSS 101.10fF
C6005 sky130_fd_sc_hd__clkinv_4_10/w_82_21# VSS 0.00fF
C6006 p2_b VSS 15.65fF
C6007 sky130_fd_sc_hd__clkinv_4_10/Y VSS 29.02fF
C6008 sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VSS 1.52fF
C6009 sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VSS 12.53fF
C6010 sky130_fd_sc_hd__clkinv_1_0/Y VSS 32.90fF
C6011 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VSS 0.19fF
C6012 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VSS 0.27fF
C6013 sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VSS 0.49fF
C6014 p2d VSS 15.07fF
C6015 sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VSS 1.51fF
C6016 p2d_b VSS 23.55fF
C6017 sky130_fd_sc_hd__clkinv_4_9/Y VSS 75.37fF
C6018 sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VSS 1.57fF
C6019 p1d_b VSS 12.85fF
C6020 sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VSS 1.63fF
.ends

.subckt sky130_fd_pr__nfet_01v8_E56BNL_AA a_n72_n90# a_16_n90# a_n32_32# VSUBS
X0 a_16_n90# a_n32_32# a_n72_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=150000u
C0 a_n32_32# a_n72_n90# 0.01fF
C1 a_16_n90# a_n72_n90# 0.14fF
C2 a_16_n90# a_n32_32# 0.01fF
C3 a_16_n90# VSUBS 0.02fF
C4 a_n72_n90# VSUBS 0.02fF
C5 a_n32_32# VSUBS 0.15fF
.ends

.subckt switch_5t_AA out en_b transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD in en VSS transmission_gate_1/in
Xtransmission_gate_0 en VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in transmission_gate_1/in VSS en_b transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_1/in out VSS en_b transmission_gate
Xsky130_fd_pr__nfet_01v8_E56BNL_0 VSS transmission_gate_1/in en_b VSS sky130_fd_pr__nfet_01v8_E56BNL_AA
C0 transmission_gate_1/in in 0.68fF
C1 VDD out 0.16fF
C2 VDD en_b 0.57fF
C3 out en_b 0.02fF
C4 en in 0.13fF
C5 VDD transmission_gate_1/in 0.42fF
C6 transmission_gate_1/in out 0.72fF
C7 transmission_gate_1/in en_b 0.23fF
C8 en en_b 0.06fF
C9 en transmission_gate_1/in 0.09fF
C10 VDD in 0.10fF
C11 out in 0.43fF
C12 en_b in 0.12fF
C13 en VSS 3.45fF
C14 out VSS 0.90fF
C15 en_b VSS 0.55fF
C16 VDD VSS 10.85fF
C17 transmission_gate_1/in VSS 2.10fF
C18 in VSS 1.01fF
.ends

.subckt a_mux4_en sky130_fd_sc_hd__nand2_1_2/a_113_47# switch_5t_1/transmission_gate_1/in
+ switch_5t_3/en sky130_fd_sc_hd__inv_1_0/Y switch_5t_2/en_b switch_5t_0/en sky130_fd_sc_hd__nand2_1_3/a_113_47#
+ sky130_fd_sc_hd__inv_1_1/Y switch_5t_2/in switch_5t_0/transmission_gate_1/in switch_5t_2/transmission_gate_1/in
+ switch_5t_3/transmission_gate_1/in sky130_fd_sc_hd__nand2_1_0/a_113_47# transmission_gate_3/en_b
+ switch_5t_1/en_b in3 switch_5t_2/en switch_5t_3/in in2 en s0 in0 switch_5t_0/en_b
+ s1 switch_5t_0/in switch_5t_1/in out in1 VDD switch_5t_3/en_b sky130_fd_sc_hd__nand2_1_1/a_113_47#
+ switch_5t_1/en VSS
Xsky130_fd_sc_hd__inv_1_4 switch_5t_0/en switch_5t_0/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_5 switch_5t_2/en switch_5t_2/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_0 out switch_5t_0/en_b switch_5t_0/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD switch_5t_0/in switch_5t_0/en VSS switch_5t_0/transmission_gate_1/in switch_5t_AA
Xsky130_fd_sc_hd__inv_1_6 switch_5t_3/en switch_5t_3/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_1 out switch_5t_1/en_b switch_5t_1/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD switch_5t_1/in switch_5t_1/en VSS switch_5t_1/transmission_gate_1/in switch_5t_AA
Xsky130_fd_sc_hd__inv_1_8 transmission_gate_3/en_b en VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xswitch_5t_2 out switch_5t_2/en_b switch_5t_2/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD switch_5t_2/in switch_5t_2/en VSS switch_5t_2/transmission_gate_1/in switch_5t_AA
Xswitch_5t_3 out switch_5t_3/en_b switch_5t_3/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ VDD switch_5t_3/in switch_5t_3/en VSS switch_5t_3/transmission_gate_1/in switch_5t_AA
Xtransmission_gate_0 en VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in0 switch_5t_0/in VSS transmission_gate_3/en_b transmission_gate
Xtransmission_gate_1 en VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in1 switch_5t_1/in VSS transmission_gate_3/en_b transmission_gate
Xtransmission_gate_2 en VDD transmission_gate_2/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in2 switch_5t_2/in VSS transmission_gate_3/en_b transmission_gate
Xtransmission_gate_3 en VDD transmission_gate_3/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in3 switch_5t_3/in VSS transmission_gate_3/en_b transmission_gate
Xsky130_fd_sc_hd__nand2_1_0 s0 s1 VSS VDD switch_5t_3/en_b VSS VDD sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_1 s0 sky130_fd_sc_hd__inv_1_0/Y VSS VDD switch_5t_2/en_b
+ VSS VDD sky130_fd_sc_hd__nand2_1_1/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_2 s1 sky130_fd_sc_hd__inv_1_1/Y VSS VDD switch_5t_1/en_b
+ VSS VDD sky130_fd_sc_hd__nand2_1_2/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_3 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_1/Y
+ VSS VDD switch_5t_0/en_b VSS VDD sky130_fd_sc_hd__nand2_1_3/a_113_47# sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/Y s0 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/Y s1 VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 switch_5t_1/en switch_5t_1/en_b VSS VDD VSS VDD sky130_fd_sc_hd__inv_1
C0 switch_5t_2/transmission_gate_1/in switch_5t_2/en 0.00fF
C1 transmission_gate_3/en_b in1 0.10fF
C2 VDD in1 -0.02fF
C3 en switch_5t_3/en_b 0.06fF
C4 switch_5t_1/en_b switch_5t_0/in 0.05fF
C5 switch_5t_2/in in2 0.00fF
C6 switch_5t_0/in in0 0.02fF
C7 sky130_fd_sc_hd__inv_1_1/Y switch_5t_1/in 0.07fF
C8 switch_5t_2/transmission_gate_1/in switch_5t_1/en 0.02fF
C9 switch_5t_2/transmission_gate_1/in switch_5t_3/en 0.09fF
C10 switch_5t_0/en switch_5t_1/en_b 0.02fF
C11 switch_5t_2/in switch_5t_2/en_b 0.15fF
C12 switch_5t_1/en_b s0 0.10fF
C13 s0 switch_5t_3/in 0.01fF
C14 sky130_fd_sc_hd__inv_1_0/Y switch_5t_0/in 0.02fF
C15 sky130_fd_sc_hd__nand2_1_0/a_113_47# switch_5t_3/en_b 0.01fF
C16 s1 switch_5t_2/in 0.30fF
C17 switch_5t_2/in switch_5t_2/en 0.09fF
C18 switch_5t_0/en sky130_fd_sc_hd__inv_1_0/Y 0.01fF
C19 s0 sky130_fd_sc_hd__inv_1_0/Y 0.98fF
C20 switch_5t_0/en_b switch_5t_2/in 0.00fF
C21 switch_5t_1/transmission_gate_1/in switch_5t_2/en_b 0.02fF
C22 transmission_gate_3/en_b switch_5t_1/in 0.41fF
C23 in3 switch_5t_2/in 0.07fF
C24 VDD switch_5t_1/in 0.60fF
C25 VDD switch_5t_3/transmission_gate_1/in 0.07fF
C26 switch_5t_1/en_b switch_5t_2/transmission_gate_1/in 0.09fF
C27 switch_5t_1/en switch_5t_2/in 0.01fF
C28 switch_5t_0/transmission_gate_1/in switch_5t_1/in 0.06fF
C29 switch_5t_2/transmission_gate_1/in switch_5t_3/in 0.06fF
C30 switch_5t_1/transmission_gate_1/in switch_5t_2/en 0.09fF
C31 switch_5t_2/in switch_5t_3/en 0.07fF
C32 en in1 0.06fF
C33 switch_5t_0/en_b switch_5t_1/transmission_gate_1/in 0.12fF
C34 switch_5t_2/transmission_gate_1/in sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C35 switch_5t_0/en switch_5t_0/in 0.11fF
C36 s0 switch_5t_0/in 0.04fF
C37 switch_5t_1/transmission_gate_1/in switch_5t_1/en 0.00fF
C38 sky130_fd_sc_hd__inv_1_1/Y switch_5t_2/en_b 0.00fF
C39 out switch_5t_3/transmission_gate_1/in 0.14fF
C40 switch_5t_0/en s0 0.03fF
C41 switch_5t_3/en_b switch_5t_3/transmission_gate_1/in 0.01fF
C42 sky130_fd_sc_hd__inv_1_1/Y s1 0.31fF
C43 switch_5t_1/en_b switch_5t_2/in 0.06fF
C44 switch_5t_3/in switch_5t_2/in 0.35fF
C45 switch_5t_0/en_b sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C46 transmission_gate_3/en_b in2 0.11fF
C47 sky130_fd_sc_hd__nand2_1_2/a_113_47# s1 0.01fF
C48 VDD in2 0.00fF
C49 en switch_5t_1/in 0.12fF
C50 sky130_fd_sc_hd__inv_1_0/Y switch_5t_2/in 0.08fF
C51 switch_5t_1/en sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C52 transmission_gate_3/en_b switch_5t_2/en_b 0.04fF
C53 VDD switch_5t_2/en_b 0.33fF
C54 switch_5t_1/en_b switch_5t_1/transmission_gate_1/in 0.04fF
C55 s1 transmission_gate_3/en_b 1.15fF
C56 switch_5t_2/transmission_gate_1/in s0 0.02fF
C57 s1 VDD 0.75fF
C58 switch_5t_0/en_b sky130_fd_sc_hd__nand2_1_3/a_113_47# -0.00fF
C59 s1 switch_5t_2/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# 0.00fF
C60 transmission_gate_3/en_b switch_5t_2/en 0.04fF
C61 VDD switch_5t_2/en 0.20fF
C62 switch_5t_0/en_b transmission_gate_3/en_b 0.06fF
C63 switch_5t_1/transmission_gate_1/in sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C64 switch_5t_0/en_b VDD 0.02fF
C65 switch_5t_0/en_b switch_5t_0/transmission_gate_1/in 0.03fF
C66 in3 transmission_gate_3/en_b 0.04fF
C67 switch_5t_1/in in1 0.14fF
C68 in3 VDD -0.12fF
C69 switch_5t_1/en transmission_gate_3/en_b 0.01fF
C70 switch_5t_1/en VDD 0.23fF
C71 switch_5t_2/en_b out 0.08fF
C72 transmission_gate_3/en_b switch_5t_3/en 0.00fF
C73 switch_5t_1/en_b sky130_fd_sc_hd__inv_1_1/Y 0.15fF
C74 switch_5t_2/en_b switch_5t_3/en_b 0.38fF
C75 switch_5t_0/transmission_gate_1/in switch_5t_1/en 0.11fF
C76 VDD switch_5t_3/en 0.21fF
C77 s1 switch_5t_3/en_b 0.03fF
C78 s0 switch_5t_2/in 0.46fF
C79 en in2 0.07fF
C80 out switch_5t_2/en 0.07fF
C81 switch_5t_1/en_b sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.01fF
C82 switch_5t_3/en_b switch_5t_2/en 0.19fF
C83 switch_5t_0/en_b out 0.07fF
C84 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__inv_1_0/Y 0.42fF
C85 switch_5t_0/en_b switch_5t_3/en_b 0.00fF
C86 switch_5t_1/transmission_gate_1/in switch_5t_0/in 0.10fF
C87 en switch_5t_2/en_b 0.03fF
C88 s1 en 0.66fF
C89 switch_5t_1/en out 0.08fF
C90 switch_5t_0/en switch_5t_1/transmission_gate_1/in 0.03fF
C91 switch_5t_1/en_b transmission_gate_3/en_b 0.04fF
C92 switch_5t_3/in transmission_gate_3/en_b 0.07fF
C93 switch_5t_3/en out 0.06fF
C94 en switch_5t_2/en 0.03fF
C95 switch_5t_1/en_b VDD 0.30fF
C96 switch_5t_3/in VDD 0.17fF
C97 switch_5t_3/en switch_5t_3/en_b 0.15fF
C98 transmission_gate_3/en_b in0 0.16fF
C99 switch_5t_0/en_b en 0.07fF
C100 switch_5t_0/transmission_gate_1/in switch_5t_1/en_b 0.03fF
C101 switch_5t_2/transmission_gate_1/in switch_5t_2/in 0.02fF
C102 VDD in0 0.07fF
C103 in2 in1 0.23fF
C104 en in3 0.04fF
C105 sky130_fd_sc_hd__inv_1_0/Y transmission_gate_3/en_b 0.10fF
C106 sky130_fd_sc_hd__inv_1_1/Y switch_5t_0/in 0.02fF
C107 sky130_fd_sc_hd__inv_1_0/Y VDD 0.77fF
C108 sky130_fd_sc_hd__inv_1_0/Y switch_5t_2/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# 0.00fF
C109 switch_5t_2/transmission_gate_1/in switch_5t_1/transmission_gate_1/in 0.30fF
C110 sky130_fd_sc_hd__inv_1_1/Y s0 0.29fF
C111 switch_5t_1/en_b out 0.08fF
C112 switch_5t_1/en_b switch_5t_3/en_b 0.01fF
C113 switch_5t_3/in switch_5t_3/en_b 0.09fF
C114 transmission_gate_3/en_b switch_5t_0/in 0.32fF
C115 sky130_fd_sc_hd__inv_1_0/Y switch_5t_3/en_b 0.00fF
C116 VDD switch_5t_0/in -0.19fF
C117 in2 switch_5t_1/in 0.07fF
C118 switch_5t_0/transmission_gate_1/in switch_5t_0/in 0.10fF
C119 switch_5t_1/en_b en 0.03fF
C120 en switch_5t_3/in 0.08fF
C121 switch_5t_0/en transmission_gate_3/en_b 0.07fF
C122 en in0 0.06fF
C123 s0 transmission_gate_3/en_b 0.47fF
C124 sky130_fd_sc_hd__nand2_1_1/a_113_47# switch_5t_2/en_b -0.00fF
C125 switch_5t_0/en VDD 0.08fF
C126 switch_5t_1/in switch_5t_2/en_b 0.02fF
C127 switch_5t_2/en_b switch_5t_3/transmission_gate_1/in 0.09fF
C128 s0 VDD 0.90fF
C129 switch_5t_1/transmission_gate_1/in switch_5t_2/in 0.06fF
C130 switch_5t_0/transmission_gate_1/in switch_5t_0/en 0.06fF
C131 s1 switch_5t_1/in 0.08fF
C132 sky130_fd_sc_hd__inv_1_0/Y en 0.07fF
C133 switch_5t_1/in switch_5t_2/en 0.05fF
C134 switch_5t_3/transmission_gate_1/in switch_5t_2/en 0.02fF
C135 switch_5t_0/en_b switch_5t_1/in 0.13fF
C136 in1 in0 0.33fF
C137 switch_5t_0/en out 0.02fF
C138 switch_5t_1/en switch_5t_1/in 0.14fF
C139 switch_5t_2/transmission_gate_1/in VDD 0.31fF
C140 sky130_fd_sc_hd__inv_1_1/Y switch_5t_2/in 0.02fF
C141 s0 switch_5t_3/en_b 0.10fF
C142 switch_5t_3/en switch_5t_3/transmission_gate_1/in 0.01fF
C143 en switch_5t_0/in 0.14fF
C144 switch_5t_0/en en 0.07fF
C145 s0 en 0.55fF
C146 s1 in2 0.00fF
C147 switch_5t_1/transmission_gate_1/in sky130_fd_sc_hd__inv_1_1/Y 0.02fF
C148 switch_5t_2/transmission_gate_1/in out 0.34fF
C149 switch_5t_2/transmission_gate_1/in switch_5t_3/en_b 0.06fF
C150 transmission_gate_3/en_b switch_5t_2/in 0.17fF
C151 switch_5t_1/en_b switch_5t_1/in 0.28fF
C152 VDD switch_5t_2/in 1.04fF
C153 s1 switch_5t_2/en_b 0.07fF
C154 switch_5t_3/in switch_5t_3/transmission_gate_1/in 0.02fF
C155 switch_5t_1/in in0 0.09fF
C156 in1 switch_5t_0/in 0.07fF
C157 switch_5t_2/en_b switch_5t_2/en 0.61fF
C158 in3 in2 0.23fF
C159 switch_5t_0/en_b switch_5t_2/en_b 0.01fF
C160 s1 switch_5t_2/en 0.03fF
C161 sky130_fd_sc_hd__inv_1_0/Y switch_5t_1/in 0.08fF
C162 switch_5t_0/en_b s1 0.07fF
C163 s0 in1 0.00fF
C164 switch_5t_1/transmission_gate_1/in VDD 0.36fF
C165 switch_5t_1/en switch_5t_2/en_b 0.01fF
C166 switch_5t_0/transmission_gate_1/in switch_5t_1/transmission_gate_1/in 0.41fF
C167 switch_5t_2/en_b switch_5t_3/en 0.46fF
C168 switch_5t_1/en s1 0.02fF
C169 switch_5t_2/in switch_5t_3/en_b 0.09fF
C170 switch_5t_1/en switch_5t_2/en 0.16fF
C171 switch_5t_0/en_b switch_5t_1/en 0.67fF
C172 switch_5t_3/en switch_5t_2/en 0.25fF
C173 switch_5t_1/in switch_5t_0/in 0.54fF
C174 switch_5t_3/in in2 0.06fF
C175 sky130_fd_sc_hd__inv_1_1/Y transmission_gate_3/en_b 0.04fF
C176 switch_5t_1/transmission_gate_1/in out 0.34fF
C177 en switch_5t_2/in 0.09fF
C178 sky130_fd_sc_hd__inv_1_1/Y VDD 0.66fF
C179 switch_5t_0/en switch_5t_1/in 0.01fF
C180 switch_5t_1/en_b switch_5t_2/en_b 0.23fF
C181 s0 sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C182 switch_5t_3/in switch_5t_2/en_b 0.09fF
C183 s0 switch_5t_1/in 0.06fF
C184 sky130_fd_sc_hd__inv_1_0/Y in2 0.01fF
C185 switch_5t_1/en_b s1 0.31fF
C186 s1 switch_5t_3/in 0.02fF
C187 switch_5t_1/en_b switch_5t_2/en 0.42fF
C188 switch_5t_3/in switch_5t_2/en 0.04fF
C189 sky130_fd_sc_hd__inv_1_0/Y switch_5t_2/en_b 0.04fF
C190 switch_5t_0/en_b switch_5t_1/en_b 0.47fF
C191 sky130_fd_sc_hd__inv_1_0/Y s1 0.46fF
C192 switch_5t_2/in in1 0.06fF
C193 transmission_gate_3/en_b VDD 0.47fF
C194 switch_5t_3/in in3 0.00fF
C195 sky130_fd_sc_hd__inv_1_0/Y switch_5t_2/en 0.01fF
C196 switch_5t_0/transmission_gate_1/in transmission_gate_3/en_b 0.02fF
C197 VDD switch_5t_2/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# 0.00fF
C198 switch_5t_1/en_b switch_5t_1/en 0.23fF
C199 switch_5t_2/transmission_gate_1/in switch_5t_1/in 0.07fF
C200 switch_5t_0/transmission_gate_1/in VDD 0.16fF
C201 switch_5t_0/en_b sky130_fd_sc_hd__inv_1_0/Y 0.10fF
C202 switch_5t_2/transmission_gate_1/in switch_5t_3/transmission_gate_1/in 0.30fF
C203 switch_5t_3/in switch_5t_3/en 0.14fF
C204 switch_5t_1/en sky130_fd_sc_hd__inv_1_0/Y 0.02fF
C205 sky130_fd_sc_hd__inv_1_1/Y en 0.03fF
C206 s0 in2 0.00fF
C207 s1 switch_5t_0/in 0.06fF
C208 transmission_gate_3/en_b switch_5t_3/en_b 0.04fF
C209 VDD out 0.97fF
C210 VDD switch_5t_3/en_b 0.28fF
C211 switch_5t_0/transmission_gate_1/in out 0.23fF
C212 s0 switch_5t_2/en_b 0.34fF
C213 switch_5t_0/en_b switch_5t_0/in 0.09fF
C214 switch_5t_0/en s1 0.03fF
C215 switch_5t_2/in switch_5t_1/in 0.30fF
C216 switch_5t_2/in switch_5t_3/transmission_gate_1/in 0.07fF
C217 s0 s1 2.16fF
C218 s0 switch_5t_2/en 0.09fF
C219 switch_5t_0/en_b switch_5t_0/en 0.15fF
C220 en transmission_gate_3/en_b 2.71fF
C221 sky130_fd_sc_hd__inv_1_1/Y in1 0.01fF
C222 switch_5t_1/en switch_5t_0/in 0.13fF
C223 switch_5t_0/en_b s0 0.08fF
C224 en VDD 0.17fF
C225 switch_5t_1/en_b sky130_fd_sc_hd__inv_1_0/Y 0.19fF
C226 switch_5t_0/transmission_gate_1/in en 0.00fF
C227 switch_5t_1/transmission_gate_1/in switch_5t_1/in 0.06fF
C228 switch_5t_0/en switch_5t_1/en 0.20fF
C229 out switch_5t_3/en_b 0.01fF
C230 switch_5t_2/transmission_gate_1/in switch_5t_2/en_b 0.05fF
C231 switch_5t_1/en s0 0.02fF
C232 s0 switch_5t_3/en 0.01fF
C233 switch_5t_2/transmission_gate_1/in s1 0.01fF
C234 sky130_fd_sc_hd__nand2_1_3/a_113_47# VSS 0.01fF
C235 sky130_fd_sc_hd__inv_1_1/Y VSS 24.03fF
C236 sky130_fd_sc_hd__nand2_1_2/a_113_47# VSS -0.00fF
C237 s0 VSS 54.12fF
C238 sky130_fd_sc_hd__inv_1_0/Y VSS 18.63fF
C239 sky130_fd_sc_hd__nand2_1_1/a_113_47# VSS 0.01fF
C240 s1 VSS 33.39fF
C241 sky130_fd_sc_hd__nand2_1_0/a_113_47# VSS -0.00fF
C242 en VSS 8.18fF
C243 switch_5t_3/in VSS 1.04fF
C244 in3 VSS 0.44fF
C245 transmission_gate_3/en_b VSS 7.83fF
C246 VDD VSS -226.82fF
C247 switch_5t_2/in VSS 0.26fF
C248 in2 VSS 0.19fF
C249 switch_5t_1/in VSS 0.85fF
C250 in1 VSS 0.17fF
C251 switch_5t_0/in VSS 2.76fF
C252 in0 VSS 0.84fF
C253 switch_5t_3/en VSS 3.47fF
C254 out VSS 1.82fF
C255 switch_5t_3/en_b VSS 8.83fF
C256 switch_5t_3/transmission_gate_1/in VSS 1.64fF
C257 switch_5t_2/en VSS 4.99fF
C258 switch_5t_2/en_b VSS 11.60fF
C259 switch_5t_2/transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262# VSS 0.00fF
C260 switch_5t_2/transmission_gate_1/in VSS 1.77fF
C261 switch_5t_1/en VSS 12.86fF
C262 switch_5t_1/en_b VSS -2.59fF
C263 switch_5t_1/transmission_gate_1/in VSS 1.77fF
C264 switch_5t_0/en VSS 4.74fF
C265 switch_5t_0/en_b VSS 8.70fF
C266 switch_5t_0/transmission_gate_1/in VSS 1.93fF
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TABSMU c1_n1210_n1160# m3_n1310_n1260# VSUBS
X0 c1_n1210_n1160# m3_n1310_n1260# sky130_fd_pr__cap_mim_m3_1 l=1.16e+07u w=1.16e+07u
C0 c1_n1210_n1160# m3_n1310_n1260# 13.72fF
C1 m3_n1310_n1260# VSUBS 4.03fF
.ends

.subckt sky130_fd_pr__pfet_01v8_VCQUSW a_n810_n632# a_1802_n632# a_n4080_n100# a_2640_n100#
+ a_2010_n100# a_3852_131# a_n3750_n632# a_n3120_n632# a_3600_n632# a_2594_n401# a_n88_n632#
+ a_n2866_n401# a_n2912_n100# a_n718_n632# a_n556_n729# a_2548_n100# a_n182_n100#
+ a_n3658_n632# a_n3028_n632# a_n3496_n729# a_2012_n632# a_2642_n632# a_n1140_n100#
+ a_n1770_n100# a_n1398_n197# a_2172_131# a_n812_n100# a_n4128_131# a_3224_n729# a_n766_n401#
+ a_3480_n100# a_n3122_n100# a_n3752_n100# a_240_n632# a_870_n632# a_n2448_131# a_3388_n100#
+ a_3434_n401# a_n3706_n401# a_3482_n632# a_492_131# a_1500_n632# a_4064_n729# a_n1650_n632#
+ a_n1020_n632# a_n768_131# a_n2238_n197# a_n1558_n632# a_n2610_n100# a_n1396_n729#
+ w_n4520_n851# a_750_n100# a_120_n100# a_1124_n729# a_n2490_n632# a_2340_n632# a_2970_n632#
+ a_1380_n100# a_658_n100# a_n510_n100# a_n1022_n100# a_n1652_n100# a_n138_n197# a_1288_n100#
+ a_n3450_n100# a_n3078_n197# a_n2398_n632# a_122_n632# a_752_n632# a_1334_n401# a_74_n401#
+ a_702_n197# a_1382_n632# a_n1606_n401# a_1962_n197# a_3012_131# a_n390_n632# a_1918_n100#
+ a_28_n100# a_3180_n632# a_n2492_n100# a_1332_131# a_n2236_n729# a_n298_n632# a_3810_n632#
+ a_2850_n100# a_2220_n100# a_n3960_n632# a_n3330_n632# a_2174_n401# a_n1608_131#
+ a_n928_n632# a_n2446_n401# a_n136_n729# a_n3868_n632# a_n3238_n632# a_2758_n100#
+ a_2128_n100# a_n392_n100# a_n3076_n729# a_2802_n197# a_2222_n632# a_2852_n632# a_n1350_n100#
+ a_n1980_n100# a_n4170_n632# a_4020_n632# a_n346_n401# a_3690_n100# a_3060_n100#
+ a_n3332_n100# a_n3962_n100# a_2592_131# a_450_n632# a_n3286_n401# a_3598_n100# a_n4078_n632#
+ a_1080_n632# a_3014_n401# a_n2868_131# a_3062_n632# a_3692_n632# a_n2190_n100# a_3642_n197#
+ a_n1860_n632# a_n1230_n632# a_1710_n632# a_n4172_n100# a_n2820_n100# a_n1768_n632#
+ a_n1138_n632# a_n1188_131# a_704_n729# a_n4126_n401# a_960_n100# a_330_n100# a_1964_n729#
+ a_1590_n100# a_282_n197# a_n2070_n632# a_2550_n632# a_n90_n100# a_n978_n197# a_n1186_n401#
+ a_868_n100# a_238_n100# a_n720_n100# a_n1232_n100# a_n1862_n100# a_914_n401# a_1498_n100#
+ a_n3030_n100# a_n3660_n100# a_n2700_n632# a_332_n632# a_962_n632# a_1542_n197# a_1592_n632#
+ a_n3918_n197# a_n2608_n632# a_3390_n632# a_n2072_n100# a_3432_131# a_n600_n632#
+ a_1752_131# a_2804_n729# a_n3540_n632# a_2430_n100# a_n2702_n100# a_n3708_131# a_n508_n632#
+ a_n2026_n401# a_2382_n197# a_2968_n100# a_2338_n100# a_n976_n729# a_n3448_n632#
+ a_n1560_n100# a_2432_n632# a_3644_n729# a_3270_n100# a_n602_n100# a_n2028_131# a_n3916_n729#
+ a_n3542_n100# a_660_n632# a_n1818_n197# a_3178_n100# a_1290_n632# a_3900_n100# a_3854_n401#
+ a_3222_n197# a_3272_n632# a_n348_131# a_30_n632# a_3808_n100# a_n1440_n632# a_1920_n632#
+ a_284_n729# a_n2658_n197# a_3902_n632# a_n2400_n100# a_n1978_n632# a_n1348_n632#
+ a_n3288_131# a_4110_n100# a_494_n401# a_540_n100# a_4062_n197# a_4018_n100# a_1544_n729#
+ a_n2280_n632# a_2130_n632# a_2760_n632# a_1170_n100# a_72_131# a_n300_n100# a_n930_n100#
+ a_n1442_n100# a_n558_n197# a_n1816_n729# a_448_n100# a_n3240_n100# a_n3870_n100#
+ a_n3498_n197# a_n2188_n632# a_4112_n632# a_1078_n100# a_1754_n401# a_1800_n100#
+ a_n2910_n632# a_542_n632# a_1122_n197# a_n180_n632# a_1172_n632# a_2384_n729# a_n2818_n632#
+ a_1708_n100# a_912_131# VSUBS a_n2656_n729# a_n2282_n100#
X0 a_n90_n100# a_n138_n197# a_n182_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_330_n100# a_282_n197# a_238_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2 a_n3868_n632# a_n3916_n729# a_n3960_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X3 a_n1348_n632# a_n1396_n729# a_n1440_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X4 a_n3450_n100# a_n3498_n197# a_n3542_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X5 a_3480_n100# a_3432_131# a_3388_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X6 a_3062_n632# a_3014_n401# a_2970_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X7 a_542_n632# a_494_n401# a_450_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X8 a_2432_n632# a_2384_n729# a_2340_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X9 a_n1770_n100# a_n1818_n197# a_n1862_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X10 a_1800_n100# a_1752_131# a_1708_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X11 a_n508_n632# a_n556_n729# a_n600_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X12 a_1592_n632# a_1544_n729# a_1500_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X13 a_2222_n632# a_2174_n401# a_2130_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X14 a_540_n100# a_492_131# a_448_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X15 a_2220_n100# a_2172_131# a_2128_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X16 a_n3660_n100# a_n3708_131# a_n3752_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X17 a_n300_n100# a_n348_131# a_n392_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X18 a_3690_n100# a_3642_n197# a_3598_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X19 a_n3028_n632# a_n3076_n729# a_n3120_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X20 a_n2398_n632# a_n2446_n401# a_n2490_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X21 a_4110_n100# a_4062_n197# a_4018_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X22 a_n1558_n632# a_n1606_n401# a_n1650_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X23 a_n1980_n100# a_n2028_131# a_n2072_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X24 a_2010_n100# a_1962_n197# a_1918_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X25 a_3272_n632# a_3224_n729# a_3180_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X26 a_n510_n100# a_n558_n197# a_n602_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X27 a_750_n100# a_702_n197# a_658_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X28 a_752_n632# a_704_n729# a_660_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X29 a_2642_n632# a_2594_n401# a_2550_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X30 a_n3870_n100# a_n3918_n197# a_n3962_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X31 a_3900_n100# a_3852_131# a_3808_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X32 a_n4078_n632# a_n4126_n401# a_n4170_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X33 a_n718_n632# a_n766_n401# a_n810_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X34 a_1802_n632# a_1754_n401# a_1710_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X35 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=2.48e+12p pd=2.096e+07u as=0p ps=0u w=1e+06u l=150000u
X36 a_n3238_n632# a_n3286_n401# a_n3330_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X37 a_n2608_n632# a_n2656_n729# a_n2700_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X38 a_n2190_n100# a_n2238_n197# a_n2282_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X39 a_n720_n100# a_n768_131# a_n812_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X40 a_960_n100# a_912_131# a_868_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X41 a_n1768_n632# a_n1816_n729# a_n1860_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X42 a_4112_n632# a_4064_n729# a_4020_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X43 a_n4080_n100# a_n4128_131# a_n4172_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X44 a_2852_n632# a_2804_n729# a_2760_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X45 a_3482_n632# a_3434_n401# a_3390_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X46 a_962_n632# a_914_n401# a_870_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X47 a_n2400_n100# a_n2448_131# a_n2492_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X48 a_2430_n100# a_2382_n197# a_2338_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X49 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n928_n632# a_n976_n729# a_n1020_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X51 a_122_n632# a_74_n401# a_30_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X52 a_2012_n632# a_1964_n729# a_1920_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X53 a_n3448_n632# a_n3496_n729# a_n3540_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X54 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_n930_n100# a_n978_n197# a_n1022_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X56 a_n2818_n632# a_n2866_n401# a_n2910_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X57 a_n1140_n100# a_n1188_131# a_n1232_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X58 a_1170_n100# a_1122_n197# a_1078_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X59 a_n88_n632# a_n136_n729# a_n180_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X60 w_n4520_n851# w_n4520_n851# w_n4520_n851# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_n2610_n100# a_n2658_n197# a_n2702_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X62 a_2640_n100# a_2592_131# a_2548_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X63 a_1172_n632# a_1124_n729# a_1080_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X64 a_3692_n632# a_3644_n729# a_3600_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X65 a_n3030_n100# a_n3078_n197# a_n3122_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X66 a_3060_n100# a_3012_131# a_2968_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X67 a_n1978_n632# a_n2026_n401# a_n2070_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X68 a_n3658_n632# a_n3706_n401# a_n3750_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X69 a_n1138_n632# a_n1186_n401# a_n1230_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X70 a_n1350_n100# a_n1398_n197# a_n1442_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X71 a_1380_n100# a_1332_131# a_1288_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X72 a_n2820_n100# a_n2868_131# a_n2912_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X73 a_2850_n100# a_2802_n197# a_2758_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X74 a_332_n632# a_284_n729# a_240_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X75 a_n3240_n100# a_n3288_131# a_n3332_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X76 a_3270_n100# a_3222_n197# a_3178_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X77 a_n298_n632# a_n346_n401# a_n390_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X78 a_1382_n632# a_1334_n401# a_1290_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X79 a_3902_n632# a_3854_n401# a_3810_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X80 a_n1560_n100# a_n1608_131# a_n1652_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X81 a_120_n100# a_72_131# a_28_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X82 a_1590_n100# a_1542_n197# a_1498_n100# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X83 a_n2188_n632# a_n2236_n729# a_n2280_n632# w_n4520_n851# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
C0 a_n1186_n401# a_n1188_131# 0.01fF
C1 a_752_n632# a_660_n632# 0.09fF
C2 a_542_n632# a_2130_n632# 0.00fF
C3 a_1172_n632# a_660_n632# 0.01fF
C4 a_n348_131# a_1122_n197# 0.00fF
C5 a_3480_n100# a_2758_n100# 0.01fF
C6 a_n2280_n632# a_n1558_n632# 0.01fF
C7 a_914_n401# a_704_n729# 0.00fF
C8 a_238_n100# a_330_n100# 0.09fF
C9 a_240_n632# a_n600_n632# 0.01fF
C10 a_n4080_n100# a_n4126_n401# 0.00fF
C11 a_n1978_n632# a_n3330_n632# 0.00fF
C12 a_n1978_n632# a_n2188_n632# 0.03fF
C13 a_n1140_n100# a_n1862_n100# 0.01fF
C14 a_n2280_n632# a_n3750_n632# 0.00fF
C15 a_3600_n632# a_2222_n632# 0.00fF
C16 a_n138_n197# a_n348_131# 0.00fF
C17 a_n136_n729# a_n1606_n401# 0.00fF
C18 a_n1770_n100# a_n2702_n100# 0.01fF
C19 a_3600_n632# a_2642_n632# 0.01fF
C20 a_1288_n100# a_1332_131# 0.00fF
C21 a_120_n100# a_868_n100# 0.01fF
C22 a_n3030_n100# a_n3542_n100# 0.01fF
C23 w_n4520_n851# a_122_n632# 0.01fF
C24 a_2852_n632# a_4020_n632# 0.01fF
C25 a_2384_n729# a_1124_n729# 0.00fF
C26 a_1288_n100# a_1498_n100# 0.03fF
C27 a_n2070_n632# a_n928_n632# 0.01fF
C28 a_n2026_n401# a_n1980_n100# 0.00fF
C29 w_n4520_n851# a_n1232_n100# 0.02fF
C30 a_n346_n401# a_n1816_n729# 0.00fF
C31 a_3902_n632# a_3692_n632# 0.03fF
C32 a_n3870_n100# a_n3542_n100# 0.02fF
C33 a_3480_n100# a_3900_n100# 0.02fF
C34 a_n3496_n729# a_n3076_n729# 0.01fF
C35 a_912_131# a_2172_131# 0.00fF
C36 a_n3540_n632# a_n1978_n632# 0.00fF
C37 a_n3030_n100# a_n1980_n100# 0.01fF
C38 a_450_n632# a_492_131# 0.00fF
C39 a_n1396_n729# a_n766_n401# 0.00fF
C40 a_n602_n100# a_n90_n100# 0.01fF
C41 a_1544_n729# a_1754_n401# 0.00fF
C42 a_752_n632# a_122_n632# 0.01fF
C43 a_2012_n632# a_1920_n632# 0.09fF
C44 a_1590_n100# a_2010_n100# 0.02fF
C45 a_914_n401# a_960_n100# 0.00fF
C46 w_n4520_n851# a_n3918_n197# 0.11fF
C47 a_n1020_n632# a_n298_n632# 0.01fF
C48 a_1172_n632# a_122_n632# 0.01fF
C49 a_n2910_n632# a_n3868_n632# 0.01fF
C50 a_n976_n729# a_74_n401# 0.00fF
C51 a_n2490_n632# a_n1650_n632# 0.01fF
C52 a_2172_131# a_2174_n401# 0.01fF
C53 a_n1978_n632# a_n1980_n100# 0.00fF
C54 a_2384_n729# a_2174_n401# 0.00fF
C55 a_1332_131# a_1752_131# 0.01fF
C56 a_n3122_n100# a_n3660_n100# 0.01fF
C57 a_n2700_n632# a_n3868_n632# 0.01fF
C58 a_n1140_n100# a_n1188_131# 0.00fF
C59 a_n4080_n100# a_n4172_n100# 0.09fF
C60 a_2968_n100# a_3270_n100# 0.02fF
C61 a_n3240_n100# a_n3660_n100# 0.02fF
C62 a_n558_n197# a_n348_131# 0.00fF
C63 a_120_n100# a_540_n100# 0.02fF
C64 a_74_n401# a_1334_n401# 0.00fF
C65 a_28_n100# a_1170_n100# 0.01fF
C66 a_1332_131# a_1122_n197# 0.00fF
C67 a_870_n632# a_1802_n632# 0.01fF
C68 a_n1020_n632# a_n508_n632# 0.01fF
C69 a_n930_n100# a_n1770_n100# 0.01fF
C70 a_n4172_n100# a_n3752_n100# 0.02fF
C71 a_n2070_n632# a_n2818_n632# 0.01fF
C72 a_n2070_n632# a_n3120_n632# 0.01fF
C73 a_2338_n100# a_2850_n100# 0.01fF
C74 a_1080_n632# a_1710_n632# 0.01fF
C75 w_n4520_n851# a_1964_n729# 0.12fF
C76 a_868_n100# a_1078_n100# 0.03fF
C77 a_n3658_n632# a_n3028_n632# 0.01fF
C78 a_658_n100# a_868_n100# 0.03fF
C79 a_3852_131# a_3222_n197# 0.00fF
C80 a_n138_n197# a_1332_131# 0.00fF
C81 a_n1650_n632# a_n2188_n632# 0.01fF
C82 a_1802_n632# a_3180_n632# 0.00fF
C83 a_870_n632# a_n180_n632# 0.01fF
C84 a_n1442_n100# a_n2610_n100# 0.01fF
C85 a_2550_n632# a_1592_n632# 0.01fF
C86 a_332_n632# a_1710_n632# 0.00fF
C87 a_4062_n197# a_3222_n197# 0.01fF
C88 a_1802_n632# a_660_n632# 0.01fF
C89 a_1708_n100# a_2548_n100# 0.01fF
C90 w_n4520_n851# a_3690_n100# 0.04fF
C91 a_n1348_n632# a_n2608_n632# 0.00fF
C92 a_238_n100# a_1708_n100# 0.00fF
C93 a_4112_n632# a_3692_n632# 0.02fF
C94 a_3270_n100# a_3178_n100# 0.09fF
C95 a_n1440_n632# a_n298_n632# 0.01fF
C96 a_n3030_n100# a_n1652_n100# 0.00fF
C97 a_n90_n100# a_28_n100# 0.07fF
C98 a_120_n100# a_1288_n100# 0.01fF
C99 a_2222_n632# a_3390_n632# 0.01fF
C100 a_n3330_n632# a_n3288_131# 0.00fF
C101 a_2760_n632# a_3180_n632# 0.02fF
C102 a_n180_n632# a_660_n632# 0.01fF
C103 a_2642_n632# a_3390_n632# 0.01fF
C104 a_n300_n100# a_n1140_n100# 0.01fF
C105 a_n1348_n632# a_n810_n632# 0.01fF
C106 a_450_n632# a_1382_n632# 0.01fF
C107 w_n4520_n851# a_n2492_n100# 0.02fF
C108 a_540_n100# a_1078_n100# 0.01fF
C109 a_658_n100# a_540_n100# 0.07fF
C110 a_n2026_n401# a_n766_n401# 0.00fF
C111 a_n1440_n632# a_n508_n632# 0.01fF
C112 a_n390_n632# a_n1138_n632# 0.01fF
C113 a_4018_n100# a_2850_n100# 0.01fF
C114 a_n2400_n100# a_n812_n100# 0.00fF
C115 a_3180_n632# a_3482_n632# 0.02fF
C116 a_3642_n197# a_2172_131# 0.00fF
C117 a_2968_n100# a_2010_n100# 0.01fF
C118 a_2432_n632# a_962_n632# 0.00fF
C119 w_n4520_n851# a_1170_n100# 0.02fF
C120 a_1918_n100# a_1920_n632# 0.00fF
C121 a_3600_n632# a_3810_n632# 0.03fF
C122 a_3062_n632# a_2130_n632# 0.01fF
C123 a_1592_n632# a_1290_n632# 0.02fF
C124 a_2852_n632# w_n4520_n851# 0.03fF
C125 a_n3870_n100# a_n3916_n729# 0.00fF
C126 a_3642_n197# a_3012_131# 0.00fF
C127 a_n2070_n632# a_n1768_n632# 0.02fF
C128 a_n3120_n632# a_n3122_n100# 0.00fF
C129 a_2384_n729# a_2430_n100# 0.00fF
C130 a_n1020_n632# w_n4520_n851# 0.01fF
C131 a_2802_n197# a_2172_131# 0.00fF
C132 a_n3448_n632# a_n4078_n632# 0.01fF
C133 a_2802_n197# a_3012_131# 0.00fF
C134 a_n2190_n100# a_n1232_n100# 0.01fF
C135 a_3060_n100# a_2758_n100# 0.02fF
C136 a_2338_n100# a_1590_n100# 0.01fF
C137 a_3600_n632# a_2550_n632# 0.01fF
C138 a_n2912_n100# a_n1442_n100# 0.00fF
C139 a_n2608_n632# a_n4078_n632# 0.00fF
C140 a_1172_n632# a_1170_n100# 0.00fF
C141 a_870_n632# a_542_n632# 0.02fF
C142 a_750_n100# a_1170_n100# 0.02fF
C143 a_2432_n632# a_2222_n632# 0.03fF
C144 a_120_n100# a_n182_n100# 0.02fF
C145 a_n180_n632# a_122_n632# 0.02fF
C146 a_4018_n100# a_4110_n100# 0.09fF
C147 a_2340_n632# a_3692_n632# 0.00fF
C148 a_1288_n100# a_1078_n100# 0.03fF
C149 a_1288_n100# a_658_n100# 0.01fF
C150 a_n3448_n632# a_n4170_n632# 0.01fF
C151 a_2432_n632# a_2642_n632# 0.03fF
C152 a_n1608_131# a_n1398_n197# 0.00fF
C153 a_n1442_n100# a_n2282_n100# 0.01fF
C154 a_n90_n100# w_n4520_n851# 0.02fF
C155 a_n510_n100# a_n1862_n100# 0.00fF
C156 a_n88_n632# a_n928_n632# 0.01fF
C157 a_2850_n100# a_1800_n100# 0.01fF
C158 a_2010_n100# a_3178_n100# 0.01fF
C159 a_n1978_n632# a_n1558_n632# 0.02fF
C160 a_n2070_n632# a_n718_n632# 0.00fF
C161 a_n3708_131# w_n4520_n851# 0.13fF
C162 a_n2608_n632# a_n4170_n632# 0.00fF
C163 a_238_n100# a_n1232_n100# 0.00fF
C164 a_n1022_n100# a_n1862_n100# 0.01fF
C165 a_494_n401# a_704_n729# 0.00fF
C166 a_n3658_n632# a_n2490_n632# 0.01fF
C167 a_2804_n729# a_2850_n100# 0.00fF
C168 a_3060_n100# a_3900_n100# 0.01fF
C169 a_n1020_n632# a_n2398_n632# 0.00fF
C170 a_542_n632# a_660_n632# 0.07fF
C171 a_450_n632# a_n600_n632# 0.01fF
C172 a_n768_131# a_702_n197# 0.00fF
C173 a_n1818_n197# a_n2028_131# 0.00fF
C174 a_n1978_n632# a_n2280_n632# 0.02fF
C175 a_n3332_n100# a_n3330_n632# 0.00fF
C176 a_n1650_n632# a_n1652_n100# 0.00fF
C177 a_2382_n197# a_2592_131# 0.00fF
C178 a_2128_n100# a_2850_n100# 0.01fF
C179 a_n2656_n729# a_n2236_n729# 0.01fF
C180 a_120_n100# a_n1442_n100# 0.00fF
C181 a_1498_n100# a_330_n100# 0.01fF
C182 w_n4520_n851# a_492_131# 0.12fF
C183 a_1962_n197# a_1332_131# 0.00fF
C184 a_n1440_n632# w_n4520_n851# 0.01fF
C185 a_n4172_n100# a_n2610_n100# 0.00fF
C186 a_n3918_n197# a_n3078_n197# 0.01fF
C187 a_n928_n632# a_n1230_n632# 0.02fF
C188 a_n3918_n197# a_n2448_131# 0.00fF
C189 a_750_n100# a_n90_n100# 0.01fF
C190 a_332_n632# a_1080_n632# 0.01fF
C191 a_30_n632# a_962_n632# 0.01fF
C192 a_n136_n729# a_1124_n729# 0.00fF
C193 a_1918_n100# a_2220_n100# 0.02fF
C194 a_n720_n100# a_n1862_n100# 0.01fF
C195 a_1122_n197# a_1078_n100# 0.00fF
C196 a_n3330_n632# a_n3658_n632# 0.02fF
C197 a_3014_n401# a_2384_n729# 0.00fF
C198 a_n3658_n632# a_n2188_n632# 0.00fF
C199 a_n1862_n100# a_n1980_n100# 0.07fF
C200 a_n602_n100# a_n600_n632# 0.00fF
C201 a_1288_n100# a_2758_n100# 0.00fF
C202 a_n2072_n100# a_n812_n100# 0.00fF
C203 a_n720_n100# a_n768_131# 0.00fF
C204 a_n2070_n632# a_n1860_n632# 0.03fF
C205 a_n3332_n100# a_n3542_n100# 0.03fF
C206 a_1754_n401# a_2594_n401# 0.01fF
C207 a_3014_n401# a_3012_131# 0.01fF
C208 a_n3448_n632# a_n3450_n100# 0.00fF
C209 a_n182_n100# a_1078_n100# 0.00fF
C210 a_658_n100# a_n182_n100# 0.01fF
C211 a_1380_n100# a_2010_n100# 0.01fF
C212 a_2970_n632# a_4020_n632# 0.01fF
C213 a_2640_n100# w_n4520_n851# 0.02fF
C214 a_2850_n100# a_3808_n100# 0.01fF
C215 w_n4520_n851# a_n1398_n197# 0.10fF
C216 a_3390_n632# a_3810_n632# 0.02fF
C217 a_3014_n401# a_4064_n729# 0.00fF
C218 a_3222_n197# a_3432_131# 0.00fF
C219 a_n2026_n401# a_n1396_n729# 0.00fF
C220 w_n4520_n851# a_1542_n197# 0.10fF
C221 a_3272_n632# a_2130_n632# 0.01fF
C222 a_1500_n632# a_2130_n632# 0.01fF
C223 a_n3332_n100# a_n1980_n100# 0.00fF
C224 a_448_n100# a_2010_n100# 0.00fF
C225 a_542_n632# a_122_n632# 0.02fF
C226 a_1544_n729# a_74_n401# 0.00fF
C227 a_2968_n100# a_2338_n100# 0.01fF
C228 a_30_n632# a_n390_n632# 0.02fF
C229 a_n3540_n632# a_n3658_n632# 0.07fF
C230 a_3690_n100# a_2548_n100# 0.01fF
C231 a_n2398_n632# a_n1440_n632# 0.01fF
C232 a_n2912_n100# a_n2910_n632# 0.00fF
C233 a_450_n632# a_1920_n632# 0.00fF
C234 a_n1650_n632# a_n1558_n632# 0.09fF
C235 a_n298_n632# a_n600_n632# 0.02fF
C236 a_n2190_n100# a_n2492_n100# 0.02fF
C237 a_2430_n100# a_3270_n100# 0.01fF
C238 a_n2818_n632# a_n1230_n632# 0.00fF
C239 a_2550_n632# a_3390_n632# 0.01fF
C240 a_1590_n100# a_1800_n100# 0.03fF
C241 a_n1350_n100# a_n182_n100# 0.01fF
C242 a_3222_n197# w_n4520_n851# 0.10fF
C243 a_n3660_n100# a_n3706_n401# 0.00fF
C244 a_1544_n729# a_1500_n632# 0.00fF
C245 a_2852_n632# a_1802_n632# 0.01fF
C246 a_n1348_n632# a_n1138_n632# 0.03fF
C247 a_n1650_n632# a_n2280_n632# 0.01fF
C248 a_3902_n632# a_3600_n632# 0.02fF
C249 a_n508_n632# a_n600_n632# 0.09fF
C250 a_4110_n100# a_3808_n100# 0.02fF
C251 a_n976_n729# a_284_n729# 0.00fF
C252 a_2128_n100# a_1590_n100# 0.01fF
C253 a_1382_n632# w_n4520_n851# 0.01fF
C254 a_n2912_n100# a_n4172_n100# 0.00fF
C255 a_450_n632# a_2012_n632# 0.00fF
C256 a_n300_n100# a_n510_n100# 0.03fF
C257 a_n2492_n100# a_n2448_131# 0.00fF
C258 a_120_n100# a_330_n100# 0.03fF
C259 a_n1022_n100# a_n978_n197# 0.00fF
C260 a_2548_n100# a_1170_n100# 0.00fF
C261 a_2338_n100# a_3178_n100# 0.01fF
C262 a_n1862_n100# a_n1652_n100# 0.03fF
C263 a_284_n729# a_1334_n401# 0.00fF
C264 a_238_n100# a_1170_n100# 0.01fF
C265 a_n2070_n632# a_n2910_n632# 0.01fF
C266 a_n1020_n632# a_n180_n632# 0.01fF
C267 a_2432_n632# a_3810_n632# 0.00fF
C268 a_n300_n100# a_n1022_n100# 0.01fF
C269 a_n1350_n100# a_n1442_n100# 0.09fF
C270 a_1708_n100# a_1498_n100# 0.03fF
C271 a_2760_n632# a_2852_n632# 0.09fF
C272 a_4018_n100# a_2968_n100# 0.01fF
C273 a_450_n632# a_240_n632# 0.03fF
C274 a_n2072_n100# a_n602_n100# 0.00fF
C275 a_n4080_n100# a_n2492_n100# 0.00fF
C276 a_960_n100# a_1590_n100# 0.01fF
C277 a_n2070_n632# a_n2700_n632# 0.01fF
C278 a_n3330_n632# a_n3286_n401# 0.00fF
C279 a_n3448_n632# a_n3960_n632# 0.01fF
C280 a_n136_n729# a_n766_n401# 0.00fF
C281 a_2172_131# a_3012_131# 0.01fF
C282 a_752_n632# a_1382_n632# 0.01fF
C283 a_1172_n632# a_1382_n632# 0.03fF
C284 a_3598_n100# a_2758_n100# 0.01fF
C285 a_n2608_n632# a_n3960_n632# 0.00fF
C286 a_n3752_n100# a_n2492_n100# 0.00fF
C287 a_n392_n100# a_n812_n100# 0.02fF
C288 a_n4078_n632# a_n3028_n632# 0.01fF
C289 a_2852_n632# a_3482_n632# 0.01fF
C290 a_2432_n632# a_2550_n632# 0.07fF
C291 a_492_131# a_72_131# 0.01fF
C292 a_n1230_n632# a_n1768_n632# 0.01fF
C293 a_n3706_n401# a_n2236_n729# 0.00fF
C294 a_n300_n100# a_n720_n100# 0.02fF
C295 a_2222_n632# a_2174_n401# 0.00fF
C296 a_3062_n632# a_3180_n632# 0.07fF
C297 a_n2446_n401# a_n2656_n729# 0.00fF
C298 a_n1770_n100# a_n1768_n632# 0.00fF
C299 a_n88_n632# a_n718_n632# 0.01fF
C300 a_2010_n100# a_2430_n100# 0.02fF
C301 a_1754_n401# a_1964_n729# 0.00fF
C302 a_n766_n401# a_n768_131# 0.01fF
C303 a_238_n100# a_n90_n100# 0.02fF
C304 a_2850_n100# a_3388_n100# 0.01fF
C305 a_n1560_n100# a_n1140_n100# 0.02fF
C306 a_n3028_n632# a_n4170_n632# 0.01fF
C307 a_n2400_n100# w_n4520_n851# 0.02fF
C308 a_n3708_131# a_n3078_n197# 0.00fF
C309 a_4018_n100# a_3178_n100# 0.01fF
C310 a_3600_n632# a_4112_n632# 0.01fF
C311 a_n3708_131# a_n2448_131# 0.00fF
C312 a_3598_n100# a_3900_n100# 0.02fF
C313 a_2338_n100# a_1380_n100# 0.01fF
C314 a_2340_n632# a_1592_n632# 0.01fF
C315 w_n4520_n851# a_n3076_n729# 0.12fF
C316 a_3014_n401# a_3854_n401# 0.01fF
C317 a_n1978_n632# a_n2026_n401# 0.00fF
C318 a_2968_n100# a_1800_n100# 0.01fF
C319 a_n3870_n100# a_n3030_n100# 0.01fF
C320 a_330_n100# a_1078_n100# 0.01fF
C321 a_n1232_n100# a_n2610_n100# 0.00fF
C322 a_658_n100# a_330_n100# 0.02fF
C323 a_72_131# a_n1398_n197# 0.00fF
C324 a_n180_n632# a_n1440_n632# 0.00fF
C325 a_2970_n632# w_n4520_n851# 0.03fF
C326 w_n4520_n851# a_n600_n632# 0.01fF
C327 a_n3542_n100# a_n3962_n100# 0.02fF
C328 a_1542_n197# a_72_131# 0.00fF
C329 a_n1560_n100# a_n1606_n401# 0.00fF
C330 a_240_n632# a_n298_n632# 0.01fF
C331 a_n1770_n100# a_n182_n100# 0.00fF
C332 a_n1348_n632# a_n2490_n632# 0.01fF
C333 a_n718_n632# a_n1230_n632# 0.01fF
C334 a_2432_n632# a_1290_n632# 0.01fF
C335 a_n1140_n100# a_n2702_n100# 0.00fF
C336 a_n3708_131# a_n3752_n100# 0.00fF
C337 a_2968_n100# a_2128_n100# 0.01fF
C338 a_n300_n100# a_448_n100# 0.01fF
C339 a_3902_n632# a_3390_n632# 0.01fF
C340 a_n1816_n729# a_n2656_n729# 0.01fF
C341 a_542_n632# a_n1020_n632# 0.00fF
C342 a_962_n632# a_1710_n632# 0.01fF
C343 a_704_n729# a_702_n197# 0.01fF
C344 a_4110_n100# a_3388_n100# 0.01fF
C345 a_752_n632# a_n600_n632# 0.00fF
C346 a_240_n632# a_n508_n632# 0.01fF
C347 a_120_n100# a_1708_n100# 0.00fF
C348 a_n2398_n632# a_n2400_n100# 0.00fF
C349 a_n2238_n197# a_n1608_131# 0.00fF
C350 a_2640_n100# a_2548_n100# 0.09fF
C351 a_n392_n100# a_n602_n100# 0.03fF
C352 a_n3122_n100# a_n4172_n100# 0.01fF
C353 a_n1348_n632# a_30_n632# 0.00fF
C354 a_1800_n100# a_3178_n100# 0.00fF
C355 a_3390_n632# a_3388_n100# 0.00fF
C356 a_n1348_n632# a_n2188_n632# 0.01fF
C357 a_n1770_n100# a_n1442_n100# 0.02fF
C358 a_914_n401# a_1334_n401# 0.01fF
C359 a_n3240_n100# a_n4172_n100# 0.01fF
C360 a_n2448_131# a_n1398_n197# 0.00fF
C361 a_n300_n100# a_n1652_n100# 0.00fF
C362 a_n2820_n100# a_n3542_n100# 0.01fF
C363 a_n3658_n632# a_n3750_n632# 0.09fF
C364 a_3480_n100# a_2850_n100# 0.01fF
C365 a_n1860_n632# a_n1230_n632# 0.01fF
C366 a_n1816_n729# a_n1770_n100# 0.00fF
C367 a_2968_n100# a_3808_n100# 0.01fF
C368 a_2222_n632# a_1710_n632# 0.01fF
C369 a_n3658_n632# a_n2280_n632# 0.00fF
C370 a_1382_n632# a_1802_n632# 0.02fF
C371 w_n4520_n851# a_1920_n632# 0.01fF
C372 a_n510_n100# a_960_n100# 0.00fF
C373 a_2642_n632# a_1710_n632# 0.01fF
C374 a_870_n632# a_1500_n632# 0.01fF
C375 a_2592_131# a_1752_131# 0.01fF
C376 a_2128_n100# a_3178_n100# 0.01fF
C377 a_3600_n632# a_2340_n632# 0.00fF
C378 a_n2820_n100# a_n1980_n100# 0.01fF
C379 a_n136_n729# a_n1396_n729# 0.00fF
C380 a_1124_n729# a_704_n729# 0.01fF
C381 a_2592_131# a_1122_n197# 0.00fF
C382 a_n2490_n632# a_n4078_n632# 0.00fF
C383 a_n1140_n100# a_n930_n100# 0.03fF
C384 a_282_n197# a_702_n197# 0.01fF
C385 a_n390_n632# a_n1558_n632# 0.01fF
C386 a_3224_n729# a_2174_n401# 0.00fF
C387 a_3854_n401# a_2384_n729# 0.00fF
C388 a_4112_n632# a_4110_n100# 0.00fF
C389 a_n2656_n729# a_n4126_n401# 0.00fF
C390 a_3902_n632# a_2432_n632# 0.00fF
C391 a_n180_n632# a_1382_n632# 0.00fF
C392 a_3272_n632# a_3180_n632# 0.09fF
C393 a_n2072_n100# w_n4520_n851# 0.02fF
C394 a_752_n632# a_1920_n632# 0.01fF
C395 a_2760_n632# a_1382_n632# 0.00fF
C396 a_30_n632# a_1290_n632# 0.00fF
C397 a_1172_n632# a_1920_n632# 0.01fF
C398 a_3854_n401# a_4064_n729# 0.00fF
C399 a_n1232_n100# a_n2282_n100# 0.01fF
C400 a_660_n632# a_1500_n632# 0.01fF
C401 a_2594_n401# a_3434_n401# 0.01fF
C402 a_3692_n632# a_2130_n632# 0.00fF
C403 a_4112_n632# a_3390_n632# 0.01fF
C404 w_n4520_n851# a_2012_n632# 0.01fF
C405 w_n4520_n851# a_n2238_n197# 0.10fF
C406 a_n3916_n729# a_n3286_n401# 0.00fF
C407 a_2338_n100# a_2430_n100# 0.09fF
C408 a_3480_n100# a_4110_n100# 0.01fF
C409 a_1380_n100# a_1800_n100# 0.02fF
C410 a_1708_n100# a_1078_n100# 0.01fF
C411 a_658_n100# a_1708_n100# 0.01fF
C412 a_704_n729# a_2174_n401# 0.00fF
C413 a_n2610_n100# a_n2492_n100# 0.07fF
C414 a_n392_n100# a_28_n100# 0.02fF
C415 a_n1978_n632# a_n1650_n632# 0.02fF
C416 a_3178_n100# a_3808_n100# 0.01fF
C417 a_n2700_n632# a_n2656_n729# 0.00fF
C418 a_n2446_n401# a_n3706_n401# 0.00fF
C419 a_448_n100# a_1800_n100# 0.00fF
C420 a_3644_n729# w_n4520_n851# 0.10fF
C421 a_n3330_n632# a_n4078_n632# 0.01fF
C422 a_4062_n197# a_3852_131# 0.00fF
C423 a_n810_n632# a_n928_n632# 0.07fF
C424 a_240_n632# w_n4520_n851# 0.01fF
C425 a_120_n100# a_122_n632# 0.00fF
C426 a_2804_n729# a_2174_n401# 0.00fF
C427 a_n3238_n632# w_n4520_n851# 0.03fF
C428 a_n3028_n632# a_n3960_n632# 0.01fF
C429 a_120_n100# a_n1232_n100# 0.00fF
C430 a_2128_n100# a_1380_n100# 0.01fF
C431 a_n2190_n100# a_n2400_n100# 0.03fF
C432 a_n602_n100# a_n812_n100# 0.03fF
C433 a_752_n632# a_2012_n632# 0.00fF
C434 a_658_n100# a_660_n632# 0.00fF
C435 a_1172_n632# a_2012_n632# 0.01fF
C436 a_74_n401# a_122_n632# 0.00fF
C437 a_n3330_n632# a_n4170_n632# 0.01fF
C438 a_284_n729# a_1544_n729# 0.00fF
C439 a_912_131# a_960_n100# 0.00fF
C440 a_n348_131# a_492_131# 0.01fF
C441 a_912_131# a_282_n197# 0.00fF
C442 a_n3448_n632# a_n2818_n632# 0.01fF
C443 a_2970_n632# a_1802_n632# 0.01fF
C444 a_n2700_n632# a_n1230_n632# 0.00fF
C445 a_n3448_n632# a_n3120_n632# 0.02fF
C446 a_n3540_n632# a_n4078_n632# 0.01fF
C447 a_752_n632# a_240_n632# 0.01fF
C448 a_n2820_n100# a_n1652_n100# 0.01fF
C449 a_240_n632# a_1172_n632# 0.01fF
C450 a_n556_n729# a_n600_n632# 0.00fF
C451 a_960_n100# a_1380_n100# 0.02fF
C452 a_2220_n100# w_n4520_n851# 0.02fF
C453 a_962_n632# a_1080_n632# 0.07fF
C454 a_n2818_n632# a_n2608_n632# 0.03fF
C455 a_1498_n100# a_1170_n100# 0.02fF
C456 a_n3120_n632# a_n2608_n632# 0.01fF
C457 a_4018_n100# a_2430_n100# 0.00fF
C458 a_448_n100# a_960_n100# 0.01fF
C459 a_1500_n632# a_122_n632# 0.00fF
C460 a_n3496_n729# w_n4520_n851# 0.12fF
C461 a_1708_n100# a_2758_n100# 0.01fF
C462 a_n2400_n100# a_n2448_131# 0.00fF
C463 a_n510_n100# a_n1560_n100# 0.01fF
C464 a_n3540_n632# a_n4170_n632# 0.01fF
C465 a_n180_n632# a_n600_n632# 0.02fF
C466 a_332_n632# a_962_n632# 0.01fF
C467 a_2968_n100# a_3388_n100# 0.02fF
C468 a_542_n632# a_1382_n632# 0.01fF
C469 a_n3076_n729# a_n3078_n197# 0.01fF
C470 a_n3238_n632# a_n2398_n632# 0.01fF
C471 a_2970_n632# a_2760_n632# 0.03fF
C472 a_n1560_n100# a_n1022_n100# 0.01fF
C473 a_704_n729# a_n766_n401# 0.00fF
C474 a_n348_131# a_n1398_n197# 0.00fF
C475 a_2852_n632# a_3062_n632# 0.03fF
C476 a_3390_n632# a_2340_n632# 0.01fF
C477 a_n976_n729# a_n1186_n401# 0.00fF
C478 a_n1818_n197# a_n1816_n729# 0.01fF
C479 a_2220_n100# a_750_n100# 0.00fF
C480 a_4062_n197# a_4020_n632# 0.00fF
C481 a_2222_n632# a_1080_n632# 0.01fF
C482 a_n1860_n632# a_n1818_n197# 0.00fF
C483 a_n392_n100# w_n4520_n851# 0.02fF
C484 a_n1186_n401# a_n2236_n729# 0.00fF
C485 a_n2912_n100# a_n2492_n100# 0.02fF
C486 a_n1818_n197# a_n558_n197# 0.00fF
C487 a_n2400_n100# a_n3752_n100# 0.00fF
C488 a_28_n100# a_n812_n100# 0.01fF
C489 a_n3030_n100# a_n1862_n100# 0.01fF
C490 a_2642_n632# a_1080_n632# 0.00fF
C491 a_n390_n632# a_1080_n632# 0.00fF
C492 a_2970_n632# a_3482_n632# 0.01fF
C493 a_284_n729# a_330_n100# 0.00fF
C494 a_n90_n100# a_1498_n100# 0.00fF
C495 a_870_n632# a_n88_n632# 0.01fF
C496 a_1918_n100# w_n4520_n851# 0.02fF
C497 a_n2282_n100# a_n2492_n100# 0.03fF
C498 a_1802_n632# a_1920_n632# 0.07fF
C499 a_n720_n100# a_n1560_n100# 0.01fF
C500 a_n390_n632# a_332_n632# 0.01fF
C501 a_1800_n100# a_2430_n100# 0.01fF
C502 a_3388_n100# a_3178_n100# 0.03fF
C503 a_1964_n729# a_3434_n401# 0.00fF
C504 a_n3332_n100# a_n3030_n100# 0.02fF
C505 a_n1560_n100# a_n1980_n100# 0.02fF
C506 a_450_n632# a_n298_n632# 0.01fF
C507 a_1332_131# a_492_131# 0.01fF
C508 a_n3706_n401# a_n4126_n401# 0.01fF
C509 a_n392_n100# a_750_n100# 0.01fF
C510 a_2550_n632# a_1710_n632# 0.01fF
C511 a_n3332_n100# a_n3870_n100# 0.01fF
C512 a_n2608_n632# a_n1768_n632# 0.01fF
C513 a_n1350_n100# a_n1232_n100# 0.07fF
C514 a_2804_n729# a_2802_n197# 0.01fF
C515 a_n88_n632# a_660_n632# 0.01fF
C516 a_2850_n100# a_3060_n100# 0.03fF
C517 a_n2190_n100# a_n2072_n100# 0.07fF
C518 a_1962_n197# a_2592_131# 0.00fF
C519 a_n3542_n100# a_n3450_n100# 0.09fF
C520 a_n1348_n632# a_n1558_n632# 0.03fF
C521 a_2128_n100# a_2430_n100# 0.02fF
C522 a_1918_n100# a_750_n100# 0.01fF
C523 a_n3542_n100# a_n2702_n100# 0.01fF
C524 a_494_n401# a_n976_n729# 0.00fF
C525 a_2760_n632# a_1920_n632# 0.01fF
C526 a_450_n632# a_n508_n632# 0.01fF
C527 a_2432_n632# a_2340_n632# 0.09fF
C528 a_n2490_n632# a_n3960_n632# 0.00fF
C529 a_2968_n100# a_3480_n100# 0.01fF
C530 a_1802_n632# a_2012_n632# 0.03fF
C531 a_n2190_n100# a_n2238_n197# 0.00fF
C532 a_n810_n632# a_n1768_n632# 0.01fF
C533 a_120_n100# a_1170_n100# 0.01fF
C534 a_n1980_n100# a_n3450_n100# 0.00fF
C535 a_914_n401# a_1544_n729# 0.00fF
C536 a_n1980_n100# a_n2702_n100# 0.01fF
C537 a_n2656_n729# a_n2866_n401# 0.00fF
C538 a_494_n401# a_1334_n401# 0.01fF
C539 a_542_n632# a_n600_n632# 0.01fF
C540 a_n1348_n632# a_n2280_n632# 0.01fF
C541 a_960_n100# a_2430_n100# 0.00fF
C542 a_1332_131# a_1542_n197# 0.00fF
C543 a_1920_n632# a_3482_n632# 0.00fF
C544 a_2640_n100# a_1498_n100# 0.01fF
C545 a_n2070_n632# a_n1020_n632# 0.01fF
C546 a_240_n632# a_1802_n632# 0.00fF
C547 a_n510_n100# a_n930_n100# 0.02fF
C548 a_3014_n401# a_3224_n729# 0.00fF
C549 a_n2658_n197# a_n3288_131# 0.00fF
C550 a_1498_n100# a_1542_n197# 0.00fF
C551 a_494_n401# a_540_n100# 0.00fF
C552 a_2010_n100# a_3270_n100# 0.00fF
C553 a_n1022_n100# a_n930_n100# 0.09fF
C554 a_2760_n632# a_2012_n632# 0.01fF
C555 w_n4520_n851# a_n812_n100# 0.02fF
C556 a_1290_n632# a_1710_n632# 0.02fF
C557 a_n602_n100# a_28_n100# 0.01fF
C558 a_2430_n100# a_3808_n100# 0.00fF
C559 a_3852_131# a_3432_131# 0.01fF
C560 a_n2238_n197# a_n3078_n197# 0.01fF
C561 a_4110_n100# a_3060_n100# 0.01fF
C562 a_n976_n729# a_n1606_n401# 0.00fF
C563 a_n3330_n632# a_n3960_n632# 0.01fF
C564 a_n2238_n197# a_n2448_131# 0.00fF
C565 a_n180_n632# a_240_n632# 0.02fF
C566 a_n928_n632# a_n1138_n632# 0.03fF
C567 a_n1606_n401# a_n2236_n729# 0.00fF
C568 a_n718_n632# a_n810_n632# 0.09fF
C569 a_1592_n632# a_2130_n632# 0.01fF
C570 a_4062_n197# a_3432_131# 0.00fF
C571 a_n88_n632# a_122_n632# 0.03fF
C572 a_2852_n632# a_3272_n632# 0.02fF
C573 a_2852_n632# a_1500_n632# 0.00fF
C574 a_240_n632# a_238_n100# 0.00fF
C575 a_3480_n100# a_3178_n100# 0.02fF
C576 a_n1560_n100# a_n1652_n100# 0.09fF
C577 a_n1978_n632# a_n390_n632# 0.00fF
C578 a_120_n100# a_n90_n100# 0.03fF
C579 a_2012_n632# a_3482_n632# 0.00fF
C580 a_1590_n100# a_868_n100# 0.01fF
C581 a_1288_n100# a_2850_n100# 0.00fF
C582 a_n720_n100# a_n930_n100# 0.03fF
C583 a_3852_131# w_n4520_n851# 0.11fF
C584 a_n3448_n632# a_n1860_n632# 0.00fF
C585 a_n508_n632# a_n298_n632# 0.03fF
C586 a_n3540_n632# a_n3960_n632# 0.02fF
C587 a_n3122_n100# a_n2492_n100# 0.01fF
C588 a_3014_n401# a_2804_n729# 0.00fF
C589 a_750_n100# a_n812_n100# 0.00fF
C590 a_3692_n632# a_3180_n632# 0.01fF
C591 a_n930_n100# a_n1980_n100# 0.01fF
C592 a_n4078_n632# a_n3750_n632# 0.02fF
C593 a_542_n632# a_1920_n632# 0.00fF
C594 a_4062_n197# w_n4520_n851# 0.10fF
C595 a_1170_n100# a_1078_n100# 0.09fF
C596 a_n3240_n100# a_n2492_n100# 0.01fF
C597 a_n1860_n632# a_n2608_n632# 0.01fF
C598 a_658_n100# a_1170_n100# 0.01fF
C599 a_2220_n100# a_2548_n100# 0.02fF
C600 a_1544_n729# a_1592_n632# 0.00fF
C601 a_n2026_n401# a_n3286_n401# 0.00fF
C602 a_1590_n100# a_3060_n100# 0.00fF
C603 a_n1230_n632# a_122_n632# 0.00fF
C604 a_n2818_n632# a_n3028_n632# 0.03fF
C605 a_n3120_n632# a_n3028_n632# 0.09fF
C606 a_n2070_n632# a_n1440_n632# 0.01fF
C607 a_450_n632# w_n4520_n851# 0.01fF
C608 a_n1232_n100# a_n1230_n632# 0.00fF
C609 a_n1348_n632# a_n1396_n729# 0.00fF
C610 a_n2702_n100# a_n1652_n100# 0.01fF
C611 a_n1980_n100# a_n2028_131# 0.00fF
C612 a_2758_n100# a_3690_n100# 0.01fF
C613 a_n2446_n401# a_n1186_n401# 0.00fF
C614 a_n1232_n100# a_n1770_n100# 0.01fF
C615 a_n1350_n100# a_n2492_n100# 0.01fF
C616 a_n3750_n632# a_n4170_n632# 0.02fF
C617 a_n1860_n632# a_n810_n632# 0.01fF
C618 a_n3238_n632# a_n3868_n632# 0.01fF
C619 a_n2400_n100# a_n2610_n100# 0.03fF
C620 a_1590_n100# a_540_n100# 0.01fF
C621 a_2550_n632# a_1080_n632# 0.00fF
C622 a_2384_n729# a_3224_n729# 0.01fF
C623 a_n3332_n100# a_n3288_131# 0.00fF
C624 a_542_n632# a_2012_n632# 0.00fF
C625 a_448_n100# a_n930_n100# 0.00fF
C626 a_n1560_n100# a_n1558_n632# 0.00fF
C627 a_450_n632# a_752_n632# 0.02fF
C628 a_3598_n100# a_3600_n632# 0.00fF
C629 a_450_n632# a_1172_n632# 0.01fF
C630 a_n602_n100# w_n4520_n851# 0.02fF
C631 a_n3030_n100# a_n3962_n100# 0.01fF
C632 a_238_n100# a_n392_n100# 0.01fF
C633 a_n90_n100# a_1078_n100# 0.01fF
C634 a_658_n100# a_n90_n100# 0.01fF
C635 a_2594_n401# a_2592_131# 0.01fF
C636 a_3600_n632# a_2130_n632# 0.00fF
C637 a_n3870_n100# a_n3962_n100# 0.09fF
C638 a_3900_n100# a_3690_n100# 0.03fF
C639 a_542_n632# a_240_n632# 0.02fF
C640 a_3224_n729# a_4064_n729# 0.01fF
C641 a_1918_n100# a_2548_n100# 0.01fF
C642 w_n4520_n851# a_4020_n632# 0.08fF
C643 a_2758_n100# a_1170_n100# 0.00fF
C644 a_n390_n632# a_n1650_n632# 0.00fF
C645 a_n1816_n729# a_n1186_n401# 0.00fF
C646 a_n3448_n632# a_n2910_n632# 0.01fF
C647 a_3388_n100# a_2430_n100# 0.01fF
C648 a_n2490_n632# a_n928_n632# 0.00fF
C649 a_n3706_n401# a_n2866_n401# 0.01fF
C650 a_n1188_131# a_n2658_n197# 0.00fF
C651 a_n930_n100# a_n1652_n100# 0.01fF
C652 a_750_n100# a_n602_n100# 0.00fF
C653 a_n3448_n632# a_n2700_n632# 0.01fF
C654 a_n2910_n632# a_n2608_n632# 0.02fF
C655 a_912_131# a_2382_n197# 0.00fF
C656 w_n4520_n851# a_n298_n632# 0.01fF
C657 a_1288_n100# a_1590_n100# 0.02fF
C658 a_2338_n100# a_3270_n100# 0.01fF
C659 a_2804_n729# a_2384_n729# 0.01fF
C660 a_n1350_n100# a_n90_n100# 0.00fF
C661 a_n1768_n632# a_n3028_n632# 0.00fF
C662 a_n1140_n100# a_n182_n100# 0.01fF
C663 a_1500_n632# a_1542_n197# 0.00fF
C664 a_3598_n100# a_2850_n100# 0.01fF
C665 a_n2700_n632# a_n2608_n632# 0.09fF
C666 a_1080_n632# a_1290_n632# 0.03fF
C667 a_2128_n100# a_2172_131# 0.00fF
C668 a_n2820_n100# a_n3030_n100# 0.03fF
C669 a_870_n632# a_914_n401# 0.00fF
C670 a_2804_n729# a_4064_n729# 0.00fF
C671 a_n3660_n100# a_n3542_n100# 0.07fF
C672 a_2970_n632# a_3062_n632# 0.09fF
C673 a_n1138_n632# a_n1768_n632# 0.01fF
C674 a_n2820_n100# a_n3870_n100# 0.01fF
C675 a_n510_n100# a_868_n100# 0.00fF
C676 a_332_n632# a_1290_n632# 0.01fF
C677 a_n508_n632# w_n4520_n851# 0.01fF
C678 a_n2190_n100# a_n812_n100# 0.00fF
C679 a_2968_n100# a_3060_n100# 0.09fF
C680 a_30_n632# a_n928_n632# 0.01fF
C681 a_n3332_n100# a_n1862_n100# 0.00fF
C682 a_752_n632# a_n298_n632# 0.01fF
C683 a_n928_n632# a_n2188_n632# 0.00fF
C684 a_1172_n632# a_n298_n632# 0.00fF
C685 w_n4520_n851# a_28_n100# 0.02fF
C686 a_2640_n100# a_1078_n100# 0.00fF
C687 a_n2912_n100# a_n2400_n100# 0.01fF
C688 a_n1020_n632# a_n88_n632# 0.01fF
C689 a_n2446_n401# a_n1606_n401# 0.01fF
C690 a_n3916_n729# a_n3960_n632# 0.00fF
C691 a_n1140_n100# a_n1442_n100# 0.02fF
C692 w_n4520_n851# a_n1608_131# 0.12fF
C693 a_n2818_n632# a_n2490_n632# 0.02fF
C694 a_n2400_n100# a_n2282_n100# 0.07fF
C695 a_n3120_n632# a_n2490_n632# 0.01fF
C696 a_n1770_n100# a_n2492_n100# 0.01fF
C697 a_1382_n632# a_1500_n632# 0.07fF
C698 a_752_n632# a_n508_n632# 0.00fF
C699 a_n2188_n632# a_n2236_n729# 0.00fF
C700 a_n2072_n100# a_n2610_n100# 0.01fF
C701 a_3598_n100# a_4110_n100# 0.01fF
C702 a_238_n100# a_n812_n100# 0.01fF
C703 a_n1348_n632# a_n1978_n632# 0.01fF
C704 a_4018_n100# a_3270_n100# 0.01fF
C705 a_494_n401# a_1544_n729# 0.00fF
C706 a_n718_n632# a_n1138_n632# 0.02fF
C707 a_750_n100# a_28_n100# 0.01fF
C708 a_n720_n100# a_868_n100# 0.00fF
C709 a_n1350_n100# a_n1398_n197# 0.00fF
C710 a_3480_n100# a_2430_n100# 0.01fF
C711 a_n1020_n632# a_n1230_n632# 0.03fF
C712 a_n1188_131# a_n768_131# 0.01fF
C713 a_n88_n632# a_n90_n100# 0.00fF
C714 a_3692_n632# a_3690_n100# 0.00fF
C715 a_n510_n100# a_540_n100# 0.01fF
C716 a_n3286_n401# a_n3288_131# 0.01fF
C717 a_3060_n100# a_3178_n100# 0.07fF
C718 a_450_n632# a_1802_n632# 0.00fF
C719 a_3224_n729# a_3270_n100# 0.00fF
C720 a_3390_n632# a_2130_n632# 0.00fF
C721 a_n1022_n100# a_540_n100# 0.00fF
C722 w_n4520_n851# a_3432_131# 0.12fF
C723 a_n1816_n729# a_n1606_n401# 0.00fF
C724 a_n3330_n632# a_n2818_n632# 0.01fF
C725 a_3062_n632# a_1920_n632# 0.01fF
C726 a_n3120_n632# a_n3330_n632# 0.03fF
C727 a_n2818_n632# a_n2188_n632# 0.01fF
C728 a_n3120_n632# a_n2188_n632# 0.01fF
C729 a_870_n632# a_1592_n632# 0.01fF
C730 a_n3750_n632# a_n3960_n632# 0.03fF
C731 a_2338_n100# a_2010_n100# 0.02fF
C732 a_2640_n100# a_2758_n100# 0.07fF
C733 a_3854_n401# a_3224_n729# 0.00fF
C734 a_n1860_n632# a_n3028_n632# 0.01fF
C735 a_912_131# a_868_n100# 0.00fF
C736 a_n2070_n632# a_n600_n632# 0.00fF
C737 a_450_n632# a_n180_n632# 0.01fF
C738 a_n88_n632# a_n1440_n632# 0.00fF
C739 a_n392_n100# a_n348_131# 0.00fF
C740 a_n2868_131# a_n3288_131# 0.01fF
C741 a_1592_n632# a_3180_n632# 0.00fF
C742 a_1380_n100# a_868_n100# 0.01fF
C743 a_n2190_n100# a_n602_n100# 0.00fF
C744 a_n2868_131# a_n2658_n197# 0.00fF
C745 a_2340_n632# a_1710_n632# 0.01fF
C746 a_2382_n197# a_3642_n197# 0.00fF
C747 a_n1860_n632# a_n1138_n632# 0.01fF
C748 a_1800_n100# a_3270_n100# 0.00fF
C749 a_n3540_n632# a_n2818_n632# 0.01fF
C750 a_n720_n100# a_540_n100# 0.00fF
C751 a_448_n100# a_868_n100# 0.02fF
C752 a_n3540_n632# a_n3120_n632# 0.02fF
C753 a_660_n632# a_1592_n632# 0.01fF
C754 a_1124_n729# a_1334_n401# 0.00fF
C755 a_2222_n632# a_962_n632# 0.00fF
C756 a_3062_n632# a_2012_n632# 0.01fF
C757 a_2852_n632# a_3692_n632# 0.01fF
C758 a_2382_n197# a_2430_n100# 0.00fF
C759 a_n2490_n632# a_n1768_n632# 0.01fF
C760 a_n390_n632# a_962_n632# 0.00fF
C761 a_2382_n197# a_2802_n197# 0.01fF
C762 a_2640_n100# a_3900_n100# 0.00fF
C763 a_n300_n100# a_n1862_n100# 0.00fF
C764 a_3854_n401# a_3810_n632# 0.00fF
C765 a_n768_131# a_n978_n197# 0.00fF
C766 a_2970_n632# a_1500_n632# 0.00fF
C767 a_n1440_n632# a_n1230_n632# 0.03fF
C768 a_2970_n632# a_3272_n632# 0.02fF
C769 a_n1140_n100# a_330_n100# 0.00fF
C770 a_n2912_n100# a_n2072_n100# 0.01fF
C771 a_2128_n100# a_3270_n100# 0.01fF
C772 a_238_n100# a_n602_n100# 0.01fF
C773 a_1544_n729# a_1590_n100# 0.00fF
C774 a_752_n632# w_n4520_n851# 0.01fF
C775 a_2804_n729# a_3854_n401# 0.00fF
C776 a_n1348_n632# a_n1650_n632# 0.02fF
C777 a_1172_n632# w_n4520_n851# 0.01fF
C778 a_1380_n100# a_1334_n401# 0.00fF
C779 a_750_n100# w_n4520_n851# 0.02fF
C780 a_2432_n632# a_2130_n632# 0.02fF
C781 a_n810_n632# a_660_n632# 0.00fF
C782 a_2220_n100# a_1498_n100# 0.01fF
C783 a_1334_n401# a_2174_n401# 0.01fF
C784 a_n2072_n100# a_n2282_n100# 0.03fF
C785 a_n3122_n100# a_n2400_n100# 0.01fF
C786 a_2760_n632# a_4020_n632# 0.00fF
C787 a_1380_n100# a_540_n100# 0.01fF
C788 a_n3330_n632# a_n1768_n632# 0.00fF
C789 a_n2188_n632# a_n1768_n632# 0.02fF
C790 a_28_n100# a_72_131# 0.00fF
C791 a_n1560_n100# a_n3030_n100# 0.00fF
C792 a_n2490_n632# a_n2446_n401# 0.00fF
C793 a_n2398_n632# w_n4520_n851# 0.01fF
C794 a_n3240_n100# a_n2400_n100# 0.01fF
C795 a_2222_n632# a_2642_n632# 0.02fF
C796 a_448_n100# a_540_n100# 0.09fF
C797 a_n180_n632# a_n298_n632# 0.07fF
C798 a_n2282_n100# a_n2238_n197# 0.00fF
C799 a_752_n632# a_1172_n632# 0.02fF
C800 a_n2910_n632# a_n3028_n632# 0.07fF
C801 a_n556_n729# a_n508_n632# 0.00fF
C802 a_n1188_131# a_n978_n197# 0.00fF
C803 a_752_n632# a_750_n100# 0.00fF
C804 a_1752_131# a_702_n197# 0.00fF
C805 a_914_n401# a_1964_n729# 0.00fF
C806 a_4020_n632# a_3482_n632# 0.01fF
C807 a_1592_n632# a_122_n632# 0.00fF
C808 a_n1350_n100# a_n2400_n100# 0.01fF
C809 a_3270_n100# a_3808_n100# 0.01fF
C810 a_n2700_n632# a_n3028_n632# 0.02fF
C811 a_3600_n632# a_3180_n632# 0.02fF
C812 a_n2070_n632# a_n2072_n100# 0.00fF
C813 a_n88_n632# a_1382_n632# 0.00fF
C814 a_450_n632# a_542_n632# 0.09fF
C815 a_702_n197# a_1122_n197# 0.01fF
C816 a_n180_n632# a_n508_n632# 0.02fF
C817 a_n3332_n100# a_n3962_n100# 0.01fF
C818 a_n510_n100# a_n182_n100# 0.02fF
C819 a_n136_n729# a_704_n729# 0.01fF
C820 a_n3030_n100# a_n3450_n100# 0.02fF
C821 a_2968_n100# a_3598_n100# 0.01fF
C822 a_1500_n632# a_1920_n632# 0.02fF
C823 a_30_n632# a_n718_n632# 0.01fF
C824 a_n3030_n100# a_n2702_n100# 0.02fF
C825 a_1920_n632# a_3272_n632# 0.00fF
C826 a_n2700_n632# a_n1138_n632# 0.00fF
C827 a_1590_n100# a_330_n100# 0.00fF
C828 a_2010_n100# a_1800_n100# 0.03fF
C829 a_1918_n100# a_1498_n100# 0.02fF
C830 a_n718_n632# a_n2188_n632# 0.00fF
C831 a_n1022_n100# a_n182_n100# 0.01fF
C832 a_238_n100# a_28_n100# 0.03fF
C833 a_n976_n729# a_n766_n401# 0.00fF
C834 a_n3870_n100# a_n3450_n100# 0.02fF
C835 a_n138_n197# a_702_n197# 0.01fF
C836 a_n3870_n100# a_n2702_n100# 0.01fF
C837 a_1288_n100# a_1380_n100# 0.09fF
C838 a_n810_n632# a_122_n632# 0.01fF
C839 a_n3708_131# a_n3706_n401# 0.01fF
C840 a_n766_n401# a_n2236_n729# 0.00fF
C841 a_n1860_n632# a_n2490_n632# 0.01fF
C842 a_2850_n100# a_1708_n100# 0.01fF
C843 a_1288_n100# a_448_n100# 0.01fF
C844 a_2430_n100# a_868_n100# 0.00fF
C845 a_n2070_n632# a_n3238_n632# 0.01fF
C846 a_n2820_n100# a_n1862_n100# 0.01fF
C847 a_n928_n632# a_n1558_n632# 0.01fF
C848 a_2128_n100# a_2010_n100# 0.07fF
C849 a_n3078_n197# a_n1608_131# 0.00fF
C850 a_n1608_131# a_n2448_131# 0.01fF
C851 a_n510_n100# a_n1442_n100# 0.01fF
C852 a_2012_n632# a_3272_n632# 0.00fF
C853 a_1500_n632# a_2012_n632# 0.01fF
C854 a_n720_n100# a_n182_n100# 0.01fF
C855 a_4112_n632# a_4064_n729# 0.00fF
C856 a_1124_n729# a_1122_n197# 0.01fF
C857 a_n1022_n100# a_n1442_n100# 0.02fF
C858 a_912_131# a_1752_131# 0.01fF
C859 a_3644_n729# a_3434_n401# 0.00fF
C860 a_n928_n632# a_n2280_n632# 0.00fF
C861 a_2340_n632# a_1080_n632# 0.00fF
C862 w_n4520_n851# a_72_131# 0.12fF
C863 a_n3332_n100# a_n2820_n100# 0.01fF
C864 a_n718_n632# a_n720_n100# 0.00fF
C865 a_3060_n100# a_2430_n100# 0.01fF
C866 a_960_n100# a_2010_n100# 0.01fF
C867 a_3598_n100# a_3178_n100# 0.02fF
C868 a_n3540_n632# a_n3498_n197# 0.00fF
C869 a_n3542_n100# a_n3498_n197# 0.00fF
C870 a_912_131# a_1122_n197# 0.00fF
C871 a_n1860_n632# a_n3330_n632# 0.00fF
C872 a_240_n632# a_1500_n632# 0.00fF
C873 a_n1860_n632# a_n2188_n632# 0.02fF
C874 a_542_n632# a_n298_n632# 0.01fF
C875 a_n510_n100# a_n558_n197# 0.00fF
C876 a_1802_n632# w_n4520_n851# 0.01fF
C877 a_n2190_n100# w_n4520_n851# 0.02fF
C878 a_n556_n729# w_n4520_n851# 0.12fF
C879 a_n3122_n100# a_n2072_n100# 0.01fF
C880 a_2640_n100# a_2592_131# 0.00fF
C881 a_n2656_n729# a_n3076_n729# 0.01fF
C882 a_n2280_n632# a_n2236_n729# 0.00fF
C883 a_1542_n197# a_2592_131# 0.00fF
C884 a_n558_n197# a_702_n197# 0.00fF
C885 a_n2026_n401# a_n2028_131# 0.01fF
C886 a_n3240_n100# a_n2072_n100# 0.01fF
C887 a_n88_n632# a_n600_n632# 0.01fF
C888 a_912_131# a_n138_n197# 0.00fF
C889 a_n720_n100# a_n1442_n100# 0.01fF
C890 a_1380_n100# a_n182_n100# 0.00fF
C891 a_n2818_n632# a_n1558_n632# 0.00fF
C892 a_n180_n632# w_n4520_n851# 0.01fF
C893 a_3902_n632# a_3854_n401# 0.00fF
C894 a_542_n632# a_n508_n632# 0.01fF
C895 a_n1442_n100# a_n1980_n100# 0.01fF
C896 a_n3120_n632# a_n1558_n632# 0.00fF
C897 a_n768_131# a_282_n197# 0.00fF
C898 a_n346_n401# a_n298_n632# 0.00fF
C899 a_120_n100# a_n392_n100# 0.01fF
C900 w_n4520_n851# a_2548_n100# 0.02fF
C901 a_752_n632# a_1802_n632# 0.01fF
C902 a_448_n100# a_n182_n100# 0.01fF
C903 a_n1350_n100# a_n2072_n100# 0.01fF
C904 a_2550_n632# a_962_n632# 0.00fF
C905 a_1172_n632# a_1802_n632# 0.01fF
C906 a_238_n100# w_n4520_n851# 0.02fF
C907 a_2760_n632# w_n4520_n851# 0.02fF
C908 a_n2818_n632# a_n3750_n632# 0.01fF
C909 a_n3120_n632# a_n3750_n632# 0.01fF
C910 a_3388_n100# a_3270_n100# 0.07fF
C911 a_n2400_n100# a_n1770_n100# 0.01fF
C912 a_n2490_n632# a_n2910_n632# 0.02fF
C913 a_3222_n197# a_2592_131# 0.00fF
C914 w_n4520_n851# a_n3078_n197# 0.10fF
C915 w_n4520_n851# a_n2448_131# 0.12fF
C916 a_2382_n197# a_2172_131# 0.00fF
C917 a_2382_n197# a_2384_n729# 0.01fF
C918 a_n2818_n632# a_n2280_n632# 0.01fF
C919 a_3390_n632# a_3180_n632# 0.03fF
C920 a_2222_n632# a_3810_n632# 0.00fF
C921 a_n3120_n632# a_n2280_n632# 0.01fF
C922 a_n1818_n197# a_n1398_n197# 0.01fF
C923 a_2384_n729# a_2340_n632# 0.00fF
C924 a_n2700_n632# a_n2490_n632# 0.03fF
C925 a_n1230_n632# a_n600_n632# 0.01fF
C926 a_2382_n197# a_3012_131# 0.00fF
C927 a_2642_n632# a_3810_n632# 0.01fF
C928 a_n3238_n632# a_n3240_n100# 0.00fF
C929 a_752_n632# a_n180_n632# 0.01fF
C930 a_960_n100# a_962_n632# 0.00fF
C931 a_1590_n100# a_1708_n100# 0.07fF
C932 a_n4080_n100# w_n4520_n851# 0.08fF
C933 a_n180_n632# a_1172_n632# 0.00fF
C934 w_n4520_n851# a_3482_n632# 0.03fF
C935 a_2852_n632# a_1592_n632# 0.00fF
C936 a_2220_n100# a_1078_n100# 0.01fF
C937 a_2220_n100# a_658_n100# 0.00fF
C938 a_2760_n632# a_1172_n632# 0.00fF
C939 a_n2866_n401# a_n1606_n401# 0.00fF
C940 a_1288_n100# a_2430_n100# 0.01fF
C941 a_238_n100# a_750_n100# 0.01fF
C942 a_n182_n100# a_n1652_n100# 0.00fF
C943 w_n4520_n851# a_n3752_n100# 0.04fF
C944 a_2222_n632# a_2550_n632# 0.02fF
C945 a_2338_n100# a_1800_n100# 0.01fF
C946 a_1544_n729# a_1124_n729# 0.01fF
C947 a_2174_n401# a_2130_n632# 0.00fF
C948 a_n1188_131# a_282_n197# 0.00fF
C949 a_n510_n100# a_330_n100# 0.01fF
C950 a_912_131# a_n558_n197# 0.00fF
C951 a_n3330_n632# a_n2910_n632# 0.02fF
C952 a_2642_n632# a_2550_n632# 0.09fF
C953 a_n2910_n632# a_n2188_n632# 0.01fF
C954 a_n1348_n632# a_n390_n632# 0.01fF
C955 a_n976_n729# a_n1396_n729# 0.01fF
C956 a_n1020_n632# a_n2608_n632# 0.00fF
C957 a_3014_n401# a_3060_n100# 0.00fF
C958 w_n4520_n851# a_n3868_n632# 0.05fF
C959 a_n1022_n100# a_330_n100# 0.00fF
C960 a_n1140_n100# a_n1232_n100# 0.09fF
C961 a_n2700_n632# a_n3330_n632# 0.01fF
C962 a_n2700_n632# a_n2188_n632# 0.01fF
C963 a_962_n632# a_1290_n632# 0.02fF
C964 a_n1396_n729# a_n2236_n729# 0.01fF
C965 a_870_n632# a_2432_n632# 0.00fF
C966 a_n2702_n100# a_n2658_n197# 0.00fF
C967 a_n2282_n100# a_n812_n100# 0.00fF
C968 a_1962_n197# a_702_n197# 0.00fF
C969 a_2338_n100# a_2128_n100# 0.03fF
C970 a_1710_n632# a_1752_131# 0.00fF
C971 a_n1768_n632# a_n1558_n632# 0.03fF
C972 a_n1020_n632# a_n810_n632# 0.03fF
C973 a_658_n100# a_n392_n100# 0.01fF
C974 a_n392_n100# a_1078_n100# 0.00fF
C975 a_332_n632# a_n928_n632# 0.00fF
C976 a_n348_131# a_n1608_131# 0.00fF
C977 a_1544_n729# a_2174_n401# 0.00fF
C978 a_n3916_n729# a_n2446_n401# 0.00fF
C979 a_n1442_n100# a_n1652_n100# 0.03fF
C980 a_n3540_n632# a_n2910_n632# 0.01fF
C981 a_2970_n632# a_3692_n632# 0.01fF
C982 a_2432_n632# a_3180_n632# 0.01fF
C983 a_n718_n632# a_n766_n401# 0.00fF
C984 a_542_n632# w_n4520_n851# 0.01fF
C985 a_3480_n100# a_3270_n100# 0.03fF
C986 a_n3658_n632# a_n4078_n632# 0.02fF
C987 a_2802_n197# a_1752_131# 0.00fF
C988 a_1918_n100# a_1078_n100# 0.01fF
C989 a_n3540_n632# a_n2700_n632# 0.01fF
C990 a_n720_n100# a_330_n100# 0.01fF
C991 a_1918_n100# a_658_n100# 0.00fF
C992 a_n2280_n632# a_n1768_n632# 0.01fF
C993 a_2338_n100# a_960_n100# 0.00fF
C994 a_n1560_n100# a_n1862_n100# 0.02fF
C995 a_120_n100# a_n812_n100# 0.01fF
C996 a_2220_n100# a_2758_n100# 0.01fF
C997 a_2010_n100# a_3388_n100# 0.00fF
C998 a_2222_n632# a_1290_n632# 0.01fF
C999 a_n3660_n100# a_n3030_n100# 0.01fF
C1000 a_n1138_n632# a_122_n632# 0.00fF
C1001 a_2642_n632# a_1290_n632# 0.00fF
C1002 a_n2398_n632# a_n3868_n632# 0.00fF
C1003 a_494_n401# a_1964_n729# 0.00fF
C1004 a_n978_n197# a_282_n197# 0.00fF
C1005 a_n88_n632# a_240_n632# 0.02fF
C1006 a_n1350_n100# a_n392_n100# 0.01fF
C1007 a_n2820_n100# a_n3962_n100# 0.01fF
C1008 a_n3658_n632# a_n4170_n632# 0.01fF
C1009 a_2850_n100# a_3690_n100# 0.01fF
C1010 a_n3870_n100# a_n3660_n100# 0.03fF
C1011 a_n300_n100# a_960_n100# 0.00fF
C1012 a_n2820_n100# a_n2868_131# 0.00fF
C1013 a_2338_n100# a_3808_n100# 0.00fF
C1014 a_2852_n632# a_3600_n632# 0.01fF
C1015 a_1754_n401# w_n4520_n851# 0.10fF
C1016 a_n346_n401# w_n4520_n851# 0.10fF
C1017 a_n718_n632# a_n1558_n632# 0.01fF
C1018 a_542_n632# a_752_n632# 0.03fF
C1019 a_n2072_n100# a_n1770_n100# 0.02fF
C1020 a_542_n632# a_1172_n632# 0.01fF
C1021 a_n1440_n632# a_n2608_n632# 0.01fF
C1022 a_n3542_n100# a_n4172_n100# 0.01fF
C1023 a_3062_n632# a_4020_n632# 0.01fF
C1024 a_n3706_n401# a_n3076_n729# 0.00fF
C1025 a_n1862_n100# a_n3450_n100# 0.00fF
C1026 a_n1816_n729# a_n766_n401# 0.00fF
C1027 a_n1862_n100# a_n2702_n100# 0.01fF
C1028 a_2968_n100# a_1708_n100# 0.00fF
C1029 a_912_131# a_1962_n197# 0.00fF
C1030 a_3598_n100# a_3642_n197# 0.00fF
C1031 a_1380_n100# a_330_n100# 0.01fF
C1032 a_n718_n632# a_n2280_n632# 0.00fF
C1033 a_1710_n632# a_2130_n632# 0.02fF
C1034 a_n3288_131# a_n2028_131# 0.00fF
C1035 a_n810_n632# a_n1440_n632# 0.01fF
C1036 a_2804_n729# a_3224_n729# 0.01fF
C1037 a_3598_n100# a_2430_n100# 0.01fF
C1038 a_448_n100# a_330_n100# 0.07fF
C1039 a_240_n632# a_n1230_n632# 0.00fF
C1040 w_n4520_n851# a_n348_131# 0.12fF
C1041 a_n2658_n197# a_n2028_131# 0.00fF
C1042 a_870_n632# a_30_n632# 0.01fF
C1043 a_n976_n729# a_n2026_n401# 0.00fF
C1044 a_3060_n100# a_3012_131# 0.00fF
C1045 a_1918_n100# a_2758_n100# 0.01fF
C1046 a_n3332_n100# a_n3450_n100# 0.07fF
C1047 a_28_n100# a_1498_n100# 0.00fF
C1048 a_2384_n729# a_1334_n401# 0.00fF
C1049 a_n3496_n729# a_n2656_n729# 0.01fF
C1050 a_n3332_n100# a_n2702_n100# 0.01fF
C1051 a_2760_n632# a_1802_n632# 0.01fF
C1052 a_n2026_n401# a_n2236_n729# 0.00fF
C1053 a_4110_n100# a_3690_n100# 0.02fF
C1054 a_2852_n632# a_2850_n100# 0.00fF
C1055 a_n1978_n632# a_n928_n632# 0.01fF
C1056 a_658_n100# a_n812_n100# 0.00fF
C1057 a_n1860_n632# a_n1558_n632# 0.02fF
C1058 a_n1140_n100# a_n2492_n100# 0.00fF
C1059 a_4018_n100# a_3808_n100# 0.03fF
C1060 a_3480_n100# a_2010_n100# 0.00fF
C1061 a_3902_n632# a_2642_n632# 0.00fF
C1062 a_120_n100# a_n602_n100# 0.01fF
C1063 a_30_n632# a_660_n632# 0.01fF
C1064 a_1708_n100# a_3178_n100# 0.00fF
C1065 a_2128_n100# a_1800_n100# 0.02fF
C1066 a_2550_n632# a_3810_n632# 0.00fF
C1067 a_n1860_n632# a_n2280_n632# 0.02fF
C1068 a_450_n632# a_1500_n632# 0.01fF
C1069 a_n3916_n729# a_n4126_n401# 0.00fF
C1070 a_660_n632# a_702_n197# 0.00fF
C1071 a_n2190_n100# a_n3752_n100# 0.00fF
C1072 a_n930_n100# a_n1862_n100# 0.01fF
C1073 a_3178_n100# a_3180_n632# 0.00fF
C1074 a_1382_n632# a_1592_n632# 0.03fF
C1075 a_n3078_n197# a_n2448_131# 0.00fF
C1076 a_3644_n729# a_3692_n632# 0.00fF
C1077 w_n4520_n851# a_n2610_n100# 0.02fF
C1078 a_n1350_n100# a_n812_n100# 0.01fF
C1079 a_2760_n632# a_3482_n632# 0.01fF
C1080 a_960_n100# a_1800_n100# 0.01fF
C1081 a_284_n729# a_240_n632# 0.00fF
C1082 a_n2446_n401# a_n1396_n729# 0.00fF
C1083 a_1080_n632# a_1122_n197# 0.00fF
C1084 a_n300_n100# a_n1560_n100# 0.00fF
C1085 a_n1978_n632# a_n2818_n632# 0.01fF
C1086 a_n392_n100# a_n1770_n100# 0.00fF
C1087 a_n1978_n632# a_n3120_n632# 0.01fF
C1088 a_n768_131# a_n2028_131# 0.00fF
C1089 a_870_n632# a_912_131# 0.00fF
C1090 a_2338_n100# a_3388_n100# 0.01fF
C1091 w_n4520_n851# a_1332_131# 0.12fF
C1092 a_3810_n632# a_3808_n100# 0.00fF
C1093 a_2852_n632# a_3390_n632# 0.01fF
C1094 a_n1140_n100# a_n90_n100# 0.01fF
C1095 a_2128_n100# a_960_n100# 0.01fF
C1096 w_n4520_n851# a_1498_n100# 0.02fF
C1097 a_542_n632# a_1802_n632# 0.00fF
C1098 a_3272_n632# a_4020_n632# 0.01fF
C1099 a_1380_n100# a_1708_n100# 0.02fF
C1100 a_30_n632# a_122_n632# 0.09fF
C1101 a_n4080_n100# a_n3752_n100# 0.02fF
C1102 a_n2070_n632# a_n508_n632# 0.00fF
C1103 a_n2910_n632# a_n1558_n632# 0.00fF
C1104 a_494_n401# a_492_131# 0.01fF
C1105 a_120_n100# a_28_n100# 0.09fF
C1106 a_n1020_n632# a_n1138_n632# 0.07fF
C1107 a_1590_n100# a_1170_n100# 0.02fF
C1108 a_n1650_n632# a_n928_n632# 0.01fF
C1109 a_n510_n100# a_n1232_n100# 0.01fF
C1110 a_448_n100# a_1708_n100# 0.00fF
C1111 a_658_n100# a_n602_n100# 0.00fF
C1112 a_n718_n632# a_332_n632# 0.01fF
C1113 a_1124_n729# a_2594_n401# 0.00fF
C1114 a_n2700_n632# a_n1558_n632# 0.01fF
C1115 a_n1818_n197# a_n2238_n197# 0.01fF
C1116 a_3062_n632# w_n4520_n851# 0.03fF
C1117 a_542_n632# a_n180_n632# 0.01fF
C1118 a_n2910_n632# a_n3750_n632# 0.01fF
C1119 a_n1816_n729# a_n1396_n729# 0.01fF
C1120 a_n3658_n632# a_n3960_n632# 0.02fF
C1121 a_4112_n632# a_2642_n632# 0.00fF
C1122 a_2172_131# a_1752_131# 0.01fF
C1123 a_n1022_n100# a_n1232_n100# 0.03fF
C1124 a_2802_n197# a_1962_n197# 0.01fF
C1125 a_1802_n632# a_1754_n401# 0.00fF
C1126 a_n2910_n632# a_n2280_n632# 0.01fF
C1127 a_n1188_131# a_n2028_131# 0.01fF
C1128 a_n2700_n632# a_n3750_n632# 0.01fF
C1129 a_1752_131# a_3012_131# 0.00fF
C1130 a_n556_n729# a_n346_n401# 0.00fF
C1131 a_2550_n632# a_1290_n632# 0.00fF
C1132 a_750_n100# a_1498_n100# 0.01fF
C1133 a_1080_n632# a_2130_n632# 0.01fF
C1134 a_2640_n100# a_2850_n100# 0.03fF
C1135 a_3060_n100# a_3270_n100# 0.03fF
C1136 a_2172_131# a_1122_n197# 0.00fF
C1137 a_3014_n401# a_1544_n729# 0.00fF
C1138 a_n2700_n632# a_n2280_n632# 0.02fF
C1139 a_n348_131# a_72_131# 0.01fF
C1140 a_2970_n632# a_1592_n632# 0.00fF
C1141 a_4018_n100# a_3388_n100# 0.01fF
C1142 a_n1350_n100# a_n602_n100# 0.01fF
C1143 a_2594_n401# a_2174_n401# 0.01fF
C1144 a_n2912_n100# w_n4520_n851# 0.03fF
C1145 a_n3496_n729# a_n3706_n401# 0.00fF
C1146 a_3852_131# a_3900_n100# 0.00fF
C1147 a_2852_n632# a_2432_n632# 0.02fF
C1148 a_n720_n100# a_n1232_n100# 0.01fF
C1149 a_n1440_n632# a_n3028_n632# 0.00fF
C1150 a_n1978_n632# a_n1768_n632# 0.03fF
C1151 a_2340_n632# a_962_n632# 0.00fF
C1152 a_n3450_n100# a_n3962_n100# 0.01fF
C1153 a_n2702_n100# a_n3962_n100# 0.00fF
C1154 a_n1232_n100# a_n1980_n100# 0.01fF
C1155 w_n4520_n851# a_n2282_n100# 0.02fF
C1156 a_2338_n100# a_3480_n100# 0.01fF
C1157 a_2968_n100# a_3690_n100# 0.01fF
C1158 a_n2446_n401# a_n2026_n401# 0.01fF
C1159 a_n2818_n632# a_n1650_n632# 0.01fF
C1160 a_n3120_n632# a_n1650_n632# 0.00fF
C1161 a_n930_n100# a_n978_n197# 0.00fF
C1162 a_n810_n632# a_n600_n632# 0.03fF
C1163 a_n1770_n100# a_n812_n100# 0.01fF
C1164 a_n1440_n632# a_n1138_n632# 0.02fF
C1165 a_n2820_n100# a_n1560_n100# 0.00fF
C1166 a_3902_n632# a_3810_n632# 0.09fF
C1167 a_n300_n100# a_n930_n100# 0.01fF
C1168 a_2640_n100# a_4110_n100# 0.00fF
C1169 a_28_n100# a_1078_n100# 0.01fF
C1170 a_658_n100# a_28_n100# 0.01fF
C1171 a_n2490_n632# a_n2492_n100# 0.00fF
C1172 a_450_n632# a_n88_n632# 0.01fF
C1173 a_2172_131# a_2130_n632# 0.00fF
C1174 a_n978_n197# a_n2028_131# 0.00fF
C1175 a_2010_n100# a_868_n100# 0.01fF
C1176 a_120_n100# w_n4520_n851# 0.02fF
C1177 a_870_n632# a_1710_n632# 0.01fF
C1178 a_3434_n401# a_3432_131# 0.01fF
C1179 a_2222_n632# a_2340_n632# 0.07fF
C1180 a_n2070_n632# w_n4520_n851# 0.01fF
C1181 a_n3332_n100# a_n3660_n100# 0.02fF
C1182 a_1708_n100# a_1710_n632# 0.00fF
C1183 a_3902_n632# a_2550_n632# 0.00fF
C1184 a_n1978_n632# a_n718_n632# 0.00fF
C1185 a_3388_n100# a_1800_n100# 0.00fF
C1186 a_2642_n632# a_2340_n632# 0.02fF
C1187 a_1592_n632# a_1920_n632# 0.02fF
C1188 w_n4520_n851# a_74_n401# 0.10fF
C1189 a_n2820_n100# a_n3450_n100# 0.01fF
C1190 a_n976_n729# a_n136_n729# 0.01fF
C1191 a_n2190_n100# a_n2610_n100# 0.02fF
C1192 a_n3030_n100# a_n1442_n100# 0.00fF
C1193 a_n1020_n632# a_n2490_n632# 0.00fF
C1194 a_n2820_n100# a_n2702_n100# 0.07fF
C1195 a_n1350_n100# a_28_n100# 0.00fF
C1196 a_1710_n632# a_3180_n632# 0.00fF
C1197 a_n2026_n401# a_n1816_n729# 0.00fF
C1198 a_1708_n100# a_2430_n100# 0.01fF
C1199 a_3690_n100# a_3178_n100# 0.01fF
C1200 a_2010_n100# a_3060_n100# 0.01fF
C1201 a_2970_n632# a_3600_n632# 0.01fF
C1202 a_2338_n100# a_2382_n197# 0.00fF
C1203 a_1544_n729# a_2384_n729# 0.01fF
C1204 a_1332_131# a_72_131# 0.00fF
C1205 a_2640_n100# a_1590_n100# 0.01fF
C1206 a_4018_n100# a_3480_n100# 0.01fF
C1207 w_n4520_n851# a_3434_n401# 0.09fF
C1208 a_2338_n100# a_2340_n632# 0.00fF
C1209 a_2128_n100# a_3388_n100# 0.00fF
C1210 a_n3658_n632# a_n3660_n100# 0.00fF
C1211 a_n3916_n729# a_n2866_n401# 0.00fF
C1212 a_1590_n100# a_1542_n197# 0.00fF
C1213 a_n136_n729# a_1334_n401# 0.00fF
C1214 a_660_n632# a_1710_n632# 0.01fF
C1215 a_120_n100# a_750_n100# 0.01fF
C1216 a_1500_n632# w_n4520_n851# 0.01fF
C1217 w_n4520_n851# a_3272_n632# 0.03fF
C1218 a_n1022_n100# a_n2492_n100# 0.00fF
C1219 a_1124_n729# a_1964_n729# 0.01fF
C1220 a_n3962_n100# a_n3960_n632# 0.00fF
C1221 a_332_n632# a_330_n100# 0.00fF
C1222 a_2010_n100# a_540_n100# 0.00fF
C1223 a_n1232_n100# a_n1652_n100# 0.02fF
C1224 a_n4078_n632# a_n4170_n632# 0.09fF
C1225 a_2012_n632# a_1592_n632# 0.02fF
C1226 a_n1650_n632# a_n1768_n632# 0.07fF
C1227 a_n2868_131# a_n2028_131# 0.01fF
C1228 a_30_n632# a_n1020_n632# 0.01fF
C1229 a_n2070_n632# a_n2398_n632# 0.02fF
C1230 a_n1020_n632# a_n2188_n632# 0.01fF
C1231 a_n1860_n632# a_n1978_n632# 0.07fF
C1232 a_n88_n632# a_n298_n632# 0.03fF
C1233 a_n3542_n100# a_n2492_n100# 0.01fF
C1234 a_4112_n632# a_3810_n632# 0.02fF
C1235 a_n602_n100# a_n1770_n100# 0.01fF
C1236 a_n1020_n632# a_n1022_n100# 0.00fF
C1237 a_240_n632# a_1592_n632# 0.00fF
C1238 a_n4080_n100# a_n2610_n100# 0.00fF
C1239 a_752_n632# a_1500_n632# 0.01fF
C1240 a_1172_n632# a_1500_n632# 0.02fF
C1241 a_1802_n632# a_3062_n632# 0.00fF
C1242 w_n4520_n851# a_1078_n100# 0.02fF
C1243 a_n3238_n632# a_n3448_n632# 0.03fF
C1244 a_658_n100# w_n4520_n851# 0.02fF
C1245 a_3388_n100# a_3808_n100# 0.02fF
C1246 a_1964_n729# a_2174_n401# 0.00fF
C1247 a_1498_n100# a_2548_n100# 0.01fF
C1248 a_n3122_n100# w_n4520_n851# 0.03fF
C1249 a_238_n100# a_1498_n100# 0.00fF
C1250 a_n1980_n100# a_n2492_n100# 0.01fF
C1251 a_n2610_n100# a_n3752_n100# 0.01fF
C1252 a_n1140_n100# a_n2400_n100# 0.00fF
C1253 a_n3238_n632# a_n2608_n632# 0.01fF
C1254 a_n1440_n632# a_n2490_n632# 0.01fF
C1255 a_n3240_n100# w_n4520_n851# 0.03fF
C1256 a_n88_n632# a_n508_n632# 0.02fF
C1257 a_4112_n632# a_2550_n632# 0.00fF
C1258 a_n510_n100# a_n90_n100# 0.02fF
C1259 a_n718_n632# a_n1650_n632# 0.01fF
C1260 a_n298_n632# a_n1230_n632# 0.01fF
C1261 a_122_n632# a_1710_n632# 0.00fF
C1262 a_3852_131# a_2592_131# 0.00fF
C1263 a_240_n632# a_n810_n632# 0.01fF
C1264 a_1962_n197# a_2172_131# 0.00fF
C1265 a_n346_n401# a_n348_131# 0.01fF
C1266 a_1288_n100# a_2010_n100# 0.01fF
C1267 a_n1022_n100# a_n90_n100# 0.01fF
C1268 a_n3916_n729# a_n3918_n197# 0.01fF
C1269 a_n2190_n100# a_n2912_n100# 0.01fF
C1270 a_2760_n632# a_3062_n632# 0.02fF
C1271 a_n1350_n100# w_n4520_n851# 0.02fF
C1272 a_750_n100# a_1078_n100# 0.02fF
C1273 a_658_n100# a_750_n100# 0.09fF
C1274 a_1962_n197# a_3012_131# 0.00fF
C1275 a_1124_n729# a_1170_n100# 0.00fF
C1276 a_n3448_n632# a_n3496_n729# 0.00fF
C1277 a_n390_n632# a_n928_n632# 0.01fF
C1278 a_4062_n197# a_2592_131# 0.00fF
C1279 a_2128_n100# a_3480_n100# 0.00fF
C1280 a_3598_n100# a_3270_n100# 0.02fF
C1281 a_30_n632# a_n1440_n632# 0.00fF
C1282 a_n2190_n100# a_n2282_n100# 0.09fF
C1283 a_n1606_n401# a_n3076_n729# 0.00fF
C1284 a_n508_n632# a_n1230_n632# 0.01fF
C1285 a_1382_n632# a_2432_n632# 0.01fF
C1286 a_n1440_n632# a_n2188_n632# 0.01fF
C1287 a_n3028_n632# a_n3076_n729# 0.00fF
C1288 a_3062_n632# a_3482_n632# 0.02fF
C1289 a_2338_n100# a_868_n100# 0.00fF
C1290 a_3600_n632# a_2012_n632# 0.00fF
C1291 a_492_131# a_702_n197# 0.00fF
C1292 a_2968_n100# a_2640_n100# 0.02fF
C1293 a_1380_n100# a_1170_n100# 0.03fF
C1294 w_n4520_n851# a_2758_n100# 0.02fF
C1295 a_120_n100# a_72_131# 0.00fF
C1296 a_n2818_n632# a_n3658_n632# 0.01fF
C1297 a_870_n632# a_1080_n632# 0.03fF
C1298 a_n3120_n632# a_n3658_n632# 0.01fF
C1299 a_n720_n100# a_n90_n100# 0.01fF
C1300 a_3692_n632# a_4020_n632# 0.02fF
C1301 a_n1978_n632# a_n2910_n632# 0.01fF
C1302 a_2970_n632# a_3390_n632# 0.02fF
C1303 a_448_n100# a_1170_n100# 0.01fF
C1304 a_3600_n632# a_3644_n729# 0.00fF
C1305 a_n3498_n197# a_n3288_131# 0.00fF
C1306 a_n300_n100# a_868_n100# 0.01fF
C1307 a_n1860_n632# a_n1650_n632# 0.03fF
C1308 a_n1978_n632# a_n2700_n632# 0.01fF
C1309 a_2340_n632# a_3810_n632# 0.00fF
C1310 a_3014_n401# a_2594_n401# 0.01fF
C1311 a_74_n401# a_72_131# 0.01fF
C1312 a_870_n632# a_332_n632# 0.01fF
C1313 a_n3660_n100# a_n3962_n100# 0.02fF
C1314 a_n2658_n197# a_n3498_n197# 0.01fF
C1315 a_2338_n100# a_3060_n100# 0.01fF
C1316 a_n600_n632# a_n1138_n632# 0.01fF
C1317 a_n2912_n100# a_n4080_n100# 0.01fF
C1318 a_3480_n100# a_3808_n100# 0.02fF
C1319 a_n3030_n100# a_n4172_n100# 0.01fF
C1320 a_n976_n729# a_n978_n197# 0.01fF
C1321 a_n2492_n100# a_n1652_n100# 0.01fF
C1322 a_n4128_131# a_n3288_131# 0.01fF
C1323 a_n3870_n100# a_n4172_n100# 0.02fF
C1324 a_n556_n729# a_74_n401# 0.00fF
C1325 a_n2866_n401# a_n1396_n729# 0.00fF
C1326 a_n2912_n100# a_n3752_n100# 0.01fF
C1327 a_660_n632# a_1080_n632# 0.02fF
C1328 w_n4520_n851# a_3900_n100# 0.06fF
C1329 a_n4128_131# a_n2658_n197# 0.00fF
C1330 a_n1560_n100# a_n2702_n100# 0.01fF
C1331 a_1542_n197# a_702_n197# 0.01fF
C1332 a_2550_n632# a_2340_n632# 0.03fF
C1333 a_n88_n632# w_n4520_n851# 0.01fF
C1334 a_n90_n100# a_1380_n100# 0.00fF
C1335 w_n4520_n851# a_n2656_n729# 0.12fF
C1336 a_n136_n729# a_n138_n197# 0.01fF
C1337 a_120_n100# a_238_n100# 0.07fF
C1338 a_2640_n100# a_3178_n100# 0.01fF
C1339 a_332_n632# a_660_n632# 0.02fF
C1340 a_n2282_n100# a_n3752_n100# 0.00fF
C1341 a_448_n100# a_n90_n100# 0.01fF
C1342 a_1802_n632# a_3272_n632# 0.00fF
C1343 a_1802_n632# a_1500_n632# 0.02fF
C1344 a_n1140_n100# a_n2072_n100# 0.01fF
C1345 a_3642_n197# a_3690_n100# 0.00fF
C1346 a_n3286_n401# a_n2236_n729# 0.00fF
C1347 a_n300_n100# a_540_n100# 0.01fF
C1348 a_912_131# a_492_131# 0.01fF
C1349 a_n4078_n632# a_n3960_n632# 0.07fF
C1350 a_2430_n100# a_3690_n100# 0.00fF
C1351 a_3598_n100# a_2010_n100# 0.00fF
C1352 a_n2820_n100# a_n3660_n100# 0.01fF
C1353 a_2970_n632# a_2432_n632# 0.01fF
C1354 a_752_n632# a_n88_n632# 0.01fF
C1355 a_3390_n632# a_1920_n632# 0.00fF
C1356 a_n88_n632# a_1172_n632# 0.00fF
C1357 a_30_n632# a_1382_n632# 0.00fF
C1358 a_n2702_n100# a_n3450_n100# 0.01fF
C1359 w_n4520_n851# a_n1230_n632# 0.01fF
C1360 a_n138_n197# a_n768_131# 0.00fF
C1361 a_4018_n100# a_3060_n100# 0.01fF
C1362 a_3222_n197# a_3178_n100# 0.00fF
C1363 a_448_n100# a_492_131# 0.00fF
C1364 w_n4520_n851# a_n1770_n100# 0.02fF
C1365 a_3902_n632# a_4112_n632# 0.03fF
C1366 a_n4170_n632# a_n3960_n632# 0.03fF
C1367 a_2760_n632# a_3272_n632# 0.01fF
C1368 a_2760_n632# a_1500_n632# 0.00fF
C1369 a_n90_n100# a_n1652_n100# 0.00fF
C1370 a_n2910_n632# a_n1650_n632# 0.00fF
C1371 a_2220_n100# a_2850_n100# 0.01fF
C1372 a_2340_n632# a_1290_n632# 0.01fF
C1373 a_n2190_n100# a_n3122_n100# 0.01fF
C1374 a_1080_n632# a_122_n632# 0.01fF
C1375 a_1288_n100# a_2338_n100# 0.01fF
C1376 a_n1442_n100# a_n1862_n100# 0.02fF
C1377 a_3434_n401# a_3482_n632# 0.00fF
C1378 a_n1560_n100# a_n930_n100# 0.01fF
C1379 a_n2700_n632# a_n1650_n632# 0.01fF
C1380 a_2852_n632# a_1710_n632# 0.01fF
C1381 a_912_131# a_1542_n197# 0.00fF
C1382 a_2384_n729# a_2594_n401# 0.00fF
C1383 a_n3240_n100# a_n2190_n100# 0.01fF
C1384 a_2640_n100# a_1380_n100# 0.00fF
C1385 a_3390_n632# a_2012_n632# 0.00fF
C1386 a_3272_n632# a_3482_n632# 0.03fF
C1387 a_1800_n100# a_868_n100# 0.01fF
C1388 a_n390_n632# a_n1768_n632# 0.00fF
C1389 a_2430_n100# a_1170_n100# 0.00fF
C1390 a_332_n632# a_122_n632# 0.03fF
C1391 a_2548_n100# a_1078_n100# 0.00fF
C1392 a_n300_n100# a_1288_n100# 0.00fF
C1393 a_238_n100# a_1078_n100# 0.01fF
C1394 a_658_n100# a_238_n100# 0.02fF
C1395 a_n1020_n632# a_n1558_n632# 0.01fF
C1396 a_n1860_n632# a_n1862_n100# 0.00fF
C1397 a_n2190_n100# a_n1350_n100# 0.01fF
C1398 a_n138_n197# a_n1188_131# 0.00fF
C1399 a_4064_n729# a_2594_n401# 0.00fF
C1400 a_n3238_n632# a_n3028_n632# 0.03fF
C1401 a_n810_n632# a_n812_n100# 0.00fF
C1402 a_n2398_n632# a_n1230_n632# 0.01fF
C1403 a_n2026_n401# a_n2866_n401# 0.01fF
C1404 a_n3122_n100# a_n3078_n197# 0.00fF
C1405 a_2128_n100# a_868_n100# 0.00fF
C1406 a_3480_n100# a_3388_n100# 0.09fF
C1407 a_2970_n632# a_2968_n100# 0.00fF
C1408 a_n558_n197# a_n768_131# 0.00fF
C1409 a_3014_n401# a_1964_n729# 0.00fF
C1410 a_3060_n100# a_1800_n100# 0.00fF
C1411 a_n1020_n632# a_n2280_n632# 0.00fF
C1412 w_n4520_n851# a_3692_n632# 0.04fF
C1413 a_2432_n632# a_1920_n632# 0.01fF
C1414 a_704_n729# a_1334_n401# 0.00fF
C1415 a_n1818_n197# a_n1608_131# 0.00fF
C1416 a_962_n632# a_2130_n632# 0.01fF
C1417 a_240_n632# a_n1138_n632# 0.00fF
C1418 a_n1348_n632# a_n928_n632# 0.02fF
C1419 a_n2700_n632# a_n2658_n197# 0.00fF
C1420 a_3432_131# a_2592_131# 0.01fF
C1421 a_n4080_n100# a_n3122_n100# 0.01fF
C1422 a_284_n729# w_n4520_n851# 0.12fF
C1423 a_1918_n100# a_2850_n100# 0.01fF
C1424 a_238_n100# a_n1350_n100# 0.00fF
C1425 a_450_n632# a_1592_n632# 0.01fF
C1426 a_n1022_n100# a_n2400_n100# 0.00fF
C1427 a_n390_n632# a_n718_n632# 0.02fF
C1428 a_n3240_n100# a_n4080_n100# 0.01fF
C1429 a_960_n100# a_868_n100# 0.09fF
C1430 a_2804_n729# a_1334_n401# 0.00fF
C1431 a_30_n632# a_n600_n632# 0.01fF
C1432 a_1800_n100# a_540_n100# 0.00fF
C1433 a_n3122_n100# a_n3752_n100# 0.01fF
C1434 a_2128_n100# a_3060_n100# 0.01fF
C1435 a_n392_n100# a_n1140_n100# 0.01fF
C1436 a_n2188_n632# a_n600_n632# 0.00fF
C1437 a_1382_n632# a_1380_n100# 0.00fF
C1438 a_3902_n632# a_2340_n632# 0.00fF
C1439 a_542_n632# a_1500_n632# 0.01fF
C1440 a_n3240_n100# a_n3752_n100# 0.01fF
C1441 a_n3708_131# a_n3750_n632# 0.00fF
C1442 a_n2820_n100# a_n2818_n632# 0.00fF
C1443 a_n346_n401# a_74_n401# 0.01fF
C1444 w_n4520_n851# a_2592_131# 0.12fF
C1445 a_2758_n100# a_2548_n100# 0.03fF
C1446 a_n2400_n100# a_n3542_n100# 0.01fF
C1447 a_2432_n632# a_2012_n632# 0.02fF
C1448 a_2760_n632# a_2758_n100# 0.00fF
C1449 a_2222_n632# a_2130_n632# 0.09fF
C1450 a_n558_n197# a_n1188_131# 0.00fF
C1451 a_450_n632# a_n810_n632# 0.00fF
C1452 a_2128_n100# a_540_n100# 0.00fF
C1453 a_2010_n100# a_1962_n197# 0.00fF
C1454 a_n300_n100# a_n182_n100# 0.07fF
C1455 a_n138_n197# a_n978_n197# 0.01fF
C1456 w_n4520_n851# a_n3706_n401# 0.10fF
C1457 a_2642_n632# a_2130_n632# 0.01fF
C1458 a_n1440_n632# a_n1558_n632# 0.07fF
C1459 a_2220_n100# a_1590_n100# 0.01fF
C1460 a_n2400_n100# a_n1980_n100# 0.02fF
C1461 a_n2912_n100# a_n2610_n100# 0.02fF
C1462 a_1708_n100# a_3270_n100# 0.00fF
C1463 a_2338_n100# a_3598_n100# 0.00fF
C1464 a_n1348_n632# a_n2818_n632# 0.00fF
C1465 a_3060_n100# a_3808_n100# 0.01fF
C1466 a_n1440_n632# a_n2280_n632# 0.01fF
C1467 a_960_n100# a_540_n100# 0.02fF
C1468 a_n1860_n632# a_n390_n632# 0.00fF
C1469 a_n1818_n197# w_n4520_n851# 0.10fF
C1470 a_n2610_n100# a_n2282_n100# 0.02fF
C1471 a_n2446_n401# a_n3286_n401# 0.01fF
C1472 a_3900_n100# a_2548_n100# 0.00fF
C1473 a_1288_n100# a_1800_n100# 0.01fF
C1474 a_n88_n632# a_n180_n632# 0.09fF
C1475 a_n3870_n100# a_n3918_n197# 0.00fF
C1476 a_n300_n100# a_n1442_n100# 0.01fF
C1477 a_2640_n100# a_2430_n100# 0.03fF
C1478 a_1334_n401# a_1290_n632# 0.00fF
C1479 a_2384_n729# a_1964_n729# 0.01fF
C1480 a_2802_n197# a_1542_n197# 0.00fF
C1481 a_n2190_n100# a_n1770_n100# 0.02fF
C1482 a_1288_n100# a_2128_n100# 0.01fF
C1483 a_1918_n100# a_1590_n100# 0.02fF
C1484 a_n558_n197# a_n978_n197# 0.01fF
C1485 a_3854_n401# a_2594_n401# 0.00fF
C1486 a_n180_n632# a_n1230_n632# 0.01fF
C1487 a_n3238_n632# a_n2490_n632# 0.01fF
C1488 a_n3658_n632# a_n2910_n632# 0.01fF
C1489 a_3222_n197# a_3642_n197# 0.01fF
C1490 a_n510_n100# a_n2072_n100# 0.00fF
C1491 a_n810_n632# a_n298_n632# 0.01fF
C1492 a_n1140_n100# a_n812_n100# 0.02fF
C1493 a_1800_n100# a_1752_131# 0.00fF
C1494 a_4018_n100# a_3598_n100# 0.02fF
C1495 a_n1816_n729# a_n3286_n401# 0.00fF
C1496 a_n1020_n632# a_332_n632# 0.00fF
C1497 a_n3332_n100# a_n4172_n100# 0.01fF
C1498 a_n3660_n100# a_n3450_n100# 0.03fF
C1499 a_n2868_131# a_n3498_n197# 0.00fF
C1500 a_n2700_n632# a_n3658_n632# 0.01fF
C1501 a_1288_n100# a_960_n100# 0.02fF
C1502 a_n3660_n100# a_n2702_n100# 0.01fF
C1503 a_n1022_n100# a_n2072_n100# 0.01fF
C1504 a_1382_n632# a_1710_n632# 0.02fF
C1505 a_3222_n197# a_2802_n197# 0.01fF
C1506 a_914_n401# w_n4520_n851# 0.10fF
C1507 a_n2818_n632# a_n4078_n632# 0.00fF
C1508 a_n3120_n632# a_n4078_n632# 0.01fF
C1509 a_n1348_n632# a_n1768_n632# 0.02fF
C1510 a_120_n100# a_1498_n100# 0.00fF
C1511 a_n2400_n100# a_n1652_n100# 0.01fF
C1512 a_n4128_131# a_n2868_131# 0.00fF
C1513 a_n810_n632# a_n508_n632# 0.02fF
C1514 a_30_n632# a_240_n632# 0.03fF
C1515 a_3600_n632# a_4020_n632# 0.02fF
C1516 a_2010_n100# a_1708_n100# 0.02fF
C1517 a_n2072_n100# a_n3542_n100# 0.00fF
C1518 a_n1440_n632# a_n1396_n729# 0.00fF
C1519 a_n3238_n632# a_n3330_n632# 0.09fF
C1520 a_n3238_n632# a_n2188_n632# 0.01fF
C1521 a_2968_n100# a_2220_n100# 0.01fF
C1522 a_494_n401# a_450_n632# 0.00fF
C1523 a_n2818_n632# a_n4170_n632# 0.00fF
C1524 a_1288_n100# a_1290_n632# 0.00fF
C1525 a_n3120_n632# a_n4170_n632# 0.01fF
C1526 a_n720_n100# a_n2072_n100# 0.00fF
C1527 a_n2912_n100# a_n2282_n100# 0.01fF
C1528 a_n556_n729# a_284_n729# 0.01fF
C1529 a_n3030_n100# a_n2492_n100# 0.01fF
C1530 a_n2072_n100# a_n1980_n100# 0.09fF
C1531 a_542_n632# a_n88_n632# 0.01fF
C1532 a_282_n197# a_1752_131# 0.00fF
C1533 a_n3870_n100# a_n2492_n100# 0.00fF
C1534 a_n3916_n729# a_n3076_n729# 0.01fF
C1535 a_1500_n632# a_1498_n100# 0.00fF
C1536 a_3388_n100# a_3060_n100# 0.02fF
C1537 a_4062_n197# a_4110_n100# 0.00fF
C1538 a_n1348_n632# a_n718_n632# 0.01fF
C1539 a_282_n197# a_1122_n197# 0.01fF
C1540 a_n3122_n100# a_n2610_n100# 0.01fF
C1541 a_2760_n632# a_3692_n632# 0.01fF
C1542 a_n3540_n632# a_n3238_n632# 0.02fF
C1543 a_n2820_n100# a_n1442_n100# 0.00fF
C1544 a_n1396_n729# a_n1398_n197# 0.01fF
C1545 a_n300_n100# a_330_n100# 0.01fF
C1546 a_n3286_n401# a_n4126_n401# 0.01fF
C1547 a_2382_n197# a_2340_n632# 0.00fF
C1548 a_n3240_n100# a_n2610_n100# 0.01fF
C1549 a_960_n100# a_n182_n100# 0.01fF
C1550 a_3062_n632# a_1500_n632# 0.00fF
C1551 a_3062_n632# a_3272_n632# 0.03fF
C1552 w_n4520_n851# a_1592_n632# 0.01fF
C1553 a_n3448_n632# w_n4520_n851# 0.03fF
C1554 a_2128_n100# a_3598_n100# 0.00fF
C1555 a_n1140_n100# a_n602_n100# 0.01fF
C1556 a_870_n632# a_962_n632# 0.09fF
C1557 a_2220_n100# a_3178_n100# 0.01fF
C1558 a_n138_n197# a_282_n197# 0.01fF
C1559 a_3692_n632# a_3482_n632# 0.03fF
C1560 a_2968_n100# a_1918_n100# 0.01fF
C1561 a_n1020_n632# a_n1978_n632# 0.01fF
C1562 a_n1350_n100# a_n2610_n100# 0.00fF
C1563 a_2970_n632# a_1710_n632# 0.00fF
C1564 a_1498_n100# a_1078_n100# 0.02fF
C1565 a_2128_n100# a_2130_n632# 0.00fF
C1566 a_n2608_n632# w_n4520_n851# 0.01fF
C1567 a_658_n100# a_1498_n100# 0.01fF
C1568 a_2548_n100# a_2592_131# 0.00fF
C1569 a_2550_n632# a_2130_n632# 0.02fF
C1570 a_n3918_n197# a_n3288_131# 0.00fF
C1571 a_1544_n729# a_704_n729# 0.01fF
C1572 a_n510_n100# a_n392_n100# 0.07fF
C1573 a_n3540_n632# a_n3496_n729# 0.00fF
C1574 a_450_n632# a_n1138_n632# 0.00fF
C1575 a_n2658_n197# a_n3918_n197# 0.00fF
C1576 a_n600_n632# a_n1558_n632# 0.01fF
C1577 a_n1022_n100# a_n392_n100# 0.01fF
C1578 a_752_n632# a_1592_n632# 0.01fF
C1579 a_1172_n632# a_1592_n632# 0.02fF
C1580 a_n810_n632# w_n4520_n851# 0.01fF
C1581 a_n928_n632# a_n930_n100# 0.00fF
C1582 a_2804_n729# a_1544_n729# 0.00fF
C1583 a_n1348_n632# a_n1860_n632# 0.01fF
C1584 a_660_n632# a_962_n632# 0.02fF
C1585 a_3644_n729# a_2174_n401# 0.00fF
C1586 a_n2910_n632# a_n2868_131# 0.00fF
C1587 a_3690_n100# a_3270_n100# 0.02fF
C1588 a_870_n632# a_2222_n632# 0.00fF
C1589 a_3598_n100# a_3808_n100# 0.03fF
C1590 a_n976_n729# a_n930_n100# 0.00fF
C1591 a_n2072_n100# a_n1652_n100# 0.02fF
C1592 a_870_n632# a_n390_n632# 0.00fF
C1593 a_120_n100# a_74_n401# 0.00fF
C1594 a_n3448_n632# a_n2398_n632# 0.01fF
C1595 a_1918_n100# a_3178_n100# 0.00fF
C1596 a_3390_n632# a_4020_n632# 0.01fF
C1597 a_3480_n100# a_3060_n100# 0.02fF
C1598 a_n1818_n197# a_n3078_n197# 0.00fF
C1599 a_752_n632# a_n810_n632# 0.00fF
C1600 a_1382_n632# a_1080_n632# 0.02fF
C1601 a_n1818_n197# a_n2448_131# 0.00fF
C1602 a_n558_n197# a_282_n197# 0.01fF
C1603 a_2222_n632# a_3180_n632# 0.01fF
C1604 a_n2398_n632# a_n2608_n632# 0.03fF
C1605 a_n720_n100# a_n392_n100# 0.02fF
C1606 a_n1232_n100# a_n1862_n100# 0.01fF
C1607 a_2220_n100# a_1380_n100# 0.01fF
C1608 a_1290_n632# a_2130_n632# 0.01fF
C1609 a_n2912_n100# a_n3122_n100# 0.03fF
C1610 a_2642_n632# a_3180_n632# 0.01fF
C1611 a_2172_131# a_1542_n197# 0.00fF
C1612 a_n4172_n100# a_n3962_n100# 0.03fF
C1613 a_1498_n100# a_2758_n100# 0.00fF
C1614 a_n392_n100# a_n1980_n100# 0.00fF
C1615 a_n1140_n100# a_28_n100# 0.01fF
C1616 a_2222_n632# a_660_n632# 0.00fF
C1617 a_2220_n100# a_2174_n401# 0.00fF
C1618 a_2338_n100# a_1708_n100# 0.01fF
C1619 a_n1978_n632# a_n1440_n632# 0.01fF
C1620 a_1382_n632# a_332_n632# 0.01fF
C1621 a_n3240_n100# a_n2912_n100# 0.02fF
C1622 a_1920_n632# a_1710_n632# 0.03fF
C1623 a_n930_n100# a_540_n100# 0.00fF
C1624 a_1542_n197# a_3012_131# 0.00fF
C1625 a_3600_n632# w_n4520_n851# 0.04fF
C1626 a_n556_n729# a_914_n401# 0.00fF
C1627 w_n4520_n851# a_n1186_n401# 0.10fF
C1628 a_n390_n632# a_660_n632# 0.01fF
C1629 a_n2656_n729# a_n2610_n100# 0.00fF
C1630 a_1800_n100# a_330_n100# 0.00fF
C1631 a_n2398_n632# a_n810_n632# 0.00fF
C1632 a_n3122_n100# a_n2282_n100# 0.01fF
C1633 a_n298_n632# a_n1138_n632# 0.01fF
C1634 a_2642_n632# a_2594_n401# 0.00fF
C1635 a_n3240_n100# a_n2282_n100# 0.01fF
C1636 a_n2912_n100# a_n1350_n100# 0.00fF
C1637 a_n1020_n632# a_n1650_n632# 0.01fF
C1638 a_3222_n197# a_2172_131# 0.00fF
C1639 a_n1560_n100# a_n182_n100# 0.00fF
C1640 a_n346_n401# a_284_n729# 0.00fF
C1641 a_284_n729# a_1754_n401# 0.00fF
C1642 a_962_n632# a_122_n632# 0.01fF
C1643 a_n2818_n632# a_n3960_n632# 0.01fF
C1644 a_2010_n100# a_1964_n729# 0.00fF
C1645 a_3222_n197# a_3012_131# 0.00fF
C1646 a_n3120_n632# a_n3960_n632# 0.01fF
C1647 a_120_n100# a_1078_n100# 0.01fF
C1648 a_120_n100# a_658_n100# 0.01fF
C1649 a_n4128_131# a_n4170_n632# 0.00fF
C1650 a_n510_n100# a_n812_n100# 0.02fF
C1651 a_n1348_n632# a_n2910_n632# 0.00fF
C1652 a_2970_n632# a_3014_n401# 0.00fF
C1653 a_n1350_n100# a_n2282_n100# 0.01fF
C1654 a_2012_n632# a_1710_n632# 0.02fF
C1655 a_448_n100# a_n392_n100# 0.01fF
C1656 a_n1606_n401# a_n1608_131# 0.01fF
C1657 a_n508_n632# a_n1138_n632# 0.01fF
C1658 a_1918_n100# a_1380_n100# 0.01fF
C1659 a_n1022_n100# a_n812_n100# 0.03fF
C1660 a_n1232_n100# a_n1188_131# 0.00fF
C1661 a_n1348_n632# a_n2700_n632# 0.00fF
C1662 a_n2820_n100# a_n4172_n100# 0.00fF
C1663 a_n1770_n100# a_n2610_n100# 0.01fF
C1664 a_2432_n632# a_4020_n632# 0.00fF
C1665 a_2850_n100# w_n4520_n851# 0.03fF
C1666 a_1918_n100# a_448_n100# 0.00fF
C1667 a_960_n100# a_330_n100# 0.01fF
C1668 a_240_n632# a_1710_n632# 0.00fF
C1669 a_330_n100# a_282_n197# 0.00fF
C1670 a_3644_n729# a_3642_n197# 0.01fF
C1671 a_n1560_n100# a_n1442_n100# 0.07fF
C1672 a_1590_n100# a_28_n100# 0.00fF
C1673 a_494_n401# w_n4520_n851# 0.10fF
C1674 a_120_n100# a_n1350_n100# 0.00fF
C1675 a_n2280_n632# a_n2238_n197# 0.00fF
C1676 a_n390_n632# a_122_n632# 0.01fF
C1677 a_1802_n632# a_1592_n632# 0.03fF
C1678 a_n3916_n729# a_n3496_n729# 0.01fF
C1679 a_n392_n100# a_n1652_n100# 0.00fF
C1680 a_n720_n100# a_n812_n100# 0.09fF
C1681 a_n1140_n100# w_n4520_n851# 0.02fF
C1682 a_3598_n100# a_3388_n100# 0.03fF
C1683 a_n3450_n100# a_n3498_n197# 0.00fF
C1684 a_450_n632# a_30_n632# 0.02fF
C1685 a_n3238_n632# a_n3750_n632# 0.01fF
C1686 a_n1980_n100# a_n812_n100# 0.01fF
C1687 a_332_n632# a_n600_n632# 0.01fF
C1688 a_n2866_n401# a_n3286_n401# 0.01fF
C1689 a_n4078_n632# a_n4126_n401# 0.00fF
C1690 a_n1440_n632# a_n1650_n632# 0.03fF
C1691 a_3390_n632# a_3432_131# 0.00fF
C1692 a_n3238_n632# a_n2280_n632# 0.01fF
C1693 a_n3708_131# a_n3288_131# 0.01fF
C1694 a_2010_n100# a_1170_n100# 0.01fF
C1695 a_3224_n729# a_3180_n632# 0.00fF
C1696 a_4110_n100# w_n4520_n851# 0.14fF
C1697 a_n1442_n100# a_n2702_n100# 0.00fF
C1698 a_n3708_131# a_n2658_n197# 0.00fF
C1699 a_n1862_n100# a_n2492_n100# 0.01fF
C1700 a_2220_n100# a_2430_n100# 0.03fF
C1701 a_2760_n632# a_1592_n632# 0.01fF
C1702 a_658_n100# a_1078_n100# 0.02fF
C1703 w_n4520_n851# a_n1606_n401# 0.10fF
C1704 a_n2910_n632# a_n4078_n632# 0.01fF
C1705 a_n4170_n632# a_n4126_n401# 0.00fF
C1706 w_n4520_n851# a_n3028_n632# 0.03fF
C1707 a_n300_n100# a_n1232_n100# 0.01fF
C1708 a_n1818_n197# a_n348_131# 0.00fF
C1709 a_n2866_n401# a_n2868_131# 0.01fF
C1710 a_1708_n100# a_1800_n100# 0.09fF
C1711 a_n2700_n632# a_n4078_n632# 0.00fF
C1712 a_2640_n100# a_3270_n100# 0.01fF
C1713 a_3390_n632# w_n4520_n851# 0.03fF
C1714 a_3224_n729# a_2594_n401# 0.00fF
C1715 a_n510_n100# a_n602_n100# 0.09fF
C1716 a_n3332_n100# a_n2492_n100# 0.01fF
C1717 a_n930_n100# a_n182_n100# 0.01fF
C1718 a_n180_n632# a_n810_n632# 0.01fF
C1719 a_n3240_n100# a_n3122_n100# 0.07fF
C1720 a_3810_n632# a_3180_n632# 0.01fF
C1721 a_448_n100# a_n812_n100# 0.00fF
C1722 a_n1022_n100# a_n602_n100# 0.02fF
C1723 a_n2910_n632# a_n4170_n632# 0.00fF
C1724 w_n4520_n851# a_n1138_n632# 0.01fF
C1725 a_n2026_n401# a_n3076_n729# 0.00fF
C1726 a_2970_n632# a_3012_131# 0.00fF
C1727 a_n2912_n100# a_n1770_n100# 0.01fF
C1728 a_n2400_n100# a_n3030_n100# 0.01fF
C1729 a_1920_n632# a_1080_n632# 0.01fF
C1730 a_n976_n729# a_n928_n632# 0.00fF
C1731 a_660_n632# a_704_n729# 0.00fF
C1732 a_2128_n100# a_1708_n100# 0.02fF
C1733 a_n2700_n632# a_n4170_n632# 0.00fF
C1734 a_n136_n729# a_n90_n100# 0.00fF
C1735 a_914_n401# a_1754_n401# 0.01fF
C1736 a_n3030_n100# a_n3076_n729# 0.00fF
C1737 a_n346_n401# a_914_n401# 0.00fF
C1738 a_n3870_n100# a_n2400_n100# 0.00fF
C1739 a_1590_n100# w_n4520_n851# 0.02fF
C1740 a_n1770_n100# a_n2282_n100# 0.01fF
C1741 a_332_n632# a_1920_n632# 0.00fF
C1742 a_n3448_n632# a_n3868_n632# 0.02fF
C1743 a_3222_n197# a_3270_n100# 0.00fF
C1744 a_30_n632# a_n298_n632# 0.02fF
C1745 a_2550_n632# a_3180_n632# 0.01fF
C1746 a_n556_n729# a_n1186_n401# 0.00fF
C1747 a_3062_n632# a_3692_n632# 0.01fF
C1748 a_3014_n401# a_3644_n729# 0.00fF
C1749 a_1918_n100# a_2430_n100# 0.01fF
C1750 a_2382_n197# a_1752_131# 0.00fF
C1751 a_n976_n729# a_n2236_n729# 0.00fF
C1752 a_3598_n100# a_3480_n100# 0.07fF
C1753 a_540_n100# a_868_n100# 0.02fF
C1754 a_1332_131# a_2592_131# 0.00fF
C1755 a_n2608_n632# a_n3868_n632# 0.00fF
C1756 a_n930_n100# a_n1442_n100# 0.01fF
C1757 a_n720_n100# a_n602_n100# 0.07fF
C1758 a_960_n100# a_1708_n100# 0.01fF
C1759 a_n2398_n632# a_n3028_n632# 0.01fF
C1760 a_n2820_n100# a_n2866_n401# 0.00fF
C1761 a_n2658_n197# a_n1398_n197# 0.00fF
C1762 a_n812_n100# a_n1652_n100# 0.01fF
C1763 a_2804_n729# a_2594_n401# 0.00fF
C1764 a_n3498_n197# a_n2028_131# 0.00fF
C1765 a_n4172_n100# a_n4170_n632# 0.00fF
C1766 a_2382_n197# a_1122_n197# 0.00fF
C1767 a_n602_n100# a_n1980_n100# 0.00fF
C1768 a_2012_n632# a_1080_n632# 0.01fF
C1769 a_n1978_n632# a_n600_n632# 0.00fF
C1770 a_n2070_n632# a_n1230_n632# 0.01fF
C1771 a_2338_n100# a_3690_n100# 0.00fF
C1772 a_n88_n632# a_1500_n632# 0.00fF
C1773 a_2550_n632# a_2594_n401# 0.00fF
C1774 a_30_n632# a_n508_n632# 0.01fF
C1775 a_750_n100# a_1590_n100# 0.01fF
C1776 a_n510_n100# a_n508_n632# 0.00fF
C1777 a_n2398_n632# a_n1138_n632# 0.00fF
C1778 a_n3962_n100# a_n3918_n197# 0.00fF
C1779 a_450_n632# a_448_n100# 0.00fF
C1780 a_542_n632# a_1592_n632# 0.01fF
C1781 a_2432_n632# w_n4520_n851# 0.01fF
C1782 a_30_n632# a_28_n100# 0.00fF
C1783 a_2760_n632# a_3600_n632# 0.01fF
C1784 a_n2868_131# a_n3918_n197# 0.00fF
C1785 a_n510_n100# a_28_n100# 0.01fF
C1786 a_240_n632# a_1080_n632# 0.01fF
C1787 a_870_n632# a_1290_n632# 0.02fF
C1788 a_n1022_n100# a_28_n100# 0.01fF
C1789 a_2852_n632# a_2222_n632# 0.01fF
C1790 a_n768_131# a_492_131# 0.00fF
C1791 a_240_n632# a_332_n632# 0.09fF
C1792 a_2852_n632# a_2642_n632# 0.03fF
C1793 a_n558_n197# a_n2028_131# 0.00fF
C1794 a_3600_n632# a_3482_n632# 0.07fF
C1795 a_2640_n100# a_2010_n100# 0.01fF
C1796 a_n2700_n632# a_n2702_n100# 0.00fF
C1797 a_n2820_n100# a_n1232_n100# 0.00fF
C1798 a_n1020_n632# a_n390_n632# 0.01fF
C1799 a_448_n100# a_n602_n100# 0.01fF
C1800 a_1172_n632# a_2432_n632# 0.00fF
C1801 a_1288_n100# a_868_n100# 0.02fF
C1802 a_542_n632# a_n810_n632# 0.00fF
C1803 a_n556_n729# a_494_n401# 0.00fF
C1804 a_2338_n100# a_1170_n100# 0.01fF
C1805 a_660_n632# a_1290_n632# 0.01fF
C1806 a_2850_n100# a_2548_n100# 0.02fF
C1807 a_n2190_n100# a_n1140_n100# 0.01fF
C1808 a_2340_n632# a_2130_n632# 0.03fF
C1809 a_n1348_n632# a_122_n632# 0.00fF
C1810 a_n720_n100# a_28_n100# 0.01fF
C1811 a_n2490_n632# w_n4520_n851# 0.01fF
C1812 a_n4172_n100# a_n3450_n100# 0.01fF
C1813 a_4018_n100# a_3690_n100# 0.02fF
C1814 a_n4172_n100# a_n2702_n100# 0.00fF
C1815 a_n3120_n632# a_n2818_n632# 0.02fF
C1816 a_3224_n729# a_1964_n729# 0.00fF
C1817 a_n2072_n100# a_n3030_n100# 0.01fF
C1818 a_n768_131# a_n1398_n197# 0.00fF
C1819 a_n300_n100# a_1170_n100# 0.00fF
C1820 a_2384_n729# a_3644_n729# 0.00fF
C1821 a_n1020_n632# a_n978_n197# 0.00fF
C1822 a_2968_n100# w_n4520_n851# 0.03fF
C1823 a_n602_n100# a_n1652_n100# 0.01fF
C1824 a_n928_n632# a_n1768_n632# 0.01fF
C1825 a_284_n729# a_74_n401# 0.00fF
C1826 a_3852_131# a_3642_n197# 0.00fF
C1827 a_n3122_n100# a_n1770_n100# 0.00fF
C1828 a_238_n100# a_n1140_n100# 0.00fF
C1829 a_n1650_n632# a_n600_n632# 0.01fF
C1830 a_n556_n729# a_n1606_n401# 0.00fF
C1831 a_n930_n100# a_330_n100# 0.00fF
C1832 a_3900_n100# a_2758_n100# 0.01fF
C1833 a_4064_n729# a_3644_n729# 0.01fF
C1834 a_1288_n100# a_540_n100# 0.01fF
C1835 a_n3240_n100# a_n1770_n100# 0.00fF
C1836 a_1802_n632# a_3390_n632# 0.00fF
C1837 a_4062_n197# a_3642_n197# 0.01fF
C1838 a_30_n632# w_n4520_n851# 0.01fF
C1839 a_1964_n729# a_704_n729# 0.00fF
C1840 a_3852_131# a_2802_n197# 0.00fF
C1841 a_n3962_n100# a_n2492_n100# 0.00fF
C1842 a_n3330_n632# w_n4520_n851# 0.03fF
C1843 w_n4520_n851# a_n2188_n632# 0.01fF
C1844 a_n510_n100# w_n4520_n851# 0.02fF
C1845 a_3692_n632# a_3272_n632# 0.02fF
C1846 a_450_n632# a_1710_n632# 0.00fF
C1847 a_4110_n100# a_2548_n100# 0.00fF
C1848 a_1380_n100# a_28_n100# 0.00fF
C1849 a_n2910_n632# a_n3960_n632# 0.01fF
C1850 a_n390_n632# a_n1440_n632# 0.01fF
C1851 a_2220_n100# a_2172_131# 0.00fF
C1852 w_n4520_n851# a_702_n197# 0.10fF
C1853 a_n1022_n100# w_n4520_n851# 0.02fF
C1854 a_n182_n100# a_868_n100# 0.01fF
C1855 a_4062_n197# a_2802_n197# 0.00fF
C1856 a_448_n100# a_28_n100# 0.02fF
C1857 a_3902_n632# a_3180_n632# 0.01fF
C1858 a_n1350_n100# a_n1770_n100# 0.02fF
C1859 a_n1188_131# a_n1398_n197# 0.00fF
C1860 a_1290_n632# a_122_n632# 0.01fF
C1861 a_n2398_n632# a_n2490_n632# 0.09fF
C1862 a_2804_n729# a_1964_n729# 0.01fF
C1863 a_n300_n100# a_n90_n100# 0.03fF
C1864 a_n2700_n632# a_n3960_n632# 0.00fF
C1865 a_n346_n401# a_n1186_n401# 0.01fF
C1866 w_n4520_n851# a_3178_n100# 0.03fF
C1867 a_n3238_n632# a_n1978_n632# 0.00fF
C1868 a_30_n632# a_752_n632# 0.01fF
C1869 a_n718_n632# a_n928_n632# 0.03fF
C1870 a_30_n632# a_1172_n632# 0.01fF
C1871 a_2760_n632# a_3390_n632# 0.01fF
C1872 a_n180_n632# a_n1138_n632# 0.01fF
C1873 a_n3540_n632# w_n4520_n851# 0.03fF
C1874 a_n3496_n729# a_n2026_n401# 0.00fF
C1875 a_n3542_n100# w_n4520_n851# 0.04fF
C1876 a_n510_n100# a_750_n100# 0.00fF
C1877 a_n2608_n632# a_n2610_n100# 0.00fF
C1878 a_n978_n197# a_492_131# 0.00fF
C1879 a_n976_n729# a_n2446_n401# 0.00fF
C1880 a_n2818_n632# a_n1768_n632# 0.01fF
C1881 a_2640_n100# a_2642_n632# 0.00fF
C1882 a_n3120_n632# a_n1768_n632# 0.00fF
C1883 a_750_n100# a_702_n197# 0.00fF
C1884 a_n720_n100# w_n4520_n851# 0.02fF
C1885 a_2128_n100# a_3690_n100# 0.00fF
C1886 a_n2446_n401# a_n2236_n729# 0.00fF
C1887 a_1590_n100# a_2548_n100# 0.01fF
C1888 a_3390_n632# a_3482_n632# 0.09fF
C1889 a_1382_n632# a_962_n632# 0.02fF
C1890 a_n2820_n100# a_n2492_n100# 0.02fF
C1891 w_n4520_n851# a_n1980_n100# 0.02fF
C1892 a_n2398_n632# a_n3330_n632# 0.01fF
C1893 a_238_n100# a_1590_n100# 0.00fF
C1894 a_n2398_n632# a_n2188_n632# 0.03fF
C1895 a_494_n401# a_542_n632# 0.00fF
C1896 a_2382_n197# a_1962_n197# 0.01fF
C1897 a_2640_n100# a_2338_n100# 0.02fF
C1898 a_2432_n632# a_1802_n632# 0.01fF
C1899 a_540_n100# a_n182_n100# 0.01fF
C1900 a_1124_n729# w_n4520_n851# 0.12fF
C1901 a_n1652_n100# a_n1608_131# 0.00fF
C1902 a_n3028_n632# a_n3868_n632# 0.01fF
C1903 a_1800_n100# a_1170_n100# 0.01fF
C1904 a_n3708_131# a_n2868_131# 0.01fF
C1905 a_3598_n100# a_3060_n100# 0.01fF
C1906 a_2852_n632# a_3810_n632# 0.01fF
C1907 a_912_131# w_n4520_n851# 0.12fF
C1908 a_n2400_n100# a_n1862_n100# 0.01fF
C1909 a_n978_n197# a_n1398_n197# 0.01fF
C1910 a_n88_n632# a_n1230_n632# 0.01fF
C1911 a_n1860_n632# a_n928_n632# 0.01fF
C1912 a_n720_n100# a_750_n100# 0.00fF
C1913 a_3062_n632# a_1592_n632# 0.00fF
C1914 a_494_n401# a_n346_n401# 0.01fF
C1915 a_494_n401# a_1754_n401# 0.00fF
C1916 a_2804_n729# a_2852_n632# 0.00fF
C1917 a_n298_n632# a_n1558_n632# 0.00fF
C1918 a_n3540_n632# a_n2398_n632# 0.01fF
C1919 a_n976_n729# a_n1816_n729# 0.01fF
C1920 a_1380_n100# w_n4520_n851# 0.02fF
C1921 a_3690_n100# a_3808_n100# 0.07fF
C1922 a_1382_n632# a_2222_n632# 0.01fF
C1923 a_2128_n100# a_1170_n100# 0.01fF
C1924 a_n1560_n100# a_n1232_n100# 0.02fF
C1925 a_1172_n632# a_1124_n729# 0.00fF
C1926 a_4112_n632# a_3180_n632# 0.01fF
C1927 a_2760_n632# a_2432_n632# 0.02fF
C1928 w_n4520_n851# a_2174_n401# 0.10fF
C1929 a_n1816_n729# a_n2236_n729# 0.01fF
C1930 a_1382_n632# a_2642_n632# 0.00fF
C1931 a_2852_n632# a_2550_n632# 0.02fF
C1932 a_448_n100# w_n4520_n851# 0.02fF
C1933 a_n3332_n100# a_n2400_n100# 0.01fF
C1934 a_914_n401# a_74_n401# 0.01fF
C1935 a_n1348_n632# a_n1020_n632# 0.02fF
C1936 a_n508_n632# a_n1558_n632# 0.01fF
C1937 a_n3238_n632# a_n1650_n632# 0.00fF
C1938 a_960_n100# a_1170_n100# 0.03fF
C1939 a_2432_n632# a_3482_n632# 0.01fF
C1940 a_3854_n401# a_3644_n729# 0.00fF
C1941 a_1288_n100# a_n182_n100# 0.00fF
C1942 a_750_n100# a_1380_n100# 0.01fF
C1943 a_4018_n100# a_2640_n100# 0.00fF
C1944 a_1544_n729# a_1334_n401# 0.00fF
C1945 a_n2238_n197# a_n3288_131# 0.00fF
C1946 a_n346_n401# a_n1606_n401# 0.00fF
C1947 a_n1232_n100# a_n2702_n100# 0.00fF
C1948 w_n4520_n851# a_n1652_n100# 0.02fF
C1949 a_30_n632# a_72_131# 0.00fF
C1950 a_n2238_n197# a_n2658_n197# 0.01fF
C1951 a_448_n100# a_750_n100# 0.02fF
C1952 a_n2868_131# a_n1398_n197# 0.00fF
C1953 a_962_n632# a_n600_n632# 0.00fF
C1954 a_450_n632# a_1080_n632# 0.01fF
C1955 a_n1860_n632# a_n2818_n632# 0.01fF
C1956 a_n1860_n632# a_n3120_n632# 0.00fF
C1957 a_2220_n100# a_3270_n100# 0.01fF
C1958 a_1752_131# a_1122_n197# 0.00fF
C1959 a_72_131# a_702_n197# 0.00fF
C1960 a_330_n100# a_868_n100# 0.01fF
C1961 a_n2490_n632# a_n2448_131# 0.00fF
C1962 a_2968_n100# a_2548_n100# 0.02fF
C1963 a_n3660_n100# a_n4172_n100# 0.01fF
C1964 a_n2190_n100# a_n2188_n632# 0.00fF
C1965 a_450_n632# a_332_n632# 0.07fF
C1966 a_n556_n729# a_n510_n100# 0.00fF
C1967 a_2852_n632# a_1290_n632# 0.00fF
C1968 a_870_n632# a_2340_n632# 0.00fF
C1969 a_n718_n632# a_n1768_n632# 0.01fF
C1970 a_n2070_n632# a_n3448_n632# 0.00fF
C1971 a_n2190_n100# a_n1022_n100# 0.01fF
C1972 a_3600_n632# a_3062_n632# 0.01fF
C1973 a_960_n100# a_n90_n100# 0.01fF
C1974 a_n3916_n729# w_n4520_n851# 0.13fF
C1975 a_3642_n197# a_3432_131# 0.00fF
C1976 w_n4520_n851# a_n766_n401# 0.10fF
C1977 a_30_n632# a_n180_n632# 0.03fF
C1978 a_n1348_n632# a_n1440_n632# 0.09fF
C1979 a_n2070_n632# a_n2608_n632# 0.01fF
C1980 a_2970_n632# a_2222_n632# 0.01fF
C1981 a_2010_n100# a_2012_n632# 0.00fF
C1982 a_2340_n632# a_3180_n632# 0.01fF
C1983 a_3852_131# a_3012_131# 0.01fF
C1984 a_n138_n197# a_1122_n197# 0.00fF
C1985 a_2970_n632# a_2642_n632# 0.02fF
C1986 a_2802_n197# a_3432_131# 0.00fF
C1987 a_3222_n197# a_3224_n729# 0.01fF
C1988 a_2640_n100# a_1800_n100# 0.01fF
C1989 a_n510_n100# a_238_n100# 0.01fF
C1990 a_n390_n632# a_n600_n632# 0.03fF
C1991 a_n1140_n100# a_n2610_n100# 0.00fF
C1992 a_n2072_n100# a_n1862_n100# 0.03fF
C1993 a_n2190_n100# a_n3542_n100# 0.00fF
C1994 w_n4520_n851# a_1710_n632# 0.01fF
C1995 a_n3706_n401# a_n2656_n729# 0.00fF
C1996 a_2850_n100# a_1498_n100# 0.00fF
C1997 a_n2490_n632# a_n3868_n632# 0.00fF
C1998 a_238_n100# a_n1022_n100# 0.00fF
C1999 a_4062_n197# a_3012_131# 0.00fF
C2000 a_n930_n100# a_n1232_n100# 0.02fF
C2001 a_1918_n100# a_3270_n100# 0.00fF
C2002 a_n2070_n632# a_n810_n632# 0.00fF
C2003 w_n4520_n851# a_3642_n197# 0.09fF
C2004 a_n138_n197# a_n182_n100# 0.00fF
C2005 a_492_131# a_282_n197# 0.00fF
C2006 a_n720_n100# a_n2190_n100# 0.00fF
C2007 w_n4520_n851# a_n1558_n632# 0.01fF
C2008 a_540_n100# a_330_n100# 0.03fF
C2009 a_1500_n632# a_1592_n632# 0.09fF
C2010 a_2548_n100# a_3178_n100# 0.01fF
C2011 a_962_n632# a_1920_n632# 0.01fF
C2012 a_3388_n100# a_3690_n100# 0.02fF
C2013 w_n4520_n851# a_2430_n100# 0.02fF
C2014 a_4062_n197# a_4064_n729# 0.01fF
C2015 a_n2190_n100# a_n1980_n100# 0.03fF
C2016 a_2640_n100# a_2128_n100# 0.01fF
C2017 a_n1816_n729# a_n1768_n632# 0.00fF
C2018 a_n1560_n100# a_n2492_n100# 0.01fF
C2019 a_n298_n632# a_1080_n632# 0.00fF
C2020 a_2802_n197# w_n4520_n851# 0.10fF
C2021 a_n3332_n100# a_n2072_n100# 0.00fF
C2022 a_n2238_n197# a_n768_131# 0.00fF
C2023 a_912_131# a_72_131# 0.01fF
C2024 w_n4520_n851# a_n3750_n632# 0.04fF
C2025 a_n1860_n632# a_n1768_n632# 0.09fF
C2026 a_n2818_n632# a_n2910_n632# 0.09fF
C2027 a_n3120_n632# a_n2910_n632# 0.03fF
C2028 a_752_n632# a_1710_n632# 0.01fF
C2029 a_1172_n632# a_1710_n632# 0.01fF
C2030 a_n2280_n632# w_n4520_n851# 0.01fF
C2031 a_332_n632# a_n298_n632# 0.01fF
C2032 a_n2700_n632# a_n2818_n632# 0.07fF
C2033 a_n1442_n100# a_n182_n100# 0.00fF
C2034 a_n720_n100# a_238_n100# 0.01fF
C2035 a_n3120_n632# a_n2700_n632# 0.02fF
C2036 a_3902_n632# a_2852_n632# 0.01fF
C2037 a_2220_n100# a_2010_n100# 0.03fF
C2038 a_n3330_n632# a_n3868_n632# 0.01fF
C2039 a_n3286_n401# a_n3076_n729# 0.00fF
C2040 a_n508_n632# a_1080_n632# 0.00fF
C2041 a_n3960_n632# a_n3918_n197# 0.00fF
C2042 a_1542_n197# a_282_n197# 0.00fF
C2043 a_n4080_n100# a_n3542_n100# 0.01fF
C2044 a_962_n632# a_2012_n632# 0.01fF
C2045 a_2222_n632# a_1920_n632# 0.02fF
C2046 a_n3450_n100# a_n2492_n100# 0.01fF
C2047 a_n2702_n100# a_n2492_n100# 0.03fF
C2048 a_n508_n632# a_332_n632# 0.01fF
C2049 a_2642_n632# a_1920_n632# 0.01fF
C2050 a_n2446_n401# a_n1816_n729# 0.00fF
C2051 a_n2400_n100# a_n3962_n100# 0.00fF
C2052 a_2640_n100# a_3808_n100# 0.01fF
C2053 a_n2398_n632# a_n1558_n632# 0.01fF
C2054 a_n3542_n100# a_n3752_n100# 0.03fF
C2055 a_n1818_n197# a_n1770_n100# 0.00fF
C2056 a_870_n632# a_868_n100# 0.00fF
C2057 a_n2238_n197# a_n1188_131# 0.00fF
C2058 a_1288_n100# a_330_n100# 0.01fF
C2059 a_n4128_131# a_n3498_n197# 0.00fF
C2060 a_74_n401# a_n1186_n401# 0.00fF
C2061 a_n1860_n632# a_n718_n632# 0.01fF
C2062 a_240_n632# a_962_n632# 0.01fF
C2063 a_n138_n197# a_n558_n197# 0.01fF
C2064 a_1708_n100# a_868_n100# 0.01fF
C2065 a_1382_n632# a_2550_n632# 0.01fF
C2066 a_30_n632# a_542_n632# 0.01fF
C2067 a_n3540_n632# a_n3868_n632# 0.02fF
C2068 a_n2398_n632# a_n3750_n632# 0.00fF
C2069 a_1380_n100# a_2548_n100# 0.01fF
C2070 a_4064_n729# a_4020_n632# 0.00fF
C2071 a_238_n100# a_1380_n100# 0.01fF
C2072 a_n1560_n100# a_n90_n100# 0.00fF
C2073 a_n2398_n632# a_n2280_n632# 0.07fF
C2074 a_n3238_n632# a_n3658_n632# 0.02fF
C2075 a_2222_n632# a_2012_n632# 0.03fF
C2076 a_448_n100# a_238_n100# 0.03fF
C2077 a_3062_n632# a_3390_n632# 0.02fF
C2078 a_3600_n632# a_3272_n632# 0.02fF
C2079 a_1918_n100# a_2010_n100# 0.09fF
C2080 a_1590_n100# a_1498_n100# 0.09fF
C2081 a_3480_n100# a_3690_n100# 0.03fF
C2082 a_2642_n632# a_2012_n632# 0.01fF
C2083 a_n2190_n100# a_n1652_n100# 0.01fF
C2084 a_n1140_n100# a_n2282_n100# 0.01fF
C2085 a_1708_n100# a_3060_n100# 0.00fF
C2086 a_n392_n100# a_n1862_n100# 0.00fF
C2087 a_n2910_n632# a_n1768_n632# 0.01fF
C2088 a_3014_n401# w_n4520_n851# 0.10fF
C2089 a_n928_n632# a_660_n632# 0.00fF
C2090 w_n4520_n851# a_n1396_n729# 0.12fF
C2091 a_n2820_n100# a_n2400_n100# 0.02fF
C2092 a_n2700_n632# a_n1768_n632# 0.01fF
C2093 a_n390_n632# a_240_n632# 0.01fF
C2094 a_n1860_n632# a_n1816_n729# 0.00fF
C2095 a_n930_n100# a_n2492_n100# 0.00fF
C2096 a_1962_n197# a_1752_131# 0.00fF
C2097 a_2852_n632# a_4112_n632# 0.00fF
C2098 a_1708_n100# a_540_n100# 0.01fF
C2099 a_120_n100# a_n1140_n100# 0.00fF
C2100 a_494_n401# a_74_n401# 0.01fF
C2101 a_1382_n632# a_1290_n632# 0.09fF
C2102 a_3852_131# a_3854_n401# 0.01fF
C2103 a_n2238_n197# a_n978_n197# 0.00fF
C2104 a_2970_n632# a_3810_n632# 0.01fF
C2105 a_1962_n197# a_1122_n197# 0.01fF
C2106 w_n4520_n851# a_1080_n632# 0.01fF
C2107 a_n556_n729# a_n766_n401# 0.00fF
C2108 a_330_n100# a_n182_n100# 0.01fF
C2109 a_2220_n100# a_2222_n632# 0.00fF
C2110 a_n348_131# a_702_n197# 0.00fF
C2111 a_2594_n401# a_1334_n401# 0.00fF
C2112 a_n1978_n632# a_n508_n632# 0.00fF
C2113 a_332_n632# w_n4520_n851# 0.01fF
C2114 a_1802_n632# a_1710_n632# 0.09fF
C2115 a_n2866_n401# a_n2236_n729# 0.00fF
C2116 a_2970_n632# a_2550_n632# 0.02fF
C2117 a_2432_n632# a_3062_n632# 0.01fF
C2118 a_n1348_n632# a_n600_n632# 0.01fF
C2119 a_n4128_131# a_n4126_n401# 0.01fF
C2120 a_n2608_n632# a_n2656_n729# 0.00fF
C2121 a_n2070_n632# a_n3028_n632# 0.01fF
C2122 a_752_n632# a_1080_n632# 0.02fF
C2123 a_2172_131# a_3432_131# 0.00fF
C2124 a_1172_n632# a_1080_n632# 0.09fF
C2125 a_n346_n401# a_1124_n729# 0.00fF
C2126 a_1754_n401# a_1124_n729# 0.00fF
C2127 a_n928_n632# a_122_n632# 0.01fF
C2128 a_2220_n100# a_2338_n100# 0.07fF
C2129 a_3432_131# a_3012_131# 0.01fF
C2130 a_2640_n100# a_3388_n100# 0.01fF
C2131 a_1288_n100# a_1708_n100# 0.02fF
C2132 a_752_n632# a_332_n632# 0.02fF
C2133 a_n3238_n632# a_n3286_n401# 0.00fF
C2134 a_1172_n632# a_332_n632# 0.01fF
C2135 a_n88_n632# a_n810_n632# 0.01fF
C2136 a_914_n401# a_284_n729# 0.00fF
C2137 a_2760_n632# a_1710_n632# 0.01fF
C2138 a_n90_n100# a_n930_n100# 0.01fF
C2139 a_n2070_n632# a_n1138_n632# 0.01fF
C2140 a_n180_n632# a_n1558_n632# 0.00fF
C2141 a_n2818_n632# a_n2866_n401# 0.00fF
C2142 a_n2868_131# a_n2238_n197# 0.00fF
C2143 a_n390_n632# a_n392_n100# 0.00fF
C2144 a_2430_n100# a_2548_n100# 0.07fF
C2145 a_120_n100# a_1590_n100# 0.00fF
C2146 w_n4520_n851# a_2172_131# 0.12fF
C2147 a_n2608_n632# a_n1230_n632# 0.00fF
C2148 a_n1862_n100# a_n812_n100# 0.01fF
C2149 a_2384_n729# w_n4520_n851# 0.12fF
C2150 a_2968_n100# a_1498_n100# 0.00fF
C2151 a_3390_n632# a_3434_n401# 0.00fF
C2152 a_1754_n401# a_2174_n401# 0.01fF
C2153 a_n1022_n100# a_n2610_n100# 0.00fF
C2154 w_n4520_n851# a_3012_131# 0.13fF
C2155 a_n1860_n632# a_n2910_n632# 0.01fF
C2156 a_2760_n632# a_2802_n197# 0.00fF
C2157 a_n3916_n729# a_n3868_n632# 0.00fF
C2158 a_2852_n632# a_2340_n632# 0.01fF
C2159 a_n812_n100# a_n768_131# 0.00fF
C2160 a_n2026_n401# w_n4520_n851# 0.10fF
C2161 a_912_131# a_n348_131# 0.00fF
C2162 a_3390_n632# a_3272_n632# 0.07fF
C2163 a_n1650_n632# a_n298_n632# 0.00fF
C2164 a_n1860_n632# a_n2700_n632# 0.01fF
C2165 a_4064_n729# w_n4520_n851# 0.11fF
C2166 a_3224_n729# a_3644_n729# 0.01fF
C2167 a_n810_n632# a_n1230_n632# 0.02fF
C2168 a_n3496_n729# a_n3286_n401# 0.00fF
C2169 a_n4128_131# a_n4172_n100# 0.00fF
C2170 a_n3030_n100# w_n4520_n851# 0.03fF
C2171 a_1708_n100# a_1752_131# 0.00fF
C2172 a_n2820_n100# a_n2072_n100# 0.01fF
C2173 a_2550_n632# a_1920_n632# 0.01fF
C2174 a_1918_n100# a_2338_n100# 0.02fF
C2175 a_n3542_n100# a_n2610_n100# 0.01fF
C2176 a_1332_131# a_702_n197# 0.00fF
C2177 a_n300_n100# a_n392_n100# 0.09fF
C2178 a_n3870_n100# w_n4520_n851# 0.05fF
C2179 a_n2656_n729# a_n1186_n401# 0.00fF
C2180 a_2850_n100# a_2758_n100# 0.09fF
C2181 a_n1350_n100# a_n1140_n100# 0.03fF
C2182 a_n508_n632# a_n1650_n632# 0.01fF
C2183 a_n1978_n632# w_n4520_n851# 0.01fF
C2184 a_n3750_n632# a_n3752_n100# 0.00fF
C2185 a_n1980_n100# a_n2610_n100# 0.01fF
C2186 a_n3660_n100# a_n2492_n100# 0.01fF
C2187 a_870_n632# a_n718_n632# 0.00fF
C2188 a_n3750_n632# a_n3868_n632# 0.07fF
C2189 a_2640_n100# a_3480_n100# 0.01fF
C2190 a_n1650_n632# a_n1608_131# 0.00fF
C2191 a_n2280_n632# a_n3868_n632# 0.00fF
C2192 a_2550_n632# a_2012_n632# 0.01fF
C2193 a_2804_n729# a_3644_n729# 0.01fF
C2194 a_n556_n729# a_n1396_n729# 0.01fF
C2195 a_542_n632# a_1710_n632# 0.01fF
C2196 a_n1230_n632# a_n1186_n401# 0.00fF
C2197 a_n1560_n100# a_n2400_n100# 0.01fF
C2198 a_1590_n100# a_1078_n100# 0.01fF
C2199 a_658_n100# a_1590_n100# 0.01fF
C2200 a_1964_n729# a_1334_n401# 0.00fF
C2201 a_n2028_131# a_n1398_n197# 0.00fF
C2202 a_2850_n100# a_3900_n100# 0.01fF
C2203 a_n346_n401# a_n766_n401# 0.01fF
C2204 a_2432_n632# a_3272_n632# 0.01fF
C2205 a_2432_n632# a_1500_n632# 0.01fF
C2206 a_3060_n100# a_3690_n100# 0.01fF
C2207 a_1920_n632# a_1290_n632# 0.01fF
C2208 a_n1348_n632# a_240_n632# 0.00fF
C2209 a_n602_n100# a_n1862_n100# 0.00fF
C2210 a_870_n632# a_2130_n632# 0.00fF
C2211 a_4110_n100# a_2758_n100# 0.00fF
C2212 a_n718_n632# a_660_n632# 0.00fF
C2213 a_1802_n632# a_1080_n632# 0.01fF
C2214 a_2970_n632# a_3902_n632# 0.01fF
C2215 a_n2070_n632# a_n2490_n632# 0.02fF
C2216 a_2220_n100# a_1800_n100# 0.02fF
C2217 a_n2700_n632# a_n2910_n632# 0.03fF
C2218 a_450_n632# a_962_n632# 0.01fF
C2219 a_n1978_n632# a_n2398_n632# 0.02fF
C2220 a_1754_n401# a_1710_n632# 0.00fF
C2221 a_912_131# a_1332_131# 0.01fF
C2222 a_868_n100# a_1170_n100# 0.02fF
C2223 a_n2658_n197# a_n1608_131# 0.00fF
C2224 a_1802_n632# a_332_n632# 0.00fF
C2225 a_2130_n632# a_3180_n632# 0.01fF
C2226 a_n2446_n401# a_n2866_n401# 0.01fF
C2227 a_n2400_n100# a_n3450_n100# 0.01fF
C2228 a_1380_n100# a_1332_131# 0.00fF
C2229 a_n1022_n100# a_n2282_n100# 0.00fF
C2230 a_n2400_n100# a_n2702_n100# 0.02fF
C2231 a_240_n632# a_282_n197# 0.00fF
C2232 a_n180_n632# a_1080_n632# 0.00fF
C2233 a_n3660_n100# a_n3708_131# 0.00fF
C2234 a_1380_n100# a_1498_n100# 0.07fF
C2235 a_n2912_n100# a_n3542_n100# 0.01fF
C2236 a_2220_n100# a_2128_n100# 0.09fF
C2237 a_n1020_n632# a_n928_n632# 0.09fF
C2238 a_2382_n197# a_1542_n197# 0.01fF
C2239 a_660_n632# a_2130_n632# 0.00fF
C2240 a_2012_n632# a_1290_n632# 0.01fF
C2241 a_4110_n100# a_3900_n100# 0.03fF
C2242 a_448_n100# a_1498_n100# 0.01fF
C2243 a_n300_n100# a_n812_n100# 0.01fF
C2244 a_n180_n632# a_332_n632# 0.01fF
C2245 a_120_n100# a_n510_n100# 0.01fF
C2246 a_n2610_n100# a_n1652_n100# 0.01fF
C2247 w_n4520_n851# a_3270_n100# 0.03fF
C2248 a_n2070_n632# a_n3330_n632# 0.00fF
C2249 a_n2070_n632# a_n2188_n632# 0.07fF
C2250 a_n1650_n632# w_n4520_n851# 0.01fF
C2251 a_1590_n100# a_2758_n100# 0.01fF
C2252 a_3600_n632# a_3692_n632# 0.09fF
C2253 a_n3542_n100# a_n2282_n100# 0.00fF
C2254 a_n2912_n100# a_n1980_n100# 0.01fF
C2255 a_n976_n729# a_n1020_n632# 0.00fF
C2256 a_120_n100# a_n1022_n100# 0.01fF
C2257 a_2220_n100# a_960_n100# 0.00fF
C2258 a_450_n632# a_n390_n632# 0.01fF
C2259 a_240_n632# a_1290_n632# 0.01fF
C2260 a_30_n632# a_74_n401# 0.00fF
C2261 a_284_n729# a_n1186_n401# 0.00fF
C2262 a_n2656_n729# a_n1606_n401# 0.00fF
C2263 a_n720_n100# a_n2282_n100# 0.00fF
C2264 a_3854_n401# w_n4520_n851# 0.08fF
C2265 a_1918_n100# a_1800_n100# 0.07fF
C2266 a_2382_n197# a_3222_n197# 0.01fF
C2267 a_n1232_n100# a_n182_n100# 0.01fF
C2268 a_n90_n100# a_868_n100# 0.01fF
C2269 a_n1980_n100# a_n2282_n100# 0.02fF
C2270 a_n718_n632# a_122_n632# 0.01fF
C2271 a_540_n100# a_1170_n100# 0.01fF
C2272 a_n1140_n100# a_n1770_n100# 0.01fF
C2273 a_n1816_n729# a_n2866_n401# 0.00fF
C2274 a_2220_n100# a_3808_n100# 0.00fF
C2275 a_n3540_n632# a_n2070_n632# 0.00fF
C2276 a_n88_n632# a_n1138_n632# 0.01fF
C2277 a_n3238_n632# a_n4078_n632# 0.01fF
C2278 a_1544_n729# a_2594_n401# 0.00fF
C2279 a_n298_n632# a_962_n632# 0.00fF
C2280 a_n556_n729# a_n2026_n401# 0.00fF
C2281 a_30_n632# a_1500_n632# 0.00fF
C2282 w_n4520_n851# a_n3288_131# 0.13fF
C2283 a_1918_n100# a_2128_n100# 0.03fF
C2284 a_120_n100# a_n720_n100# 0.01fF
C2285 a_1382_n632# a_2340_n632# 0.01fF
C2286 a_2970_n632# a_4112_n632# 0.01fF
C2287 w_n4520_n851# a_n2658_n197# 0.10fF
C2288 a_n2400_n100# a_n930_n100# 0.00fF
C2289 a_n2190_n100# a_n3030_n100# 0.01fF
C2290 a_n392_n100# a_960_n100# 0.00fF
C2291 a_n1560_n100# a_n2072_n100# 0.01fF
C2292 a_n768_131# a_n1608_131# 0.01fF
C2293 a_n2398_n632# a_n1650_n632# 0.01fF
C2294 a_n3238_n632# a_n4170_n632# 0.01fF
C2295 a_n1232_n100# a_n1442_n100# 0.03fF
C2296 a_n1440_n632# a_n928_n632# 0.01fF
C2297 a_2642_n632# a_4020_n632# 0.00fF
C2298 a_1708_n100# a_330_n100# 0.00fF
C2299 a_n508_n632# a_962_n632# 0.00fF
C2300 a_1918_n100# a_960_n100# 0.01fF
C2301 a_n3918_n197# a_n3498_n197# 0.01fF
C2302 a_n1230_n632# a_n1138_n632# 0.09fF
C2303 a_n90_n100# a_540_n100# 0.01fF
C2304 a_3014_n401# a_1754_n401# 0.00fF
C2305 a_494_n401# a_284_n729# 0.00fF
C2306 a_n510_n100# a_1078_n100# 0.00fF
C2307 a_542_n632# a_1080_n632# 0.01fF
C2308 a_n510_n100# a_658_n100# 0.01fF
C2309 a_1124_n729# a_74_n401# 0.00fF
C2310 a_1288_n100# a_1170_n100# 0.07fF
C2311 a_n346_n401# a_n1396_n729# 0.00fF
C2312 a_4018_n100# a_4062_n197# 0.00fF
C2313 a_n390_n632# a_n298_n632# 0.09fF
C2314 a_658_n100# a_702_n197# 0.00fF
C2315 a_n3030_n100# a_n3078_n197# 0.00fF
C2316 a_n300_n100# a_n602_n100# 0.02fF
C2317 a_n2912_n100# a_n1652_n100# 0.00fF
C2318 a_n4128_131# a_n3918_n197# 0.00fF
C2319 a_120_n100# a_1380_n100# 0.00fF
C2320 a_n2072_n100# a_n3450_n100# 0.00fF
C2321 a_n136_n729# w_n4520_n851# 0.12fF
C2322 a_2010_n100# w_n4520_n851# 0.02fF
C2323 a_542_n632# a_332_n632# 0.03fF
C2324 a_n2072_n100# a_n2702_n100# 0.01fF
C2325 a_n2866_n401# a_n4126_n401# 0.00fF
C2326 a_120_n100# a_448_n100# 0.02fF
C2327 a_n1188_131# a_n1608_131# 0.01fF
C2328 a_n4080_n100# a_n3030_n100# 0.01fF
C2329 a_2802_n197# a_1332_131# 0.00fF
C2330 a_540_n100# a_492_131# 0.00fF
C2331 a_1498_n100# a_2430_n100# 0.01fF
C2332 a_n2282_n100# a_n1652_n100# 0.01fF
C2333 a_n390_n632# a_n508_n632# 0.07fF
C2334 a_n510_n100# a_n1350_n100# 0.01fF
C2335 a_2968_n100# a_2758_n100# 0.03fF
C2336 a_3062_n632# a_1710_n632# 0.00fF
C2337 a_n3870_n100# a_n4080_n100# 0.03fF
C2338 w_n4520_n851# a_n1862_n100# 0.02fF
C2339 a_n2910_n632# a_n2866_n401# 0.00fF
C2340 a_n3122_n100# a_n3542_n100# 0.02fF
C2341 a_n3030_n100# a_n3752_n100# 0.01fF
C2342 a_2640_n100# a_3060_n100# 0.02fF
C2343 a_n1440_n632# a_n2818_n632# 0.00fF
C2344 a_n1350_n100# a_n1022_n100# 0.02fF
C2345 a_n720_n100# a_658_n100# 0.00fF
C2346 a_3390_n632# a_3692_n632# 0.02fF
C2347 a_n3240_n100# a_n3542_n100# 0.02fF
C2348 a_n300_n100# a_n298_n632# 0.00fF
C2349 a_n3870_n100# a_n3752_n100# 0.07fF
C2350 w_n4520_n851# a_n768_131# 0.12fF
C2351 a_n1020_n632# a_n1768_n632# 0.01fF
C2352 a_750_n100# a_2010_n100# 0.00fF
C2353 a_3434_n401# a_2174_n401# 0.00fF
C2354 a_3852_131# a_3810_n632# 0.00fF
C2355 a_1288_n100# a_n90_n100# 0.00fF
C2356 a_2970_n632# a_2340_n632# 0.01fF
C2357 a_n3122_n100# a_n1980_n100# 0.01fF
C2358 a_n3448_n632# a_n2608_n632# 0.01fF
C2359 a_3598_n100# a_3690_n100# 0.09fF
C2360 a_1170_n100# a_1122_n197# 0.00fF
C2361 a_n3332_n100# w_n4520_n851# 0.03fF
C2362 a_n3870_n100# a_n3868_n632# 0.00fF
C2363 a_n3240_n100# a_n1980_n100# 0.00fF
C2364 a_4018_n100# a_4020_n632# 0.00fF
C2365 a_2220_n100# a_3388_n100# 0.01fF
C2366 a_2968_n100# a_3900_n100# 0.01fF
C2367 a_n182_n100# a_1170_n100# 0.00fF
C2368 a_n720_n100# a_n1350_n100# 0.01fF
C2369 w_n4520_n851# a_962_n632# 0.01fF
C2370 a_n300_n100# a_28_n100# 0.02fF
C2371 a_n2072_n100# a_n930_n100# 0.01fF
C2372 a_n1232_n100# a_330_n100# 0.00fF
C2373 a_n1560_n100# a_n392_n100# 0.01fF
C2374 a_2758_n100# a_3178_n100# 0.02fF
C2375 a_1544_n729# a_1964_n729# 0.01fF
C2376 a_n1350_n100# a_n1980_n100# 0.01fF
C2377 a_1380_n100# a_1078_n100# 0.02fF
C2378 a_658_n100# a_1380_n100# 0.01fF
C2379 a_n978_n197# a_n1608_131# 0.00fF
C2380 a_n3496_n729# a_n3450_n100# 0.00fF
C2381 a_n3658_n632# w_n4520_n851# 0.04fF
C2382 a_2384_n729# a_1754_n401# 0.00fF
C2383 w_n4520_n851# a_n1188_131# 0.12fF
C2384 a_n2400_n100# a_n3660_n100# 0.00fF
C2385 a_448_n100# a_1078_n100# 0.01fF
C2386 a_658_n100# a_448_n100# 0.03fF
C2387 a_n1020_n632# a_n718_n632# 0.02fF
C2388 a_n1442_n100# a_n2492_n100# 0.01fF
C2389 a_n2072_n100# a_n2028_131# 0.00fF
C2390 a_n2490_n632# a_n1230_n632# 0.00fF
C2391 a_n180_n632# a_n1650_n632# 0.00fF
C2392 a_30_n632# a_n88_n632# 0.07fF
C2393 a_1382_n632# a_1334_n401# 0.00fF
C2394 a_2548_n100# a_3270_n100# 0.01fF
C2395 a_752_n632# a_962_n632# 0.03fF
C2396 a_1172_n632# a_962_n632# 0.03fF
C2397 a_74_n401# a_n766_n401# 0.01fF
C2398 a_n2238_n197# a_n2028_131# 0.00fF
C2399 a_2432_n632# a_3692_n632# 0.00fF
C2400 a_n2280_n632# a_n2282_n100# 0.00fF
C2401 a_2222_n632# w_n4520_n851# 0.01fF
C2402 a_2640_n100# a_1288_n100# 0.00fF
C2403 a_870_n632# a_660_n632# 0.03fF
C2404 a_494_n401# a_914_n401# 0.01fF
C2405 a_n1440_n632# a_n1768_n632# 0.02fF
C2406 a_3852_131# a_3808_n100# 0.00fF
C2407 a_2852_n632# a_2130_n632# 0.01fF
C2408 a_3900_n100# a_3178_n100# 0.01fF
C2409 a_2340_n632# a_1920_n632# 0.02fF
C2410 a_n90_n100# a_n182_n100# 0.09fF
C2411 a_n390_n632# w_n4520_n851# 0.01fF
C2412 a_2642_n632# w_n4520_n851# 0.02fF
C2413 a_1918_n100# a_3388_n100# 0.00fF
C2414 a_492_131# a_1752_131# 0.00fF
C2415 a_3810_n632# a_4020_n632# 0.03fF
C2416 a_n2070_n632# a_n1558_n632# 0.01fF
C2417 a_n138_n197# a_n90_n100# 0.00fF
C2418 a_n3238_n632# a_n3960_n632# 0.01fF
C2419 a_30_n632# a_n1230_n632# 0.00fF
C2420 a_492_131# a_1122_n197# 0.00fF
C2421 a_n3122_n100# a_n1652_n100# 0.00fF
C2422 a_n1230_n632# a_n2188_n632# 0.01fF
C2423 a_3014_n401# a_3062_n632# 0.00fF
C2424 a_n2398_n632# a_n3658_n632# 0.00fF
C2425 a_n2868_131# a_n1608_131# 0.00fF
C2426 a_2338_n100# w_n4520_n851# 0.02fF
C2427 a_752_n632# a_2222_n632# 0.00fF
C2428 a_n2070_n632# a_n2280_n632# 0.03fF
C2429 a_n3240_n100# a_n1652_n100# 0.00fF
C2430 a_1380_n100# a_2758_n100# 0.00fF
C2431 a_n510_n100# a_n1770_n100# 0.00fF
C2432 a_1172_n632# a_2222_n632# 0.01fF
C2433 a_n1860_n632# a_n1020_n632# 0.01fF
C2434 a_n3078_n197# a_n3288_131# 0.00fF
C2435 a_n3708_131# a_n3498_n197# 0.00fF
C2436 a_2550_n632# a_4020_n632# 0.00fF
C2437 a_2220_n100# a_3480_n100# 0.00fF
C2438 a_n3288_131# a_n2448_131# 0.01fF
C2439 a_752_n632# a_n390_n632# 0.01fF
C2440 a_1172_n632# a_2642_n632# 0.00fF
C2441 a_3272_n632# a_1710_n632# 0.00fF
C2442 a_1500_n632# a_1710_n632# 0.03fF
C2443 a_n390_n632# a_1172_n632# 0.00fF
C2444 a_960_n100# a_n602_n100# 0.00fF
C2445 a_n1022_n100# a_n1770_n100# 0.01fF
C2446 w_n4520_n851# a_n978_n197# 0.10fF
C2447 a_450_n632# a_1290_n632# 0.01fF
C2448 a_n2658_n197# a_n3078_n197# 0.01fF
C2449 a_n928_n632# a_n600_n632# 0.02fF
C2450 a_1964_n729# a_1962_n197# 0.01fF
C2451 a_n138_n197# a_492_131# 0.00fF
C2452 a_2340_n632# a_2012_n632# 0.02fF
C2453 a_n2658_n197# a_n2448_131# 0.00fF
C2454 a_n90_n100# a_n1442_n100# 0.00fF
C2455 a_n718_n632# a_n1440_n632# 0.01fF
C2456 a_n300_n100# w_n4520_n851# 0.02fF
C2457 a_n1350_n100# a_n1652_n100# 0.02fF
C2458 a_1542_n197# a_1752_131# 0.00fF
C2459 a_n4128_131# a_n3708_131# 0.01fF
C2460 a_n556_n729# a_n136_n729# 0.01fF
C2461 a_n2236_n729# a_n3076_n729# 0.01fF
C2462 a_n1348_n632# a_n298_n632# 0.01fF
C2463 a_n1560_n100# a_n812_n100# 0.01fF
C2464 a_1542_n197# a_1122_n197# 0.01fF
C2465 a_2338_n100# a_750_n100# 0.00fF
C2466 a_870_n632# a_122_n632# 0.01fF
C2467 w_n4520_n851# a_n3286_n401# 0.10fF
C2468 a_n768_131# a_72_131# 0.01fF
C2469 a_n392_n100# a_n930_n100# 0.01fF
C2470 a_n136_n729# a_n180_n632# 0.00fF
C2471 a_n2190_n100# a_n1862_n100# 0.02fF
C2472 a_n720_n100# a_n1770_n100# 0.01fF
C2473 a_n1440_n632# a_n1442_n100# 0.00fF
C2474 a_2010_n100# a_2548_n100# 0.01fF
C2475 a_3222_n197# a_1752_131# 0.00fF
C2476 a_n1770_n100# a_n1980_n100# 0.03fF
C2477 a_n138_n197# a_n1398_n197# 0.00fF
C2478 a_n1348_n632# a_n508_n632# 0.01fF
C2479 a_n3030_n100# a_n2610_n100# 0.02fF
C2480 a_n300_n100# a_750_n100# 0.01fF
C2481 a_2172_131# a_1332_131# 0.01fF
C2482 a_2430_n100# a_1078_n100# 0.00fF
C2483 a_n2072_n100# a_n3660_n100# 0.00fF
C2484 a_1918_n100# a_3480_n100# 0.00fF
C2485 a_4018_n100# w_n4520_n851# 0.08fF
C2486 a_n3120_n632# a_n3076_n729# 0.00fF
C2487 a_n3870_n100# a_n2610_n100# 0.00fF
C2488 w_n4520_n851# a_n3962_n100# 0.06fF
C2489 a_330_n100# a_1170_n100# 0.01fF
C2490 a_n3332_n100# a_n2190_n100# 0.01fF
C2491 w_n4520_n851# a_n2868_131# 0.12fF
C2492 a_660_n632# a_122_n632# 0.01fF
C2493 a_n1860_n632# a_n1440_n632# 0.02fF
C2494 a_n558_n197# a_492_131# 0.00fF
C2495 a_2640_n100# a_3598_n100# 0.01fF
C2496 a_960_n100# a_28_n100# 0.01fF
C2497 a_n298_n632# a_1290_n632# 0.00fF
C2498 a_n1188_131# a_72_131# 0.00fF
C2499 a_1802_n632# a_962_n632# 0.01fF
C2500 a_3224_n729# w_n4520_n851# 0.12fF
C2501 a_n1442_n100# a_n1398_n197# 0.00fF
C2502 a_n3448_n632# a_n3028_n632# 0.02fF
C2503 a_74_n401# a_n1396_n729# 0.00fF
C2504 a_3014_n401# a_3434_n401# 0.01fF
C2505 a_n2608_n632# a_n3028_n632# 0.02fF
C2506 a_n180_n632# a_962_n632# 0.01fF
C2507 a_n558_n197# a_n1398_n197# 0.01fF
C2508 w_n4520_n851# a_704_n729# 0.12fF
C2509 a_n90_n100# a_330_n100# 0.02fF
C2510 a_2758_n100# a_2430_n100# 0.02fF
C2511 a_n1560_n100# a_n602_n100# 0.01fF
C2512 w_n4520_n851# a_3810_n632# 0.05fF
C2513 w_n4520_n851# a_1800_n100# 0.02fF
C2514 a_n2820_n100# w_n4520_n851# 0.02fF
C2515 a_n3332_n100# a_n4080_n100# 0.01fF
C2516 a_1544_n729# a_1542_n197# 0.01fF
C2517 a_1802_n632# a_2222_n632# 0.02fF
C2518 a_2802_n197# a_2758_n100# 0.00fF
C2519 a_n2608_n632# a_n1138_n632# 0.00fF
C2520 a_n3916_n729# a_n2656_n729# 0.00fF
C2521 a_1590_n100# a_1592_n632# 0.00fF
C2522 a_284_n729# a_1124_n729# 0.01fF
C2523 a_1802_n632# a_2642_n632# 0.01fF
C2524 a_2804_n729# w_n4520_n851# 0.12fF
C2525 a_n930_n100# a_n812_n100# 0.07fF
C2526 a_n3332_n100# a_n3752_n100# 0.02fF
C2527 a_n1770_n100# a_n1652_n100# 0.07fF
C2528 a_240_n632# a_n928_n632# 0.01fF
C2529 a_3902_n632# a_4020_n632# 0.07fF
C2530 a_n1188_131# a_n2448_131# 0.00fF
C2531 a_1382_n632# a_2130_n632# 0.01fF
C2532 a_n2236_n729# a_n2238_n197# 0.01fF
C2533 a_2128_n100# w_n4520_n851# 0.02fF
C2534 a_n2912_n100# a_n3030_n100# 0.07fF
C2535 a_n1140_n100# a_n1186_n401# 0.00fF
C2536 a_752_n632# a_704_n729# 0.00fF
C2537 a_2550_n632# w_n4520_n851# 0.01fF
C2538 a_1500_n632# a_1080_n632# 0.02fF
C2539 a_n1348_n632# w_n4520_n851# 0.01fF
C2540 a_n810_n632# a_n1138_n632# 0.02fF
C2541 a_n978_n197# a_72_131# 0.00fF
C2542 a_n600_n632# a_n1768_n632# 0.01fF
C2543 a_750_n100# a_704_n729# 0.00fF
C2544 a_n1440_n632# a_n2910_n632# 0.00fF
C2545 a_n390_n632# a_n180_n632# 0.03fF
C2546 a_n3870_n100# a_n2912_n100# 0.01fF
C2547 a_1964_n729# a_2594_n401# 0.00fF
C2548 a_750_n100# a_1800_n100# 0.01fF
C2549 a_2760_n632# a_2222_n632# 0.01fF
C2550 a_3900_n100# a_2430_n100# 0.00fF
C2551 a_1962_n197# a_492_131# 0.00fF
C2552 a_n3030_n100# a_n2282_n100# 0.01fF
C2553 a_n2700_n632# a_n1440_n632# 0.00fF
C2554 a_n88_n632# a_n1558_n632# 0.00fF
C2555 a_332_n632# a_1500_n632# 0.01fF
C2556 a_2760_n632# a_2642_n632# 0.07fF
C2557 a_n346_n401# a_n136_n729# 0.00fF
C2558 a_2220_n100# a_868_n100# 0.00fF
C2559 a_960_n100# w_n4520_n851# 0.02fF
C2560 a_2432_n632# a_1592_n632# 0.01fF
C2561 w_n4520_n851# a_282_n197# 0.10fF
C2562 a_n3870_n100# a_n2282_n100# 0.00fF
C2563 a_n1186_n401# a_n1606_n401# 0.01fF
C2564 a_n2446_n401# a_n2400_n100# 0.00fF
C2565 a_n3658_n632# a_n3868_n632# 0.03fF
C2566 a_1172_n632# a_2550_n632# 0.00fF
C2567 a_1080_n632# a_1078_n100# 0.00fF
C2568 a_2222_n632# a_3482_n632# 0.00fF
C2569 a_2128_n100# a_750_n100# 0.00fF
C2570 a_2338_n100# a_2548_n100# 0.03fF
C2571 a_1708_n100# a_1170_n100# 0.01fF
C2572 a_n2446_n401# a_n3076_n729# 0.00fF
C2573 a_n2070_n632# a_n2026_n401# 0.00fF
C2574 a_3600_n632# a_3390_n632# 0.03fF
C2575 a_2642_n632# a_3482_n632# 0.01fF
C2576 w_n4520_n851# a_3808_n100# 0.05fF
C2577 a_n1560_n100# a_28_n100# 0.00fF
C2578 a_n1350_n100# a_n1396_n729# 0.00fF
C2579 a_2220_n100# a_3060_n100# 0.01fF
C2580 a_n718_n632# a_n600_n632# 0.07fF
C2581 a_n1230_n632# a_n1558_n632# 0.02fF
C2582 a_2384_n729# a_3434_n401# 0.00fF
C2583 a_n1138_n632# a_n1186_n401# 0.00fF
C2584 a_n1348_n632# a_n2398_n632# 0.01fF
C2585 a_2852_n632# a_3180_n632# 0.02fF
C2586 a_542_n632# a_962_n632# 0.02fF
C2587 a_1962_n197# a_1542_n197# 0.01fF
C2588 a_n3238_n632# a_n2818_n632# 0.02fF
C2589 w_n4520_n851# a_1290_n632# 0.01fF
C2590 a_n3238_n632# a_n3120_n632# 0.07fF
C2591 a_n300_n100# a_238_n100# 0.01fF
C2592 a_n978_n197# a_n2448_131# 0.00fF
C2593 a_n3496_n729# a_n2236_n729# 0.00fF
C2594 a_750_n100# a_960_n100# 0.03fF
C2595 a_n1560_n100# a_n1608_131# 0.00fF
C2596 a_n2400_n100# a_n1442_n100# 0.01fF
C2597 a_n392_n100# a_868_n100# 0.00fF
C2598 a_n2610_n100# a_n2658_n197# 0.00fF
C2599 a_n2070_n632# a_n1978_n632# 0.09fF
C2600 a_4110_n100# a_2850_n100# 0.00fF
C2601 a_4064_n729# a_3434_n401# 0.00fF
C2602 a_n2280_n632# a_n1230_n632# 0.01fF
C2603 a_1918_n100# a_868_n100# 0.01fF
C2604 a_n3448_n632# a_n2490_n632# 0.01fF
C2605 w_n4520_n851# a_n4078_n632# 0.08fF
C2606 a_n602_n100# a_n930_n100# 0.02fF
C2607 a_4112_n632# a_4020_n632# 0.09fF
C2608 a_2970_n632# a_2130_n632# 0.01fF
C2609 a_n768_131# a_n348_131# 0.01fF
C2610 a_3222_n197# a_1962_n197# 0.00fF
C2611 a_3852_131# a_2382_n197# 0.00fF
C2612 a_n1816_n729# a_n3076_n729# 0.00fF
C2613 a_n2490_n632# a_n2608_n632# 0.07fF
C2614 a_752_n632# a_1290_n632# 0.01fF
C2615 a_1172_n632# a_1290_n632# 0.07fF
C2616 a_284_n729# a_n766_n401# 0.00fF
C2617 a_4018_n100# a_2548_n100# 0.00fF
C2618 w_n4520_n851# a_n4170_n632# 0.14fF
C2619 a_542_n632# a_n390_n632# 0.01fF
C2620 a_1918_n100# a_3060_n100# 0.01fF
C2621 a_n1860_n632# a_n600_n632# 0.00fF
C2622 a_914_n401# a_1124_n729# 0.00fF
C2623 a_n558_n197# a_n600_n632# 0.00fF
C2624 a_2432_n632# a_3600_n632# 0.01fF
C2625 a_30_n632# a_1592_n632# 0.00fF
C2626 a_n392_n100# a_540_n100# 0.01fF
C2627 a_1590_n100# a_2850_n100# 0.00fF
C2628 a_n3448_n632# a_n3330_n632# 0.07fF
C2629 a_n2868_131# a_n3078_n197# 0.00fF
C2630 a_n3448_n632# a_n2188_n632# 0.00fF
C2631 a_n2868_131# a_n2448_131# 0.01fF
C2632 a_n2656_n729# a_n1396_n729# 0.00fF
C2633 a_n1232_n100# a_n2492_n100# 0.00fF
C2634 a_912_131# a_914_n401# 0.01fF
C2635 a_n3330_n632# a_n2608_n632# 0.01fF
C2636 a_n556_n729# a_704_n729# 0.00fF
C2637 a_n2608_n632# a_n2188_n632# 0.02fF
C2638 a_n3122_n100# a_n3030_n100# 0.09fF
C2639 a_1918_n100# a_540_n100# 0.00fF
C2640 a_n3916_n729# a_n3706_n401# 0.00fF
C2641 a_n1140_n100# a_n1138_n632# 0.00fF
C2642 a_2220_n100# a_1288_n100# 0.01fF
C2643 a_1802_n632# a_1800_n100# 0.00fF
C2644 a_n4080_n100# a_n3962_n100# 0.07fF
C2645 a_3388_n100# a_3432_131# 0.00fF
C2646 a_n1188_131# a_n348_131# 0.01fF
C2647 a_n2820_n100# a_n2190_n100# 0.01fF
C2648 a_n1862_n100# a_n2610_n100# 0.01fF
C2649 a_n1560_n100# w_n4520_n851# 0.02fF
C2650 a_n346_n401# a_n390_n632# 0.00fF
C2651 a_3902_n632# w_n4520_n851# 0.06fF
C2652 a_n3238_n632# a_n1768_n632# 0.00fF
C2653 a_n3240_n100# a_n3030_n100# 0.03fF
C2654 a_n3870_n100# a_n3122_n100# 0.01fF
C2655 a_914_n401# a_2174_n401# 0.00fF
C2656 a_n1020_n632# a_122_n632# 0.01fF
C2657 a_n3752_n100# a_n3962_n100# 0.03fF
C2658 a_2010_n100# a_1498_n100# 0.01fF
C2659 a_n88_n632# a_1080_n632# 0.01fF
C2660 a_30_n632# a_n810_n632# 0.01fF
C2661 a_3642_n197# a_2592_131# 0.00fF
C2662 a_n3240_n100# a_n3870_n100# 0.01fF
C2663 a_n3540_n632# a_n3448_n632# 0.09fF
C2664 a_n810_n632# a_n2188_n632# 0.00fF
C2665 a_n930_n100# a_28_n100# 0.01fF
C2666 a_1920_n632# a_2130_n632# 0.03fF
C2667 a_2640_n100# a_1708_n100# 0.01fF
C2668 a_n3076_n729# a_n4126_n401# 0.00fF
C2669 a_1802_n632# a_2550_n632# 0.01fF
C2670 a_n3332_n100# a_n2610_n100# 0.01fF
C2671 a_1800_n100# a_2548_n100# 0.01fF
C2672 a_n3540_n632# a_n2608_n632# 0.01fF
C2673 a_n88_n632# a_332_n632# 0.02fF
C2674 a_n2070_n632# a_n1650_n632# 0.02fF
C2675 a_238_n100# a_1800_n100# 0.00fF
C2676 a_2802_n197# a_2592_131# 0.00fF
C2677 w_n4520_n851# a_3388_n100# 0.03fF
C2678 a_2760_n632# a_3810_n632# 0.01fF
C2679 a_n390_n632# a_n348_131# 0.00fF
C2680 a_282_n197# a_72_131# 0.00fF
C2681 w_n4520_n851# a_n3450_n100# 0.03fF
C2682 w_n4520_n851# a_n2702_n100# 0.02fF
C2683 a_n2238_n197# a_n3498_n197# 0.00fF
C2684 a_n2072_n100# a_n1442_n100# 0.01fF
C2685 a_n300_n100# a_n346_n401# 0.00fF
C2686 a_2760_n632# a_2804_n729# 0.00fF
C2687 a_240_n632# a_n718_n632# 0.01fF
C2688 a_n3706_n401# a_n3750_n632# 0.00fF
C2689 a_n1348_n632# a_n180_n632# 0.01fF
C2690 a_2128_n100# a_2548_n100# 0.02fF
C2691 a_2550_n632# a_2548_n100# 0.00fF
C2692 a_n2820_n100# a_n4080_n100# 0.00fF
C2693 a_n90_n100# a_n1232_n100# 0.01fF
C2694 a_3810_n632# a_3482_n632# 0.02fF
C2695 a_n2028_131# a_n1608_131# 0.01fF
C2696 a_1918_n100# a_1288_n100# 0.01fF
C2697 a_2760_n632# a_2550_n632# 0.03fF
C2698 a_2012_n632# a_2130_n632# 0.07fF
C2699 a_2640_n100# a_2594_n401# 0.00fF
C2700 a_332_n632# a_n1230_n632# 0.00fF
C2701 a_n978_n197# a_n348_131# 0.00fF
C2702 a_n2820_n100# a_n3752_n100# 0.01fF
C2703 a_3272_n632# a_3270_n100# 0.00fF
C2704 a_3854_n401# a_3434_n401# 0.01fF
C2705 a_3222_n197# a_3180_n632# 0.00fF
C2706 a_870_n632# a_1382_n632# 0.01fF
C2707 a_n300_n100# a_n348_131# 0.00fF
C2708 a_960_n100# a_2548_n100# 0.00fF
C2709 a_540_n100# a_n812_n100# 0.00fF
C2710 a_238_n100# a_960_n100# 0.01fF
C2711 a_n1440_n632# a_122_n632# 0.00fF
C2712 a_2550_n632# a_3482_n632# 0.01fF
C2713 a_n3708_131# a_n3918_n197# 0.00fF
C2714 a_3480_n100# a_3432_131# 0.00fF
C2715 a_1802_n632# a_1290_n632# 0.01fF
C2716 a_238_n100# a_282_n197# 0.00fF
C2717 a_n3496_n729# a_n2446_n401# 0.00fF
C2718 a_450_n632# a_n928_n632# 0.00fF
C2719 a_4112_n632# w_n4520_n851# 0.14fF
C2720 a_n2026_n401# a_n2656_n729# 0.00fF
C2721 a_2968_n100# a_2850_n100# 0.07fF
C2722 a_n2912_n100# a_n1862_n100# 0.01fF
C2723 a_2548_n100# a_3808_n100# 0.00fF
C2724 a_2432_n632# a_3390_n632# 0.01fF
C2725 a_2220_n100# a_3598_n100# 0.00fF
C2726 a_n180_n632# a_1290_n632# 0.00fF
C2727 a_n3238_n632# a_n1860_n632# 0.00fF
C2728 a_n3496_n729# a_n3498_n197# 0.01fF
C2729 a_1382_n632# a_660_n632# 0.01fF
C2730 w_n4520_n851# a_n930_n100# 0.02fF
C2731 a_1754_n401# a_3224_n729# 0.00fF
C2732 a_n1862_n100# a_n2282_n100# 0.02fF
C2733 a_n392_n100# a_n182_n100# 0.03fF
C2734 a_3480_n100# w_n4520_n851# 0.04fF
C2735 a_n3332_n100# a_n2912_n100# 0.02fF
C2736 a_n602_n100# a_868_n100# 0.00fF
C2737 a_2760_n632# a_1290_n632# 0.00fF
C2738 w_n4520_n851# a_n3960_n632# 0.06fF
C2739 w_n4520_n851# a_n2028_131# 0.12fF
C2740 a_1920_n632# a_1962_n197# 0.00fF
C2741 a_n3332_n100# a_n2282_n100# 0.01fF
C2742 a_n136_n729# a_74_n401# 0.00fF
C2743 a_284_n729# a_332_n632# 0.00fF
C2744 a_1754_n401# a_704_n729# 0.00fF
C2745 a_3062_n632# a_2222_n632# 0.01fF
C2746 a_2382_n197# a_3432_131# 0.00fF
C2747 a_n346_n401# a_704_n729# 0.00fF
C2748 a_n2490_n632# a_n3028_n632# 0.01fF
C2749 a_2968_n100# a_4110_n100# 0.01fF
C2750 a_2850_n100# a_3178_n100# 0.02fF
C2751 a_n3030_n100# a_n1770_n100# 0.00fF
C2752 a_1754_n401# a_1800_n100# 0.00fF
C2753 a_2338_n100# a_1498_n100# 0.01fF
C2754 a_n510_n100# a_n1140_n100# 0.01fF
C2755 a_3062_n632# a_2642_n632# 0.02fF
C2756 a_n392_n100# a_n1442_n100# 0.01fF
C2757 a_n3240_n100# a_n3288_131# 0.00fF
C2758 a_n4080_n100# a_n4078_n632# 0.00fF
C2759 a_n1978_n632# a_n1230_n632# 0.01fF
C2760 a_2804_n729# a_1754_n401# 0.00fF
C2761 a_n1022_n100# a_n1140_n100# 0.07fF
C2762 a_n2190_n100# a_n1560_n100# 0.01fF
C2763 a_870_n632# a_n600_n632# 0.00fF
C2764 a_n928_n632# a_n298_n632# 0.01fF
C2765 a_n2490_n632# a_n1138_n632# 0.00fF
C2766 a_2758_n100# a_3270_n100# 0.01fF
C2767 a_n602_n100# a_540_n100# 0.01fF
C2768 a_2382_n197# w_n4520_n851# 0.10fF
C2769 a_1382_n632# a_122_n632# 0.00fF
C2770 a_2340_n632# w_n4520_n851# 0.01fF
C2771 a_n2398_n632# a_n3960_n632# 0.00fF
C2772 a_n2610_n100# a_n3962_n100# 0.00fF
C2773 a_1592_n632# a_1710_n632# 0.07fF
C2774 a_2970_n632# a_3180_n632# 0.03fF
C2775 a_n3330_n632# a_n3028_n632# 0.02fF
C2776 a_n2188_n632# a_n3028_n632# 0.01fF
C2777 a_n4078_n632# a_n3868_n632# 0.03fF
C2778 a_n3238_n632# a_n2910_n632# 0.02fF
C2779 a_n508_n632# a_n928_n632# 0.02fF
C2780 a_28_n100# a_868_n100# 0.01fF
C2781 a_n90_n100# a_1170_n100# 0.00fF
C2782 a_2968_n100# a_1590_n100# 0.00fF
C2783 a_2010_n100# a_1078_n100# 0.01fF
C2784 a_658_n100# a_2010_n100# 0.00fF
C2785 a_2760_n632# a_3902_n632# 0.01fF
C2786 a_n810_n632# a_n766_n401# 0.00fF
C2787 a_n720_n100# a_n1140_n100# 0.02fF
C2788 a_4110_n100# a_3178_n100# 0.01fF
C2789 a_n2070_n632# a_n3658_n632# 0.00fF
C2790 a_660_n632# a_n600_n632# 0.00fF
C2791 a_n2190_n100# a_n3450_n100# 0.00fF
C2792 a_n3238_n632# a_n2700_n632# 0.01fF
C2793 a_494_n401# a_1124_n729# 0.00fF
C2794 a_n2190_n100# a_n2702_n100# 0.01fF
C2795 a_30_n632# a_n1138_n632# 0.01fF
C2796 a_542_n632# a_1290_n632# 0.01fF
C2797 a_n1140_n100# a_n1980_n100# 0.01fF
C2798 a_n2188_n632# a_n1138_n632# 0.01fF
C2799 a_n3448_n632# a_n3750_n632# 0.02fF
C2800 a_n2608_n632# a_n1558_n632# 0.01fF
C2801 a_3900_n100# a_3270_n100# 0.01fF
C2802 a_n3496_n729# a_n4126_n401# 0.00fF
C2803 a_752_n632# a_2340_n632# 0.00fF
C2804 a_n812_n100# a_n182_n100# 0.01fF
C2805 a_n4170_n632# a_n3868_n632# 0.02fF
C2806 a_1172_n632# a_2340_n632# 0.01fF
C2807 a_2640_n100# a_3690_n100# 0.01fF
C2808 a_n2866_n401# a_n3076_n729# 0.00fF
C2809 a_1380_n100# a_2850_n100# 0.00fF
C2810 a_2172_131# a_2592_131# 0.01fF
C2811 a_n3448_n632# a_n2280_n632# 0.01fF
C2812 a_n88_n632# a_n1650_n632# 0.00fF
C2813 a_3388_n100# a_2548_n100# 0.01fF
C2814 a_n2608_n632# a_n3750_n632# 0.01fF
C2815 a_n3540_n632# a_n3028_n632# 0.01fF
C2816 a_3902_n632# a_3482_n632# 0.02fF
C2817 a_2592_131# a_3012_131# 0.01fF
C2818 a_3854_n401# a_3900_n100# 0.00fF
C2819 a_n2608_n632# a_n2280_n632# 0.02fF
C2820 a_n3122_n100# a_n1862_n100# 0.00fF
C2821 a_1500_n632# a_962_n632# 0.01fF
C2822 a_n810_n632# a_n1558_n632# 0.01fF
C2823 a_n348_131# a_282_n197# 0.00fF
C2824 a_870_n632# a_1920_n632# 0.01fF
C2825 a_n3240_n100# a_n1862_n100# 0.00fF
C2826 a_n1020_n632# a_n1440_n632# 0.02fF
C2827 a_n2820_n100# a_n2610_n100# 0.03fF
C2828 a_n3660_n100# w_n4520_n851# 0.04fF
C2829 a_28_n100# a_540_n100# 0.01fF
C2830 a_1590_n100# a_3178_n100# 0.00fF
C2831 a_n810_n632# a_n2280_n632# 0.00fF
C2832 a_n3332_n100# a_n3122_n100# 0.03fF
C2833 a_n1186_n401# a_n766_n401# 0.01fF
C2834 a_n1442_n100# a_n812_n100# 0.01fF
C2835 a_n2400_n100# a_n1232_n100# 0.01fF
C2836 a_n1650_n632# a_n1230_n632# 0.02fF
C2837 a_448_n100# a_n1140_n100# 0.00fF
C2838 a_n4080_n100# a_n3450_n100# 0.01fF
C2839 a_n1350_n100# a_n1862_n100# 0.01fF
C2840 a_1920_n632# a_3180_n632# 0.00fF
C2841 a_n4080_n100# a_n2702_n100# 0.00fF
C2842 a_n3332_n100# a_n3240_n100# 0.09fF
C2843 a_2010_n100# a_2758_n100# 0.01fF
C2844 a_n392_n100# a_330_n100# 0.01fF
C2845 a_2640_n100# a_1170_n100# 0.00fF
C2846 a_n2656_n729# a_n2658_n197# 0.01fF
C2847 a_n600_n632# a_122_n632# 0.01fF
C2848 a_2222_n632# a_1500_n632# 0.01fF
C2849 a_2222_n632# a_3272_n632# 0.01fF
C2850 a_660_n632# a_1920_n632# 0.00fF
C2851 a_n3752_n100# a_n3450_n100# 0.02fF
C2852 a_n2190_n100# a_n930_n100# 0.00fF
C2853 a_n2702_n100# a_n3752_n100# 0.01fF
C2854 a_870_n632# a_2012_n632# 0.01fF
C2855 a_1800_n100# a_1498_n100# 0.02fF
C2856 a_1918_n100# a_330_n100# 0.00fF
C2857 a_n2912_n100# a_n3962_n100# 0.01fF
C2858 a_n300_n100# a_120_n100# 0.02fF
C2859 a_2642_n632# a_1500_n632# 0.01fF
C2860 a_3600_n632# a_3642_n197# 0.00fF
C2861 a_2642_n632# a_3272_n632# 0.01fF
C2862 a_450_n632# a_n718_n632# 0.01fF
C2863 a_n2912_n100# a_n2868_131# 0.00fF
C2864 w_n4520_n851# a_868_n100# 0.02fF
C2865 a_2760_n632# a_4112_n632# 0.00fF
C2866 a_1918_n100# a_1962_n197# 0.00fF
C2867 a_n928_n632# w_n4520_n851# 0.01fF
C2868 a_n1140_n100# a_n1652_n100# 0.01fF
C2869 a_870_n632# a_240_n632# 0.01fF
C2870 a_2012_n632# a_3180_n632# 0.01fF
C2871 a_3062_n632# a_3810_n632# 0.01fF
C2872 a_2128_n100# a_1498_n100# 0.01fF
C2873 a_238_n100# a_n930_n100# 0.01fF
C2874 a_n976_n729# w_n4520_n851# 0.12fF
C2875 a_1288_n100# a_28_n100# 0.00fF
C2876 a_n602_n100# a_n182_n100# 0.02fF
C2877 a_3480_n100# a_2548_n100# 0.01fF
C2878 a_n298_n632# a_n1768_n632# 0.00fF
C2879 a_660_n632# a_2012_n632# 0.00fF
C2880 a_4112_n632# a_3482_n632# 0.01fF
C2881 a_n88_n632# a_n136_n729# 0.00fF
C2882 w_n4520_n851# a_3060_n100# 0.03fF
C2883 w_n4520_n851# a_n2236_n729# 0.12fF
C2884 a_914_n401# a_2384_n729# 0.00fF
C2885 a_1380_n100# a_1590_n100# 0.03fF
C2886 a_494_n401# a_n766_n401# 0.00fF
C2887 a_n3330_n632# a_n2490_n632# 0.01fF
C2888 a_n2490_n632# a_n2188_n632# 0.02fF
C2889 w_n4520_n851# a_1334_n401# 0.10fF
C2890 a_750_n100# a_868_n100# 0.07fF
C2891 a_1332_131# a_282_n197# 0.00fF
C2892 a_448_n100# a_1590_n100# 0.01fF
C2893 a_2852_n632# a_1382_n632# 0.00fF
C2894 a_3062_n632# a_2550_n632# 0.01fF
C2895 a_960_n100# a_1498_n100# 0.01fF
C2896 a_1592_n632# a_1080_n632# 0.01fF
C2897 a_240_n632# a_660_n632# 0.02fF
C2898 a_n3078_n197# a_n2028_131# 0.00fF
C2899 a_n2028_131# a_n2448_131# 0.01fF
C2900 a_n2820_n100# a_n2912_n100# 0.09fF
C2901 a_2338_n100# a_1078_n100# 0.00fF
C2902 a_3480_n100# a_3482_n632# 0.00fF
C2903 a_n508_n632# a_n1768_n632# 0.00fF
C2904 w_n4520_n851# a_540_n100# 0.02fF
C2905 a_2220_n100# a_1708_n100# 0.01fF
C2906 a_2850_n100# a_2430_n100# 0.02fF
C2907 a_3644_n729# a_2594_n401# 0.00fF
C2908 a_1802_n632# a_2340_n632# 0.01fF
C2909 a_2802_n197# a_2850_n100# 0.00fF
C2910 a_n2398_n632# a_n928_n632# 0.00fF
C2911 a_332_n632# a_1592_n632# 0.00fF
C2912 a_n602_n100# a_n1442_n100# 0.01fF
C2913 a_n1440_n632# a_n1398_n197# 0.00fF
C2914 a_1542_n197# a_492_131# 0.00fF
C2915 a_n2820_n100# a_n2282_n100# 0.01fF
C2916 a_n2818_n632# w_n4520_n851# 0.02fF
C2917 a_n3120_n632# w_n4520_n851# 0.03fF
C2918 a_n3540_n632# a_n2490_n632# 0.01fF
C2919 a_n718_n632# a_n298_n632# 0.02fF
C2920 a_n300_n100# a_1078_n100# 0.00fF
C2921 a_1290_n632# a_1332_131# 0.00fF
C2922 a_n300_n100# a_658_n100# 0.01fF
C2923 a_2968_n100# a_3178_n100# 0.03fF
C2924 a_n812_n100# a_330_n100# 0.01fF
C2925 a_n3330_n632# a_n2188_n632# 0.01fF
C2926 a_n1606_n401# a_n766_n401# 0.01fF
C2927 a_n2072_n100# a_n1232_n100# 0.01fF
C2928 a_n510_n100# a_n1022_n100# 0.01fF
C2929 a_n3960_n632# a_n3868_n632# 0.09fF
C2930 a_n602_n100# a_n558_n197# 0.00fF
C2931 a_2760_n632# a_2340_n632# 0.02fF
C2932 a_750_n100# a_540_n100# 0.03fF
C2933 a_n2400_n100# a_n2492_n100# 0.09fF
C2934 a_n88_n632# a_962_n632# 0.01fF
C2935 a_28_n100# a_n182_n100# 0.03fF
C2936 a_3224_n729# a_3434_n401# 0.00fF
C2937 a_n810_n632# a_332_n632# 0.01fF
C2938 a_n1770_n100# a_n1862_n100# 0.09fF
C2939 a_n718_n632# a_n508_n632# 0.03fF
C2940 a_n1396_n729# a_n1186_n401# 0.00fF
C2941 a_3224_n729# a_3272_n632# 0.00fF
C2942 a_n3240_n100# a_n3286_n401# 0.00fF
C2943 a_n300_n100# a_n1350_n100# 0.01fF
C2944 a_n3540_n632# a_n3330_n632# 0.03fF
C2945 a_n3540_n632# a_n2188_n632# 0.00fF
C2946 a_1918_n100# a_1708_n100# 0.03fF
C2947 a_704_n729# a_74_n401# 0.00fF
C2948 a_1288_n100# w_n4520_n851# 0.02fF
C2949 a_n1606_n401# a_n1558_n632# 0.00fF
C2950 a_240_n632# a_122_n632# 0.07fF
C2951 a_2340_n632# a_3482_n632# 0.01fF
C2952 a_n3028_n632# a_n1558_n632# 0.00fF
C2953 a_n3496_n729# a_n2866_n401# 0.00fF
C2954 a_2338_n100# a_2758_n100# 0.02fF
C2955 a_n3332_n100# a_n1770_n100# 0.00fF
C2956 a_n2190_n100# a_n3660_n100# 0.00fF
C2957 a_n1560_n100# a_n2610_n100# 0.01fF
C2958 a_n138_n197# a_n1608_131# 0.00fF
C2959 a_n2398_n632# a_n2818_n632# 0.02fF
C2960 a_n3120_n632# a_n2398_n632# 0.01fF
C2961 a_n720_n100# a_n510_n100# 0.03fF
C2962 a_n3750_n632# a_n3028_n632# 0.01fF
C2963 a_n3122_n100# a_n3962_n100# 0.01fF
C2964 a_n1860_n632# a_n298_n632# 0.00fF
C2965 a_1964_n729# a_1920_n632# 0.00fF
C2966 a_n2070_n632# a_n1348_n632# 0.01fF
C2967 a_2970_n632# a_2852_n632# 0.07fF
C2968 a_n510_n100# a_n1980_n100# 0.00fF
C2969 a_n720_n100# a_n1022_n100# 0.02fF
C2970 a_n2280_n632# a_n3028_n632# 0.01fF
C2971 a_n3240_n100# a_n3962_n100# 0.01fF
C2972 a_n136_n729# a_284_n729# 0.01fF
C2973 a_n1138_n632# a_n1558_n632# 0.02fF
C2974 a_n1442_n100# a_28_n100# 0.00fF
C2975 a_n1020_n632# a_n600_n632# 0.02fF
C2976 a_3272_n632# a_3810_n632# 0.01fF
C2977 a_n1022_n100# a_n1980_n100# 0.01fF
C2978 a_2968_n100# a_1380_n100# 0.00fF
C2979 a_n88_n632# a_n390_n632# 0.02fF
C2980 a_2804_n729# a_3434_n401# 0.00fF
C2981 a_n1230_n632# a_n1188_131# 0.00fF
C2982 a_n3540_n632# a_n3542_n100# 0.00fF
C2983 a_120_n100# a_960_n100# 0.01fF
C2984 w_n4520_n851# a_n1768_n632# 0.01fF
C2985 a_1288_n100# a_750_n100# 0.01fF
C2986 a_n1818_n197# a_n3288_131# 0.00fF
C2987 a_1590_n100# a_2430_n100# 0.01fF
C2988 a_n1860_n632# a_n508_n632# 0.00fF
C2989 a_n3448_n632# a_n1978_n632# 0.00fF
C2990 a_2338_n100# a_3900_n100# 0.00fF
C2991 a_n2280_n632# a_n1138_n632# 0.01fF
C2992 w_n4520_n851# a_1752_131# 0.12fF
C2993 a_n2610_n100# a_n3450_n100# 0.01fF
C2994 a_n1818_n197# a_n2658_n197# 0.01fF
C2995 a_n2702_n100# a_n2610_n100# 0.09fF
C2996 a_n1978_n632# a_n2608_n632# 0.01fF
C2997 a_912_131# a_702_n197# 0.00fF
C2998 a_n3542_n100# a_n1980_n100# 0.00fF
C2999 a_n602_n100# a_330_n100# 0.01fF
C3000 a_2012_n632# a_1964_n729# 0.00fF
C3001 a_2550_n632# a_3272_n632# 0.01fF
C3002 a_2550_n632# a_1500_n632# 0.01fF
C3003 w_n4520_n851# a_1122_n197# 0.10fF
C3004 a_n4080_n100# a_n3660_n100# 0.02fF
C3005 a_1800_n100# a_1078_n100# 0.01fF
C3006 a_658_n100# a_1800_n100# 0.01fF
C3007 a_n720_n100# a_n1980_n100# 0.00fF
C3008 a_n390_n632# a_n1230_n632# 0.01fF
C3009 a_4018_n100# a_2758_n100# 0.00fF
C3010 a_n510_n100# a_448_n100# 0.01fF
C3011 a_3902_n632# a_3062_n632# 0.01fF
C3012 a_n558_n197# a_n1608_131# 0.00fF
C3013 a_2432_n632# a_1710_n632# 0.01fF
C3014 a_n2820_n100# a_n3122_n100# 0.02fF
C3015 a_n556_n729# a_n976_n729# 0.01fF
C3016 w_n4520_n851# a_n182_n100# 0.02fF
C3017 a_n1978_n632# a_n810_n632# 0.01fF
C3018 a_n180_n632# a_n928_n632# 0.01fF
C3019 a_n3660_n100# a_n3752_n100# 0.09fF
C3020 a_448_n100# a_n1022_n100# 0.00fF
C3021 a_n2820_n100# a_n3240_n100# 0.02fF
C3022 a_n2190_n100# a_n2236_n729# 0.00fF
C3023 a_238_n100# a_868_n100# 0.01fF
C3024 a_n2446_n401# w_n4520_n851# 0.10fF
C3025 a_n138_n197# w_n4520_n851# 0.10fF
C3026 a_n718_n632# w_n4520_n851# 0.01fF
C3027 a_2432_n632# a_2430_n100# 0.00fF
C3028 a_n392_n100# a_n1232_n100# 0.01fF
C3029 a_2128_n100# a_1078_n100# 0.01fF
C3030 a_658_n100# a_2128_n100# 0.00fF
C3031 a_2852_n632# a_1920_n632# 0.01fF
C3032 a_n2398_n632# a_n1768_n632# 0.01fF
C3033 a_3644_n729# a_3690_n100# 0.00fF
C3034 a_n2656_n729# a_n3286_n401# 0.00fF
C3035 a_n2072_n100# a_n2492_n100# 0.02fF
C3036 a_n2026_n401# a_n1186_n401# 0.01fF
C3037 a_n2820_n100# a_n1350_n100# 0.00fF
C3038 a_n1440_n632# a_n600_n632# 0.01fF
C3039 w_n4520_n851# a_n3498_n197# 0.11fF
C3040 a_n1560_n100# a_n2912_n100# 0.00fF
C3041 a_n1396_n729# a_n1606_n401# 0.00fF
C3042 a_n510_n100# a_n1652_n100# 0.01fF
C3043 a_3060_n100# a_2548_n100# 0.01fF
C3044 a_3598_n100# w_n4520_n851# 0.04fF
C3045 a_4018_n100# a_3900_n100# 0.07fF
C3046 a_750_n100# a_n182_n100# 0.01fF
C3047 a_752_n632# a_n718_n632# 0.00fF
C3048 a_n720_n100# a_448_n100# 0.01fF
C3049 a_960_n100# a_1078_n100# 0.07fF
C3050 w_n4520_n851# a_n1442_n100# 0.02fF
C3051 a_658_n100# a_960_n100# 0.02fF
C3052 a_n1022_n100# a_n1652_n100# 0.01fF
C3053 a_1500_n632# a_1290_n632# 0.03fF
C3054 a_n300_n100# a_n1770_n100# 0.00fF
C3055 w_n4520_n851# a_2130_n632# 0.01fF
C3056 a_n1818_n197# a_n1862_n100# 0.00fF
C3057 a_n1560_n100# a_n2282_n100# 0.01fF
C3058 a_n4128_131# w_n4520_n851# 0.14fF
C3059 a_2222_n632# a_3692_n632# 0.00fF
C3060 a_n1348_n632# a_n1350_n100# 0.00fF
C3061 a_28_n100# a_330_n100# 0.02fF
C3062 a_1800_n100# a_2758_n100# 0.01fF
C3063 a_n1818_n197# a_n768_131# 0.00fF
C3064 a_2852_n632# a_2012_n632# 0.01fF
C3065 a_n1816_n729# w_n4520_n851# 0.12fF
C3066 a_2642_n632# a_3692_n632# 0.01fF
C3067 a_1124_n729# a_2174_n401# 0.00fF
C3068 a_2220_n100# a_3690_n100# 0.00fF
C3069 a_870_n632# a_450_n632# 0.02fF
C3070 a_238_n100# a_540_n100# 0.02fF
C3071 a_n2490_n632# a_n1558_n632# 0.01fF
C3072 a_n2398_n632# a_n2446_n401# 0.00fF
C3073 a_n2912_n100# a_n3450_n100# 0.01fF
C3074 a_n1860_n632# w_n4520_n851# 0.01fF
C3075 a_n2912_n100# a_n2702_n100# 0.03fF
C3076 a_n558_n197# w_n4520_n851# 0.10fF
C3077 a_n3658_n632# a_n3706_n401# 0.00fF
C3078 a_n2490_n632# a_n3750_n632# 0.00fF
C3079 a_n2608_n632# a_n1650_n632# 0.01fF
C3080 a_752_n632# a_2130_n632# 0.00fF
C3081 a_1172_n632# a_2130_n632# 0.01fF
C3082 a_2968_n100# a_2430_n100# 0.01fF
C3083 a_n720_n100# a_n1652_n100# 0.01fF
C3084 a_n136_n729# a_914_n401# 0.00fF
C3085 a_1544_n729# w_n4520_n851# 0.12fF
C3086 a_2128_n100# a_2758_n100# 0.01fF
C3087 a_n2490_n632# a_n2280_n632# 0.03fF
C3088 a_n3120_n632# a_n3078_n197# 0.00fF
C3089 a_n2282_n100# a_n3450_n100# 0.01fF
C3090 a_4112_n632# a_3062_n632# 0.01fF
C3091 a_n1020_n632# a_240_n632# 0.00fF
C3092 a_n1980_n100# a_n1652_n100# 0.02fF
C3093 a_n2702_n100# a_n2282_n100# 0.02fF
C3094 a_448_n100# a_1380_n100# 0.01fF
C3095 a_450_n632# a_660_n632# 0.03fF
C3096 a_n810_n632# a_n1650_n632# 0.01fF
C3097 a_332_n632# a_n1138_n632# 0.00fF
C3098 a_30_n632# a_n1558_n632# 0.00fF
C3099 a_542_n632# a_n928_n632# 0.00fF
C3100 a_n2188_n632# a_n1558_n632# 0.01fF
C3101 a_n1818_n197# a_n1188_131# 0.00fF
C3102 a_n3708_131# a_n2238_n197# 0.00fF
C3103 a_2220_n100# a_1170_n100# 0.01fF
C3104 a_n1232_n100# a_n812_n100# 0.02fF
C3105 a_1288_n100# a_2548_n100# 0.00fF
C3106 a_n3330_n632# a_n3750_n632# 0.02fF
C3107 a_n2188_n632# a_n3750_n632# 0.00fF
C3108 a_n720_n100# a_n766_n401# 0.00fF
C3109 a_2970_n632# a_1382_n632# 0.00fF
C3110 a_1288_n100# a_238_n100# 0.01fF
C3111 a_n3330_n632# a_n2280_n632# 0.01fF
C3112 a_n1860_n632# a_n2398_n632# 0.01fF
C3113 a_3902_n632# a_3272_n632# 0.01fF
C3114 a_n2280_n632# a_n2188_n632# 0.09fF
C3115 a_n2818_n632# a_n3868_n632# 0.01fF
C3116 a_n3120_n632# a_n3868_n632# 0.01fF
C3117 w_n4520_n851# a_n4126_n401# 0.12fF
C3118 a_1962_n197# a_3432_131# 0.00fF
C3119 a_2758_n100# a_3808_n100# 0.01fF
C3120 a_72_131# a_1122_n197# 0.00fF
C3121 a_2430_n100# a_3178_n100# 0.01fF
C3122 a_4110_n100# a_4064_n729# 0.00fF
C3123 a_n1348_n632# a_n88_n632# 0.00fF
C3124 a_870_n632# a_n298_n632# 0.01fF
C3125 a_n2026_n401# a_n1606_n401# 0.01fF
C3126 a_4020_n632# a_3180_n632# 0.01fF
C3127 a_2382_n197# a_1332_131# 0.00fF
C3128 a_2432_n632# a_1080_n632# 0.00fF
C3129 a_n976_n729# a_n346_n401# 0.00fF
C3130 a_914_n401# a_962_n632# 0.00fF
C3131 a_n180_n632# a_n1768_n632# 0.00fF
C3132 w_n4520_n851# a_330_n100# 0.02fF
C3133 a_542_n632# a_540_n100# 0.00fF
C3134 a_n2820_n100# a_n1770_n100# 0.01fF
C3135 a_n3540_n632# a_n3750_n632# 0.03fF
C3136 a_n392_n100# a_1170_n100# 0.00fF
C3137 a_n2910_n632# w_n4520_n851# 0.03fF
C3138 a_n3030_n100# a_n3028_n632# 0.00fF
C3139 a_n138_n197# a_72_131# 0.00fF
C3140 a_n930_n100# a_n2282_n100# 0.00fF
C3141 a_n3540_n632# a_n2280_n632# 0.00fF
C3142 w_n4520_n851# a_1962_n197# 0.10fF
C3143 a_n2700_n632# w_n4520_n851# 0.02fF
C3144 a_870_n632# a_n508_n632# 0.00fF
C3145 a_450_n632# a_122_n632# 0.02fF
C3146 a_n1560_n100# a_n3122_n100# 0.00fF
C3147 a_1754_n401# a_1334_n401# 0.01fF
C3148 a_1918_n100# a_1170_n100# 0.01fF
C3149 a_n1348_n632# a_n1230_n632# 0.07fF
C3150 a_3900_n100# a_3808_n100# 0.09fF
C3151 a_n1818_n197# a_n978_n197# 0.01fF
C3152 a_660_n632# a_n298_n632# 0.01fF
C3153 a_n1978_n632# a_n3028_n632# 0.01fF
C3154 a_3062_n632# a_2340_n632# 0.01fF
C3155 a_n3706_n401# a_n3286_n401# 0.01fF
C3156 a_n3660_n100# a_n2610_n100# 0.01fF
C3157 a_n2238_n197# a_n1398_n197# 0.01fF
C3158 a_n180_n632# a_n182_n100# 0.00fF
C3159 a_120_n100# a_n930_n100# 0.01fF
C3160 a_750_n100# a_330_n100# 0.02fF
C3161 w_n4520_n851# a_n4172_n100# 0.14fF
C3162 a_n88_n632# a_1290_n632# 0.00fF
C3163 a_1382_n632# a_1920_n632# 0.01fF
C3164 a_n1560_n100# a_n1350_n100# 0.03fF
C3165 a_n180_n632# a_n138_n197# 0.00fF
C3166 a_n1978_n632# a_n1138_n632# 0.01fF
C3167 a_n180_n632# a_n718_n632# 0.01fF
C3168 a_238_n100# a_n182_n100# 0.02fF
C3169 a_n508_n632# a_660_n632# 0.01fF
C3170 a_2850_n100# a_3270_n100# 0.02fF
C3171 a_1380_n100# a_2430_n100# 0.01fF
C3172 a_n3122_n100# a_n3450_n100# 0.02fF
C3173 a_n392_n100# a_n90_n100# 0.02fF
C3174 a_n3122_n100# a_n2702_n100# 0.02fF
C3175 a_n2190_n100# a_n1442_n100# 0.01fF
C3176 a_n602_n100# a_n1232_n100# 0.01fF
C3177 a_2432_n632# a_2384_n729# 0.00fF
C3178 a_1802_n632# a_2130_n632# 0.02fF
C3179 a_3692_n632# a_3810_n632# 0.07fF
C3180 a_n2398_n632# a_n2910_n632# 0.01fF
C3181 a_n2446_n401# a_n2448_131# 0.01fF
C3182 a_n3240_n100# a_n3450_n100# 0.03fF
C3183 a_n2070_n632# a_n2028_131# 0.00fF
C3184 a_284_n729# a_704_n729# 0.01fF
C3185 a_4112_n632# a_3272_n632# 0.01fF
C3186 a_n3240_n100# a_n2702_n100# 0.01fF
C3187 a_n558_n197# a_72_131# 0.00fF
C3188 a_n2398_n632# a_n2700_n632# 0.02fF
C3189 a_n556_n729# a_n1816_n729# 0.00fF
C3190 a_3598_n100# a_2548_n100# 0.01fF
C3191 a_962_n632# a_1592_n632# 0.01fF
C3192 a_3480_n100# a_3434_n401# 0.00fF
C3193 a_n810_n632# a_n768_131# 0.00fF
C3194 a_n3498_n197# a_n3078_n197# 0.01fF
C3195 a_2220_n100# a_2640_n100# 0.02fF
C3196 a_n3498_n197# a_n2448_131# 0.00fF
C3197 a_1382_n632# a_2012_n632# 0.01fF
C3198 a_30_n632# a_1080_n632# 0.01fF
C3199 a_n1818_n197# a_n2868_131# 0.00fF
C3200 a_n1350_n100# a_n2702_n100# 0.00fF
C3201 a_n556_n729# a_n558_n197# 0.01fF
C3202 a_2550_n632# a_3692_n632# 0.01fF
C3203 a_n3448_n632# a_n3658_n632# 0.03fF
C3204 a_n298_n632# a_122_n632# 0.02fF
C3205 a_2760_n632# a_2130_n632# 0.01fF
C3206 a_n136_n729# a_n1186_n401# 0.00fF
C3207 a_n3658_n632# a_n2608_n632# 0.01fF
C3208 a_n4128_131# a_n3078_n197# 0.00fF
C3209 a_30_n632# a_332_n632# 0.02fF
C3210 a_3388_n100# a_2758_n100# 0.01fF
C3211 a_240_n632# a_1382_n632# 0.01fF
C3212 a_4110_n100# a_3270_n100# 0.01fF
C3213 a_1498_n100# a_868_n100# 0.01fF
C3214 a_870_n632# w_n4520_n851# 0.01fF
C3215 a_n1650_n632# a_n1606_n401# 0.00fF
C3216 a_3902_n632# a_3900_n100# 0.00fF
C3217 a_n4128_131# a_n4080_n100# 0.00fF
C3218 a_2130_n632# a_3482_n632# 0.00fF
C3219 a_n508_n632# a_122_n632# 0.01fF
C3220 a_658_n100# a_n930_n100# 0.00fF
C3221 a_2222_n632# a_1592_n632# 0.01fF
C3222 w_n4520_n851# a_1708_n100# 0.02fF
C3223 a_n1650_n632# a_n3028_n632# 0.00fF
C3224 a_n2912_n100# a_n3660_n100# 0.01fF
C3225 a_284_n729# a_282_n197# 0.01fF
C3226 a_2550_n632# a_2592_131# 0.00fF
C3227 a_2642_n632# a_1592_n632# 0.01fF
C3228 a_n1232_n100# a_28_n100# 0.00fF
C3229 a_2968_n100# a_3012_131# 0.00fF
C3230 a_2970_n632# a_1920_n632# 0.01fF
C3231 w_n4520_n851# a_3180_n632# 0.03fF
C3232 a_1754_n401# a_1752_131# 0.01fF
C3233 a_3060_n100# a_1498_n100# 0.00fF
C3234 a_1334_n401# a_1332_131# 0.01fF
C3235 a_1918_n100# a_2640_n100# 0.01fF
C3236 a_n3660_n100# a_n2282_n100# 0.00fF
C3237 a_n1650_n632# a_n1138_n632# 0.01fF
C3238 a_n2072_n100# a_n2400_n100# 0.02fF
C3239 a_870_n632# a_752_n632# 0.07fF
C3240 a_3388_n100# a_3900_n100# 0.01fF
C3241 a_542_n632# a_n718_n632# 0.00fF
C3242 a_870_n632# a_1172_n632# 0.02fF
C3243 a_2010_n100# a_2850_n100# 0.01fF
C3244 a_660_n632# w_n4520_n851# 0.01fF
C3245 a_n90_n100# a_n812_n100# 0.01fF
C3246 a_2340_n632# a_3272_n632# 0.01fF
C3247 a_2340_n632# a_1500_n632# 0.01fF
C3248 a_n1350_n100# a_n930_n100# 0.02fF
C3249 a_1124_n729# a_1080_n632# 0.00fF
C3250 a_n1978_n632# a_n2490_n632# 0.01fF
C3251 a_750_n100# a_1708_n100# 0.01fF
C3252 a_3014_n401# a_2174_n401# 0.01fF
C3253 a_n390_n632# a_n810_n632# 0.02fF
C3254 w_n4520_n851# a_2594_n401# 0.10fF
C3255 a_3062_n632# a_3060_n100# 0.00fF
C3256 a_1498_n100# a_540_n100# 0.01fF
C3257 a_2172_131# a_702_n197# 0.00fF
C3258 a_494_n401# a_n136_n729# 0.00fF
C3259 a_n1560_n100# a_n1770_n100# 0.03fF
C3260 w_n4520_n851# a_n2866_n401# 0.10fF
C3261 a_450_n632# a_n1020_n632# 0.00fF
C3262 a_2970_n632# a_2012_n632# 0.01fF
C3263 a_2802_n197# a_3642_n197# 0.01fF
C3264 w_n4520_n851# VSUBS 31.73fF
.ends

.subckt latch_pmos_pair sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n632#
+ VSUBS sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
Xsky130_fd_pr__pfet_01v8_VCQUSW_0 sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1802_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4080_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2640_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2010_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3852_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3750_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3120_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3600_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2594_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n88_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2866_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2912_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n718_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n556_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2548_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n182_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3658_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3028_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3496_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2012_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2642_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1140_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1770_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1398_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2172_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n812_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4128_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3224_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n766_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3480_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3122_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3752_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_240_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_870_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2448_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3388_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3434_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3706_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3482_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_492_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1500_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4064_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1650_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n768_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2238_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1558_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2610_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1396_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_750_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_120_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1124_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2490_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2340_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2970_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1380_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_658_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n510_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1022_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1652_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n138_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1288_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3450_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3078_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2398_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_122_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_752_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1334_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_74_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_702_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1382_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1606_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1962_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3012_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1918_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_28_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2492_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1332_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2236_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n298_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3810_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2850_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2220_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3960_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3330_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2174_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1608_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n928_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2446_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n136_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3868_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3238_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2758_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2128_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n392_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3076_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2802_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2222_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2852_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1350_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1980_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4170_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4020_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n346_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3690_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3060_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3332_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3962_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2592_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_450_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3286_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3598_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4078_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1080_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3014_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2868_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3062_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3692_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2190_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3642_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1860_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1230_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1710_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4172_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2820_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1768_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1138_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1188_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_704_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n4126_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_960_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_330_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1964_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1590_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_282_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2070_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2550_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n90_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n978_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1186_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_868_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_238_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n720_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1232_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1862_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_914_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1498_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3030_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3660_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2700_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_332_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_962_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1542_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1592_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3918_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2608_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3390_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2072_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3432_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n600_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1752_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2804_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3540_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2430_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2702_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3708_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n508_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2026_n401#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2382_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2968_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2338_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n976_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3448_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1560_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2432_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3644_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3270_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n602_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2028_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3916_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3542_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_660_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1818_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3178_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1290_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3900_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3854_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3222_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3272_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n348_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_30_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3808_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1440_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1920_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_284_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2658_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_3902_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2400_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1978_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1348_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3288_131# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4110_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_494_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_540_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4062_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4018_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1544_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2280_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2130_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2760_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1170_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_72_131#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n300_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n930_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1442_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n558_n197#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n1816_n729# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_448_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3240_n100# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3870_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n3498_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2188_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_4112_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1078_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1754_n401# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1800_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2910_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_542_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1122_n197# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n180_n632#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1172_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_2384_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2818_n632# sky130_fd_pr__pfet_01v8_VCQUSW_0/a_1708_n100#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_912_131# VSUBS sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2656_n729#
+ sky130_fd_pr__pfet_01v8_VCQUSW_0/a_n2282_n100# sky130_fd_pr__pfet_01v8_VCQUSW
C0 sky130_fd_pr__pfet_01v8_VCQUSW_0/w_n4520_n851# VSUBS 31.73fF
.ends

.subckt sky130_fd_pr__pfet_01v8_VCG74W a_543_n100# a_159_n100# a_n609_n100# a_495_n197#
+ a_n705_n100# a_255_n100# a_n657_n197# a_n369_131# a_351_n100# a_n417_n100# a_n801_n100#
+ a_303_n197# a_n129_n100# a_n513_n100# a_n465_n197# a_n561_131# a_63_n100# a_n225_n100#
+ a_399_131# a_111_n197# a_n321_n100# a_n273_n197# a_15_131# a_n753_131# a_639_n100#
+ w_n1031_n319# a_591_131# a_207_131# a_735_n100# a_n33_n100# a_687_n197# a_447_n100#
+ a_n81_n197# a_n177_131# VSUBS
X0 a_63_n100# a_15_131# a_n33_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n197# a_n129_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_255_n100# a_207_131# a_159_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_351_n100# a_303_n197# a_255_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_543_n100# a_495_n197# a_447_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 w_n1031_n319# w_n1031_n319# a_735_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=6.2e+11p pd=5.24e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_159_n100# a_111_n197# a_63_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_447_n100# a_399_131# a_351_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_639_n100# a_591_131# a_543_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_735_n100# a_687_n197# a_639_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n801_n100# w_n1031_n319# w_n1031_n319# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_n513_n100# a_n561_131# a_n609_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_n321_n100# a_n369_131# a_n417_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_n225_n100# a_n273_n197# a_n321_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_n705_n100# a_n753_131# a_n801_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_n609_n100# a_n657_n197# a_n705_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n417_n100# a_n465_n197# a_n513_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n129_n100# a_n177_131# a_n225_n100# w_n1031_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n513_n100# a_63_n100# 0.01fF
C1 a_n417_n100# a_n33_n100# 0.02fF
C2 a_n417_n100# a_639_n100# 0.01fF
C3 a_735_n100# a_447_n100# 0.02fF
C4 a_n657_n197# a_207_131# 0.00fF
C5 a_207_131# a_n753_131# 0.01fF
C6 a_591_131# a_15_131# 0.01fF
C7 a_735_n100# a_63_n100# 0.01fF
C8 a_n177_131# a_n225_n100# 0.00fF
C9 a_447_n100# a_63_n100# 0.02fF
C10 a_207_131# w_n1031_n319# 0.12fF
C11 a_495_n197# a_303_n197# 0.04fF
C12 a_111_n197# a_n561_131# 0.00fF
C13 a_399_131# a_n273_n197# 0.00fF
C14 a_n321_n100# a_255_n100# 0.01fF
C15 a_111_n197# a_63_n100# 0.00fF
C16 a_351_n100# a_n33_n100# 0.02fF
C17 a_255_n100# a_n225_n100# 0.01fF
C18 a_351_n100# a_639_n100# 0.02fF
C19 a_n33_n100# w_n1031_n319# 0.04fF
C20 a_639_n100# w_n1031_n319# 0.08fF
C21 a_n81_n197# a_399_131# 0.00fF
C22 a_n417_n100# a_n801_n100# 0.02fF
C23 a_207_131# a_687_n197# 0.00fF
C24 a_255_n100# a_n609_n100# 0.01fF
C25 a_255_n100# a_n513_n100# 0.01fF
C26 a_303_n197# a_n465_n197# 0.01fF
C27 a_n561_131# a_n177_131# 0.01fF
C28 a_n273_n197# a_15_131# 0.00fF
C29 a_639_n100# a_687_n197# 0.00fF
C30 a_111_n197# a_n177_131# 0.00fF
C31 a_n801_n100# a_n753_131# 0.00fF
C32 a_735_n100# a_255_n100# 0.01fF
C33 a_159_n100# a_543_n100# 0.02fF
C34 a_n81_n197# a_15_131# 0.01fF
C35 a_255_n100# a_447_n100# 0.04fF
C36 a_n705_n100# a_543_n100# 0.00fF
C37 a_351_n100# a_n801_n100# 0.01fF
C38 a_n801_n100# w_n1031_n319# 0.15fF
C39 a_n273_n197# a_591_131# 0.00fF
C40 a_255_n100# a_63_n100# 0.04fF
C41 a_n81_n197# a_591_131# 0.00fF
C42 a_543_n100# a_591_131# 0.00fF
C43 a_n129_n100# a_n33_n100# 0.09fF
C44 a_n129_n100# a_639_n100# 0.01fF
C45 a_495_n197# a_447_n100# 0.00fF
C46 a_n369_131# a_207_131# 0.01fF
C47 a_495_n197# a_n561_131# 0.00fF
C48 a_n513_n100# a_n465_n197# 0.00fF
C49 a_495_n197# a_111_n197# 0.01fF
C50 a_n657_n197# a_399_131# 0.00fF
C51 a_399_131# a_n753_131# 0.00fF
C52 a_n417_n100# a_159_n100# 0.01fF
C53 a_n417_n100# a_n705_n100# 0.02fF
C54 a_351_n100# a_399_131# 0.00fF
C55 a_399_131# w_n1031_n319# 0.12fF
C56 a_n561_131# a_n465_n197# 0.01fF
C57 a_n81_n197# a_n273_n197# 0.04fF
C58 a_111_n197# a_n465_n197# 0.01fF
C59 a_n801_n100# a_n129_n100# 0.01fF
C60 a_495_n197# a_n177_131# 0.00fF
C61 a_n657_n197# a_15_131# 0.00fF
C62 a_15_131# a_n753_131# 0.01fF
C63 a_n705_n100# a_n657_n197# 0.00fF
C64 a_n705_n100# a_n753_131# 0.00fF
C65 a_399_131# a_687_n197# 0.00fF
C66 a_159_n100# a_351_n100# 0.04fF
C67 a_159_n100# w_n1031_n319# 0.04fF
C68 a_n705_n100# a_351_n100# 0.01fF
C69 a_15_131# w_n1031_n319# 0.12fF
C70 a_n705_n100# w_n1031_n319# 0.08fF
C71 a_n657_n197# a_591_131# 0.00fF
C72 a_591_131# a_n753_131# 0.00fF
C73 a_n177_131# a_n465_n197# 0.00fF
C74 a_303_n197# a_207_131# 0.01fF
C75 a_591_131# w_n1031_n319# 0.12fF
C76 a_15_131# a_687_n197# 0.00fF
C77 a_591_131# a_687_n197# 0.01fF
C78 a_n417_n100# a_543_n100# 0.01fF
C79 a_399_131# a_n369_131# 0.01fF
C80 a_n657_n197# a_n273_n197# 0.01fF
C81 a_n273_n197# a_n753_131# 0.00fF
C82 a_495_n197# a_n465_n197# 0.01fF
C83 a_159_n100# a_n129_n100# 0.02fF
C84 a_n705_n100# a_n129_n100# 0.01fF
C85 a_n657_n197# a_n81_n197# 0.01fF
C86 a_n81_n197# a_n753_131# 0.00fF
C87 a_n321_n100# a_n33_n100# 0.02fF
C88 a_n321_n100# a_639_n100# 0.01fF
C89 a_n273_n197# w_n1031_n319# 0.13fF
C90 a_n33_n100# a_n225_n100# 0.04fF
C91 a_639_n100# a_n225_n100# 0.01fF
C92 a_n81_n197# w_n1031_n319# 0.13fF
C93 a_543_n100# a_351_n100# 0.04fF
C94 a_543_n100# w_n1031_n319# 0.06fF
C95 a_n369_131# a_15_131# 0.01fF
C96 a_n609_n100# a_n33_n100# 0.01fF
C97 a_n513_n100# a_n33_n100# 0.01fF
C98 a_639_n100# a_n609_n100# 0.00fF
C99 a_n513_n100# a_639_n100# 0.01fF
C100 a_n273_n197# a_687_n197# 0.01fF
C101 a_n561_131# a_207_131# 0.01fF
C102 a_735_n100# a_n33_n100# 0.01fF
C103 a_n81_n197# a_687_n197# 0.01fF
C104 a_735_n100# a_639_n100# 0.09fF
C105 a_n369_131# a_591_131# 0.01fF
C106 a_111_n197# a_207_131# 0.01fF
C107 a_n801_n100# a_n321_n100# 0.01fF
C108 a_447_n100# a_n33_n100# 0.01fF
C109 a_447_n100# a_639_n100# 0.04fF
C110 a_n801_n100# a_n225_n100# 0.01fF
C111 a_n33_n100# a_63_n100# 0.09fF
C112 a_639_n100# a_63_n100# 0.01fF
C113 a_399_131# a_303_n197# 0.01fF
C114 a_n801_n100# a_n609_n100# 0.04fF
C115 a_n801_n100# a_n513_n100# 0.02fF
C116 a_n417_n100# a_351_n100# 0.01fF
C117 a_n417_n100# w_n1031_n319# 0.05fF
C118 a_n177_131# a_207_131# 0.01fF
C119 a_n81_n197# a_n129_n100# 0.00fF
C120 a_735_n100# a_n801_n100# 0.00fF
C121 a_543_n100# a_n129_n100# 0.01fF
C122 a_n657_n197# a_n753_131# 0.01fF
C123 a_n273_n197# a_n369_131# 0.01fF
C124 a_n801_n100# a_447_n100# 0.00fF
C125 a_n657_n197# w_n1031_n319# 0.16fF
C126 a_255_n100# a_207_131# 0.00fF
C127 w_n1031_n319# a_n753_131# 0.17fF
C128 a_303_n197# a_15_131# 0.00fF
C129 a_n81_n197# a_n369_131# 0.00fF
C130 a_n801_n100# a_63_n100# 0.01fF
C131 a_351_n100# w_n1031_n319# 0.05fF
C132 a_255_n100# a_n33_n100# 0.02fF
C133 a_255_n100# a_639_n100# 0.02fF
C134 a_591_131# a_303_n197# 0.00fF
C135 a_n657_n197# a_687_n197# 0.00fF
C136 a_n753_131# a_687_n197# 0.00fF
C137 a_495_n197# a_207_131# 0.00fF
C138 a_159_n100# a_n321_n100# 0.01fF
C139 w_n1031_n319# a_687_n197# 0.13fF
C140 a_159_n100# a_n225_n100# 0.02fF
C141 a_n705_n100# a_n321_n100# 0.02fF
C142 a_n417_n100# a_n129_n100# 0.02fF
C143 a_n705_n100# a_n225_n100# 0.01fF
C144 a_399_131# a_447_n100# 0.00fF
C145 a_159_n100# a_n609_n100# 0.01fF
C146 a_159_n100# a_n513_n100# 0.01fF
C147 a_399_131# a_n561_131# 0.01fF
C148 a_n801_n100# a_255_n100# 0.01fF
C149 a_n705_n100# a_n609_n100# 0.09fF
C150 a_n705_n100# a_n513_n100# 0.04fF
C151 a_111_n197# a_399_131# 0.00fF
C152 a_n465_n197# a_207_131# 0.00fF
C153 a_n417_n100# a_n369_131# 0.00fF
C154 a_735_n100# a_159_n100# 0.01fF
C155 a_n273_n197# a_303_n197# 0.01fF
C156 a_n705_n100# a_735_n100# 0.00fF
C157 a_159_n100# a_447_n100# 0.02fF
C158 a_351_n100# a_n129_n100# 0.01fF
C159 a_n129_n100# w_n1031_n319# 0.04fF
C160 a_n705_n100# a_447_n100# 0.01fF
C161 a_n81_n197# a_303_n197# 0.01fF
C162 a_n657_n197# a_n369_131# 0.00fF
C163 a_n369_131# a_n753_131# 0.01fF
C164 a_159_n100# a_111_n197# 0.00fF
C165 a_n561_131# a_15_131# 0.01fF
C166 a_159_n100# a_63_n100# 0.09fF
C167 a_111_n197# a_15_131# 0.01fF
C168 a_15_131# a_63_n100# 0.00fF
C169 a_399_131# a_n177_131# 0.01fF
C170 a_n705_n100# a_63_n100# 0.01fF
C171 a_n369_131# w_n1031_n319# 0.13fF
C172 a_n321_n100# a_n273_n197# 0.00fF
C173 a_591_131# a_n561_131# 0.00fF
C174 a_n273_n197# a_n225_n100# 0.00fF
C175 a_111_n197# a_591_131# 0.00fF
C176 a_543_n100# a_n321_n100# 0.01fF
C177 a_n369_131# a_687_n197# 0.00fF
C178 a_15_131# a_n177_131# 0.04fF
C179 a_543_n100# a_n225_n100# 0.01fF
C180 a_543_n100# a_n609_n100# 0.01fF
C181 a_543_n100# a_n513_n100# 0.01fF
C182 a_159_n100# a_255_n100# 0.09fF
C183 a_495_n197# a_399_131# 0.01fF
C184 a_591_131# a_n177_131# 0.01fF
C185 a_n705_n100# a_255_n100# 0.01fF
C186 a_n273_n197# a_n561_131# 0.00fF
C187 a_735_n100# a_543_n100# 0.04fF
C188 a_111_n197# a_n273_n197# 0.01fF
C189 a_n657_n197# a_303_n197# 0.01fF
C190 a_303_n197# a_n753_131# 0.00fF
C191 a_543_n100# a_447_n100# 0.09fF
C192 a_n81_n197# a_n561_131# 0.00fF
C193 a_n81_n197# a_111_n197# 0.04fF
C194 a_399_131# a_n465_n197# 0.00fF
C195 a_495_n197# a_15_131# 0.00fF
C196 a_351_n100# a_303_n197# 0.00fF
C197 a_n417_n100# a_n321_n100# 0.09fF
C198 a_543_n100# a_63_n100# 0.01fF
C199 a_303_n197# w_n1031_n319# 0.11fF
C200 a_n417_n100# a_n225_n100# 0.04fF
C201 a_n273_n197# a_n177_131# 0.01fF
C202 a_n417_n100# a_n609_n100# 0.04fF
C203 a_495_n197# a_591_131# 0.01fF
C204 a_n417_n100# a_n513_n100# 0.09fF
C205 a_303_n197# a_687_n197# 0.01fF
C206 a_15_131# a_n465_n197# 0.00fF
C207 a_n81_n197# a_n177_131# 0.01fF
C208 a_351_n100# a_n321_n100# 0.01fF
C209 a_n417_n100# a_735_n100# 0.01fF
C210 a_n321_n100# w_n1031_n319# 0.05fF
C211 a_351_n100# a_n225_n100# 0.01fF
C212 a_n657_n197# a_n609_n100# 0.00fF
C213 a_n225_n100# w_n1031_n319# 0.04fF
C214 a_n417_n100# a_447_n100# 0.01fF
C215 a_639_n100# a_n33_n100# 0.01fF
C216 a_591_131# a_n465_n197# 0.00fF
C217 a_543_n100# a_255_n100# 0.02fF
C218 a_351_n100# a_n609_n100# 0.01fF
C219 a_n417_n100# a_63_n100# 0.01fF
C220 a_351_n100# a_n513_n100# 0.01fF
C221 a_n609_n100# w_n1031_n319# 0.06fF
C222 a_n513_n100# w_n1031_n319# 0.05fF
C223 a_495_n197# a_n273_n197# 0.01fF
C224 a_735_n100# a_351_n100# 0.02fF
C225 a_n657_n197# a_n561_131# 0.01fF
C226 a_n561_131# a_n753_131# 0.04fF
C227 a_735_n100# w_n1031_n319# 0.15fF
C228 a_n657_n197# a_111_n197# 0.01fF
C229 a_111_n197# a_n753_131# 0.00fF
C230 a_351_n100# a_447_n100# 0.09fF
C231 a_n81_n197# a_495_n197# 0.01fF
C232 a_447_n100# w_n1031_n319# 0.05fF
C233 a_543_n100# a_495_n197# 0.00fF
C234 a_n369_131# a_303_n197# 0.00fF
C235 a_n561_131# w_n1031_n319# 0.14fF
C236 a_n801_n100# a_n33_n100# 0.01fF
C237 a_n801_n100# a_639_n100# 0.00fF
C238 a_351_n100# a_63_n100# 0.02fF
C239 a_111_n197# w_n1031_n319# 0.12fF
C240 w_n1031_n319# a_63_n100# 0.04fF
C241 a_735_n100# a_687_n197# 0.00fF
C242 a_n273_n197# a_n465_n197# 0.04fF
C243 a_n321_n100# a_n129_n100# 0.04fF
C244 a_n129_n100# a_n225_n100# 0.09fF
C245 a_n417_n100# a_255_n100# 0.01fF
C246 a_n81_n197# a_n465_n197# 0.01fF
C247 a_n561_131# a_687_n197# 0.00fF
C248 a_n657_n197# a_n177_131# 0.00fF
C249 a_n177_131# a_n753_131# 0.01fF
C250 a_111_n197# a_687_n197# 0.01fF
C251 a_n321_n100# a_n369_131# 0.00fF
C252 a_n129_n100# a_n609_n100# 0.01fF
C253 a_n513_n100# a_n129_n100# 0.02fF
C254 a_n177_131# w_n1031_n319# 0.13fF
C255 a_399_131# a_207_131# 0.04fF
C256 a_735_n100# a_n129_n100# 0.01fF
C257 a_351_n100# a_255_n100# 0.09fF
C258 a_255_n100# w_n1031_n319# 0.05fF
C259 a_447_n100# a_n129_n100# 0.01fF
C260 a_n177_131# a_687_n197# 0.00fF
C261 a_159_n100# a_207_131# 0.00fF
C262 a_n129_n100# a_63_n100# 0.04fF
C263 a_n657_n197# a_495_n197# 0.00fF
C264 a_15_131# a_207_131# 0.04fF
C265 a_495_n197# a_n753_131# 0.00fF
C266 a_n417_n100# a_n465_n197# 0.00fF
C267 a_159_n100# a_n33_n100# 0.04fF
C268 a_159_n100# a_639_n100# 0.01fF
C269 a_n369_131# a_n561_131# 0.04fF
C270 a_495_n197# w_n1031_n319# 0.11fF
C271 a_15_131# a_n33_n100# 0.00fF
C272 a_n705_n100# a_n33_n100# 0.01fF
C273 a_111_n197# a_n369_131# 0.00fF
C274 a_n705_n100# a_639_n100# 0.00fF
C275 a_591_131# a_207_131# 0.01fF
C276 a_n129_n100# a_n177_131# 0.00fF
C277 a_n657_n197# a_n465_n197# 0.04fF
C278 a_n465_n197# a_n753_131# 0.00fF
C279 a_591_131# a_639_n100# 0.00fF
C280 a_495_n197# a_687_n197# 0.04fF
C281 a_n465_n197# w_n1031_n319# 0.14fF
C282 a_255_n100# a_n129_n100# 0.02fF
C283 a_n369_131# a_n177_131# 0.04fF
C284 a_159_n100# a_n801_n100# 0.01fF
C285 a_n705_n100# a_n801_n100# 0.09fF
C286 a_n465_n197# a_687_n197# 0.00fF
C287 a_n273_n197# a_207_131# 0.00fF
C288 a_n321_n100# a_n225_n100# 0.09fF
C289 a_n81_n197# a_207_131# 0.00fF
C290 a_n561_131# a_303_n197# 0.00fF
C291 a_111_n197# a_303_n197# 0.04fF
C292 a_n321_n100# a_n609_n100# 0.02fF
C293 a_n81_n197# a_n33_n100# 0.00fF
C294 a_n321_n100# a_n513_n100# 0.04fF
C295 a_495_n197# a_n369_131# 0.00fF
C296 a_543_n100# a_n33_n100# 0.01fF
C297 a_543_n100# a_639_n100# 0.09fF
C298 a_n609_n100# a_n225_n100# 0.02fF
C299 a_n513_n100# a_n225_n100# 0.02fF
C300 a_735_n100# a_n321_n100# 0.01fF
C301 a_399_131# a_15_131# 0.01fF
C302 a_n513_n100# a_n609_n100# 0.09fF
C303 a_735_n100# a_n225_n100# 0.01fF
C304 a_n321_n100# a_447_n100# 0.01fF
C305 a_447_n100# a_n225_n100# 0.01fF
C306 a_303_n197# a_n177_131# 0.00fF
C307 a_n369_131# a_n465_n197# 0.01fF
C308 a_n321_n100# a_63_n100# 0.02fF
C309 a_735_n100# a_n609_n100# 0.00fF
C310 a_735_n100# a_n513_n100# 0.00fF
C311 a_399_131# a_591_131# 0.04fF
C312 a_n225_n100# a_63_n100# 0.02fF
C313 a_447_n100# a_n609_n100# 0.01fF
C314 a_n513_n100# a_447_n100# 0.01fF
C315 a_n705_n100# a_159_n100# 0.01fF
C316 a_543_n100# a_n801_n100# 0.00fF
C317 a_n561_131# a_n609_n100# 0.00fF
C318 a_n513_n100# a_n561_131# 0.00fF
C319 a_255_n100# a_303_n197# 0.00fF
C320 a_n609_n100# a_63_n100# 0.01fF
C321 w_n1031_n319# VSUBS 3.95fF
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=5.63e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=3.6625e+11p ps=3.78e+06u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
C0 VPWR X 0.30fF
C1 VPB a_27_47# 0.12fF
C2 A VPWR 0.02fF
C3 VGND VPWR 0.06fF
C4 VPB VPWR 0.24fF
C5 VPWR a_27_47# 0.24fF
C6 A X 0.01fF
C7 VGND X 0.19fF
C8 A VGND 0.02fF
C9 VPB X 0.00fF
C10 a_27_47# X 0.26fF
C11 VPB A 0.10fF
C12 A a_27_47# 0.21fF
C13 VGND a_27_47# 0.19fF
C14 VGND VNB 0.28fF
C15 X VNB 0.00fF
C16 VPWR VNB 0.08fF
C17 A VNB 0.13fF
C18 VPB VNB 0.43fF
C19 a_27_47# VNB 0.15fF
.ends

.subckt precharge_pmos sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131#
+ VSUBS
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_pr__pfet_01v8_VCG74W_0/a_543_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_159_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n609_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_495_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n705_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_255_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n657_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n369_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_351_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n417_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n801_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_303_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n129_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n513_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n465_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n561_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_63_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n225_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_399_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_111_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n321_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n273_n197#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_15_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n753_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_639_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_591_131# sky130_fd_pr__pfet_01v8_VCG74W_0/a_207_131#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_735_n100# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n33_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_687_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_447_n100#
+ sky130_fd_pr__pfet_01v8_VCG74W_0/a_n81_n197# sky130_fd_pr__pfet_01v8_VCG74W_0/a_n177_131#
+ VSUBS sky130_fd_pr__pfet_01v8_VCG74W
C0 sky130_fd_pr__pfet_01v8_VCG74W_0/w_n1031_n319# VSUBS 3.95fF
.ends

.subckt current_tail a_543_n100# a_159_n100# a_n609_n100# a_n1569_n100# a_n705_n100#
+ a_255_n100# a_1407_n100# a_351_n100# a_n417_n100# a_n801_n100# a_1503_n100# a_1119_n100#
+ a_n1377_n100# a_n129_n100# a_n513_n100# a_1215_n100# a_63_n100# a_n1089_n100# a_n1473_n100#
+ a_n225_n100# a_1311_n100# a_927_n100# a_n1185_n100# a_n321_n100# a_1023_n100# a_639_n100#
+ a_n1281_n100# a_735_n100# a_n33_n100# a_n897_n100# a_831_n100# a_447_n100# a_n1521_122#
+ a_n993_n100# a_n1763_n274#
X0 a_n801_n100# a_n1521_122# a_n897_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n513_n100# a_n1521_122# a_n609_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n321_n100# a_n1521_122# a_n417_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n225_n100# a_n1521_122# a_n321_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_n897_n100# a_n1521_122# a_n993_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 a_n705_n100# a_n1521_122# a_n801_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n609_n100# a_n1521_122# a_n705_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n417_n100# a_n1521_122# a_n513_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n129_n100# a_n1521_122# a_n225_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_63_n100# a_n1521_122# a_n33_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_927_n100# a_n1521_122# a_831_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11 a_1023_n100# a_n1521_122# a_927_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_n1569_n100# a_n1763_n274# a_n1763_n274# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=6.2e+11p ps=5.24e+06u w=1e+06u l=150000u
X13 a_1119_n100# a_n1521_122# a_1023_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_1215_n100# a_n1521_122# a_1119_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_1311_n100# a_n1521_122# a_1215_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_1407_n100# a_n1521_122# a_1311_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_1503_n100# a_n1521_122# a_1407_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1763_n274# a_n1763_n274# a_1503_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n33_n100# a_n1521_122# a_n129_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_351_n100# a_n1521_122# a_255_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X21 a_159_n100# a_n1521_122# a_63_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22 a_255_n100# a_n1521_122# a_159_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_447_n100# a_n1521_122# a_351_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X24 a_543_n100# a_n1521_122# a_447_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X25 a_639_n100# a_n1521_122# a_543_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_735_n100# a_n1521_122# a_639_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_831_n100# a_n1521_122# a_735_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n1473_n100# a_n1521_122# a_n1569_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X29 a_n1377_n100# a_n1521_122# a_n1473_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X30 a_n1281_n100# a_n1521_122# a_n1377_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X31 a_n1185_n100# a_n1521_122# a_n1281_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X32 a_n1089_n100# a_n1521_122# a_n1185_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X33 a_n993_n100# a_n1521_122# a_n1089_n100# a_n1763_n274# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n801_n100# a_n1377_n100# 0.01fF
C1 a_735_n100# a_n609_n100# 0.00fF
C2 a_n129_n100# a_n1569_n100# 0.00fF
C3 a_447_n100# a_n993_n100# 0.00fF
C4 a_1023_n100# a_n513_n100# 0.00fF
C5 a_159_n100# a_1407_n100# 0.00fF
C6 a_n129_n100# a_n801_n100# 0.01fF
C7 a_543_n100# a_n129_n100# 0.01fF
C8 a_255_n100# a_1407_n100# 0.01fF
C9 a_n1473_n100# a_n1521_122# 0.03fF
C10 a_447_n100# a_159_n100# 0.02fF
C11 a_n129_n100# a_n1377_n100# 0.00fF
C12 a_447_n100# a_255_n100# 0.04fF
C13 a_n33_n100# a_1407_n100# 0.00fF
C14 a_1119_n100# a_1407_n100# 0.02fF
C15 a_n417_n100# a_n225_n100# 0.04fF
C16 a_831_n100# a_1503_n100# 0.01fF
C17 a_447_n100# a_n33_n100# 0.01fF
C18 a_n705_n100# a_351_n100# 0.01fF
C19 a_639_n100# a_n801_n100# 0.00fF
C20 a_447_n100# a_1119_n100# 0.01fF
C21 a_639_n100# a_543_n100# 0.09fF
C22 a_n705_n100# a_n1473_n100# 0.01fF
C23 a_831_n100# a_351_n100# 0.01fF
C24 a_1215_n100# a_1503_n100# 0.02fF
C25 a_1215_n100# a_351_n100# 0.01fF
C26 a_927_n100# a_n513_n100# 0.00fF
C27 a_159_n100# a_1023_n100# 0.01fF
C28 a_n1089_n100# a_63_n100# 0.01fF
C29 a_255_n100# a_1023_n100# 0.01fF
C30 a_639_n100# a_n129_n100# 0.01fF
C31 a_n321_n100# a_n1089_n100# 0.01fF
C32 a_n705_n100# a_n609_n100# 0.09fF
C33 a_n1185_n100# a_n1281_n100# 0.09fF
C34 a_831_n100# a_n609_n100# 0.00fF
C35 a_n33_n100# a_1023_n100# 0.01fF
C36 a_1119_n100# a_1023_n100# 0.09fF
C37 a_63_n100# a_n513_n100# 0.01fF
C38 a_n417_n100# a_447_n100# 0.01fF
C39 a_n1569_n100# a_n1281_n100# 0.02fF
C40 a_1503_n100# a_1311_n100# 0.04fF
C41 a_n801_n100# a_n1281_n100# 0.01fF
C42 a_n321_n100# a_n513_n100# 0.04fF
C43 a_1311_n100# a_351_n100# 0.01fF
C44 a_63_n100# a_n897_n100# 0.01fF
C45 a_n225_n100# a_1407_n100# 0.00fF
C46 a_159_n100# a_927_n100# 0.01fF
C47 a_n1377_n100# a_n1281_n100# 0.09fF
C48 a_n321_n100# a_n897_n100# 0.01fF
C49 a_735_n100# a_n513_n100# 0.00fF
C50 a_255_n100# a_927_n100# 0.01fF
C51 a_n129_n100# a_n1281_n100# 0.01fF
C52 a_447_n100# a_n225_n100# 0.01fF
C53 a_n993_n100# a_63_n100# 0.01fF
C54 a_n417_n100# a_1023_n100# 0.00fF
C55 a_735_n100# a_n897_n100# 0.00fF
C56 a_n1089_n100# a_n1521_122# 0.03fF
C57 a_n33_n100# a_927_n100# 0.01fF
C58 a_n321_n100# a_n993_n100# 0.01fF
C59 a_1119_n100# a_927_n100# 0.04fF
C60 a_159_n100# a_63_n100# 0.09fF
C61 a_255_n100# a_63_n100# 0.04fF
C62 a_n321_n100# a_159_n100# 0.01fF
C63 a_n1521_122# a_n513_n100# 0.03fF
C64 a_255_n100# a_n321_n100# 0.01fF
C65 a_n225_n100# a_1023_n100# 0.00fF
C66 a_447_n100# a_1407_n100# 0.01fF
C67 a_n33_n100# a_63_n100# 0.09fF
C68 a_1119_n100# a_63_n100# 0.01fF
C69 a_n705_n100# a_n1089_n100# 0.02fF
C70 a_159_n100# a_735_n100# 0.01fF
C71 a_n1185_n100# a_351_n100# 0.00fF
C72 a_n1521_122# a_n897_n100# 0.03fF
C73 a_n33_n100# a_n321_n100# 0.02fF
C74 a_n1185_n100# a_n1473_n100# 0.02fF
C75 a_n321_n100# a_1119_n100# 0.00fF
C76 a_255_n100# a_735_n100# 0.01fF
C77 a_n417_n100# a_927_n100# 0.00fF
C78 a_n1473_n100# a_n1569_n100# 0.09fF
C79 a_543_n100# a_1503_n100# 0.01fF
C80 a_n705_n100# a_n513_n100# 0.04fF
C81 a_n801_n100# a_351_n100# 0.01fF
C82 a_n33_n100# a_735_n100# 0.01fF
C83 a_543_n100# a_351_n100# 0.04fF
C84 a_735_n100# a_1119_n100# 0.02fF
C85 a_831_n100# a_n513_n100# 0.00fF
C86 a_n801_n100# a_n1473_n100# 0.01fF
C87 a_1407_n100# a_1023_n100# 0.02fF
C88 a_n1185_n100# a_n609_n100# 0.01fF
C89 a_n705_n100# a_n897_n100# 0.04fF
C90 a_n417_n100# a_63_n100# 0.01fF
C91 a_n1473_n100# a_n1377_n100# 0.09fF
C92 a_n129_n100# a_1503_n100# 0.00fF
C93 a_n225_n100# a_927_n100# 0.01fF
C94 a_447_n100# a_1023_n100# 0.01fF
C95 a_n129_n100# a_351_n100# 0.01fF
C96 a_n1569_n100# a_n609_n100# 0.01fF
C97 a_n129_n100# a_n1473_n100# 0.00fF
C98 a_n417_n100# a_n321_n100# 0.09fF
C99 a_255_n100# a_n1521_122# 0.03fF
C100 a_n801_n100# a_n609_n100# 0.04fF
C101 a_543_n100# a_n609_n100# 0.01fF
C102 a_n705_n100# a_n993_n100# 0.02fF
C103 a_n1377_n100# a_n609_n100# 0.01fF
C104 a_n417_n100# a_735_n100# 0.01fF
C105 a_n225_n100# a_63_n100# 0.02fF
C106 a_n705_n100# a_159_n100# 0.01fF
C107 a_639_n100# a_1503_n100# 0.01fF
C108 a_n129_n100# a_n609_n100# 0.01fF
C109 a_831_n100# a_159_n100# 0.01fF
C110 a_639_n100# a_351_n100# 0.02fF
C111 a_1407_n100# a_927_n100# 0.01fF
C112 a_n321_n100# a_n225_n100# 0.09fF
C113 a_n705_n100# a_255_n100# 0.01fF
C114 a_1215_n100# a_159_n100# 0.01fF
C115 a_831_n100# a_255_n100# 0.01fF
C116 a_1215_n100# a_255_n100# 0.01fF
C117 a_447_n100# a_927_n100# 0.01fF
C118 a_n705_n100# a_n33_n100# 0.01fF
C119 a_735_n100# a_n225_n100# 0.01fF
C120 a_n33_n100# a_831_n100# 0.01fF
C121 a_831_n100# a_1119_n100# 0.02fF
C122 a_1215_n100# a_n33_n100# 0.00fF
C123 a_1407_n100# a_63_n100# 0.00fF
C124 a_1215_n100# a_1119_n100# 0.09fF
C125 a_639_n100# a_n609_n100# 0.00fF
C126 a_447_n100# a_63_n100# 0.02fF
C127 a_n1185_n100# a_n1089_n100# 0.09fF
C128 a_159_n100# a_1311_n100# 0.01fF
C129 a_n1281_n100# a_351_n100# 0.00fF
C130 a_927_n100# a_1023_n100# 0.09fF
C131 a_447_n100# a_n321_n100# 0.01fF
C132 a_255_n100# a_1311_n100# 0.01fF
C133 a_n1089_n100# a_n1569_n100# 0.01fF
C134 a_n1473_n100# a_n1281_n100# 0.04fF
C135 a_735_n100# a_1407_n100# 0.01fF
C136 a_n705_n100# a_n417_n100# 0.02fF
C137 a_n801_n100# a_n1089_n100# 0.02fF
C138 a_543_n100# a_n1089_n100# 0.00fF
C139 a_n417_n100# a_831_n100# 0.00fF
C140 a_n1185_n100# a_n513_n100# 0.01fF
C141 a_n33_n100# a_1311_n100# 0.00fF
C142 a_n417_n100# a_1215_n100# 0.00fF
C143 a_1311_n100# a_1119_n100# 0.04fF
C144 a_447_n100# a_735_n100# 0.02fF
C145 a_n1377_n100# a_n1089_n100# 0.02fF
C146 a_n1569_n100# a_n513_n100# 0.01fF
C147 a_63_n100# a_1023_n100# 0.01fF
C148 a_n1185_n100# a_n897_n100# 0.02fF
C149 a_n1281_n100# a_n609_n100# 0.01fF
C150 a_n129_n100# a_n1089_n100# 0.01fF
C151 a_n801_n100# a_n513_n100# 0.02fF
C152 a_543_n100# a_n513_n100# 0.01fF
C153 a_n321_n100# a_1023_n100# 0.00fF
C154 a_n705_n100# a_n225_n100# 0.01fF
C155 a_n1569_n100# a_n897_n100# 0.01fF
C156 a_831_n100# a_n225_n100# 0.01fF
C157 a_n1377_n100# a_n513_n100# 0.01fF
C158 a_n1521_122# a_1407_n100# 0.03fF
C159 a_n801_n100# a_n897_n100# 0.09fF
C160 a_1215_n100# a_n225_n100# 0.00fF
C161 a_543_n100# a_n897_n100# 0.00fF
C162 a_n1185_n100# a_n993_n100# 0.04fF
C163 a_n129_n100# a_n513_n100# 0.02fF
C164 a_735_n100# a_1023_n100# 0.02fF
C165 a_447_n100# a_n1521_122# 0.03fF
C166 a_n1377_n100# a_n897_n100# 0.01fF
C167 a_n1569_n100# a_n993_n100# 0.01fF
C168 a_n1185_n100# a_159_n100# 0.00fF
C169 a_n801_n100# a_n993_n100# 0.04fF
C170 a_n129_n100# a_n897_n100# 0.01fF
C171 a_543_n100# a_n993_n100# 0.00fF
C172 a_n1185_n100# a_255_n100# 0.00fF
C173 a_927_n100# a_63_n100# 0.01fF
C174 a_831_n100# a_1407_n100# 0.01fF
C175 a_n1377_n100# a_n993_n100# 0.02fF
C176 a_n801_n100# a_159_n100# 0.01fF
C177 a_1503_n100# a_351_n100# 0.01fF
C178 a_543_n100# a_159_n100# 0.02fF
C179 a_n1185_n100# a_n33_n100# 0.01fF
C180 a_n321_n100# a_927_n100# 0.00fF
C181 a_1215_n100# a_1407_n100# 0.04fF
C182 a_639_n100# a_n513_n100# 0.01fF
C183 a_n705_n100# a_447_n100# 0.01fF
C184 a_n129_n100# a_n993_n100# 0.01fF
C185 a_1311_n100# a_n225_n100# 0.00fF
C186 a_n801_n100# a_255_n100# 0.01fF
C187 a_543_n100# a_255_n100# 0.02fF
C188 a_447_n100# a_831_n100# 0.02fF
C189 a_n1377_n100# a_159_n100# 0.00fF
C190 a_n1521_122# a_1023_n100# 0.03fF
C191 a_n33_n100# a_n1569_n100# 0.00fF
C192 a_1215_n100# a_447_n100# 0.01fF
C193 a_255_n100# a_n1377_n100# 0.00fF
C194 a_639_n100# a_n897_n100# 0.00fF
C195 a_n129_n100# a_159_n100# 0.02fF
C196 a_735_n100# a_927_n100# 0.04fF
C197 a_n33_n100# a_n801_n100# 0.01fF
C198 a_n33_n100# a_543_n100# 0.01fF
C199 a_543_n100# a_1119_n100# 0.01fF
C200 a_n129_n100# a_255_n100# 0.02fF
C201 a_n321_n100# a_63_n100# 0.02fF
C202 a_n1089_n100# a_n1281_n100# 0.04fF
C203 a_n33_n100# a_n1377_n100# 0.00fF
C204 a_n609_n100# a_351_n100# 0.01fF
C205 a_n1473_n100# a_n609_n100# 0.01fF
C206 a_639_n100# a_n993_n100# 0.00fF
C207 a_1311_n100# a_1407_n100# 0.09fF
C208 a_n33_n100# a_n129_n100# 0.09fF
C209 a_n417_n100# a_n1185_n100# 0.01fF
C210 a_n129_n100# a_1119_n100# 0.00fF
C211 a_831_n100# a_1023_n100# 0.04fF
C212 a_735_n100# a_63_n100# 0.01fF
C213 a_1215_n100# a_1023_n100# 0.04fF
C214 a_n1281_n100# a_n513_n100# 0.01fF
C215 a_639_n100# a_159_n100# 0.01fF
C216 a_447_n100# a_1311_n100# 0.01fF
C217 a_n417_n100# a_n1569_n100# 0.01fF
C218 a_n321_n100# a_735_n100# 0.01fF
C219 a_639_n100# a_255_n100# 0.02fF
C220 a_n417_n100# a_n801_n100# 0.02fF
C221 a_n417_n100# a_543_n100# 0.01fF
C222 a_n1281_n100# a_n897_n100# 0.02fF
C223 a_n1185_n100# a_n225_n100# 0.01fF
C224 a_639_n100# a_n33_n100# 0.01fF
C225 a_n417_n100# a_n1377_n100# 0.01fF
C226 a_639_n100# a_1119_n100# 0.01fF
C227 a_n417_n100# a_n129_n100# 0.02fF
C228 a_n1569_n100# a_n225_n100# 0.00fF
C229 a_n1521_122# a_63_n100# 0.03fF
C230 a_n1281_n100# a_n993_n100# 0.02fF
C231 a_n705_n100# a_927_n100# 0.00fF
C232 a_1311_n100# a_1023_n100# 0.02fF
C233 a_n801_n100# a_n225_n100# 0.01fF
C234 a_831_n100# a_927_n100# 0.09fF
C235 a_543_n100# a_n225_n100# 0.01fF
C236 a_n321_n100# a_n1521_122# 0.03fF
C237 a_1215_n100# a_927_n100# 0.02fF
C238 a_159_n100# a_n1281_n100# 0.00fF
C239 a_n1377_n100# a_n225_n100# 0.01fF
C240 a_255_n100# a_n1281_n100# 0.00fF
C241 a_n129_n100# a_n225_n100# 0.09fF
C242 a_n705_n100# a_63_n100# 0.01fF
C243 a_n1089_n100# a_351_n100# 0.00fF
C244 a_n417_n100# a_639_n100# 0.01fF
C245 a_n1473_n100# a_n1089_n100# 0.02fF
C246 a_831_n100# a_63_n100# 0.01fF
C247 a_n1185_n100# a_447_n100# 0.00fF
C248 a_n33_n100# a_n1281_n100# 0.00fF
C249 a_1215_n100# a_63_n100# 0.01fF
C250 a_n705_n100# a_n321_n100# 0.02fF
C251 a_831_n100# a_n321_n100# 0.01fF
C252 a_543_n100# a_1407_n100# 0.01fF
C253 a_1215_n100# a_n321_n100# 0.00fF
C254 a_1311_n100# a_927_n100# 0.02fF
C255 a_351_n100# a_n513_n100# 0.01fF
C256 a_447_n100# a_n801_n100# 0.00fF
C257 a_n1473_n100# a_n513_n100# 0.01fF
C258 a_447_n100# a_543_n100# 0.09fF
C259 a_n705_n100# a_735_n100# 0.00fF
C260 a_n1089_n100# a_n609_n100# 0.01fF
C261 a_639_n100# a_n225_n100# 0.01fF
C262 a_831_n100# a_735_n100# 0.09fF
C263 a_n129_n100# a_1407_n100# 0.00fF
C264 a_1215_n100# a_735_n100# 0.01fF
C265 a_351_n100# a_n897_n100# 0.00fF
C266 a_n1473_n100# a_n897_n100# 0.01fF
C267 a_447_n100# a_n129_n100# 0.01fF
C268 a_n417_n100# a_n1281_n100# 0.01fF
C269 a_1311_n100# a_63_n100# 0.00fF
C270 a_n609_n100# a_n513_n100# 0.09fF
C271 a_n993_n100# a_351_n100# 0.00fF
C272 a_n321_n100# a_1311_n100# 0.00fF
C273 a_n1473_n100# a_n993_n100# 0.01fF
C274 a_543_n100# a_1023_n100# 0.01fF
C275 a_639_n100# a_1407_n100# 0.01fF
C276 a_n705_n100# a_n1521_122# 0.03fF
C277 a_n609_n100# a_n897_n100# 0.02fF
C278 a_159_n100# a_1503_n100# 0.00fF
C279 a_831_n100# a_n1521_122# 0.03fF
C280 a_159_n100# a_351_n100# 0.04fF
C281 a_255_n100# a_1503_n100# 0.00fF
C282 a_n1473_n100# a_159_n100# 0.00fF
C283 a_1215_n100# a_n1521_122# 0.03fF
C284 a_735_n100# a_1311_n100# 0.01fF
C285 a_n1281_n100# a_n225_n100# 0.01fF
C286 a_447_n100# a_639_n100# 0.04fF
C287 a_255_n100# a_351_n100# 0.09fF
C288 a_n129_n100# a_1023_n100# 0.01fF
C289 a_n609_n100# a_n993_n100# 0.02fF
C290 a_n33_n100# a_1503_n100# 0.00fF
C291 a_1503_n100# a_1119_n100# 0.02fF
C292 a_n33_n100# a_351_n100# 0.02fF
C293 a_1119_n100# a_351_n100# 0.01fF
C294 a_n33_n100# a_n1473_n100# 0.00fF
C295 a_n705_n100# a_831_n100# 0.00fF
C296 a_159_n100# a_n609_n100# 0.01fF
C297 a_255_n100# a_n609_n100# 0.01fF
C298 a_1215_n100# a_831_n100# 0.02fF
C299 a_543_n100# a_927_n100# 0.02fF
C300 a_639_n100# a_1023_n100# 0.02fF
C301 a_n1185_n100# a_63_n100# 0.00fF
C302 a_n33_n100# a_n609_n100# 0.01fF
C303 a_n1185_n100# a_n321_n100# 0.01fF
C304 a_n1569_n100# a_63_n100# 0.00fF
C305 a_n129_n100# a_927_n100# 0.01fF
C306 a_n1089_n100# a_n513_n100# 0.01fF
C307 a_n801_n100# a_63_n100# 0.01fF
C308 a_n417_n100# a_351_n100# 0.01fF
C309 a_543_n100# a_63_n100# 0.01fF
C310 a_n321_n100# a_n1569_n100# 0.00fF
C311 a_n417_n100# a_n1473_n100# 0.01fF
C312 a_n801_n100# a_n321_n100# 0.01fF
C313 a_543_n100# a_n321_n100# 0.01fF
C314 a_n1377_n100# a_63_n100# 0.00fF
C315 a_831_n100# a_1311_n100# 0.01fF
C316 a_n1089_n100# a_n897_n100# 0.04fF
C317 a_1215_n100# a_1311_n100# 0.09fF
C318 a_n129_n100# a_63_n100# 0.04fF
C319 a_n321_n100# a_n1377_n100# 0.01fF
C320 a_639_n100# a_927_n100# 0.02fF
C321 a_n801_n100# a_735_n100# 0.00fF
C322 a_n225_n100# a_351_n100# 0.01fF
C323 a_n417_n100# a_n609_n100# 0.04fF
C324 a_543_n100# a_735_n100# 0.04fF
C325 a_n129_n100# a_n321_n100# 0.04fF
C326 a_n1473_n100# a_n225_n100# 0.00fF
C327 a_n1089_n100# a_n993_n100# 0.09fF
C328 a_n897_n100# a_n513_n100# 0.02fF
C329 a_n129_n100# a_735_n100# 0.01fF
C330 a_159_n100# a_n1089_n100# 0.00fF
C331 a_639_n100# a_63_n100# 0.01fF
C332 a_255_n100# a_n1089_n100# 0.00fF
C333 a_n993_n100# a_n513_n100# 0.01fF
C334 a_n225_n100# a_n609_n100# 0.02fF
C335 a_1503_n100# a_1407_n100# 0.09fF
C336 a_639_n100# a_n321_n100# 0.01fF
C337 a_1407_n100# a_351_n100# 0.01fF
C338 a_n33_n100# a_n1089_n100# 0.01fF
C339 a_n993_n100# a_n897_n100# 0.09fF
C340 a_159_n100# a_n513_n100# 0.01fF
C341 a_447_n100# a_1503_n100# 0.01fF
C342 a_n705_n100# a_n1185_n100# 0.01fF
C343 a_255_n100# a_n513_n100# 0.01fF
C344 a_447_n100# a_351_n100# 0.09fF
C345 a_639_n100# a_735_n100# 0.09fF
C346 a_159_n100# a_n897_n100# 0.01fF
C347 a_n129_n100# a_n1521_122# 0.03fF
C348 a_n705_n100# a_n1569_n100# 0.01fF
C349 a_n33_n100# a_n513_n100# 0.01fF
C350 a_255_n100# a_n897_n100# 0.01fF
C351 a_1119_n100# a_n513_n100# 0.00fF
C352 a_n705_n100# a_n801_n100# 0.09fF
C353 a_n705_n100# a_543_n100# 0.00fF
C354 a_831_n100# a_n801_n100# 0.00fF
C355 a_n1281_n100# a_63_n100# 0.00fF
C356 a_543_n100# a_831_n100# 0.02fF
C357 a_159_n100# a_n993_n100# 0.01fF
C358 a_n33_n100# a_n897_n100# 0.01fF
C359 a_n705_n100# a_n1377_n100# 0.01fF
C360 a_1215_n100# a_543_n100# 0.01fF
C361 a_447_n100# a_n609_n100# 0.01fF
C362 a_1503_n100# a_1023_n100# 0.01fF
C363 a_n321_n100# a_n1281_n100# 0.01fF
C364 a_n417_n100# a_n1089_n100# 0.01fF
C365 a_255_n100# a_n993_n100# 0.00fF
C366 a_351_n100# a_1023_n100# 0.01fF
C367 a_n705_n100# a_n129_n100# 0.01fF
C368 a_639_n100# a_n1521_122# 0.03fF
C369 a_n129_n100# a_831_n100# 0.01fF
C370 a_n33_n100# a_n993_n100# 0.01fF
C371 a_1215_n100# a_n129_n100# 0.00fF
C372 a_255_n100# a_159_n100# 0.09fF
C373 a_n417_n100# a_n513_n100# 0.09fF
C374 a_n1089_n100# a_n225_n100# 0.01fF
C375 a_n33_n100# a_159_n100# 0.04fF
C376 a_n609_n100# a_1023_n100# 0.00fF
C377 a_159_n100# a_1119_n100# 0.01fF
C378 a_543_n100# a_1311_n100# 0.01fF
C379 a_n417_n100# a_n897_n100# 0.01fF
C380 a_n33_n100# a_255_n100# 0.02fF
C381 a_n705_n100# a_639_n100# 0.00fF
C382 a_255_n100# a_1119_n100# 0.01fF
C383 a_639_n100# a_831_n100# 0.04fF
C384 a_1503_n100# a_927_n100# 0.01fF
C385 a_1215_n100# a_639_n100# 0.01fF
C386 a_351_n100# a_927_n100# 0.01fF
C387 a_n225_n100# a_n513_n100# 0.02fF
C388 a_n33_n100# a_1119_n100# 0.01fF
C389 a_n129_n100# a_1311_n100# 0.00fF
C390 a_n417_n100# a_n993_n100# 0.01fF
C391 a_n1521_122# a_n1281_n100# 0.03fF
C392 a_n225_n100# a_n897_n100# 0.01fF
C393 a_1503_n100# a_63_n100# 0.00fF
C394 a_n417_n100# a_159_n100# 0.01fF
C395 a_351_n100# a_63_n100# 0.02fF
C396 a_447_n100# a_n1089_n100# 0.00fF
C397 a_n609_n100# a_927_n100# 0.00fF
C398 a_n417_n100# a_255_n100# 0.01fF
C399 a_n1473_n100# a_63_n100# 0.00fF
C400 a_n705_n100# a_n1281_n100# 0.01fF
C401 a_n225_n100# a_n993_n100# 0.01fF
C402 a_639_n100# a_1311_n100# 0.01fF
C403 a_n321_n100# a_351_n100# 0.01fF
C404 a_n1473_n100# a_n321_n100# 0.01fF
C405 a_n417_n100# a_n33_n100# 0.02fF
C406 a_n1185_n100# a_n1569_n100# 0.02fF
C407 a_n417_n100# a_1119_n100# 0.00fF
C408 a_1503_n100# a_735_n100# 0.01fF
C409 a_159_n100# a_n225_n100# 0.02fF
C410 a_447_n100# a_n513_n100# 0.01fF
C411 a_n1185_n100# a_n801_n100# 0.02fF
C412 a_735_n100# a_351_n100# 0.02fF
C413 a_n609_n100# a_63_n100# 0.01fF
C414 a_255_n100# a_n225_n100# 0.01fF
C415 a_n801_n100# a_n1569_n100# 0.01fF
C416 a_n1185_n100# a_n1377_n100# 0.04fF
C417 a_447_n100# a_n897_n100# 0.00fF
C418 a_n321_n100# a_n609_n100# 0.02fF
C419 a_543_n100# a_n801_n100# 0.00fF
C420 a_n33_n100# a_n225_n100# 0.04fF
C421 a_n1185_n100# a_n129_n100# 0.01fF
C422 a_n225_n100# a_1119_n100# 0.00fF
C423 a_n1377_n100# a_n1569_n100# 0.04fF
C424 a_1503_n100# a_n1763_n274# 0.14fF
C425 a_1407_n100# a_n1763_n274# 0.07fF
C426 a_1311_n100# a_n1763_n274# 0.06fF
C427 a_1215_n100# a_n1763_n274# 0.05fF
C428 a_1119_n100# a_n1763_n274# 0.04fF
C429 a_1023_n100# a_n1763_n274# 0.04fF
C430 a_927_n100# a_n1763_n274# 0.03fF
C431 a_831_n100# a_n1763_n274# 0.03fF
C432 a_735_n100# a_n1763_n274# 0.03fF
C433 a_639_n100# a_n1763_n274# 0.03fF
C434 a_543_n100# a_n1763_n274# 0.03fF
C435 a_447_n100# a_n1763_n274# 0.03fF
C436 a_351_n100# a_n1763_n274# 0.03fF
C437 a_255_n100# a_n1763_n274# 0.03fF
C438 a_159_n100# a_n1763_n274# 0.03fF
C439 a_63_n100# a_n1763_n274# 0.02fF
C440 a_n33_n100# a_n1763_n274# 0.03fF
C441 a_n129_n100# a_n1763_n274# 0.02fF
C442 a_n225_n100# a_n1763_n274# 0.03fF
C443 a_n321_n100# a_n1763_n274# 0.03fF
C444 a_n417_n100# a_n1763_n274# 0.03fF
C445 a_n513_n100# a_n1763_n274# 0.03fF
C446 a_n609_n100# a_n1763_n274# 0.03fF
C447 a_n705_n100# a_n1763_n274# 0.03fF
C448 a_n801_n100# a_n1763_n274# 0.03fF
C449 a_n897_n100# a_n1763_n274# 0.03fF
C450 a_n993_n100# a_n1763_n274# 0.03fF
C451 a_n1089_n100# a_n1763_n274# 0.04fF
C452 a_n1185_n100# a_n1763_n274# 0.04fF
C453 a_n1281_n100# a_n1763_n274# 0.05fF
C454 a_n1377_n100# a_n1763_n274# 0.06fF
C455 a_n1473_n100# a_n1763_n274# 0.08fF
C456 a_n1569_n100# a_n1763_n274# 0.15fF
C457 a_n1521_122# a_n1763_n274# 3.88fF
.ends

.subckt sky130_fd_pr__nfet_01v8_J3WY8C a_n4080_n100# a_n1188_122# a_282_n188# a_n978_n188#
+ a_1542_n188# a_n3918_n188# a_3432_122# a_1752_122# a_n3708_122# a_2382_n188# a_4228_n100#
+ a_n2028_122# a_n1818_n188# a_3222_n188# a_n348_122# a_n2658_n188# a_n3288_122# a_4062_n188#
+ a_72_122# a_n558_n188# a_n3498_n188# a_1122_n188# a_912_122# a_n4172_n100# a_3852_122#
+ a_n1398_n188# a_2172_122# a_n4128_122# a_n2448_122# a_492_122# a_n768_122# a_n2238_n188#
+ a_n138_n188# a_n3078_n188# a_1962_n188# a_702_n188# a_3012_122# a_1332_122# a_n1608_122#
+ a_n4382_n100# a_2802_n188# a_2592_122# a_3642_n188# a_n2868_122# VSUBS
X0 a_n4080_n100# a_n1398_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=1.24e+13p pd=1.048e+08u as=1.24e+13p ps=1.048e+08u w=1e+06u l=150000u
X1 a_n4080_n100# a_1332_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_n4080_n100# a_n2868_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n4080_n100# a_2802_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n4080_n100# a_n3288_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n4080_n100# a_3222_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n4080_n100# a_72_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n4080_n100# a_n1608_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_n4080_n100# a_1542_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n4080_n100# a_n138_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n4080_n100# a_282_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n4080_n100# a_n3498_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_n4080_n100# a_3432_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_n4080_n100# a_n1818_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n4080_n100# a_1752_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n4080_n100# a_492_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n4080_n100# a_2172_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n4080_n100# a_n3708_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n4080_n100# a_n348_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_n4080_n100# a_3642_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_n4080_n100# a_4062_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n4080_n100# a_n2028_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_n4080_n100# a_1962_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n4080_n100# a_702_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n4080_n100# a_n3918_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_n4080_n100# a_n558_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_n4080_n100# a_3852_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_4228_n100# a_4228_n100# a_4228_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X28 a_n4080_n100# a_n2238_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_n4080_n100# a_n768_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n4080_n100# a_912_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n4080_n100# a_n4128_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_n4080_n100# a_n2448_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_n4080_n100# a_2382_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_n4080_n100# a_n978_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n4382_n100# a_n4382_n100# a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=6.2e+11p pd=5.24e+06u as=0p ps=0u w=1e+06u l=150000u
X36 a_n4080_n100# a_n1188_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_n4080_n100# a_1122_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_n4080_n100# a_n2658_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_n4080_n100# a_2592_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_n4080_n100# a_n3078_n188# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_n4080_n100# a_3012_122# a_n4172_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 a_n3708_122# a_n4128_122# 0.01fF
C1 a_n4172_n100# a_3432_122# 0.06fF
C2 a_3432_122# a_3852_122# 0.01fF
C3 a_n4172_n100# a_2382_n188# 0.02fF
C4 a_n4080_n100# a_3432_122# 0.02fF
C5 a_2382_n188# a_3852_122# 0.00fF
C6 a_n3288_122# a_n3918_n188# 0.00fF
C7 a_4228_n100# a_n4172_n100# 0.14fF
C8 a_n4080_n100# a_2382_n188# 0.06fF
C9 a_4228_n100# a_3852_122# 0.01fF
C10 a_4228_n100# a_n4080_n100# 0.21fF
C11 a_1542_n188# a_1962_n188# 0.01fF
C12 a_282_n188# a_n1188_122# 0.00fF
C13 a_n3708_122# a_n4172_n100# 0.06fF
C14 a_492_122# a_1962_n188# 0.00fF
C15 a_n2028_122# a_n1398_n188# 0.00fF
C16 a_n2658_n188# a_n4128_122# 0.00fF
C17 a_n4172_n100# a_1122_n188# 0.02fF
C18 a_1962_n188# a_1332_122# 0.00fF
C19 a_n138_n188# a_n1188_122# 0.00fF
C20 a_n3708_122# a_n4080_n100# 0.02fF
C21 a_n2238_n188# a_n3708_122# 0.00fF
C22 a_282_n188# a_n4172_n100# 0.02fF
C23 a_n4172_n100# a_912_122# 0.06fF
C24 a_n4080_n100# a_1122_n188# 0.06fF
C25 a_1542_n188# a_2382_n188# 0.01fF
C26 a_282_n188# a_n4080_n100# 0.06fF
C27 a_n138_n188# a_n4172_n100# 0.02fF
C28 a_n4080_n100# a_912_122# 0.02fF
C29 a_n1188_122# a_n2658_n188# 0.00fF
C30 a_2592_122# a_3222_n188# 0.00fF
C31 a_n1188_122# a_n558_n188# 0.00fF
C32 a_3012_122# a_1962_n188# 0.00fF
C33 a_2382_n188# a_1332_122# 0.00fF
C34 a_n3078_n188# a_n3708_122# 0.00fF
C35 a_n768_122# a_282_n188# 0.00fF
C36 a_2172_122# a_1962_n188# 0.00fF
C37 a_702_n188# a_n4172_n100# 0.02fF
C38 a_n138_n188# a_n4080_n100# 0.06fF
C39 a_n3498_n188# a_n4128_122# 0.00fF
C40 a_n1608_122# a_n1818_n188# 0.00fF
C41 a_n2028_122# a_n3288_122# 0.00fF
C42 a_3222_n188# a_1752_122# 0.00fF
C43 a_n4172_n100# a_n2658_n188# 0.02fF
C44 a_n4172_n100# a_n558_n188# 0.02fF
C45 a_n1818_n188# a_n978_n188# 0.01fF
C46 a_n768_122# a_n138_n188# 0.00fF
C47 a_3012_122# a_3432_122# 0.01fF
C48 a_n1608_122# a_n978_n188# 0.00fF
C49 a_702_n188# a_n4080_n100# 0.06fF
C50 a_2172_122# a_3432_122# 0.00fF
C51 a_n1818_n188# a_n2448_122# 0.00fF
C52 a_2592_122# a_4062_n188# 0.00fF
C53 a_n1608_122# a_n2448_122# 0.01fF
C54 a_3012_122# a_2382_n188# 0.00fF
C55 a_72_122# a_1122_n188# 0.00fF
C56 a_n768_122# a_702_n188# 0.00fF
C57 a_n4080_n100# a_n2658_n188# 0.06fF
C58 a_2172_122# a_2382_n188# 0.00fF
C59 a_n4080_n100# a_n558_n188# 0.06fF
C60 a_n2238_n188# a_n2658_n188# 0.01fF
C61 a_1542_n188# a_1122_n188# 0.01fF
C62 a_n2448_122# a_n978_n188# 0.00fF
C63 a_282_n188# a_72_122# 0.00fF
C64 a_3012_122# a_4228_n100# 0.00fF
C65 a_72_122# a_912_122# 0.01fF
C66 a_492_122# a_1122_n188# 0.00fF
C67 a_n1818_n188# a_n2868_122# 0.00fF
C68 a_2802_n188# a_1962_n188# 0.01fF
C69 a_n768_122# a_n558_n188# 0.00fF
C70 a_1542_n188# a_282_n188# 0.00fF
C71 a_n1608_122# a_n2868_122# 0.00fF
C72 a_1542_n188# a_912_122# 0.00fF
C73 a_282_n188# a_492_122# 0.00fF
C74 a_1122_n188# a_1332_122# 0.00fF
C75 a_492_122# a_912_122# 0.01fF
C76 a_72_122# a_n138_n188# 0.00fF
C77 a_282_n188# a_1332_122# 0.00fF
C78 a_n3498_n188# a_n4172_n100# 0.02fF
C79 a_n3078_n188# a_n2658_n188# 0.01fF
C80 a_n4382_n100# a_n2868_122# 0.00fF
C81 a_912_122# a_1332_122# 0.01fF
C82 a_n2448_122# a_n2868_122# 0.01fF
C83 a_n3708_122# a_n3918_n188# 0.00fF
C84 a_n348_122# a_1122_n188# 0.00fF
C85 a_2802_n188# a_3432_122# 0.00fF
C86 a_n138_n188# a_492_122# 0.00fF
C87 a_702_n188# a_72_122# 0.00fF
C88 a_n348_122# a_282_n188# 0.00fF
C89 a_1542_n188# a_702_n188# 0.01fF
C90 a_2802_n188# a_2382_n188# 0.01fF
C91 a_n3498_n188# a_n4080_n100# 0.06fF
C92 a_2592_122# a_n4172_n100# 0.06fF
C93 a_n348_122# a_912_122# 0.00fF
C94 a_n138_n188# a_1332_122# 0.00fF
C95 a_n3498_n188# a_n2238_n188# 0.00fF
C96 a_702_n188# a_492_122# 0.00fF
C97 a_72_122# a_n558_n188# 0.00fF
C98 a_2592_122# a_3852_122# 0.00fF
C99 a_2172_122# a_1122_n188# 0.00fF
C100 a_4228_n100# a_2802_n188# 0.00fF
C101 a_702_n188# a_1332_122# 0.00fF
C102 a_2592_122# a_n4080_n100# 0.02fF
C103 a_n348_122# a_n138_n188# 0.00fF
C104 a_492_122# a_n558_n188# 0.00fF
C105 a_3642_n188# a_3222_n188# 0.01fF
C106 a_n4172_n100# a_1752_122# 0.06fF
C107 a_2172_122# a_912_122# 0.00fF
C108 a_n3498_n188# a_n3078_n188# 0.01fF
C109 a_n348_122# a_702_n188# 0.00fF
C110 a_n4080_n100# a_1752_122# 0.02fF
C111 a_n348_122# a_n558_n188# 0.00fF
C112 a_n2658_n188# a_n3918_n188# 0.00fF
C113 a_3642_n188# a_4062_n188# 0.01fF
C114 a_702_n188# a_2172_122# 0.00fF
C115 a_1542_n188# a_2592_122# 0.00fF
C116 a_n138_n188# a_n1398_n188# 0.00fF
C117 a_n3708_122# a_n3288_122# 0.01fF
C118 a_2592_122# a_1332_122# 0.00fF
C119 a_1542_n188# a_1752_122# 0.00fF
C120 a_n3498_n188# a_n3918_n188# 0.01fF
C121 a_492_122# a_1752_122# 0.00fF
C122 a_n2658_n188# a_n1398_n188# 0.00fF
C123 a_3432_122# a_1962_n188# 0.00fF
C124 a_3642_n188# a_n4172_n100# 0.02fF
C125 a_n558_n188# a_n1398_n188# 0.01fF
C126 a_1752_122# a_1332_122# 0.01fF
C127 a_2382_n188# a_1962_n188# 0.01fF
C128 a_3642_n188# a_3852_122# 0.00fF
C129 a_n4382_n100# a_n4128_122# 0.00fF
C130 a_3642_n188# a_n4080_n100# 0.06fF
C131 a_3012_122# a_2592_122# 0.01fF
C132 a_n1188_122# a_n1818_n188# 0.00fF
C133 a_2592_122# a_2172_122# 0.01fF
C134 a_n1188_122# a_n1608_122# 0.01fF
C135 a_n2868_122# a_n4128_122# 0.00fF
C136 a_3432_122# a_2382_n188# 0.00fF
C137 a_n1188_122# a_n978_n188# 0.00fF
C138 a_3012_122# a_1752_122# 0.00fF
C139 a_n2028_122# a_n2658_n188# 0.00fF
C140 a_n1188_122# a_n2448_122# 0.00fF
C141 a_n2028_122# a_n558_n188# 0.00fF
C142 a_n1818_n188# a_n4172_n100# 0.02fF
C143 a_2172_122# a_1752_122# 0.01fF
C144 a_4228_n100# a_3432_122# 0.00fF
C145 a_n1608_122# a_n4172_n100# 0.06fF
C146 a_n2658_n188# a_n3288_122# 0.00fF
C147 a_n4172_n100# a_n978_n188# 0.02fF
C148 a_n1818_n188# a_n4080_n100# 0.06fF
C149 a_n2238_n188# a_n1818_n188# 0.01fF
C150 a_n4382_n100# a_n4172_n100# 0.21fF
C151 a_n1608_122# a_n4080_n100# 0.02fF
C152 a_n2448_122# a_n4172_n100# 0.06fF
C153 a_1122_n188# a_1962_n188# 0.01fF
C154 a_n2238_n188# a_n1608_122# 0.00fF
C155 a_2592_122# a_2802_n188# 0.00fF
C156 a_n768_122# a_n1818_n188# 0.00fF
C157 a_n4080_n100# a_n978_n188# 0.06fF
C158 a_n768_122# a_n1608_122# 0.01fF
C159 a_n2238_n188# a_n978_n188# 0.00fF
C160 a_912_122# a_1962_n188# 0.00fF
C161 a_n4382_n100# a_n4080_n100# 0.14fF
C162 a_n2448_122# a_n4080_n100# 0.02fF
C163 a_n4172_n100# a_n2868_122# 0.06fF
C164 a_n2238_n188# a_n2448_122# 0.00fF
C165 a_n768_122# a_n978_n188# 0.00fF
C166 a_n3498_n188# a_n2028_122# 0.00fF
C167 a_2802_n188# a_1752_122# 0.00fF
C168 a_n3078_n188# a_n1818_n188# 0.00fF
C169 a_n3078_n188# a_n1608_122# 0.00fF
C170 a_n3498_n188# a_n3288_122# 0.00fF
C171 a_1122_n188# a_2382_n188# 0.00fF
C172 a_n4080_n100# a_n2868_122# 0.02fF
C173 a_n2238_n188# a_n2868_122# 0.00fF
C174 a_702_n188# a_1962_n188# 0.00fF
C175 a_n3078_n188# a_n4382_n100# 0.00fF
C176 a_2382_n188# a_912_122# 0.00fF
C177 a_n3078_n188# a_n2448_122# 0.00fF
C178 a_3012_122# a_3642_n188# 0.00fF
C179 a_72_122# a_n978_n188# 0.00fF
C180 a_4062_n188# a_3222_n188# 0.01fF
C181 a_3642_n188# a_2172_122# 0.00fF
C182 a_n3078_n188# a_n2868_122# 0.00fF
C183 a_492_122# a_n978_n188# 0.00fF
C184 a_n348_122# a_n1818_n188# 0.00fF
C185 a_n348_122# a_n1608_122# 0.00fF
C186 a_n348_122# a_n978_n188# 0.00fF
C187 a_282_n188# a_1122_n188# 0.01fF
C188 a_1122_n188# a_912_122# 0.00fF
C189 a_3642_n188# a_2802_n188# 0.01fF
C190 a_282_n188# a_912_122# 0.00fF
C191 a_n4382_n100# a_n3918_n188# 0.01fF
C192 a_n2448_122# a_n3918_n188# 0.00fF
C193 a_n4172_n100# a_3222_n188# 0.02fF
C194 a_n138_n188# a_1122_n188# 0.00fF
C195 a_2592_122# a_1962_n188# 0.00fF
C196 a_3852_122# a_3222_n188# 0.00fF
C197 a_282_n188# a_n138_n188# 0.01fF
C198 a_n138_n188# a_912_122# 0.00fF
C199 a_702_n188# a_1122_n188# 0.01fF
C200 a_n3708_122# a_n2658_n188# 0.00fF
C201 a_n2868_122# a_n3918_n188# 0.00fF
C202 a_n4080_n100# a_3222_n188# 0.06fF
C203 a_1752_122# a_1962_n188# 0.00fF
C204 a_282_n188# a_702_n188# 0.01fF
C205 a_2592_122# a_3432_122# 0.01fF
C206 a_702_n188# a_912_122# 0.00fF
C207 a_n1818_n188# a_n1398_n188# 0.01fF
C208 a_n4172_n100# a_n4128_122# 0.06fF
C209 a_n1608_122# a_n1398_n188# 0.00fF
C210 a_n4172_n100# a_4062_n188# 0.02fF
C211 a_2592_122# a_2382_n188# 0.00fF
C212 a_282_n188# a_n558_n188# 0.01fF
C213 a_4062_n188# a_3852_122# 0.00fF
C214 a_n978_n188# a_n1398_n188# 0.01fF
C215 a_n558_n188# a_912_122# 0.00fF
C216 a_702_n188# a_n138_n188# 0.01fF
C217 a_2592_122# a_4228_n100# 0.00fF
C218 a_n2448_122# a_n1398_n188# 0.00fF
C219 a_n4080_n100# a_n4128_122# 0.02fF
C220 a_n4080_n100# a_4062_n188# 0.06fF
C221 a_2382_n188# a_1752_122# 0.00fF
C222 a_n138_n188# a_n558_n188# 0.01fF
C223 a_n1188_122# a_n4172_n100# 0.06fF
C224 a_n3498_n188# a_n3708_122# 0.00fF
C225 a_n2868_122# a_n1398_n188# 0.00fF
C226 a_n2028_122# a_n1818_n188# 0.00fF
C227 a_702_n188# a_n558_n188# 0.00fF
C228 a_n2028_122# a_n1608_122# 0.01fF
C229 a_n3078_n188# a_n4128_122# 0.00fF
C230 a_n1818_n188# a_n3288_122# 0.00fF
C231 a_n1188_122# a_n4080_n100# 0.02fF
C232 a_n2238_n188# a_n1188_122# 0.00fF
C233 a_n2028_122# a_n978_n188# 0.00fF
C234 a_n768_122# a_n1188_122# 0.01fF
C235 a_2592_122# a_1122_n188# 0.00fF
C236 a_n2028_122# a_n2448_122# 0.01fF
C237 a_n4172_n100# a_3852_122# 0.06fF
C238 a_n4382_n100# a_n3288_122# 0.00fF
C239 a_n2448_122# a_n3288_122# 0.01fF
C240 a_n4172_n100# a_n4080_n100# 15.77fF
C241 a_n2238_n188# a_n4172_n100# 0.02fF
C242 a_n2028_122# a_n2868_122# 0.01fF
C243 a_n4080_n100# a_3852_122# 0.02fF
C244 a_1122_n188# a_1752_122# 0.00fF
C245 a_n768_122# a_n4172_n100# 0.06fF
C246 a_n2868_122# a_n3288_122# 0.01fF
C247 a_282_n188# a_1752_122# 0.00fF
C248 a_n2238_n188# a_n4080_n100# 0.06fF
C249 a_912_122# a_1752_122# 0.01fF
C250 a_3012_122# a_3222_n188# 0.00fF
C251 a_n3498_n188# a_n2658_n188# 0.01fF
C252 a_2172_122# a_3222_n188# 0.00fF
C253 a_n768_122# a_n4080_n100# 0.02fF
C254 a_72_122# a_n1188_122# 0.00fF
C255 a_3642_n188# a_3432_122# 0.00fF
C256 a_n768_122# a_n2238_n188# 0.00fF
C257 a_n3078_n188# a_n4172_n100# 0.02fF
C258 a_3642_n188# a_2382_n188# 0.00fF
C259 a_n4128_122# a_n3918_n188# 0.00fF
C260 a_n3078_n188# a_n4080_n100# 0.06fF
C261 a_3642_n188# a_4228_n100# 0.00fF
C262 a_n3078_n188# a_n2238_n188# 0.01fF
C263 a_72_122# a_n4172_n100# 0.06fF
C264 a_702_n188# a_1752_122# 0.00fF
C265 a_3012_122# a_4062_n188# 0.00fF
C266 a_1542_n188# a_n4172_n100# 0.02fF
C267 a_n4172_n100# a_492_122# 0.06fF
C268 a_n348_122# a_n1188_122# 0.01fF
C269 a_72_122# a_n4080_n100# 0.02fF
C270 a_2802_n188# a_3222_n188# 0.01fF
C271 a_n4172_n100# a_1332_122# 0.06fF
C272 a_1542_n188# a_n4080_n100# 0.06fF
C273 a_n768_122# a_72_122# 0.01fF
C274 a_n4080_n100# a_492_122# 0.02fF
C275 a_n348_122# a_n4172_n100# 0.06fF
C276 a_n4080_n100# a_1332_122# 0.02fF
C277 a_n768_122# a_492_122# 0.00fF
C278 a_n4172_n100# a_n3918_n188# 0.02fF
C279 a_2802_n188# a_4062_n188# 0.00fF
C280 a_n348_122# a_n4080_n100# 0.02fF
C281 a_3012_122# a_n4172_n100# 0.06fF
C282 a_n4172_n100# a_2172_122# 0.06fF
C283 a_n4080_n100# a_n3918_n188# 0.06fF
C284 a_3012_122# a_3852_122# 0.01fF
C285 a_n348_122# a_n768_122# 0.01fF
C286 a_3012_122# a_n4080_n100# 0.02fF
C287 a_1542_n188# a_72_122# 0.00fF
C288 a_n1188_122# a_n1398_n188# 0.00fF
C289 a_2592_122# a_1752_122# 0.01fF
C290 a_n4080_n100# a_2172_122# 0.02fF
C291 a_72_122# a_492_122# 0.01fF
C292 a_1542_n188# a_492_122# 0.00fF
C293 a_72_122# a_1332_122# 0.00fF
C294 a_n4382_n100# a_n3708_122# 0.00fF
C295 a_n3288_122# a_n4128_122# 0.01fF
C296 a_n3708_122# a_n2448_122# 0.00fF
C297 a_n3078_n188# a_n3918_n188# 0.01fF
C298 a_n4172_n100# a_n1398_n188# 0.02fF
C299 a_1542_n188# a_1332_122# 0.00fF
C300 a_492_122# a_1332_122# 0.01fF
C301 a_2802_n188# a_n4172_n100# 0.02fF
C302 a_n348_122# a_72_122# 0.01fF
C303 a_282_n188# a_n978_n188# 0.00fF
C304 a_2802_n188# a_3852_122# 0.00fF
C305 a_n3708_122# a_n2868_122# 0.01fF
C306 a_n4080_n100# a_n1398_n188# 0.06fF
C307 a_n2238_n188# a_n1398_n188# 0.01fF
C308 a_n138_n188# a_n1608_122# 0.00fF
C309 a_n2028_122# a_n1188_122# 0.01fF
C310 a_n348_122# a_492_122# 0.01fF
C311 a_2802_n188# a_n4080_n100# 0.06fF
C312 a_n768_122# a_n1398_n188# 0.00fF
C313 a_n138_n188# a_n978_n188# 0.01fF
C314 a_3012_122# a_1542_n188# 0.00fF
C315 a_3222_n188# a_1962_n188# 0.00fF
C316 a_1542_n188# a_2172_122# 0.00fF
C317 a_n1818_n188# a_n2658_n188# 0.01fF
C318 a_n2028_122# a_n4172_n100# 0.06fF
C319 a_n1818_n188# a_n558_n188# 0.00fF
C320 a_n1608_122# a_n2658_n188# 0.00fF
C321 a_n1608_122# a_n558_n188# 0.00fF
C322 a_n4172_n100# a_n3288_122# 0.06fF
C323 a_2172_122# a_1332_122# 0.01fF
C324 a_n558_n188# a_n978_n188# 0.01fF
C325 a_n2028_122# a_n4080_n100# 0.02fF
C326 a_3432_122# a_3222_n188# 0.00fF
C327 a_n2238_n188# a_n2028_122# 0.00fF
C328 a_n4382_n100# a_n2658_n188# 0.00fF
C329 a_2592_122# a_3642_n188# 0.00fF
C330 a_n2448_122# a_n2658_n188# 0.00fF
C331 a_72_122# a_n1398_n188# 0.00fF
C332 a_n4080_n100# a_n3288_122# 0.02fF
C333 a_n2238_n188# a_n3288_122# 0.00fF
C334 a_2382_n188# a_3222_n188# 0.01fF
C335 a_n768_122# a_n2028_122# 0.00fF
C336 a_n2658_n188# a_n2868_122# 0.00fF
C337 a_4228_n100# a_3222_n188# 0.00fF
C338 a_1542_n188# a_2802_n188# 0.00fF
C339 a_3012_122# a_2172_122# 0.01fF
C340 a_n3078_n188# a_n2028_122# 0.00fF
C341 a_4062_n188# a_3432_122# 0.00fF
C342 a_n3078_n188# a_n3288_122# 0.00fF
C343 a_2802_n188# a_1332_122# 0.00fF
C344 a_n348_122# a_n1398_n188# 0.00fF
C345 a_n3498_n188# a_n4382_n100# 0.00fF
C346 a_n3498_n188# a_n2448_122# 0.00fF
C347 a_4228_n100# a_4062_n188# 0.00fF
C348 a_n4172_n100# a_1962_n188# 0.02fF
C349 a_n3498_n188# a_n2868_122# 0.00fF
C350 a_3012_122# a_2802_n188# 0.00fF
C351 a_2802_n188# a_2172_122# 0.00fF
C352 a_n4080_n100# a_1962_n188# 0.06fF
C353 a_n4080_n100# VSUBS 1.08fF
C354 a_n4172_n100# VSUBS 1.03fF
C355 a_4062_n188# VSUBS 0.11fF
C356 a_4228_n100# VSUBS 0.17fF
C357 a_3642_n188# VSUBS 0.10fF
C358 a_3852_122# VSUBS 0.09fF
C359 a_3222_n188# VSUBS 0.11fF
C360 a_3432_122# VSUBS 0.11fF
C361 a_2802_n188# VSUBS 0.12fF
C362 a_3012_122# VSUBS 0.11fF
C363 a_2382_n188# VSUBS 0.12fF
C364 a_2592_122# VSUBS 0.12fF
C365 a_1962_n188# VSUBS 0.12fF
C366 a_2172_122# VSUBS 0.12fF
C367 a_1542_n188# VSUBS 0.12fF
C368 a_1752_122# VSUBS 0.12fF
C369 a_1122_n188# VSUBS 0.12fF
C370 a_1332_122# VSUBS 0.12fF
C371 a_702_n188# VSUBS 0.12fF
C372 a_912_122# VSUBS 0.12fF
C373 a_282_n188# VSUBS 0.12fF
C374 a_492_122# VSUBS 0.12fF
C375 a_n138_n188# VSUBS 0.12fF
C376 a_72_122# VSUBS 0.12fF
C377 a_n558_n188# VSUBS 0.12fF
C378 a_n348_122# VSUBS 0.12fF
C379 a_n978_n188# VSUBS 0.12fF
C380 a_n768_122# VSUBS 0.12fF
C381 a_n1398_n188# VSUBS 0.12fF
C382 a_n1188_122# VSUBS 0.12fF
C383 a_n1818_n188# VSUBS 0.12fF
C384 a_n1608_122# VSUBS 0.12fF
C385 a_n2238_n188# VSUBS 0.12fF
C386 a_n2028_122# VSUBS 0.12fF
C387 a_n2658_n188# VSUBS 0.12fF
C388 a_n2448_122# VSUBS 0.12fF
C389 a_n3078_n188# VSUBS 0.12fF
C390 a_n2868_122# VSUBS 0.12fF
C391 a_n3498_n188# VSUBS 0.12fF
C392 a_n3288_122# VSUBS 0.12fF
C393 a_n3918_n188# VSUBS 0.12fF
C394 a_n3708_122# VSUBS 0.12fF
C395 a_n4382_n100# VSUBS 0.20fF
C396 a_n4128_122# VSUBS 0.13fF
.ends

.subckt latch_nmos_pair sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
C0 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C2 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C3 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C4 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C5 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C6 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C7 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C8 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C9 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C10 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# -0.00fF
C11 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C12 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C13 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C14 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C15 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C16 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C17 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C18 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C19 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.01fF
C20 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C21 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C22 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C23 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C24 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C25 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C26 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C27 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C28 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C29 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C30 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C31 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C32 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C33 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C34 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C35 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C36 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C37 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C38 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C39 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C40 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C41 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C42 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.30fF
C43 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C44 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C45 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C46 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# -0.00fF
C47 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C48 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.00fF
C49 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C50 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C51 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C52 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C53 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C54 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C55 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.02fF
C56 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C57 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C58 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# -0.00fF
C59 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C60 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C61 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C62 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.02fF
C63 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C64 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C65 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C66 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C67 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.27fF
C68 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C69 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C70 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C71 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C72 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.02fF
C73 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C74 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C75 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C76 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# -0.00fF
C77 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C78 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C79 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# -0.00fF
C80 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C81 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C82 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C83 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C84 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C85 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C86 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C87 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C88 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C89 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C90 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C91 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C92 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C93 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.02fF
C94 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C95 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C96 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C97 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C98 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C99 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C100 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# -0.00fF
C102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# -0.00fF
C103 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C105 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C106 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C107 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C108 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C109 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C110 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C112 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.02fF
C115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C116 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C118 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C119 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C121 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C122 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C123 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C125 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.02fF
C126 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C127 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C129 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.22fF
C130 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C132 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C133 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C134 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C135 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C136 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C137 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C138 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.01fF
C139 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C140 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C141 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C142 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C143 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C146 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C147 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C148 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C149 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C151 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C152 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C153 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C154 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# -0.00fF
C155 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C156 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C157 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C158 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C159 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C160 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C161 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C162 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C163 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.76fF
C164 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C165 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C166 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C167 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C168 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# -0.00fF
C169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C170 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C171 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# -0.00fF
C172 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C173 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C174 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C175 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C176 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C177 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C178 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C179 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# -0.00fF
C180 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C181 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C183 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C184 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C185 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C186 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C187 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C189 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C190 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C191 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C192 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C193 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# -0.00fF
C194 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C195 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C196 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C197 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C201 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C202 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C204 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C206 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C207 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C208 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C209 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.42fF
C210 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C211 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C212 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C213 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C214 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.01fF
C215 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C216 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C217 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C218 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C219 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C221 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.02fF
C222 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C223 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C224 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C225 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C226 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C227 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C228 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C229 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.02fF
C230 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C231 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C232 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C233 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C235 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C236 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C237 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C238 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C239 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.02fF
C240 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C241 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# -0.00fF
C242 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# -0.00fF
C243 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.93fF
C244 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C245 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# -0.00fF
C246 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C247 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.02fF
C248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C249 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C250 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C251 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C252 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C253 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C254 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C255 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C256 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.02fF
C257 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C258 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C259 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C260 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C261 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C262 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# -0.00fF
C264 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C265 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C266 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.02fF
C268 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C269 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C270 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C271 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C272 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C273 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.02fF
C274 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C275 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C276 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C277 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C278 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C279 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C281 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C282 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C283 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C284 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C285 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C286 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.02fF
C287 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C288 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C289 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C290 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C291 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C292 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C293 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C294 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# -0.00fF
C295 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C296 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C297 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C298 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C299 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C300 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C301 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C302 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C303 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C304 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# -0.00fF
C305 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# -0.01fF
C306 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C307 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C308 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C309 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C310 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C311 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C312 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C313 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C314 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C315 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C316 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.01fF
C317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C318 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# -0.00fF
C319 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C320 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C321 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C322 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C323 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.02fF
C324 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C325 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.02fF
C326 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C327 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.00fF
C329 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C330 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C331 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C332 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C333 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C334 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C335 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C336 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C337 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C338 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C339 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C340 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C341 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C342 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C343 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C344 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C345 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 1.18fF
C346 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C347 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C348 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C350 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# -0.00fF
C351 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C352 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C353 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C354 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.01fF
C355 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C356 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C357 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C358 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C359 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C360 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C361 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C362 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C363 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C364 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C365 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C366 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C367 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C368 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C369 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C371 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C372 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C373 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C374 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C376 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# -0.00fF
C377 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C378 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C379 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.02fF
C380 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C381 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C382 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C383 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C384 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C385 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C386 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C388 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C389 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C390 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C391 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C392 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.02fF
C393 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C394 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C395 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.02fF
C396 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C398 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C399 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C400 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C401 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.02fF
C402 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C405 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C406 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C407 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C408 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.27fF
C409 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C410 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C411 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# -0.00fF
C412 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.02fF
C413 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C414 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C415 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.02fF
C416 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C417 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C418 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C419 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C421 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C422 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C424 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C426 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C427 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C428 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C429 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.31fF
C430 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C431 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C432 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C433 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C434 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C435 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C436 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C437 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# -0.00fF
C438 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C439 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C440 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C441 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C442 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C443 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C444 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C445 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.02fF
C446 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C447 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C448 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C449 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# -0.00fF
C450 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.02fF
C451 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C452 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C453 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C454 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C455 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C456 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C457 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C458 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C459 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C460 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C461 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C462 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# -0.00fF
C463 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C464 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C465 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C466 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# -0.00fF
C467 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C468 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C469 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C470 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C471 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.01fF
C472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C473 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C474 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C475 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C476 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C477 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.02fF
C478 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C479 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C480 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C481 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C483 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C484 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C485 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C486 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C487 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# -0.00fF
C488 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C489 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C490 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# -0.00fF
C491 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C492 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C493 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# -0.00fF
C494 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C495 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C496 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C497 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C498 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C499 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C500 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C501 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C503 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C504 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.02fF
C505 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C506 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C507 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.02fF
C508 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C509 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C510 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# -0.01fF
C511 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C512 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C513 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C515 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C516 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C517 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.02fF
C519 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.93fF
C520 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C521 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# -0.00fF
C522 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C523 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C524 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C525 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C526 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C527 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# -0.00fF
C528 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C529 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C530 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C531 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.02fF
C532 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C533 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C534 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C535 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C536 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C537 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C538 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# -0.00fF
C539 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C541 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C542 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# -0.00fF
C543 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C544 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C545 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C546 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.02fF
C547 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C548 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.01fF
C549 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C550 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C551 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C552 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C553 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C554 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# 0.00fF
C555 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C556 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C557 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C558 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C559 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C560 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C561 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C563 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.42fF
C564 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# -0.00fF
C565 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C567 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C568 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.02fF
C569 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C570 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C571 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C572 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C573 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C574 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C575 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C576 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C577 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# -0.00fF
C579 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C580 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C581 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C582 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C583 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C585 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C586 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C587 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# -0.00fF
C588 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C589 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C590 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C591 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C592 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C593 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C594 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C595 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C596 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C597 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C598 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C599 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C600 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C601 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# -0.00fF
C602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C604 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C605 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C606 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.02fF
C607 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C608 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C609 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C610 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C611 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C612 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C613 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C615 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C616 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C617 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C618 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C619 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C620 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C621 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C622 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C623 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C624 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C625 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.02fF
C626 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C627 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C628 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C629 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C630 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C631 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C632 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C633 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C634 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C635 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C637 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 1.18fF
C638 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# -0.00fF
C639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C641 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C642 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C643 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C644 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# -0.00fF
C645 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C646 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# -0.00fF
C647 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C649 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C650 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# -0.00fF
C652 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.02fF
C653 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C654 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.02fF
C655 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C656 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C657 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C658 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C659 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C660 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C661 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.02fF
C662 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C663 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# -0.00fF
C664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C665 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C666 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C667 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C668 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C669 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C671 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C672 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C673 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C674 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C675 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C676 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C677 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C678 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C679 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C680 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C682 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C683 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C684 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C685 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C686 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C687 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C688 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C689 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# -0.00fF
C691 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C692 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C693 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C694 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C695 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C696 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C697 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C699 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# -0.00fF
C700 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C702 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C703 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C704 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C705 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.02fF
C706 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C708 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.02fF
C709 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C710 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C711 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C712 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C713 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C714 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C715 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C716 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C717 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C718 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C719 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# -0.01fF
C720 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C721 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C722 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C724 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C725 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# -0.00fF
C726 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C727 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C728 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C729 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C730 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C731 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C732 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C733 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# -0.00fF
C734 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C735 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# -0.00fF
C736 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C738 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C739 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C740 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.42fF
C741 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C742 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C743 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C744 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C745 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C746 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C747 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C748 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C749 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C750 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C751 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C752 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.02fF
C753 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C754 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C755 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C756 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C757 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C758 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C759 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C760 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C761 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C762 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C763 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C764 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C765 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C766 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C767 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.42fF
C768 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C769 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C770 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C771 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.02fF
C772 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.02fF
C773 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C774 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C775 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C776 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C777 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C778 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C779 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C780 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C781 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C782 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C783 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C784 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C785 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C786 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.02fF
C787 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C788 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C789 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# -0.00fF
C790 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C791 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C792 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C793 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C794 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C795 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.02fF
C796 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C797 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C798 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C799 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C800 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C801 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C802 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C803 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C804 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C805 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C806 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C807 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C808 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C809 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C810 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C811 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# -0.00fF
C812 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C813 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C814 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C815 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C816 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C817 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C818 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C819 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C820 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# -0.00fF
C821 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.02fF
C822 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C823 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C824 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C825 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.57fF
C826 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C827 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C828 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C830 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# -0.00fF
C831 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C832 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C833 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# -0.00fF
C834 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C835 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C836 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C838 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C839 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C840 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C841 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C842 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C843 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C844 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C845 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# -0.00fF
C846 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C847 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.02fF
C848 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C849 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C850 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# -0.00fF
C851 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C852 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C854 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C855 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C856 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# -0.00fF
C857 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C858 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C859 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.44fF
C860 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C861 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C862 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C863 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C864 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# -0.00fF
C865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C866 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C867 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C868 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C869 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.93fF
C870 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C871 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C872 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C873 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C874 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C875 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C876 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C877 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C878 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C879 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# -0.00fF
C880 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C881 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C882 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C883 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C884 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C885 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C886 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# -0.00fF
C887 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C888 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C889 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C890 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C891 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C892 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C893 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C894 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C895 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C896 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C897 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C898 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.02fF
C899 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C900 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C901 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C902 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C903 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C904 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# -0.00fF
C905 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C906 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C907 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C908 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C909 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C910 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C911 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C912 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C913 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C914 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C915 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C916 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C917 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C918 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C919 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C920 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C921 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C922 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C923 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C924 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C925 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C926 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C927 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C928 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C929 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C930 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C931 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C932 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C933 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C934 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.02fF
C935 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C936 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C937 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# -0.00fF
C938 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C939 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C940 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C941 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C942 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C943 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C944 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C945 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C946 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C947 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C948 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C949 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C950 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C951 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C952 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C953 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C954 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C955 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C956 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.24fF
C957 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C958 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C959 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C960 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C961 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C962 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C963 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C964 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C965 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C966 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C967 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.01fF
C968 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C969 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C970 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C971 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C972 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C973 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# -0.00fF
C974 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C975 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C976 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C977 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C978 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C979 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C980 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C981 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C982 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C983 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# -0.00fF
C984 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C985 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C986 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C987 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C988 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C989 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C990 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C991 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C992 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C993 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C994 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C995 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C996 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C997 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C998 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C999 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1000 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1001 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1002 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C1003 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1004 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1005 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C1006 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1007 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C1008 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1009 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1010 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C1011 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1012 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1013 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C1014 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C1015 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C1016 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1017 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1018 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1019 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C1020 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C1021 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1022 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1023 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1024 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# -0.00fF
C1025 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C1026 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1027 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1028 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1029 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1030 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C1031 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C1032 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1033 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1034 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1035 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C1036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C1037 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C1038 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1039 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1040 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1041 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1042 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C1043 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C1044 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1045 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1046 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.01fF
C1047 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1048 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C1050 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C1051 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.02fF
C1052 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1053 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1054 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# -0.00fF
C1055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1056 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C1057 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1058 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1059 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1060 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1061 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C1062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C1064 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C1065 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C1066 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# -0.00fF
C1067 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.02fF
C1068 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1069 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1070 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.00fF
C1071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C1072 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1074 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1075 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.02fF
C1076 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C1077 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1078 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1079 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1081 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1082 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1083 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C1084 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# -0.00fF
C1085 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1086 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# -0.00fF
C1087 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C1088 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1089 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1090 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.01fF
C1091 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# -0.00fF
C1092 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1093 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1094 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1095 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# -0.00fF
C1096 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# -0.00fF
C1097 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1098 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C1099 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.00fF
C1100 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1101 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C1102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1103 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1104 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C1105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C1106 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.01fF
C1107 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1108 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1109 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C1110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1111 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1112 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1113 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1114 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1115 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.02fF
C1116 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1118 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1119 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C1120 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1121 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1122 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1125 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1126 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.02fF
C1129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.31fF
C1131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# -0.00fF
C1132 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1133 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1134 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C1135 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1136 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C1137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1138 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C1139 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.17fF
C1140 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C1141 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1142 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1143 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# -0.00fF
C1145 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# -0.00fF
C1146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C1147 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# -0.00fF
C1148 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1150 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C1151 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C1152 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1153 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1154 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1155 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1156 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1158 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C1159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1161 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C1162 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C1163 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1164 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1165 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C1166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1167 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 1.18fF
C1168 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1169 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1170 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C1172 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1173 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C1175 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C1176 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C1177 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1178 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1179 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1180 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1181 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C1182 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C1183 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C1184 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1185 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1187 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C1190 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1191 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C1192 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1193 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C1194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1195 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1196 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.01fF
C1197 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C1199 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.02fF
C1201 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1202 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.02fF
C1204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C1205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1206 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C1207 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C1208 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.00fF
C1209 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1210 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.02fF
C1211 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C1212 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C1213 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.02fF
C1214 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1215 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1216 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1217 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C1218 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C1219 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C1220 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1221 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# -0.00fF
C1222 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C1223 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# -0.00fF
C1224 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# 0.00fF
C1225 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1226 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1227 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1228 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C1229 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C1230 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1231 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# -0.01fF
C1232 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# -0.00fF
C1233 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1234 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C1235 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1236 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.02fF
C1237 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1238 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C1239 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C1240 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C1241 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C1242 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1243 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1244 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1245 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1246 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1247 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C1248 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C1249 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1250 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.02fF
C1251 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1252 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1253 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1254 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1255 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# -0.00fF
C1256 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1257 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C1258 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# -0.00fF
C1259 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1260 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# -0.00fF
C1261 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1262 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C1263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1264 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1265 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1266 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1267 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1268 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1269 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# -0.00fF
C1270 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1271 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C1272 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# -0.00fF
C1273 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C1274 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C1275 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1276 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1277 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1278 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C1279 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C1281 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.01fF
C1282 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C1283 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1284 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C1285 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1286 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C1287 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1288 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1289 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C1290 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1291 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C1292 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1293 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1294 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1295 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C1296 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1297 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1298 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1299 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1300 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1301 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1302 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1303 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C1304 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C1305 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C1306 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1307 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1308 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1309 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1310 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C1311 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.01fF
C1312 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1313 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1314 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1315 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1316 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C1317 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1318 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C1319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C1320 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.02fF
C1321 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C1322 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# -0.00fF
C1323 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1324 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# -0.00fF
C1325 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1326 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1327 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1329 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.00fF
C1330 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1331 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1332 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# -0.00fF
C1333 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C1334 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1335 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C1336 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1337 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1338 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C1339 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C1340 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1341 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C1342 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1343 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C1344 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C1345 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.02fF
C1346 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1347 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1348 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C1349 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C1350 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C1352 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1353 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1354 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C1355 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C1356 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1357 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1358 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.02fF
C1359 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C1360 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C1362 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1363 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.00fF
C1364 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1365 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# -0.00fF
C1366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# -0.00fF
C1367 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C1368 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1369 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# -0.00fF
C1370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.02fF
C1371 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C1372 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1373 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1374 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C1376 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C1377 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1379 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1380 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C1381 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C1382 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C1383 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C1384 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1385 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C1386 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C1387 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1388 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C1389 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1390 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1391 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1392 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1393 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C1394 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1395 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C1396 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1397 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1398 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1399 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C1401 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1403 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1405 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1406 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1407 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# -0.00fF
C1408 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# 0.02fF
C1409 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1410 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C1411 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1412 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C1413 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1414 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1415 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C1416 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1417 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# -0.00fF
C1418 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1419 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# -0.00fF
C1420 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1421 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1422 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.01fF
C1423 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C1424 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C1425 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.00fF
C1426 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.02fF
C1427 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1428 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1429 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.00fF
C1430 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1431 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# -0.00fF
C1432 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.02fF
C1433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C1434 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1435 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C1436 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1437 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1438 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.57fF
C1439 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C1440 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1441 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C1442 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C1443 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.00fF
C1444 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C1445 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.44fF
C1446 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C1447 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1448 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1449 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1450 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C1451 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1452 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1453 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1454 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1455 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C1456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.00fF
C1457 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C1458 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C1459 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1460 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.02fF
C1461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1462 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C1463 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1464 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1465 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C1466 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.02fF
C1467 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C1468 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1469 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C1470 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1471 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C1472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1473 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1474 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C1475 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1476 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.01fF
C1477 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1478 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C1479 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1480 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C1481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1482 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1483 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1484 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C1485 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.00fF
C1486 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1487 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1488 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C1489 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1490 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1491 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1492 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# -0.00fF
C1493 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C1494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1495 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C1496 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1497 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.00fF
C1498 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1499 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1500 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# -0.00fF
C1501 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1502 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C1503 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1504 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1505 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1506 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C1507 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1508 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1509 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1510 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C1511 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1512 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C1513 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1514 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C1515 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1516 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1517 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1518 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C1519 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1520 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1521 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1522 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1523 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.01fF
C1524 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1525 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C1526 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# 0.57fF
C1527 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1528 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1529 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1530 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1531 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1532 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C1533 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1534 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.02fF
C1535 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1537 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1538 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1539 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C1541 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C1542 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C1543 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C1544 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C1545 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1546 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1547 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C1548 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1549 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1550 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C1551 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1552 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1553 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1554 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C1555 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# -0.00fF
C1556 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1557 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# -0.00fF
C1558 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1559 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C1560 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# VSUBS 1.08fF
C1561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# VSUBS 1.03fF
C1562 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# VSUBS 0.11fF
C1563 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# VSUBS 0.17fF
C1564 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# VSUBS 0.10fF
C1565 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# VSUBS 0.09fF
C1566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# VSUBS 0.11fF
C1567 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# VSUBS 0.11fF
C1568 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# VSUBS 0.12fF
C1569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# VSUBS 0.11fF
C1570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# VSUBS 0.12fF
C1571 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# VSUBS 0.12fF
C1572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# VSUBS 0.12fF
C1573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# VSUBS 0.12fF
C1574 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# VSUBS 0.12fF
C1575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# VSUBS 0.12fF
C1576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# VSUBS 0.12fF
C1577 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# VSUBS 0.12fF
C1578 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# VSUBS 0.12fF
C1579 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# VSUBS 0.12fF
C1580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# VSUBS 0.12fF
C1581 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# VSUBS 0.12fF
C1582 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# VSUBS 0.12fF
C1583 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# VSUBS 0.12fF
C1584 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# VSUBS 0.12fF
C1585 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# VSUBS 0.12fF
C1586 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# VSUBS 0.12fF
C1587 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# VSUBS 0.12fF
C1588 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# VSUBS 0.12fF
C1589 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# VSUBS 0.12fF
C1590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# VSUBS 0.12fF
C1591 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# VSUBS 0.12fF
C1592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# VSUBS 0.12fF
C1593 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# VSUBS 0.12fF
C1594 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# VSUBS 0.12fF
C1595 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# VSUBS 0.12fF
C1596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# VSUBS 0.12fF
C1597 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# VSUBS 0.12fF
C1598 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# VSUBS 0.12fF
C1599 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# VSUBS 0.12fF
C1600 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# VSUBS 0.12fF
C1601 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# VSUBS 0.12fF
C1602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# VSUBS 0.20fF
C1603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# VSUBS 0.13fF
C1604 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# VSUBS 1.08fF
C1605 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# VSUBS 1.03fF
C1606 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# VSUBS 0.11fF
C1607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# VSUBS 0.17fF
C1608 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# VSUBS 0.10fF
C1609 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# VSUBS 0.09fF
C1610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# VSUBS 0.11fF
C1611 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# VSUBS 0.11fF
C1612 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# VSUBS 0.12fF
C1613 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# VSUBS 0.11fF
C1614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# VSUBS 0.12fF
C1615 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# VSUBS 0.12fF
C1616 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# VSUBS 0.12fF
C1617 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# VSUBS 0.12fF
C1618 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# VSUBS 0.12fF
C1619 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# VSUBS 0.12fF
C1620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# VSUBS 0.12fF
C1621 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# VSUBS 0.12fF
C1622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# VSUBS 0.12fF
C1623 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# VSUBS 0.12fF
C1624 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# VSUBS 0.12fF
C1625 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# VSUBS 0.12fF
C1626 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# VSUBS 0.12fF
C1627 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# VSUBS 0.12fF
C1628 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# VSUBS 0.12fF
C1629 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# VSUBS 0.12fF
C1630 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# VSUBS 0.12fF
C1631 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# VSUBS 0.12fF
C1632 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# VSUBS 0.12fF
C1633 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# VSUBS 0.12fF
C1634 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# VSUBS 0.12fF
C1635 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# VSUBS 0.12fF
C1636 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# VSUBS 0.12fF
C1637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# VSUBS 0.12fF
C1638 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# VSUBS 0.12fF
C1639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# VSUBS 0.12fF
C1640 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# VSUBS 0.12fF
C1641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# VSUBS 0.12fF
C1642 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# VSUBS 0.12fF
C1643 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# VSUBS 0.12fF
C1644 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# VSUBS 0.12fF
C1645 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# VSUBS 0.12fF
C1646 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# VSUBS 0.20fF
C1647 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# VSUBS 0.13fF
C1648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# VSUBS 1.08fF
C1649 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# VSUBS 1.03fF
C1650 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# VSUBS 0.11fF
C1651 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# VSUBS 0.17fF
C1652 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# VSUBS 0.10fF
C1653 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# VSUBS 0.09fF
C1654 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# VSUBS 0.11fF
C1655 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# VSUBS 0.11fF
C1656 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# VSUBS 0.12fF
C1657 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# VSUBS 0.11fF
C1658 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# VSUBS 0.12fF
C1659 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# VSUBS 0.12fF
C1660 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# VSUBS 0.12fF
C1661 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# VSUBS 0.12fF
C1662 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# VSUBS 0.12fF
C1663 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# VSUBS 0.12fF
C1664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# VSUBS 0.12fF
C1665 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# VSUBS 0.12fF
C1666 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# VSUBS 0.12fF
C1667 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# VSUBS 0.12fF
C1668 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# VSUBS 0.12fF
C1669 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# VSUBS 0.12fF
C1670 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# VSUBS 0.12fF
C1671 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# VSUBS 0.12fF
C1672 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# VSUBS 0.12fF
C1673 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# VSUBS 0.12fF
C1674 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# VSUBS 0.12fF
C1675 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# VSUBS 0.12fF
C1676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# VSUBS 0.12fF
C1677 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# VSUBS 0.12fF
C1678 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# VSUBS 0.12fF
C1679 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# VSUBS 0.12fF
C1680 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# VSUBS 0.12fF
C1681 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# VSUBS 0.12fF
C1682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# VSUBS 0.12fF
C1683 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# VSUBS 0.12fF
C1684 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# VSUBS 0.12fF
C1685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# VSUBS 0.12fF
C1686 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# VSUBS 0.12fF
C1687 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# VSUBS 0.12fF
C1688 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# VSUBS 0.12fF
C1689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# VSUBS 0.12fF
C1690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# VSUBS 0.20fF
C1691 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# VSUBS 0.13fF
C1692 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# VSUBS 1.08fF
C1693 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# VSUBS 1.03fF
C1694 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# VSUBS 0.11fF
C1695 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# VSUBS 0.17fF
C1696 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# VSUBS 0.10fF
C1697 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# VSUBS 0.09fF
C1698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# VSUBS 0.11fF
C1699 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# VSUBS 0.11fF
C1700 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# VSUBS 0.12fF
C1701 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# VSUBS 0.11fF
C1702 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# VSUBS 0.12fF
C1703 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# VSUBS 0.12fF
C1704 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# VSUBS 0.12fF
C1705 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# VSUBS 0.12fF
C1706 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# VSUBS 0.12fF
C1707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# VSUBS 0.12fF
C1708 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# VSUBS 0.12fF
C1709 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# VSUBS 0.12fF
C1710 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# VSUBS 0.12fF
C1711 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# VSUBS 0.12fF
C1712 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# VSUBS 0.12fF
C1713 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# VSUBS 0.12fF
C1714 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# VSUBS 0.12fF
C1715 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# VSUBS 0.12fF
C1716 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# VSUBS 0.12fF
C1717 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# VSUBS 0.12fF
C1718 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# VSUBS 0.12fF
C1719 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# VSUBS 0.12fF
C1720 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# VSUBS 0.12fF
C1721 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# VSUBS 0.12fF
C1722 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# VSUBS 0.12fF
C1723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# VSUBS 0.12fF
C1724 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# VSUBS 0.12fF
C1725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# VSUBS 0.12fF
C1726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# VSUBS 0.12fF
C1727 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# VSUBS 0.12fF
C1728 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# VSUBS 0.12fF
C1729 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# VSUBS 0.12fF
C1730 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# VSUBS 0.12fF
C1731 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# VSUBS 0.12fF
C1732 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# VSUBS 0.12fF
C1733 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# VSUBS 0.12fF
C1734 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# VSUBS 0.20fF
C1735 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# VSUBS 0.13fF
.ends

.subckt input_diff_pair sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122#
Xsky130_fd_pr__nfet_01v8_J3WY8C_0 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_1 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_2 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_3 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_4 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_5 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_6 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
Xsky130_fd_pr__nfet_01v8_J3WY8C_7 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122#
+ sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122#
+ VSUBS sky130_fd_pr__nfet_01v8_J3WY8C
C0 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C2 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C3 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C5 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C6 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.02fF
C7 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C8 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C9 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C10 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.01fF
C11 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C12 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C13 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C14 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C15 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C16 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C17 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C18 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C19 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C20 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C21 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C22 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C23 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C24 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C25 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C26 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C27 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C28 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C29 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C30 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C31 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C32 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C33 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C34 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C35 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C36 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C37 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C38 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C39 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C40 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C41 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C42 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C43 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C44 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C45 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# -0.00fF
C46 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C47 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C48 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# -0.00fF
C49 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C50 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C51 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C52 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C53 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C54 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C55 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# -0.00fF
C56 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C57 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C58 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C59 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C60 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C61 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C62 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# -0.00fF
C63 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.02fF
C64 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C65 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C66 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C67 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C68 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C69 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C70 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C71 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C72 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C73 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C74 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C75 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C76 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C77 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C78 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C79 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C80 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C81 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C82 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C83 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C84 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C85 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C86 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C87 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C88 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C89 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C90 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C91 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.93fF
C92 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C93 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.02fF
C94 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C95 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C96 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C97 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C98 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C99 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C100 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.02fF
C101 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.02fF
C102 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C103 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C104 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C105 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.01fF
C106 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C107 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C108 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C109 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# -0.00fF
C110 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C111 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C112 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C113 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C114 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C115 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C116 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C117 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C118 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C119 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.01fF
C120 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C121 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C122 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C123 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.02fF
C124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C125 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C126 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.02fF
C127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C128 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# -0.00fF
C129 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C130 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C131 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C132 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C133 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C134 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C135 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C136 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C137 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C138 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.01fF
C139 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C140 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C142 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C143 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C147 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C148 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C149 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C151 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C152 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C153 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C155 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.02fF
C156 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C157 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C158 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C160 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C161 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C162 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# -0.00fF
C163 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C164 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C165 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.00fF
C166 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C167 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C168 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.02fF
C169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C170 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C171 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C172 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C173 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.01fF
C175 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C176 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C177 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C178 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C179 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.00fF
C180 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C181 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.02fF
C182 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C183 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C184 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C185 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C187 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C188 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C189 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.01fF
C190 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C191 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C192 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C193 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C194 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C195 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C196 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C197 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C198 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C199 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.02fF
C200 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C201 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.01fF
C202 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# -0.00fF
C203 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C204 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.02fF
C206 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C207 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C208 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C209 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C210 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# -0.01fF
C211 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C212 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C213 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C214 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C215 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# -0.00fF
C216 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C217 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C218 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C219 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C220 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C221 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C222 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C223 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C224 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.01fF
C225 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.02fF
C226 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.01fF
C227 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C228 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C229 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C230 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C231 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C232 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.02fF
C233 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C234 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C235 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C236 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C237 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C238 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# 0.01fF
C239 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# -0.00fF
C240 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C241 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C242 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C243 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C244 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C245 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C246 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C247 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# -0.00fF
C248 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C249 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C250 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C251 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C252 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C253 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C254 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C255 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# -0.00fF
C256 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C257 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# -0.00fF
C258 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C259 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C260 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C261 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C262 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C263 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C264 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.02fF
C265 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C266 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C267 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C268 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C269 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C270 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.22fF
C271 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C272 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C273 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C274 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C275 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C276 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C277 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.01fF
C278 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C279 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C280 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C281 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.02fF
C283 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C284 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C285 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C286 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C287 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.01fF
C288 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C289 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.02fF
C290 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C291 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C292 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.01fF
C293 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C294 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.02fF
C295 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C296 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C297 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.02fF
C298 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C299 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C300 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C301 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C302 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.02fF
C303 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C304 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C305 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C306 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C307 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C308 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C309 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.02fF
C310 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C311 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C312 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C313 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C314 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C315 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C316 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C317 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C318 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C320 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.00fF
C321 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C322 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C323 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C324 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C325 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C326 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C327 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C328 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C329 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C330 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.42fF
C331 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C332 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C333 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C334 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C335 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C336 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C337 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C338 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C339 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C340 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C341 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C342 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C343 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# -0.00fF
C344 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.57fF
C345 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C346 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C347 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 1.18fF
C348 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C349 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C350 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C352 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.02fF
C353 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.01fF
C354 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C355 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.02fF
C356 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C357 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C358 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C359 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C360 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C361 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C362 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C363 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C364 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C365 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C367 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C368 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C369 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.01fF
C370 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C371 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C372 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.01fF
C373 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C374 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C375 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C376 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C377 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C378 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C379 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C380 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C381 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C382 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.27fF
C383 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C384 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C385 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C386 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C387 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# 0.00fF
C388 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C389 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C390 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C391 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C392 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C393 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C394 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C395 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C396 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C397 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C398 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C399 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C400 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C401 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.78fF
C402 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C404 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C405 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C406 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C407 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C408 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C409 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C410 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C411 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C412 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C413 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C414 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C415 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C416 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C417 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C418 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C419 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.01fF
C420 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.02fF
C421 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C422 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C423 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C424 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C425 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C426 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C427 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C428 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C429 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C430 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C431 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C432 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C433 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# -0.00fF
C434 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C435 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C436 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C437 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C438 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C439 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# -0.01fF
C440 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C441 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.27fF
C442 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.01fF
C443 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C444 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.01fF
C445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C446 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C447 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# -0.00fF
C448 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C449 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C450 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.01fF
C451 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C452 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C453 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C454 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C455 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.02fF
C456 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C457 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# -0.00fF
C458 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C459 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C460 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C461 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C462 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C463 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C464 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C465 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C466 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C467 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# -0.00fF
C468 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C469 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C470 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C471 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# -0.00fF
C472 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C473 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C474 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C475 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C476 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C477 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C478 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.02fF
C479 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C480 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C481 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C483 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C484 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C485 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C486 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C487 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C488 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C489 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.02fF
C490 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C491 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C492 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.00fF
C493 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C494 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C495 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C496 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# -0.00fF
C497 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# -0.00fF
C498 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C499 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C500 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C501 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C502 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C503 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C504 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C505 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C506 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# -0.00fF
C507 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C508 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C509 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C510 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C511 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C512 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# 0.02fF
C513 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C514 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C515 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C516 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C517 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.01fF
C519 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C520 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C521 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C522 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C523 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C524 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C525 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C526 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C527 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C528 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C529 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C530 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C531 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# -0.00fF
C532 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C533 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C534 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C535 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C536 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# -0.00fF
C537 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C538 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# -0.00fF
C539 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C540 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C541 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C542 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C543 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C544 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C545 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C546 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C547 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C548 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C549 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C550 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C551 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C552 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C553 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C554 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C555 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C556 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C557 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C558 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C559 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C560 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# -0.00fF
C561 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C562 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C563 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C564 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C565 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C566 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C567 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# -0.00fF
C568 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C569 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# 0.00fF
C570 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C571 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C572 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C573 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C574 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C575 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C577 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C578 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C579 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C580 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C581 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.02fF
C582 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C583 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C584 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C585 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C586 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C587 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.01fF
C588 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C589 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C590 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C591 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.44fF
C592 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# -0.00fF
C593 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C594 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C595 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C597 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C598 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C599 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C600 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C601 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C602 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C603 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# -0.00fF
C604 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C605 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C606 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C607 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.93fF
C608 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.01fF
C609 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C610 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C611 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C612 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# -0.00fF
C613 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C614 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C615 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C616 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C617 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C618 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C619 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C620 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C621 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C622 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C623 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C624 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C625 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C626 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C627 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C628 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C629 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C630 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C631 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C632 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C633 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C634 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C635 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C636 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# -0.00fF
C637 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C638 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C639 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C640 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C641 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C642 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C643 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.02fF
C644 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# -0.30fF
C645 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C646 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C647 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C648 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C649 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C650 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C651 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# 0.00fF
C652 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C653 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C654 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C655 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C656 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C657 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C658 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.02fF
C659 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C660 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C661 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C662 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C663 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.02fF
C664 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C665 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.01fF
C666 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C667 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C668 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C669 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C670 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C671 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C672 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# 0.02fF
C673 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C674 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C675 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C677 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# 0.01fF
C678 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C679 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C680 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C681 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.01fF
C682 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# -0.00fF
C683 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C684 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C685 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C686 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C687 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C688 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C689 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.02fF
C690 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C691 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C692 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C693 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# -0.00fF
C694 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C695 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C696 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C697 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.31fF
C698 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C699 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C700 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C701 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C702 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C703 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C704 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C705 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C706 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C707 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C708 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C709 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C710 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# -0.00fF
C711 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.01fF
C712 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C713 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C714 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C715 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.02fF
C716 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C717 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.01fF
C718 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C719 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C720 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C721 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C722 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C723 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C724 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# -0.00fF
C725 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C726 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C727 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C728 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C729 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C730 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.01fF
C731 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C732 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.02fF
C733 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C734 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C735 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C736 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C737 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.01fF
C738 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.02fF
C739 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C740 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C741 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# -0.00fF
C742 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C743 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C744 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C745 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C746 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C747 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C748 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C749 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C750 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.22fF
C751 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C752 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C753 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C754 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C755 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C756 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C757 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C758 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C759 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C760 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C761 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C763 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C764 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C765 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C766 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C767 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C768 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C769 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# -0.00fF
C770 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.00fF
C771 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C772 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C773 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C774 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C775 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C776 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C777 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C778 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C779 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C780 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C781 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C782 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C783 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C784 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C785 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C786 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C787 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C788 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C789 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C790 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C791 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.01fF
C792 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C793 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.01fF
C794 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C795 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C796 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C797 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.01fF
C798 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# 0.01fF
C799 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C800 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.02fF
C801 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.01fF
C802 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C803 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C804 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.02fF
C805 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.01fF
C806 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C807 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C808 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C809 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C810 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C811 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.02fF
C812 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C813 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C814 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C815 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C816 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C817 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C818 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C819 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C820 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C821 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.02fF
C822 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C823 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C824 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C825 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# -0.00fF
C826 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C827 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C828 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C829 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C830 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C831 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C832 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C833 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# -0.00fF
C834 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C835 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C836 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C837 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C838 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C839 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C840 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C841 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C842 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C843 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C844 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C845 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C846 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C847 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C848 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C849 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C850 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C851 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C852 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C853 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C854 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.01fF
C855 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.01fF
C856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C857 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C858 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C859 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C860 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.44fF
C862 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C863 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C864 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C865 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C866 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C867 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C868 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C869 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C870 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C871 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C872 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C873 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.01fF
C874 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.02fF
C875 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C876 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.01fF
C877 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# -0.00fF
C878 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# -0.00fF
C879 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# -0.00fF
C880 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C881 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C882 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C883 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C884 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C885 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C886 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C887 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C888 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C889 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.02fF
C890 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# -0.01fF
C891 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C892 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C893 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C894 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C895 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C896 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C897 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C898 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.01fF
C899 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.02fF
C900 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C901 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C902 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C903 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C904 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.01fF
C905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C906 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C907 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.01fF
C908 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C909 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C910 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C911 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# -0.00fF
C912 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C913 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C914 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C915 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C916 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C917 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C918 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C919 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C920 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C921 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C922 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C923 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C924 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C925 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# -0.00fF
C926 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C927 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C928 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C930 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C931 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C932 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.01fF
C933 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.02fF
C934 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.42fF
C935 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C936 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C937 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# -0.00fF
C938 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C939 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C940 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C941 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C942 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C943 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C944 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C945 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C946 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C947 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C948 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C949 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C950 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C951 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C952 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C953 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.42fF
C954 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C955 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C956 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# -0.00fF
C957 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C958 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C959 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C960 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C961 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C962 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C963 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C964 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C965 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.01fF
C966 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C967 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C968 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.01fF
C969 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.02fF
C970 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C971 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.02fF
C973 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C974 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C975 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.02fF
C976 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C978 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C979 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C980 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C981 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C982 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C983 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.02fF
C984 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C985 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C986 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C987 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C988 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.01fF
C989 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.00fF
C990 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C991 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C992 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C994 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C995 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C996 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C997 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C998 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C999 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1000 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1001 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.00fF
C1002 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1003 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1004 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1006 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C1008 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1009 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1010 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C1011 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1012 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1013 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1014 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1015 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1016 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1017 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C1018 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1019 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1020 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1021 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C1022 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1023 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.01fF
C1024 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.02fF
C1025 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C1026 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.27fF
C1027 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C1028 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C1029 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.02fF
C1030 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1032 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1033 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C1034 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1035 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# -0.00fF
C1036 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1037 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1038 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C1039 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C1040 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1041 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C1042 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1043 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1044 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1045 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1046 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1047 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1048 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1049 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1050 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C1051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1052 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C1053 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C1054 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1055 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1056 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C1057 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1058 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1059 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C1060 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1061 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C1062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C1063 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# 0.01fF
C1064 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C1065 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1066 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C1067 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1068 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1069 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C1070 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1071 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1072 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1073 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1074 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1075 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1077 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.02fF
C1078 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1079 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1081 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1082 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C1083 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1084 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.93fF
C1085 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1086 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1087 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1088 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C1089 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C1090 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1091 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1092 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1093 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1094 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C1095 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1096 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C1097 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1098 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1099 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C1100 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C1101 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C1102 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.02fF
C1103 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C1104 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1105 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C1106 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1107 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1108 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C1109 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1110 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1111 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1112 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1113 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1114 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.02fF
C1115 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# 0.01fF
C1116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1117 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.01fF
C1118 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1119 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1120 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C1121 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1122 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1123 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C1124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1125 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1126 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C1128 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1129 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.01fF
C1130 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1131 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1132 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1133 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1134 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1135 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1136 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1137 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1138 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C1139 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.02fF
C1140 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1141 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C1142 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1143 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1144 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C1145 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1146 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1147 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C1148 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C1149 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C1151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1152 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1153 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# 0.01fF
C1154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1155 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C1156 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C1157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C1158 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1159 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1160 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C1161 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1162 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1163 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1164 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1165 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1166 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1167 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1168 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C1169 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1170 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1171 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1172 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C1173 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1174 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1175 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1176 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1177 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1178 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1179 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C1180 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1181 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1182 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# -0.00fF
C1183 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# -0.00fF
C1184 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1185 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1186 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# -0.00fF
C1187 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C1188 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# -0.00fF
C1189 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1190 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1191 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# -0.00fF
C1192 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C1193 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1194 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# 0.00fF
C1195 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# -0.00fF
C1196 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C1197 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.02fF
C1198 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1199 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1200 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1201 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C1202 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1204 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C1205 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C1206 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1207 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1208 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C1209 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C1210 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1211 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1212 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C1213 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.02fF
C1214 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.02fF
C1215 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1216 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C1217 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1218 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C1219 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1220 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C1221 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C1222 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C1223 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C1224 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C1225 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1226 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C1227 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1228 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C1229 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1230 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1231 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C1232 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1233 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C1234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1235 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1236 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# -0.17fF
C1237 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1238 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C1239 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C1240 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1241 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1242 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.02fF
C1243 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.01fF
C1244 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.01fF
C1245 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1246 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C1247 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1249 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C1250 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1251 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1252 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1253 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C1254 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# -0.00fF
C1255 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1256 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# 0.01fF
C1257 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C1258 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C1259 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1260 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C1261 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1262 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C1263 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1264 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1265 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1266 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.01fF
C1267 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1268 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1269 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1270 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1271 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1272 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C1273 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1274 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1275 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C1276 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C1277 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C1278 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1279 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C1280 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1281 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C1282 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C1283 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C1284 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1285 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1286 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C1287 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1288 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C1289 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1290 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1291 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C1292 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1293 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C1294 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C1295 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.02fF
C1296 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1297 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1298 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1299 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1300 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1301 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C1302 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.48fF
C1303 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# -0.00fF
C1304 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1305 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C1306 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.01fF
C1307 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1308 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1309 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C1310 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1311 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C1312 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# -0.00fF
C1313 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# -0.00fF
C1314 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C1315 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1316 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C1317 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1318 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C1319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C1320 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C1321 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.02fF
C1322 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C1323 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1324 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.02fF
C1325 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C1326 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# -0.01fF
C1327 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.02fF
C1328 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C1329 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C1330 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1331 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.02fF
C1332 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1333 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C1334 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# -0.00fF
C1335 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.02fF
C1336 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# -0.00fF
C1337 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C1338 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1339 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1340 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C1341 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C1342 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# -0.00fF
C1343 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C1344 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.02fF
C1345 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1346 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C1347 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# -0.01fF
C1348 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C1349 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C1350 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C1351 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C1352 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1353 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.01fF
C1354 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.31fF
C1355 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.57fF
C1356 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1357 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# -0.01fF
C1358 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1359 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.01fF
C1360 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C1361 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# -0.00fF
C1362 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.02fF
C1363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1364 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.02fF
C1365 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1366 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1367 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C1368 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1369 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1370 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1371 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C1372 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C1373 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.02fF
C1374 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.19fF
C1375 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C1376 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# -0.01fF
C1377 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# -0.00fF
C1378 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1379 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1380 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C1381 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1382 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# -0.00fF
C1383 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C1384 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.00fF
C1385 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C1386 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1387 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1388 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C1389 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1390 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C1391 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.02fF
C1392 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1393 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C1394 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1395 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1396 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1397 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1398 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1399 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1400 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1401 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1402 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C1403 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C1404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C1405 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C1406 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# -0.00fF
C1407 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C1408 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C1409 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.02fF
C1410 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1411 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.31fF
C1412 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C1413 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C1414 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# -0.00fF
C1415 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1416 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.02fF
C1417 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1418 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1419 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1420 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C1421 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1422 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1423 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C1424 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1425 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C1426 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C1427 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.02fF
C1428 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1429 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.01fF
C1430 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.01fF
C1431 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.01fF
C1432 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1433 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1434 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1435 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C1436 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1437 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.02fF
C1438 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1439 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1440 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C1441 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1442 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1443 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1444 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C1445 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1446 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1447 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1448 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C1449 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1450 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.01fF
C1451 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C1452 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C1453 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1454 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C1455 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.02fF
C1456 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1457 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# -0.00fF
C1458 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.02fF
C1459 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C1460 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1461 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1462 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1463 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C1464 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.02fF
C1465 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.02fF
C1466 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1467 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C1468 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C1469 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C1470 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.01fF
C1471 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1472 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C1473 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1474 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C1475 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1476 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.01fF
C1477 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C1478 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C1479 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1480 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.02fF
C1481 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C1482 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.01fF
C1483 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C1484 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# 0.00fF
C1485 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C1486 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C1487 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1488 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# -0.00fF
C1489 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C1490 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1491 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1492 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1493 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.02fF
C1494 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C1495 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1496 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1497 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.42fF
C1498 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1499 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C1500 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C1501 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C1502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1503 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1504 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C1505 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1506 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C1507 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1508 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C1509 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C1510 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# -0.00fF
C1511 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1512 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.02fF
C1513 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1514 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1515 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1516 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1517 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1518 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C1519 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# -0.01fF
C1520 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# -0.00fF
C1521 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1522 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1523 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1524 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1525 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C1526 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1527 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C1528 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C1529 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1530 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.02fF
C1531 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C1532 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.01fF
C1533 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C1534 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C1535 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C1536 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C1537 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.02fF
C1538 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1539 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C1540 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.01fF
C1541 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1542 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1543 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C1544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C1545 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C1546 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.02fF
C1547 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.02fF
C1548 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C1549 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1550 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1551 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.02fF
C1552 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1553 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1554 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C1555 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1556 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.02fF
C1557 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1558 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# -0.00fF
C1559 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.01fF
C1560 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1561 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.02fF
C1562 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1563 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C1564 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1565 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.02fF
C1566 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C1567 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1568 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C1569 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1570 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1571 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C1572 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.24fF
C1573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1574 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1576 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1577 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1578 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C1579 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1580 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# -0.00fF
C1581 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C1582 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C1583 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C1584 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1585 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1586 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C1587 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# -0.00fF
C1588 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C1589 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1590 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1591 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1592 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C1593 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C1594 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1595 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C1596 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C1597 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C1598 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C1599 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C1600 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# -0.00fF
C1601 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.01fF
C1602 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1603 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1604 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1605 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1606 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C1607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C1608 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1609 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1610 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1611 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1612 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1613 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C1614 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1615 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C1616 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1617 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1618 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1619 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1620 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1621 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.02fF
C1623 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1624 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1625 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1626 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1627 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.02fF
C1628 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C1629 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C1630 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# -0.00fF
C1631 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.01fF
C1632 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1633 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1634 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1635 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1636 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C1637 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1638 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C1639 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 1.18fF
C1640 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C1641 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1642 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# -0.00fF
C1643 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C1644 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1645 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1646 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1647 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1648 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.02fF
C1649 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# 0.02fF
C1650 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1651 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1652 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C1653 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C1654 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1655 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# -0.00fF
C1656 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1657 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1658 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1659 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C1660 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C1661 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# -0.00fF
C1662 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C1663 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1664 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1665 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1666 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C1667 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.02fF
C1668 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C1669 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.02fF
C1670 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1671 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C1672 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1673 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C1674 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1675 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C1676 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.02fF
C1677 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1678 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1679 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1680 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1681 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C1682 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C1683 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C1684 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# -0.00fF
C1685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C1686 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1687 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C1688 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1689 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1690 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1691 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C1692 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C1693 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C1694 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C1695 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C1696 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.42fF
C1697 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C1698 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C1699 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C1700 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C1701 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1702 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1703 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C1704 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C1705 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1706 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C1707 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C1708 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C1709 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C1710 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C1711 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# -0.00fF
C1712 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C1713 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.02fF
C1714 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C1715 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1716 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C1717 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C1718 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C1719 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C1720 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C1721 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1722 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.02fF
C1723 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.01fF
C1724 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C1725 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C1726 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C1727 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1728 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.01fF
C1729 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1730 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C1731 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1732 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C1733 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1734 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1735 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1736 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C1737 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1738 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C1739 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1740 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.02fF
C1741 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# -0.00fF
C1742 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1743 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1744 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1745 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C1746 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.02fF
C1747 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1748 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C1749 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C1750 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.02fF
C1751 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1752 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.02fF
C1753 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C1754 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1755 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1756 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C1757 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C1758 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.01fF
C1759 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1760 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1761 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C1762 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C1763 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C1764 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C1765 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.01fF
C1766 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1767 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C1768 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1769 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1770 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C1771 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C1772 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C1773 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# -0.00fF
C1774 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C1775 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1776 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C1777 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C1778 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.01fF
C1779 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.02fF
C1780 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.00fF
C1781 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1782 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C1783 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# -0.00fF
C1784 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C1785 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C1786 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# 0.01fF
C1787 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.00fF
C1788 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C1789 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C1790 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# -0.00fF
C1791 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C1792 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C1793 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1794 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1795 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.01fF
C1796 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C1797 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1798 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C1799 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1800 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1801 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1802 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C1803 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C1804 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.00fF
C1805 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C1806 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C1807 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# 0.00fF
C1808 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.02fF
C1809 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C1810 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1811 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.00fF
C1812 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C1813 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C1814 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1815 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C1816 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C1817 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# -0.00fF
C1818 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C1819 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C1820 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C1821 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1822 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# -0.00fF
C1823 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C1824 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1825 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1826 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1827 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1828 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1829 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1830 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C1831 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C1832 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1833 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C1834 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1835 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C1836 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C1837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C1838 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.02fF
C1839 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# -0.01fF
C1840 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C1841 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C1842 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C1843 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1844 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C1845 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C1846 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C1847 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C1848 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C1849 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C1850 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1851 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.01fF
C1852 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C1853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1854 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C1855 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1857 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.02fF
C1858 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.01fF
C1859 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1860 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1861 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C1862 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C1863 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C1864 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1865 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1866 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C1867 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C1868 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.02fF
C1869 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.01fF
C1870 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C1871 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1872 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C1873 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C1874 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C1875 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1876 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C1877 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# -0.00fF
C1878 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1879 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C1880 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1881 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1882 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C1883 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C1884 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C1885 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C1886 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C1887 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C1888 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C1889 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.02fF
C1890 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.01fF
C1891 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C1892 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# -0.01fF
C1893 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1894 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1895 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1896 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1897 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C1898 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1899 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C1900 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C1901 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C1902 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1903 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C1904 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C1905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C1906 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C1907 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C1908 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C1909 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C1910 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C1911 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C1912 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.19fF
C1913 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# -0.00fF
C1914 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C1915 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1916 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1917 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1918 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C1919 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C1920 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.01fF
C1921 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# -0.00fF
C1922 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C1923 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1924 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.01fF
C1925 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C1926 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C1927 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C1928 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C1929 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1930 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# -0.00fF
C1931 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C1932 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C1933 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1934 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1935 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1936 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C1937 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C1938 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C1939 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.02fF
C1940 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C1941 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1942 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C1943 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1944 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C1945 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C1946 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C1947 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1948 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1949 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C1950 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C1951 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1952 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C1954 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C1955 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1956 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C1957 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C1958 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# -0.00fF
C1959 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C1960 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C1961 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1962 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C1963 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# -0.00fF
C1964 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1965 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C1966 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C1967 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C1968 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.02fF
C1969 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1970 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C1971 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C1973 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C1974 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1975 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.01fF
C1976 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C1977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C1978 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C1979 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C1980 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C1981 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C1982 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C1983 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C1984 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C1985 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C1986 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C1987 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C1988 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C1989 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C1990 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C1991 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C1992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C1993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C1994 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C1995 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C1996 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C1997 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C1998 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C1999 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C2000 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.02fF
C2001 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C2002 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2003 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2004 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.02fF
C2005 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C2006 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C2007 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# -0.00fF
C2008 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C2009 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C2010 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2011 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C2012 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C2013 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C2014 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2015 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C2016 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2017 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2018 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C2019 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.01fF
C2020 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2021 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.02fF
C2022 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C2023 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2024 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2025 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C2026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# -0.00fF
C2027 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.01fF
C2028 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.02fF
C2029 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2030 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C2031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2032 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C2033 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2034 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.01fF
C2035 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2036 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C2037 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.02fF
C2038 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2039 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C2040 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C2041 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C2042 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# -0.00fF
C2043 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# -0.00fF
C2044 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C2045 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2046 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2047 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C2048 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2049 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2050 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.01fF
C2051 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C2052 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C2053 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.02fF
C2054 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C2055 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.44fF
C2056 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2057 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2058 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2059 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C2060 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C2061 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2062 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C2063 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C2064 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2065 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C2066 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2067 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.01fF
C2068 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C2069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.01fF
C2070 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# -0.00fF
C2071 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2072 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# -0.00fF
C2073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C2074 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C2075 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C2076 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2077 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C2078 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.02fF
C2079 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C2080 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C2081 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C2082 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# -0.00fF
C2083 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2084 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C2085 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C2086 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C2087 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C2088 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C2089 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.01fF
C2090 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C2091 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2092 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2093 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2094 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.44fF
C2095 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2096 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C2097 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.02fF
C2098 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2099 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2100 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C2101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C2102 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# -0.00fF
C2103 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C2104 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2105 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C2106 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C2107 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2108 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C2109 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C2110 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C2111 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C2112 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# -0.00fF
C2113 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C2114 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# -0.00fF
C2115 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C2116 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C2117 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# -0.00fF
C2118 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C2119 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2120 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C2121 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C2122 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C2123 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# -0.00fF
C2124 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C2125 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C2126 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C2127 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2128 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2129 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C2130 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.01fF
C2131 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C2132 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C2133 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2134 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2135 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C2136 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C2138 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C2139 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# -0.00fF
C2140 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C2141 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.01fF
C2142 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# -0.00fF
C2143 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C2144 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.01fF
C2145 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.01fF
C2146 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2147 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2148 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C2149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C2150 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C2151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C2152 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C2153 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.01fF
C2154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C2155 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C2156 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2157 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2158 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2159 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.01fF
C2160 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C2161 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# -0.00fF
C2162 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C2163 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2164 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C2165 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2166 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C2167 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.01fF
C2168 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2169 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C2170 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.00fF
C2171 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.01fF
C2172 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C2173 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C2174 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C2175 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2176 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# -0.00fF
C2177 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C2178 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.02fF
C2179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C2180 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C2181 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2182 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.01fF
C2183 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.01fF
C2184 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# -0.00fF
C2185 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# -0.01fF
C2186 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2187 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C2188 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C2189 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2190 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2191 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C2192 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2193 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C2194 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C2195 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C2196 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2197 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2198 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.01fF
C2199 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2200 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C2201 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# -0.00fF
C2202 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C2203 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C2204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2205 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.01fF
C2206 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C2207 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2208 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2209 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C2210 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C2211 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2212 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# -0.00fF
C2213 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2214 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2215 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2216 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C2217 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.57fF
C2218 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.02fF
C2219 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C2220 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C2221 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# -0.01fF
C2222 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.00fF
C2223 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C2224 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C2225 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C2226 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# -0.00fF
C2227 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C2228 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2229 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C2230 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.02fF
C2231 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2232 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C2233 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C2234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C2235 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C2236 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2237 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C2238 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2239 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2240 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2241 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2242 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C2243 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C2244 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2245 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C2246 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# -0.00fF
C2247 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C2248 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2249 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2250 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C2251 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2252 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2253 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C2254 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C2255 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C2256 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.01fF
C2257 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C2258 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2259 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2260 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C2261 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2262 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2263 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# -0.01fF
C2264 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2265 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C2266 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C2267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C2268 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C2269 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C2270 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2271 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2272 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C2273 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C2274 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C2275 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C2276 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C2277 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2278 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2279 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2280 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2281 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C2283 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.01fF
C2284 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2285 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.01fF
C2286 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C2287 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.02fF
C2288 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C2289 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# -0.00fF
C2290 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# -0.00fF
C2291 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C2292 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2293 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C2294 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2295 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C2296 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2297 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# -0.01fF
C2298 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C2299 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C2300 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# -0.00fF
C2301 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C2302 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C2303 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C2304 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C2305 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C2306 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2307 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2308 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2309 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C2310 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2311 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# -0.00fF
C2312 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2313 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C2314 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C2315 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2316 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C2317 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C2318 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2319 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C2320 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C2321 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C2322 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.02fF
C2323 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.02fF
C2324 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C2325 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C2326 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C2327 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.01fF
C2328 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# 0.02fF
C2329 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C2330 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2331 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2332 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C2333 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C2334 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2335 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.01fF
C2336 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2337 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C2338 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C2339 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2340 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2341 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2342 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C2343 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C2344 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C2345 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2346 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2347 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C2348 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.00fF
C2349 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C2350 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2351 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2352 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2353 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.01fF
C2354 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2355 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# -0.00fF
C2356 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C2357 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.02fF
C2358 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.02fF
C2359 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.02fF
C2360 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.02fF
C2361 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C2362 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2363 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.02fF
C2364 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2365 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2366 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.01fF
C2367 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2368 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C2369 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2370 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2371 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2372 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C2373 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C2374 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# -0.00fF
C2375 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.01fF
C2376 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C2377 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2378 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.01fF
C2379 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C2380 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2381 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.01fF
C2382 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.01fF
C2383 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2384 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2385 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C2386 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C2387 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2389 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2390 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.01fF
C2391 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2392 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2393 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2394 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2395 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2396 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2397 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C2398 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2399 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2400 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.00fF
C2401 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.02fF
C2402 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C2403 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.00fF
C2404 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.22fF
C2405 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2406 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.01fF
C2407 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.01fF
C2408 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2409 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.02fF
C2410 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C2411 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C2412 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.01fF
C2413 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2414 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C2415 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C2416 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2417 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2418 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C2419 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2420 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C2421 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C2422 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C2423 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2424 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2425 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.02fF
C2426 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C2427 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2428 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2429 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# -0.00fF
C2430 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2431 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C2432 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C2433 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C2434 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2435 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2436 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2437 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C2438 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2439 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.02fF
C2440 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# -0.00fF
C2441 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.02fF
C2442 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2443 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2444 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C2445 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2446 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 1.18fF
C2447 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C2448 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C2449 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C2450 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C2451 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2452 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C2453 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C2454 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2455 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.48fF
C2456 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2457 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C2458 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2459 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2460 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C2461 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C2462 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C2463 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2464 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.02fF
C2465 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.01fF
C2466 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2467 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C2468 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C2469 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2470 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2471 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C2472 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C2473 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C2474 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.01fF
C2475 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2476 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2477 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2478 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2479 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C2480 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C2481 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2482 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2483 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C2484 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2485 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# 0.01fF
C2486 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C2487 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.01fF
C2488 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.01fF
C2489 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C2490 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.01fF
C2491 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C2492 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2493 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C2494 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C2495 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# -0.00fF
C2496 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2497 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2498 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C2499 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C2500 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2501 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2502 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2503 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2504 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C2505 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C2506 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2507 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.44fF
C2508 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# -0.00fF
C2509 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# -0.00fF
C2510 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C2511 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2512 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C2513 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2514 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C2515 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C2516 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C2517 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2518 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C2519 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C2520 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C2521 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C2522 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2523 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2524 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# 0.01fF
C2525 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2526 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C2527 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2528 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C2529 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.01fF
C2530 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C2531 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.01fF
C2532 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2533 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2534 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2535 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# 0.01fF
C2536 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.00fF
C2537 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C2538 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# -0.00fF
C2539 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.01fF
C2540 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2541 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2542 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# 0.01fF
C2543 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C2544 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C2545 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C2546 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C2547 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.02fF
C2548 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C2549 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2550 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C2551 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# -0.00fF
C2552 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C2553 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2554 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C2555 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2556 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2557 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.01fF
C2558 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.00fF
C2559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2560 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.01fF
C2561 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2562 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2563 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C2564 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C2565 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2566 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C2567 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C2568 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C2569 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# -0.00fF
C2570 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C2571 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C2572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.01fF
C2573 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C2574 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C2575 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# 0.01fF
C2576 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C2577 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# -0.00fF
C2578 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# -0.00fF
C2579 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2580 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C2581 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C2582 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C2583 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2584 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C2585 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2586 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C2587 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# -0.00fF
C2588 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2589 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C2590 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C2591 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2592 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2593 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2594 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C2595 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2596 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2597 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C2598 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2599 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C2600 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C2601 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C2602 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.02fF
C2603 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C2604 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C2605 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2606 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C2607 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.01fF
C2608 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2609 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.01fF
C2610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2611 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# -0.00fF
C2612 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.02fF
C2613 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2614 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2615 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C2616 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C2617 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2618 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.00fF
C2619 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2620 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C2621 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C2622 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.01fF
C2623 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# -0.00fF
C2624 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2625 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2626 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C2627 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2628 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.02fF
C2629 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.02fF
C2630 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C2631 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2632 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2633 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C2634 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2635 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2636 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2637 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C2638 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2639 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C2640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C2641 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2642 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2643 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.00fF
C2644 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.01fF
C2645 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C2646 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C2647 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.57fF
C2648 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2649 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C2650 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C2651 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C2652 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C2653 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C2654 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C2655 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2656 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.02fF
C2657 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2658 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C2659 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2660 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# -0.00fF
C2661 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2662 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.01fF
C2663 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C2664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# 0.00fF
C2665 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C2666 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C2667 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2668 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2669 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C2670 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C2671 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.93fF
C2672 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2673 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.19fF
C2674 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C2675 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C2676 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.01fF
C2677 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.01fF
C2678 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C2679 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C2680 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2681 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# -0.00fF
C2682 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C2683 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2684 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.02fF
C2685 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C2686 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# -0.00fF
C2687 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C2688 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# -0.00fF
C2689 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C2690 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.02fF
C2691 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C2692 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C2693 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.02fF
C2694 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2695 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C2696 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.01fF
C2697 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2698 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C2699 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C2700 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2701 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C2702 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2703 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2704 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2705 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2706 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C2707 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# -0.00fF
C2708 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.01fF
C2709 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C2710 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C2711 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2712 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2713 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.02fF
C2714 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.01fF
C2715 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2716 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2717 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C2718 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C2719 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C2720 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2721 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C2722 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C2723 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C2724 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C2725 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2726 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C2727 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2728 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.46fF
C2729 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2730 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C2731 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C2732 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C2733 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C2734 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C2735 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2736 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C2737 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2738 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C2739 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C2740 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2741 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2742 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C2743 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C2744 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2745 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2746 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C2747 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C2748 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C2749 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2750 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C2751 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C2752 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2753 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2754 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# -0.00fF
C2755 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2756 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2757 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2758 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C2759 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C2760 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C2761 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C2762 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C2763 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C2764 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.93fF
C2765 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2766 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2767 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.01fF
C2768 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.02fF
C2769 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2770 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2771 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2772 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.01fF
C2773 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.01fF
C2774 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C2775 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2776 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2777 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C2778 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# -0.00fF
C2779 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C2780 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.02fF
C2781 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C2782 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C2783 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.02fF
C2784 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.01fF
C2785 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C2786 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# -0.00fF
C2787 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.19fF
C2788 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2789 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C2790 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.01fF
C2791 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.02fF
C2792 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2793 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2794 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.01fF
C2795 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C2796 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# 0.02fF
C2797 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C2798 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2799 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# 0.02fF
C2800 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C2801 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C2802 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2803 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C2804 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C2805 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2806 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C2807 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.01fF
C2808 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.01fF
C2809 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C2810 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.02fF
C2811 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.02fF
C2812 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2813 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C2814 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C2815 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C2816 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# -0.00fF
C2817 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.01fF
C2818 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C2819 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C2820 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2821 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2822 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2823 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.02fF
C2824 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# -0.00fF
C2825 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2826 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.01fF
C2827 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.02fF
C2828 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2830 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C2831 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# -0.00fF
C2832 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.01fF
C2833 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C2834 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C2835 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C2836 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C2838 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# -0.00fF
C2839 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.01fF
C2840 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C2841 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C2842 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C2843 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2844 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C2845 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C2846 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C2847 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2848 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C2849 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.02fF
C2850 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C2851 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C2852 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C2853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C2854 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C2855 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2856 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2857 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2858 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2859 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# -0.00fF
C2860 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# -0.00fF
C2861 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C2862 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2863 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C2864 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C2865 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C2866 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C2867 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C2868 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# -0.00fF
C2869 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C2870 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.02fF
C2871 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C2872 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2873 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2874 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2875 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C2876 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C2877 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2878 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2879 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# -0.00fF
C2880 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.00fF
C2881 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.01fF
C2882 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C2883 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C2884 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C2885 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2886 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C2887 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C2888 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C2889 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2890 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# -0.00fF
C2891 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# -0.00fF
C2892 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C2893 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C2894 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.01fF
C2895 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2896 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C2897 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.93fF
C2898 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2899 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C2900 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2901 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2902 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C2903 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C2904 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.01fF
C2905 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.02fF
C2906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C2907 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C2908 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C2909 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C2910 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.01fF
C2911 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.00fF
C2912 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C2913 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C2914 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C2915 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C2916 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C2917 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2918 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.02fF
C2919 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C2920 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C2921 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.02fF
C2922 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.02fF
C2923 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2924 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C2925 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C2926 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C2927 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.01fF
C2928 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.01fF
C2929 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C2930 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2931 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# 0.00fF
C2932 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C2933 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2934 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C2935 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2936 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C2937 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C2938 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C2939 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C2940 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C2941 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2942 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.02fF
C2943 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C2944 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.02fF
C2945 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C2946 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C2947 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C2948 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C2949 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# -0.00fF
C2950 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C2951 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C2952 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C2953 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2954 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C2955 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C2956 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2957 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# 0.00fF
C2958 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C2959 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2960 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C2961 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2962 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C2963 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2964 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.42fF
C2965 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C2966 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2967 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C2968 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2969 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.02fF
C2970 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C2971 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C2972 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2973 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C2974 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2975 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.01fF
C2976 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.02fF
C2977 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C2978 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2979 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2980 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C2981 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C2982 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.01fF
C2983 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2984 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C2985 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C2986 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C2987 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C2988 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C2989 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C2990 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C2991 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.22fF
C2992 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C2993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C2994 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C2995 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C2996 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C2997 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C2998 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C2999 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3000 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3001 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.01fF
C3002 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# 0.00fF
C3003 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.00fF
C3004 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3005 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C3006 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3008 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3009 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3010 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3011 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C3012 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C3013 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3014 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.22fF
C3015 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3016 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.01fF
C3017 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C3018 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3019 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.00fF
C3020 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.02fF
C3022 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3023 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C3024 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.01fF
C3025 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3026 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3027 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C3028 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3029 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# -0.00fF
C3030 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# -0.00fF
C3031 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3032 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C3033 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3034 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C3035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C3036 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3037 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3038 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3039 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3040 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.02fF
C3041 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C3042 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3043 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3044 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C3045 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C3046 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.01fF
C3047 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C3048 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3049 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3050 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C3051 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3052 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3053 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3054 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C3055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# -0.00fF
C3056 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3057 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.31fF
C3058 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C3059 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3060 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3061 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.02fF
C3063 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.01fF
C3064 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3065 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3066 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# -0.00fF
C3067 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3068 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.00fF
C3069 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C3070 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C3071 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C3072 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3073 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# -0.00fF
C3074 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C3075 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3076 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.02fF
C3077 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.00fF
C3078 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.42fF
C3079 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3080 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3081 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.02fF
C3082 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C3083 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C3084 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3085 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3086 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.02fF
C3087 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3088 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3089 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3090 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.00fF
C3091 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3092 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C3093 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C3094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C3095 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3096 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3097 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3098 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3099 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3100 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.01fF
C3101 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.02fF
C3102 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C3103 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C3104 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# -0.00fF
C3105 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3106 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3107 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3108 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3109 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3110 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3111 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3112 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.01fF
C3113 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3114 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3115 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.93fF
C3116 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3117 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3118 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C3119 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3120 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# -0.00fF
C3121 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C3122 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C3123 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3124 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3125 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3126 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C3127 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3128 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3129 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3130 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C3131 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C3132 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C3133 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C3134 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3135 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.44fF
C3136 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3137 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3138 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C3139 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3140 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3141 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C3142 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 1.18fF
C3143 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.02fF
C3144 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3145 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3146 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3147 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3148 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C3149 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C3150 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C3151 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3152 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3153 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3154 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.02fF
C3155 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3156 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3157 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3158 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3159 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C3160 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3161 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C3162 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C3163 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C3164 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3165 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.02fF
C3166 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.01fF
C3167 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3168 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# -0.00fF
C3170 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C3171 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.00fF
C3172 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C3173 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3174 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C3175 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3176 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C3177 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# -0.00fF
C3178 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.02fF
C3179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3180 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3181 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C3182 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3183 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C3184 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.01fF
C3185 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3186 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.02fF
C3187 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3188 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C3189 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C3190 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.02fF
C3191 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3192 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3193 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C3194 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3195 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3196 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3197 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.02fF
C3198 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3199 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C3200 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3201 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C3202 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C3203 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3204 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.01fF
C3205 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.02fF
C3206 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3207 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.00fF
C3208 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C3209 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C3210 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.01fF
C3211 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3212 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C3213 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C3214 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3215 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3216 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3217 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3218 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3219 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3220 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3221 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3222 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3223 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.01fF
C3224 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# -0.00fF
C3225 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3226 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3227 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C3228 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.01fF
C3229 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3230 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3231 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C3232 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C3233 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3234 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C3235 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.02fF
C3236 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3237 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3238 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3239 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3240 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3241 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3242 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C3243 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C3244 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# -0.00fF
C3245 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# -0.00fF
C3246 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3247 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# 0.01fF
C3248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3249 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3250 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3251 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C3252 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.01fF
C3253 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.02fF
C3254 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.00fF
C3255 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.01fF
C3256 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C3257 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C3258 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C3259 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3260 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C3261 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# -0.00fF
C3262 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3263 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C3264 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.02fF
C3265 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3266 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3267 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.01fF
C3268 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3269 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# -0.00fF
C3270 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C3271 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3272 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C3273 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C3274 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C3275 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.02fF
C3276 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C3277 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.01fF
C3278 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# -0.01fF
C3279 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3280 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C3281 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C3282 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.02fF
C3283 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3284 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C3285 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C3286 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C3287 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3288 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# -0.00fF
C3289 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# -0.00fF
C3290 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3291 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3292 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C3293 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.02fF
C3294 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3295 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C3296 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C3297 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C3298 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3299 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C3300 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3301 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3302 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.02fF
C3303 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C3304 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C3305 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3306 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C3307 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C3308 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.02fF
C3309 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C3310 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3311 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3312 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C3313 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3314 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C3315 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3316 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3317 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C3318 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3319 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3320 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C3321 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3322 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3323 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3324 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.02fF
C3325 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C3326 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3327 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C3328 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C3329 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3330 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C3331 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C3332 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C3333 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3334 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3335 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3336 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3337 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# 0.01fF
C3338 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C3339 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3340 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# 0.01fF
C3341 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3342 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C3343 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.01fF
C3344 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3345 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C3346 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3347 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C3348 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.00fF
C3349 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# -0.00fF
C3350 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3351 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# -0.00fF
C3352 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.01fF
C3353 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3354 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C3355 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3356 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C3357 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3358 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C3359 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C3360 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# 0.00fF
C3361 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.01fF
C3362 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C3363 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C3364 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# -0.00fF
C3365 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C3366 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3367 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3368 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3369 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C3370 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C3371 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3372 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3373 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C3374 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3375 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# -0.00fF
C3376 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C3377 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C3378 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C3379 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# 0.00fF
C3380 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3381 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3382 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C3383 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.01fF
C3384 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3385 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.01fF
C3386 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# 0.00fF
C3387 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3388 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C3389 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# 0.01fF
C3390 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3391 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.01fF
C3392 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C3393 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3394 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C3395 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3396 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3397 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# -0.00fF
C3398 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C3399 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3400 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3401 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3402 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.02fF
C3403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3404 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.01fF
C3405 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3406 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.02fF
C3407 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C3408 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3409 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C3410 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.02fF
C3411 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3412 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# -0.01fF
C3413 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C3414 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C3415 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.02fF
C3416 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3417 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# 0.00fF
C3418 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C3419 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3420 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C3421 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# -0.00fF
C3422 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.01fF
C3423 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3424 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C3425 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.27fF
C3426 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# 0.00fF
C3427 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3428 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3429 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3430 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# -0.00fF
C3431 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C3432 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C3433 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3434 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C3435 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C3436 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C3437 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C3438 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C3439 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C3440 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.01fF
C3441 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C3442 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C3443 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3444 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3445 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# -0.00fF
C3446 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C3447 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C3448 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C3449 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3450 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.02fF
C3451 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C3452 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3453 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3454 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3455 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C3456 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3457 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3458 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C3459 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3460 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3461 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.01fF
C3462 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3463 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3464 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C3465 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C3466 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C3467 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3468 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C3469 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# 0.00fF
C3470 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3471 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C3472 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C3473 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.00fF
C3474 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3475 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.01fF
C3476 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.01fF
C3477 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.02fF
C3478 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3479 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3480 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C3481 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3482 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.01fF
C3483 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3484 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3485 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3486 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3487 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C3488 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# 0.01fF
C3489 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.02fF
C3490 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C3491 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.00fF
C3492 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# -0.00fF
C3493 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3494 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C3495 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3496 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3497 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C3498 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3499 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# -0.00fF
C3500 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.01fF
C3501 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3502 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3503 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C3504 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3505 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3506 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.01fF
C3507 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C3508 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C3509 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# -0.00fF
C3510 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3511 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C3512 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C3513 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3514 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C3515 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3516 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3517 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C3518 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3519 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.01fF
C3520 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C3521 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3522 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C3523 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.01fF
C3524 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C3525 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C3526 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3527 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# -0.00fF
C3528 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.27fF
C3529 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C3530 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# -0.00fF
C3531 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C3532 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# -0.00fF
C3533 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3534 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# -0.00fF
C3535 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C3536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3537 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# -0.00fF
C3538 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C3539 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.01fF
C3540 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.57fF
C3541 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C3542 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# 0.00fF
C3543 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3544 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C3545 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C3546 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C3547 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C3548 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3549 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3550 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# -0.00fF
C3551 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C3552 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.02fF
C3553 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C3554 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3555 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C3556 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.01fF
C3557 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C3558 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# -0.00fF
C3559 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C3560 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C3561 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3562 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C3563 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3564 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# -0.00fF
C3565 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.01fF
C3566 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.00fF
C3567 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3568 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.01fF
C3569 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3570 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# 0.01fF
C3571 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.02fF
C3572 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# -0.00fF
C3573 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.02fF
C3574 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.02fF
C3575 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C3576 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3577 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C3578 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3579 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C3580 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3581 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.00fF
C3582 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3583 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C3584 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.02fF
C3585 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.01fF
C3586 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.01fF
C3587 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C3588 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# -0.00fF
C3589 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C3590 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C3591 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3592 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C3593 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C3594 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.02fF
C3595 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C3596 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3597 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3598 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C3599 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C3600 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C3601 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.01fF
C3602 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3603 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C3604 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.02fF
C3605 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C3606 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C3607 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# -0.00fF
C3608 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3609 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.00fF
C3610 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3611 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3612 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# -0.00fF
C3613 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C3614 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3615 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3616 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C3617 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3618 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C3619 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3620 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C3621 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C3622 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C3623 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C3624 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C3625 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C3626 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.00fF
C3627 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3628 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3629 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C3630 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C3631 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.02fF
C3632 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C3633 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# -0.00fF
C3634 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# 0.00fF
C3635 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3636 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.01fF
C3637 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C3638 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3639 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.02fF
C3640 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3641 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3642 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C3643 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# 0.02fF
C3644 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# 0.00fF
C3645 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3646 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.01fF
C3647 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3648 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C3649 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C3650 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.27fF
C3651 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3652 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3653 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3654 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.01fF
C3655 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3656 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3657 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3658 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C3659 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C3660 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3661 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.02fF
C3662 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3663 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3664 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# 0.00fF
C3665 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3666 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3667 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3668 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3669 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.01fF
C3670 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3671 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# 0.00fF
C3672 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.01fF
C3673 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C3674 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C3675 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C3676 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.02fF
C3677 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C3678 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.01fF
C3679 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# -0.00fF
C3680 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C3681 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3682 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# -0.00fF
C3683 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3684 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3685 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C3686 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.02fF
C3687 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.01fF
C3688 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.00fF
C3689 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.00fF
C3690 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C3691 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.02fF
C3692 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3693 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3694 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C3695 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.01fF
C3696 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.02fF
C3697 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C3698 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3699 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C3700 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C3701 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C3702 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3703 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.00fF
C3704 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C3705 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.01fF
C3706 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C3707 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.42fF
C3708 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3709 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C3710 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C3711 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# 0.00fF
C3712 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3713 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C3714 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.02fF
C3715 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.01fF
C3716 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3717 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C3718 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3719 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# 0.01fF
C3720 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3721 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3722 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.00fF
C3723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C3724 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C3725 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C3726 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.00fF
C3727 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C3728 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3729 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3730 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.00fF
C3731 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C3732 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.01fF
C3733 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C3734 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C3735 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C3736 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3737 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C3738 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.01fF
C3739 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3740 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C3741 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C3742 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.02fF
C3743 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.00fF
C3744 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C3745 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3746 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3747 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C3748 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# 0.00fF
C3749 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C3750 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C3751 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C3752 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# 0.02fF
C3753 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.02fF
C3754 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3755 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C3756 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 1.18fF
C3757 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C3758 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.00fF
C3759 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C3760 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C3761 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3762 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C3763 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C3764 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3765 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C3766 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C3767 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C3768 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3769 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3770 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3771 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# 0.00fF
C3772 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.02fF
C3773 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C3774 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.27fF
C3775 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C3776 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.42fF
C3777 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3778 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3779 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3780 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C3781 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.01fF
C3782 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.02fF
C3783 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.00fF
C3784 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C3785 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.02fF
C3786 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C3787 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C3788 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3789 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.00fF
C3790 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C3791 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# 0.02fF
C3792 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C3793 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.01fF
C3794 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.02fF
C3795 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3796 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3797 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3798 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3799 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# -0.00fF
C3800 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C3801 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3802 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.01fF
C3803 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3804 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.01fF
C3805 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.01fF
C3806 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C3807 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C3808 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3809 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.00fF
C3810 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# -0.00fF
C3811 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# -0.00fF
C3812 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# -0.00fF
C3813 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# 0.00fF
C3814 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C3815 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3816 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C3817 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C3818 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C3819 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C3820 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.00fF
C3821 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C3822 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3823 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.02fF
C3824 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C3825 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3826 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3827 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C3828 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# 0.00fF
C3829 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3830 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.02fF
C3831 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.00fF
C3832 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3833 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3834 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C3835 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C3836 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3837 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C3838 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3839 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3840 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C3841 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# 0.00fF
C3842 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C3843 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.02fF
C3844 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C3845 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.00fF
C3846 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C3847 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C3848 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3849 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# 0.01fF
C3850 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.02fF
C3851 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.01fF
C3852 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# 0.00fF
C3853 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C3854 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C3855 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C3856 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C3857 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C3858 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# 0.00fF
C3859 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3860 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C3861 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3862 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3863 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C3864 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# 0.02fF
C3865 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C3866 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.01fF
C3867 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.02fF
C3868 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C3869 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3870 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3871 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# -0.00fF
C3872 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C3873 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# 0.01fF
C3874 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3875 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C3876 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C3877 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C3878 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.93fF
C3879 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3880 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C3881 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.01fF
C3882 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C3883 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3884 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C3885 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3886 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C3887 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3888 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3889 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C3890 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.00fF
C3891 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3892 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.02fF
C3893 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C3894 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.01fF
C3895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3896 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C3897 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3898 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3899 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3900 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.02fF
C3901 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C3902 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C3903 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3904 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.02fF
C3905 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# 0.00fF
C3906 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C3907 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.01fF
C3908 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3909 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C3910 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C3911 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# -0.00fF
C3912 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C3913 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C3914 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# 0.00fF
C3915 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# -0.00fF
C3916 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.00fF
C3917 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.01fF
C3918 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# 0.02fF
C3919 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3920 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3921 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C3922 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.01fF
C3923 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3924 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3925 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3926 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# -0.00fF
C3927 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3928 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# 0.00fF
C3929 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C3930 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.01fF
C3931 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3932 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C3933 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3934 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C3935 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3936 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C3937 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3938 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C3939 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.42fF
C3940 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3941 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# 0.01fF
C3942 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C3943 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C3944 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C3945 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C3946 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.01fF
C3947 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# -0.00fF
C3948 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.01fF
C3949 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.42fF
C3950 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C3951 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# -0.00fF
C3952 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.00fF
C3953 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C3954 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C3955 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3956 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.02fF
C3957 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# 0.02fF
C3958 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C3959 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3960 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.00fF
C3961 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.00fF
C3962 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C3963 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3964 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.01fF
C3965 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C3966 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.01fF
C3967 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C3968 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C3969 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3970 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C3971 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.02fF
C3972 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C3973 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C3974 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.02fF
C3975 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C3976 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C3977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3978 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# 0.00fF
C3979 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# -0.01fF
C3980 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# -0.00fF
C3981 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C3982 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C3983 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.01fF
C3984 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C3985 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3986 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3987 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.01fF
C3988 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3989 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C3990 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C3991 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C3992 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C3993 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C3994 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C3995 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.01fF
C3996 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C3997 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C3998 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C3999 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4000 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4001 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4002 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C4003 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C4004 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C4006 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.27fF
C4007 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C4008 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.93fF
C4009 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4010 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4011 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4012 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C4013 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4014 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# 0.00fF
C4015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4016 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4017 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.02fF
C4018 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4019 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4020 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4021 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4022 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.00fF
C4023 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C4024 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C4025 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4027 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# -0.00fF
C4028 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4029 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# 0.00fF
C4030 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4031 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.00fF
C4032 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4033 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# -0.00fF
C4034 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4035 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4036 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C4037 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C4038 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4039 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4040 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.02fF
C4041 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C4042 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4043 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.01fF
C4044 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# -0.00fF
C4045 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.01fF
C4046 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4047 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4048 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C4049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# 0.02fF
C4050 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C4051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C4052 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C4053 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# 0.00fF
C4054 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.01fF
C4055 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.02fF
C4056 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4057 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.00fF
C4058 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4060 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4061 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# 0.01fF
C4062 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.02fF
C4063 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4064 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C4065 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# -0.00fF
C4066 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# 0.00fF
C4067 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# 0.01fF
C4068 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.00fF
C4069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4070 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C4071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4072 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4073 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C4074 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4075 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C4076 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C4077 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C4078 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C4079 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# -0.00fF
C4080 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.00fF
C4081 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.01fF
C4082 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4083 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4084 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4085 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4086 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4087 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4088 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4089 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.01fF
C4090 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# 0.00fF
C4091 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C4092 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.02fF
C4093 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C4094 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C4095 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C4096 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# 0.00fF
C4097 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.02fF
C4098 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.01fF
C4099 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4100 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C4101 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# -0.00fF
C4102 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4103 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# -0.00fF
C4104 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.02fF
C4106 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C4107 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.00fF
C4108 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# 0.00fF
C4109 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C4110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4111 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C4112 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# 0.01fF
C4113 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4114 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4115 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4116 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# 0.00fF
C4117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4118 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C4119 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C4120 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# 0.02fF
C4121 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 1.18fF
C4122 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C4123 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C4124 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# -0.00fF
C4125 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C4126 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4127 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4128 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4129 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4130 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# 0.00fF
C4131 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# -0.00fF
C4132 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.01fF
C4133 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C4134 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C4135 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.01fF
C4136 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# 0.00fF
C4137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C4138 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.01fF
C4139 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.02fF
C4140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.02fF
C4141 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.00fF
C4142 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# 0.00fF
C4143 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C4144 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C4145 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C4146 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4147 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.02fF
C4148 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C4149 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4150 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C4151 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C4152 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C4153 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.01fF
C4154 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4155 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4156 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# -0.00fF
C4157 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.01fF
C4158 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# -0.00fF
C4159 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.00fF
C4160 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# 0.01fF
C4161 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# -0.00fF
C4162 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# -0.00fF
C4163 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C4164 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.01fF
C4165 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C4166 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# 0.00fF
C4167 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.01fF
C4168 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.02fF
C4169 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.01fF
C4170 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.02fF
C4171 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# 0.00fF
C4172 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C4173 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C4174 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C4175 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.01fF
C4176 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# 0.00fF
C4177 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# 0.00fF
C4178 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# 0.00fF
C4179 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C4180 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# 0.01fF
C4181 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# 0.00fF
C4182 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4183 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# 0.01fF
C4184 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C4185 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# 0.00fF
C4186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.01fF
C4187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# 0.01fF
C4188 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4189 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C4190 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C4191 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.01fF
C4192 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4193 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.27fF
C4194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# -0.00fF
C4195 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C4196 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.00fF
C4197 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# 0.01fF
C4198 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# 0.00fF
C4199 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# -0.00fF
C4200 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# 0.00fF
C4201 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.01fF
C4202 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4203 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# 0.00fF
C4204 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4205 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C4206 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C4207 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# 0.00fF
C4208 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# 0.01fF
C4209 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4210 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C4211 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4212 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C4213 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C4214 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C4215 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# 0.00fF
C4216 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C4217 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C4218 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# 0.01fF
C4219 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# 0.02fF
C4220 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.02fF
C4221 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C4222 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4223 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C4224 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C4225 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.01fF
C4226 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4227 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.00fF
C4228 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4229 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4230 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.02fF
C4231 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.01fF
C4232 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4233 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# 0.02fF
C4234 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# -0.00fF
C4235 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C4236 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# -0.00fF
C4237 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C4238 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C4239 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C4240 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4241 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C4242 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4243 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C4244 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C4245 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.93fF
C4246 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4247 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.01fF
C4248 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.01fF
C4249 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C4250 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4251 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.01fF
C4252 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4253 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# 0.00fF
C4254 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# 0.00fF
C4255 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C4256 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# -0.00fF
C4257 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.02fF
C4258 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# 0.00fF
C4259 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.01fF
C4260 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.00fF
C4261 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.01fF
C4262 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# 0.00fF
C4263 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C4264 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C4265 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4266 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.01fF
C4267 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4268 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C4269 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C4270 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C4271 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.02fF
C4272 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4273 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# -0.00fF
C4274 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4275 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# 0.00fF
C4276 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4277 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# 0.00fF
C4278 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C4279 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4280 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C4281 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4282 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4283 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# 0.00fF
C4284 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C4285 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C4286 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.02fF
C4287 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4288 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# -0.00fF
C4289 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# 0.00fF
C4290 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4291 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# -0.00fF
C4292 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4293 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4294 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4295 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.00fF
C4296 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4297 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C4298 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# 0.00fF
C4299 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4300 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C4301 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C4302 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# 0.00fF
C4303 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C4304 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.00fF
C4305 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4306 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.01fF
C4307 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# 0.01fF
C4308 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.02fF
C4309 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4310 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# -0.00fF
C4311 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C4312 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.01fF
C4313 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4314 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C4315 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4316 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# -0.00fF
C4317 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# 0.01fF
C4318 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# 0.00fF
C4319 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C4320 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4321 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4322 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.31fF
C4323 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.02fF
C4324 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4325 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C4326 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# -0.00fF
C4327 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4328 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4329 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C4330 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# 0.01fF
C4331 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4332 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C4333 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4334 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# 0.00fF
C4335 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.00fF
C4336 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# -0.00fF
C4337 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.01fF
C4338 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# 0.00fF
C4339 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.01fF
C4340 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# 0.00fF
C4341 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# 0.00fF
C4342 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.00fF
C4343 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# 0.01fF
C4344 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# 0.00fF
C4345 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4346 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C4347 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.01fF
C4348 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# 0.01fF
C4349 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4350 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4351 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.00fF
C4352 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# 0.00fF
C4353 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.02fF
C4354 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.01fF
C4355 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4356 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.00fF
C4357 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4358 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C4359 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# 0.00fF
C4360 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4361 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.02fF
C4362 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C4363 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# 0.00fF
C4364 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C4365 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# 0.00fF
C4366 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C4367 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4368 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4369 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.01fF
C4370 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4371 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C4372 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C4373 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# 0.00fF
C4374 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4375 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C4376 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# 0.00fF
C4377 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4378 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# 0.00fF
C4379 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.01fF
C4380 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.01fF
C4381 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# 0.00fF
C4382 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C4383 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.01fF
C4384 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# -0.00fF
C4385 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4386 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4387 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4388 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C4389 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# 0.01fF
C4390 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4391 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.02fF
C4392 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.01fF
C4393 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C4394 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4395 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.00fF
C4396 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4397 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4398 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C4399 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4400 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# 0.00fF
C4401 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4402 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.01fF
C4403 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C4404 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.57fF
C4405 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C4406 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4407 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.00fF
C4408 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# 0.02fF
C4409 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# 0.00fF
C4410 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# 0.00fF
C4411 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4412 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4413 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4414 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4415 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C4416 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4417 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.00fF
C4418 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# -0.00fF
C4419 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4420 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4421 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4422 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.00fF
C4423 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# 0.00fF
C4424 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.01fF
C4425 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.02fF
C4426 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# 0.02fF
C4427 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# 0.00fF
C4428 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.01fF
C4429 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# 0.00fF
C4430 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# -0.00fF
C4431 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.00fF
C4432 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# 0.01fF
C4433 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# 0.00fF
C4434 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# 0.01fF
C4435 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.02fF
C4436 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4437 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# 0.00fF
C4438 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4439 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# 0.01fF
C4440 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# -0.00fF
C4441 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.00fF
C4442 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# -0.00fF
C4443 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.01fF
C4444 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C4445 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4446 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.02fF
C4447 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C4448 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4449 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4450 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4451 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C4452 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.01fF
C4453 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4454 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4455 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C4456 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# 0.00fF
C4457 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C4458 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# 0.00fF
C4459 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# -0.00fF
C4460 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4461 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4462 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4463 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.01fF
C4464 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4465 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4466 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# -0.00fF
C4467 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4468 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C4469 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.00fF
C4470 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# 0.00fF
C4471 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# 0.02fF
C4472 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# 0.00fF
C4473 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.01fF
C4474 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# -0.00fF
C4475 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# 0.02fF
C4476 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# 0.02fF
C4477 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# -0.00fF
C4478 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4479 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C4480 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.01fF
C4481 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4482 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.01fF
C4483 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4484 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C4485 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C4486 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# -0.00fF
C4487 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4488 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C4489 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# 0.00fF
C4490 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4491 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.00fF
C4492 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.01fF
C4493 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# 0.00fF
C4494 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4495 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4496 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C4497 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# 0.02fF
C4498 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.00fF
C4499 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# 0.01fF
C4500 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4501 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.02fF
C4502 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# 0.01fF
C4503 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# -0.00fF
C4504 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.27fF
C4505 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4506 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# 0.00fF
C4507 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C4508 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.00fF
C4509 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# 0.00fF
C4510 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4511 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 1.18fF
C4512 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4513 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# 0.00fF
C4514 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# 0.01fF
C4515 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4516 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4517 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# 0.00fF
C4518 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4519 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# 0.01fF
C4520 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.00fF
C4521 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4522 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.01fF
C4523 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C4524 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4525 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4526 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.00fF
C4527 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4528 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# 0.01fF
C4529 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4530 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C4531 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# 0.00fF
C4532 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.00fF
C4533 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.01fF
C4534 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.57fF
C4535 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# 0.00fF
C4536 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# 0.00fF
C4537 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# -0.00fF
C4538 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# 0.02fF
C4539 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4540 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# 0.01fF
C4541 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# 0.00fF
C4542 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.00fF
C4543 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4544 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C4545 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# 0.00fF
C4546 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# 0.00fF
C4547 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# 0.00fF
C4548 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# 0.00fF
C4549 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C4550 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C4551 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4552 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C4553 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4554 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4555 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4556 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.00fF
C4557 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4558 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# 0.00fF
C4559 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# 0.01fF
C4560 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4561 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# 0.01fF
C4562 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# 0.00fF
C4563 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4564 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4565 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# 0.01fF
C4566 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.00fF
C4567 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# -0.00fF
C4568 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4569 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4570 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# 0.00fF
C4571 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C4572 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4573 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# 0.00fF
C4574 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# 0.00fF
C4575 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C4576 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4577 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4578 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# 0.00fF
C4579 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# 0.01fF
C4580 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4581 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# -0.00fF
C4582 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4583 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.31fF
C4584 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# 0.02fF
C4585 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# -0.00fF
C4586 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# 0.00fF
C4587 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C4588 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# 0.01fF
C4589 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# 0.00fF
C4590 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# 0.00fF
C4591 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# -0.00fF
C4592 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# 0.00fF
C4593 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# 0.00fF
C4594 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.02fF
C4595 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4596 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# 0.00fF
C4597 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# 0.00fF
C4598 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C4599 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C4600 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4601 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# 0.01fF
C4602 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.02fF
C4603 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# 0.00fF
C4604 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.00fF
C4605 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.01fF
C4606 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4607 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4608 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.01fF
C4609 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# 0.01fF
C4610 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C4611 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C4612 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# -0.00fF
C4613 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# 0.01fF
C4614 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C4615 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# 0.00fF
C4616 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.00fF
C4617 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C4618 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C4619 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# -0.00fF
C4620 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# 0.00fF
C4621 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.00fF
C4622 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.00fF
C4623 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# 0.01fF
C4624 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# 0.01fF
C4625 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# -0.00fF
C4626 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# 0.00fF
C4627 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# 0.00fF
C4628 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4629 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4630 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4631 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.01fF
C4632 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.01fF
C4633 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4634 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# 0.01fF
C4635 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# 0.01fF
C4636 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# 0.01fF
C4637 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# 0.00fF
C4638 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4639 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C4640 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# 0.00fF
C4641 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# 0.00fF
C4642 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.00fF
C4643 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# -0.00fF
C4644 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C4645 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4646 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4647 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# -0.00fF
C4648 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4649 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# 0.00fF
C4650 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# 0.00fF
C4651 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.01fF
C4652 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# -0.00fF
C4653 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# 0.00fF
C4654 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# 0.00fF
C4655 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4656 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# 0.02fF
C4657 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4658 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# 0.00fF
C4659 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# 0.00fF
C4660 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# 0.00fF
C4661 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.01fF
C4662 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# 0.01fF
C4663 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# 0.00fF
C4664 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.01fF
C4665 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# 0.00fF
C4666 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# 0.00fF
C4667 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4668 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4669 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# 0.01fF
C4670 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# -0.01fF
C4671 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# 0.01fF
C4672 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# -0.00fF
C4673 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# 0.00fF
C4674 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# 0.00fF
C4675 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4676 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# 0.00fF
C4677 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4678 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# 0.00fF
C4679 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4680 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4681 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# 0.02fF
C4682 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.02fF
C4683 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4684 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.00fF
C4685 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4686 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# 0.00fF
C4687 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# 0.00fF
C4688 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# 0.00fF
C4689 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4690 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# 0.00fF
C4691 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4692 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4693 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# -0.00fF
C4694 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# 0.00fF
C4695 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# 0.00fF
C4696 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# 0.00fF
C4697 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4698 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# -0.00fF
C4699 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C4700 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# -0.01fF
C4701 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4702 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.01fF
C4703 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# 0.00fF
C4704 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# 0.00fF
C4705 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# -0.00fF
C4706 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4707 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# 0.00fF
C4708 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# 0.00fF
C4709 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# 0.01fF
C4710 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# 0.00fF
C4711 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# 0.01fF
C4712 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.01fF
C4713 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# -0.00fF
C4714 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.00fF
C4715 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# -0.00fF
C4716 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4717 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4718 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C4719 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# 0.00fF
C4720 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.01fF
C4721 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# 0.01fF
C4722 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# 0.00fF
C4723 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# 0.00fF
C4724 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# 0.00fF
C4725 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4726 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# 0.00fF
C4727 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# 0.00fF
C4728 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.42fF
C4729 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.01fF
C4730 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4731 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# 0.00fF
C4732 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# 0.00fF
C4733 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.00fF
C4734 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# 0.00fF
C4735 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# 0.02fF
C4736 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# 0.00fF
C4737 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4738 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# 0.00fF
C4739 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# 0.00fF
C4740 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# 0.00fF
C4741 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4742 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# 0.00fF
C4743 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# -0.01fF
C4744 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4745 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4746 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4747 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# 0.00fF
C4748 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# 0.00fF
C4749 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4750 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# 0.00fF
C4751 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4752 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.01fF
C4753 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# 0.00fF
C4754 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# 0.00fF
C4755 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# 0.01fF
C4756 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# 0.00fF
C4757 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# 0.00fF
C4758 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# 0.01fF
C4759 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# 0.00fF
C4760 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4761 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# 0.01fF
C4762 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# -0.00fF
C4763 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# 0.00fF
C4764 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# 0.00fF
C4765 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# 0.02fF
C4766 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# 0.00fF
C4767 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4768 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# 0.00fF
C4769 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4770 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.93fF
C4771 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# -0.00fF
C4772 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# 0.00fF
C4773 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4774 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4775 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4776 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# 0.00fF
C4777 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# -0.00fF
C4778 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C4779 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4780 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# 0.00fF
C4781 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# 0.02fF
C4782 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4783 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# 0.01fF
C4784 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# 0.01fF
C4785 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.00fF
C4786 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# 0.00fF
C4787 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4788 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4789 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.01fF
C4790 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# 0.00fF
C4791 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# 0.00fF
C4792 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# 0.02fF
C4793 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# 0.93fF
C4794 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4795 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# 0.00fF
C4796 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# 0.00fF
C4797 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# 0.01fF
C4798 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# 0.01fF
C4799 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# 0.00fF
C4800 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# 0.00fF
C4801 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4802 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# 0.00fF
C4803 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# 0.00fF
C4804 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.93fF
C4805 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.00fF
C4806 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# 0.02fF
C4807 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4808 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# 0.00fF
C4809 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4810 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# 0.00fF
C4811 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4812 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# 0.01fF
C4813 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4814 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# 0.00fF
C4815 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# 0.00fF
C4816 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# 0.01fF
C4817 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# -0.00fF
C4818 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# 0.00fF
C4819 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# 0.00fF
C4820 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# 0.01fF
C4821 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# 0.00fF
C4822 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# 0.00fF
C4823 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# -0.00fF
C4824 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# -0.00fF
C4825 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# 0.00fF
C4826 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# 0.01fF
C4827 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# 0.01fF
C4828 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.00fF
C4829 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# 0.00fF
C4830 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# 0.00fF
C4831 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# 0.00fF
C4832 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# 0.01fF
C4833 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# 0.00fF
C4834 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# 0.02fF
C4835 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# -0.00fF
C4836 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# -0.00fF
C4837 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# 0.02fF
C4838 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# 0.00fF
C4839 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# 0.00fF
C4840 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# 0.02fF
C4841 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# 0.00fF
C4842 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4843 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# 0.00fF
C4844 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# 0.01fF
C4845 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# 0.01fF
C4846 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# -0.00fF
C4847 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# 0.00fF
C4848 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.00fF
C4849 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# 0.00fF
C4850 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# 0.00fF
C4851 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# 0.48fF
C4852 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# 0.00fF
C4853 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# 0.00fF
C4854 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# 0.01fF
C4855 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# 0.00fF
C4856 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4080_n100# VSUBS 1.08fF
C4857 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4172_n100# VSUBS 1.03fF
C4858 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4062_n188# VSUBS 0.11fF
C4859 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_4228_n100# VSUBS 0.17fF
C4860 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3642_n188# VSUBS 0.10fF
C4861 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3852_122# VSUBS 0.09fF
C4862 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3222_n188# VSUBS 0.11fF
C4863 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3432_122# VSUBS 0.11fF
C4864 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2802_n188# VSUBS 0.12fF
C4865 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_3012_122# VSUBS 0.11fF
C4866 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2382_n188# VSUBS 0.12fF
C4867 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2592_122# VSUBS 0.12fF
C4868 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1962_n188# VSUBS 0.12fF
C4869 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_2172_122# VSUBS 0.12fF
C4870 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1542_n188# VSUBS 0.12fF
C4871 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1752_122# VSUBS 0.12fF
C4872 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1122_n188# VSUBS 0.12fF
C4873 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_1332_122# VSUBS 0.12fF
C4874 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_702_n188# VSUBS 0.12fF
C4875 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_912_122# VSUBS 0.12fF
C4876 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_282_n188# VSUBS 0.12fF
C4877 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_492_122# VSUBS 0.12fF
C4878 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n138_n188# VSUBS 0.12fF
C4879 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_72_122# VSUBS 0.12fF
C4880 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n558_n188# VSUBS 0.12fF
C4881 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n348_122# VSUBS 0.12fF
C4882 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n978_n188# VSUBS 0.12fF
C4883 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n768_122# VSUBS 0.12fF
C4884 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1398_n188# VSUBS 0.12fF
C4885 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1188_122# VSUBS 0.12fF
C4886 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1818_n188# VSUBS 0.12fF
C4887 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n1608_122# VSUBS 0.12fF
C4888 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2238_n188# VSUBS 0.12fF
C4889 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2028_122# VSUBS 0.12fF
C4890 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2658_n188# VSUBS 0.12fF
C4891 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2448_122# VSUBS 0.12fF
C4892 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3078_n188# VSUBS 0.12fF
C4893 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n2868_122# VSUBS 0.12fF
C4894 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3498_n188# VSUBS 0.12fF
C4895 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3288_122# VSUBS 0.12fF
C4896 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3918_n188# VSUBS 0.12fF
C4897 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n3708_122# VSUBS 0.12fF
C4898 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4382_n100# VSUBS 0.20fF
C4899 sky130_fd_pr__nfet_01v8_J3WY8C_7/a_n4128_122# VSUBS 0.13fF
C4900 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4080_n100# VSUBS 1.08fF
C4901 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4172_n100# VSUBS 1.03fF
C4902 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4062_n188# VSUBS 0.11fF
C4903 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_4228_n100# VSUBS 0.17fF
C4904 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3642_n188# VSUBS 0.10fF
C4905 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3852_122# VSUBS 0.09fF
C4906 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3222_n188# VSUBS 0.11fF
C4907 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3432_122# VSUBS 0.11fF
C4908 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2802_n188# VSUBS 0.12fF
C4909 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_3012_122# VSUBS 0.11fF
C4910 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2382_n188# VSUBS 0.12fF
C4911 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2592_122# VSUBS 0.12fF
C4912 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1962_n188# VSUBS 0.12fF
C4913 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_2172_122# VSUBS 0.12fF
C4914 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1542_n188# VSUBS 0.12fF
C4915 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1752_122# VSUBS 0.12fF
C4916 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1122_n188# VSUBS 0.12fF
C4917 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_1332_122# VSUBS 0.12fF
C4918 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_702_n188# VSUBS 0.12fF
C4919 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_912_122# VSUBS 0.12fF
C4920 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_282_n188# VSUBS 0.12fF
C4921 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_492_122# VSUBS 0.12fF
C4922 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n138_n188# VSUBS 0.12fF
C4923 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_72_122# VSUBS 0.12fF
C4924 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n558_n188# VSUBS 0.12fF
C4925 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n348_122# VSUBS 0.12fF
C4926 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n978_n188# VSUBS 0.12fF
C4927 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n768_122# VSUBS 0.12fF
C4928 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1398_n188# VSUBS 0.12fF
C4929 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1188_122# VSUBS 0.12fF
C4930 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1818_n188# VSUBS 0.12fF
C4931 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n1608_122# VSUBS 0.12fF
C4932 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2238_n188# VSUBS 0.12fF
C4933 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2028_122# VSUBS 0.12fF
C4934 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2658_n188# VSUBS 0.12fF
C4935 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2448_122# VSUBS 0.12fF
C4936 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3078_n188# VSUBS 0.12fF
C4937 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n2868_122# VSUBS 0.12fF
C4938 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3498_n188# VSUBS 0.12fF
C4939 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3288_122# VSUBS 0.12fF
C4940 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3918_n188# VSUBS 0.12fF
C4941 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n3708_122# VSUBS 0.12fF
C4942 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4382_n100# VSUBS 0.20fF
C4943 sky130_fd_pr__nfet_01v8_J3WY8C_6/a_n4128_122# VSUBS 0.13fF
C4944 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4080_n100# VSUBS 1.08fF
C4945 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4172_n100# VSUBS 1.03fF
C4946 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4062_n188# VSUBS 0.11fF
C4947 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_4228_n100# VSUBS 0.17fF
C4948 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3642_n188# VSUBS 0.10fF
C4949 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3852_122# VSUBS 0.09fF
C4950 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3222_n188# VSUBS 0.11fF
C4951 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3432_122# VSUBS 0.11fF
C4952 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2802_n188# VSUBS 0.12fF
C4953 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_3012_122# VSUBS 0.11fF
C4954 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2382_n188# VSUBS 0.12fF
C4955 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2592_122# VSUBS 0.12fF
C4956 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1962_n188# VSUBS 0.12fF
C4957 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_2172_122# VSUBS 0.12fF
C4958 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1542_n188# VSUBS 0.12fF
C4959 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1752_122# VSUBS 0.12fF
C4960 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1122_n188# VSUBS 0.12fF
C4961 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_1332_122# VSUBS 0.12fF
C4962 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_702_n188# VSUBS 0.12fF
C4963 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_912_122# VSUBS 0.12fF
C4964 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_282_n188# VSUBS 0.12fF
C4965 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_492_122# VSUBS 0.12fF
C4966 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n138_n188# VSUBS 0.12fF
C4967 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_72_122# VSUBS 0.12fF
C4968 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n558_n188# VSUBS 0.12fF
C4969 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n348_122# VSUBS 0.12fF
C4970 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n978_n188# VSUBS 0.12fF
C4971 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n768_122# VSUBS 0.12fF
C4972 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1398_n188# VSUBS 0.12fF
C4973 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1188_122# VSUBS 0.12fF
C4974 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1818_n188# VSUBS 0.12fF
C4975 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n1608_122# VSUBS 0.12fF
C4976 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2238_n188# VSUBS 0.12fF
C4977 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2028_122# VSUBS 0.12fF
C4978 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2658_n188# VSUBS 0.12fF
C4979 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2448_122# VSUBS 0.12fF
C4980 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3078_n188# VSUBS 0.12fF
C4981 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n2868_122# VSUBS 0.12fF
C4982 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3498_n188# VSUBS 0.12fF
C4983 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3288_122# VSUBS 0.12fF
C4984 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3918_n188# VSUBS 0.12fF
C4985 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n3708_122# VSUBS 0.12fF
C4986 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4382_n100# VSUBS 0.20fF
C4987 sky130_fd_pr__nfet_01v8_J3WY8C_5/a_n4128_122# VSUBS 0.13fF
C4988 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4080_n100# VSUBS 1.08fF
C4989 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4172_n100# VSUBS 1.03fF
C4990 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4062_n188# VSUBS 0.11fF
C4991 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_4228_n100# VSUBS 0.17fF
C4992 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3642_n188# VSUBS 0.10fF
C4993 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3852_122# VSUBS 0.09fF
C4994 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3222_n188# VSUBS 0.11fF
C4995 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3432_122# VSUBS 0.11fF
C4996 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2802_n188# VSUBS 0.12fF
C4997 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_3012_122# VSUBS 0.11fF
C4998 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2382_n188# VSUBS 0.12fF
C4999 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2592_122# VSUBS 0.12fF
C5000 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1962_n188# VSUBS 0.12fF
C5001 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_2172_122# VSUBS 0.12fF
C5002 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1542_n188# VSUBS 0.12fF
C5003 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1752_122# VSUBS 0.12fF
C5004 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1122_n188# VSUBS 0.12fF
C5005 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_1332_122# VSUBS 0.12fF
C5006 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_702_n188# VSUBS 0.12fF
C5007 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_912_122# VSUBS 0.12fF
C5008 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_282_n188# VSUBS 0.12fF
C5009 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_492_122# VSUBS 0.12fF
C5010 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n138_n188# VSUBS 0.12fF
C5011 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_72_122# VSUBS 0.12fF
C5012 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n558_n188# VSUBS 0.12fF
C5013 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n348_122# VSUBS 0.12fF
C5014 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n978_n188# VSUBS 0.12fF
C5015 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n768_122# VSUBS 0.12fF
C5016 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1398_n188# VSUBS 0.12fF
C5017 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1188_122# VSUBS 0.12fF
C5018 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1818_n188# VSUBS 0.12fF
C5019 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n1608_122# VSUBS 0.12fF
C5020 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2238_n188# VSUBS 0.12fF
C5021 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2028_122# VSUBS 0.12fF
C5022 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2658_n188# VSUBS 0.12fF
C5023 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2448_122# VSUBS 0.12fF
C5024 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3078_n188# VSUBS 0.12fF
C5025 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n2868_122# VSUBS 0.12fF
C5026 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3498_n188# VSUBS 0.12fF
C5027 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3288_122# VSUBS 0.12fF
C5028 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3918_n188# VSUBS 0.12fF
C5029 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n3708_122# VSUBS 0.12fF
C5030 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4382_n100# VSUBS 0.20fF
C5031 sky130_fd_pr__nfet_01v8_J3WY8C_4/a_n4128_122# VSUBS 0.13fF
C5032 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4080_n100# VSUBS 1.08fF
C5033 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4172_n100# VSUBS 1.03fF
C5034 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4062_n188# VSUBS 0.11fF
C5035 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_4228_n100# VSUBS 0.17fF
C5036 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3642_n188# VSUBS 0.10fF
C5037 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3852_122# VSUBS 0.09fF
C5038 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3222_n188# VSUBS 0.11fF
C5039 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3432_122# VSUBS 0.11fF
C5040 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2802_n188# VSUBS 0.12fF
C5041 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_3012_122# VSUBS 0.11fF
C5042 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2382_n188# VSUBS 0.12fF
C5043 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2592_122# VSUBS 0.12fF
C5044 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1962_n188# VSUBS 0.12fF
C5045 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_2172_122# VSUBS 0.12fF
C5046 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1542_n188# VSUBS 0.12fF
C5047 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1752_122# VSUBS 0.12fF
C5048 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1122_n188# VSUBS 0.12fF
C5049 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_1332_122# VSUBS 0.12fF
C5050 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_702_n188# VSUBS 0.12fF
C5051 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_912_122# VSUBS 0.12fF
C5052 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_282_n188# VSUBS 0.12fF
C5053 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_492_122# VSUBS 0.12fF
C5054 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n138_n188# VSUBS 0.12fF
C5055 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_72_122# VSUBS 0.12fF
C5056 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n558_n188# VSUBS 0.12fF
C5057 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n348_122# VSUBS 0.12fF
C5058 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n978_n188# VSUBS 0.12fF
C5059 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n768_122# VSUBS 0.12fF
C5060 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1398_n188# VSUBS 0.12fF
C5061 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1188_122# VSUBS 0.12fF
C5062 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1818_n188# VSUBS 0.12fF
C5063 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n1608_122# VSUBS 0.12fF
C5064 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2238_n188# VSUBS 0.12fF
C5065 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2028_122# VSUBS 0.12fF
C5066 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2658_n188# VSUBS 0.12fF
C5067 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2448_122# VSUBS 0.12fF
C5068 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3078_n188# VSUBS 0.12fF
C5069 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n2868_122# VSUBS 0.12fF
C5070 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3498_n188# VSUBS 0.12fF
C5071 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3288_122# VSUBS 0.12fF
C5072 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3918_n188# VSUBS 0.12fF
C5073 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n3708_122# VSUBS 0.12fF
C5074 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4382_n100# VSUBS 0.20fF
C5075 sky130_fd_pr__nfet_01v8_J3WY8C_3/a_n4128_122# VSUBS 0.13fF
C5076 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4080_n100# VSUBS 1.08fF
C5077 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4172_n100# VSUBS 1.03fF
C5078 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4062_n188# VSUBS 0.11fF
C5079 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_4228_n100# VSUBS 0.17fF
C5080 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3642_n188# VSUBS 0.10fF
C5081 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3852_122# VSUBS 0.09fF
C5082 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3222_n188# VSUBS 0.11fF
C5083 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3432_122# VSUBS 0.11fF
C5084 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2802_n188# VSUBS 0.12fF
C5085 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_3012_122# VSUBS 0.11fF
C5086 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2382_n188# VSUBS 0.12fF
C5087 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2592_122# VSUBS 0.12fF
C5088 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1962_n188# VSUBS 0.12fF
C5089 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_2172_122# VSUBS 0.12fF
C5090 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1542_n188# VSUBS 0.12fF
C5091 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1752_122# VSUBS 0.12fF
C5092 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1122_n188# VSUBS 0.12fF
C5093 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_1332_122# VSUBS 0.12fF
C5094 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_702_n188# VSUBS 0.12fF
C5095 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_912_122# VSUBS 0.12fF
C5096 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_282_n188# VSUBS 0.12fF
C5097 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_492_122# VSUBS 0.12fF
C5098 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n138_n188# VSUBS 0.12fF
C5099 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_72_122# VSUBS 0.12fF
C5100 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n558_n188# VSUBS 0.12fF
C5101 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n348_122# VSUBS 0.12fF
C5102 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n978_n188# VSUBS 0.12fF
C5103 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n768_122# VSUBS 0.12fF
C5104 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1398_n188# VSUBS 0.12fF
C5105 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1188_122# VSUBS 0.12fF
C5106 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1818_n188# VSUBS 0.12fF
C5107 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n1608_122# VSUBS 0.12fF
C5108 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2238_n188# VSUBS 0.12fF
C5109 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2028_122# VSUBS 0.12fF
C5110 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2658_n188# VSUBS 0.12fF
C5111 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2448_122# VSUBS 0.12fF
C5112 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3078_n188# VSUBS 0.12fF
C5113 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n2868_122# VSUBS 0.12fF
C5114 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3498_n188# VSUBS 0.12fF
C5115 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3288_122# VSUBS 0.12fF
C5116 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3918_n188# VSUBS 0.12fF
C5117 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n3708_122# VSUBS 0.12fF
C5118 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4382_n100# VSUBS 0.20fF
C5119 sky130_fd_pr__nfet_01v8_J3WY8C_2/a_n4128_122# VSUBS 0.13fF
C5120 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4080_n100# VSUBS 1.08fF
C5121 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4172_n100# VSUBS 1.03fF
C5122 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4062_n188# VSUBS 0.11fF
C5123 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_4228_n100# VSUBS 0.17fF
C5124 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3642_n188# VSUBS 0.10fF
C5125 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3852_122# VSUBS 0.09fF
C5126 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3222_n188# VSUBS 0.11fF
C5127 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3432_122# VSUBS 0.11fF
C5128 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2802_n188# VSUBS 0.12fF
C5129 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_3012_122# VSUBS 0.11fF
C5130 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2382_n188# VSUBS 0.12fF
C5131 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2592_122# VSUBS 0.12fF
C5132 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1962_n188# VSUBS 0.12fF
C5133 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_2172_122# VSUBS 0.12fF
C5134 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1542_n188# VSUBS 0.12fF
C5135 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1752_122# VSUBS 0.12fF
C5136 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1122_n188# VSUBS 0.12fF
C5137 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_1332_122# VSUBS 0.12fF
C5138 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_702_n188# VSUBS 0.12fF
C5139 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_912_122# VSUBS 0.12fF
C5140 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_282_n188# VSUBS 0.12fF
C5141 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_492_122# VSUBS 0.12fF
C5142 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n138_n188# VSUBS 0.12fF
C5143 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_72_122# VSUBS 0.12fF
C5144 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n558_n188# VSUBS 0.12fF
C5145 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n348_122# VSUBS 0.12fF
C5146 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n978_n188# VSUBS 0.12fF
C5147 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n768_122# VSUBS 0.12fF
C5148 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1398_n188# VSUBS 0.12fF
C5149 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1188_122# VSUBS 0.12fF
C5150 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1818_n188# VSUBS 0.12fF
C5151 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n1608_122# VSUBS 0.12fF
C5152 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2238_n188# VSUBS 0.12fF
C5153 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2028_122# VSUBS 0.12fF
C5154 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2658_n188# VSUBS 0.12fF
C5155 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2448_122# VSUBS 0.12fF
C5156 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3078_n188# VSUBS 0.12fF
C5157 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n2868_122# VSUBS 0.12fF
C5158 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3498_n188# VSUBS 0.12fF
C5159 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3288_122# VSUBS 0.12fF
C5160 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3918_n188# VSUBS 0.12fF
C5161 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n3708_122# VSUBS 0.12fF
C5162 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4382_n100# VSUBS 0.20fF
C5163 sky130_fd_pr__nfet_01v8_J3WY8C_1/a_n4128_122# VSUBS 0.13fF
C5164 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4080_n100# VSUBS 1.08fF
C5165 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4172_n100# VSUBS 1.03fF
C5166 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4062_n188# VSUBS 0.11fF
C5167 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_4228_n100# VSUBS 0.17fF
C5168 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3642_n188# VSUBS 0.10fF
C5169 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3852_122# VSUBS 0.09fF
C5170 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3222_n188# VSUBS 0.11fF
C5171 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3432_122# VSUBS 0.11fF
C5172 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2802_n188# VSUBS 0.12fF
C5173 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_3012_122# VSUBS 0.11fF
C5174 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2382_n188# VSUBS 0.12fF
C5175 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2592_122# VSUBS 0.12fF
C5176 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1962_n188# VSUBS 0.12fF
C5177 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_2172_122# VSUBS 0.12fF
C5178 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1542_n188# VSUBS 0.12fF
C5179 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1752_122# VSUBS 0.12fF
C5180 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1122_n188# VSUBS 0.12fF
C5181 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_1332_122# VSUBS 0.12fF
C5182 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_702_n188# VSUBS 0.12fF
C5183 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_912_122# VSUBS 0.12fF
C5184 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_282_n188# VSUBS 0.12fF
C5185 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_492_122# VSUBS 0.12fF
C5186 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n138_n188# VSUBS 0.12fF
C5187 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_72_122# VSUBS 0.12fF
C5188 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n558_n188# VSUBS 0.12fF
C5189 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n348_122# VSUBS 0.12fF
C5190 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n978_n188# VSUBS 0.12fF
C5191 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n768_122# VSUBS 0.12fF
C5192 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1398_n188# VSUBS 0.12fF
C5193 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1188_122# VSUBS 0.12fF
C5194 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1818_n188# VSUBS 0.12fF
C5195 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n1608_122# VSUBS 0.12fF
C5196 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2238_n188# VSUBS 0.12fF
C5197 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2028_122# VSUBS 0.12fF
C5198 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2658_n188# VSUBS 0.12fF
C5199 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2448_122# VSUBS 0.12fF
C5200 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3078_n188# VSUBS 0.12fF
C5201 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n2868_122# VSUBS 0.12fF
C5202 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3498_n188# VSUBS 0.12fF
C5203 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3288_122# VSUBS 0.12fF
C5204 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3918_n188# VSUBS 0.12fF
C5205 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n3708_122# VSUBS 0.12fF
C5206 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4382_n100# VSUBS 0.20fF
C5207 sky130_fd_pr__nfet_01v8_J3WY8C_0/a_n4128_122# VSUBS 0.13fF
.ends

.subckt comparator_v2 sky130_fd_sc_hd__buf_2_1/a_27_47# outp outn sky130_fd_sc_hd__buf_2_0/X
+ li_n2324_818# sky130_fd_sc_hd__nand2_4_0/a_27_47# li_940_818# sky130_fd_sc_hd__buf_2_0/a_27_47#
+ VSS sky130_fd_sc_hd__buf_2_1/X VDD clk li_940_3458# in sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__nand2_4_1/a_27_47# ip sky130_fd_sc_hd__buf_2_1/A
Xlatch_pmos_pair_0 VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD VDD VDD
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VDD sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A VDD VDD VDD VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A VDD VDD sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VDD VDD sky130_fd_sc_hd__buf_2_1/A VDD sky130_fd_sc_hd__buf_2_0/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VDD latch_pmos_pair
Xsky130_fd_sc_hd__nand2_4_0 sky130_fd_sc_hd__buf_2_1/X outp VSS VDD outn VSS VDD sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_sc_hd__nand2_4_1 sky130_fd_sc_hd__buf_2_0/X outn VSS VDD outp VSS VDD sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ sky130_fd_sc_hd__nand2_4
Xsky130_fd_pr__pfet_01v8_VCG74W_1 li_940_3458# li_940_3458# li_940_3458# clk VDD VDD
+ clk clk li_940_3458# li_940_3458# li_940_3458# clk VDD VDD clk clk VDD li_940_3458#
+ clk clk VDD clk clk clk VDD VDD clk clk li_940_3458# li_940_3458# clk VDD clk clk
+ VSS sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_pr__pfet_01v8_VCG74W_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A clk VDD VDD clk clk VDD sky130_fd_sc_hd__buf_2_1/A clk
+ clk VDD clk clk clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ clk VDD clk clk VSS sky130_fd_pr__pfet_01v8_VCG74W
Xsky130_fd_sc_hd__buf_2_0 sky130_fd_sc_hd__buf_2_0/A VSS VDD sky130_fd_sc_hd__buf_2_0/X
+ VSS VDD sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__buf_2_1 sky130_fd_sc_hd__buf_2_1/A VSS VDD sky130_fd_sc_hd__buf_2_1/X
+ VSS VDD sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__decap_12_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_0 clk sky130_fd_sc_hd__buf_2_0/A clk VDD VDD clk sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A clk sky130_fd_sc_hd__buf_2_0/A
+ VDD VDD clk VDD VDD clk clk sky130_fd_sc_hd__buf_2_0/A VDD sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A clk clk VDD VDD clk clk clk sky130_fd_sc_hd__buf_2_0/A
+ clk clk clk clk VSS precharge_pmos
Xcurrent_tail_0 li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# VSS VSS VSS
+ li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS VSS VSS li_n2324_818# li_n2324_818# li_n2324_818# li_n2324_818#
+ VSS VSS VSS VSS li_n2324_818# li_n2324_818# VSS VSS VSS clk li_n2324_818# VSS current_tail
Xsky130_fd_sc_hd__decap_12_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_12
Xprecharge_pmos_1 clk li_940_818# clk VDD VDD clk li_940_818# li_940_818# li_940_818#
+ clk li_940_818# VDD VDD clk VDD VDD clk clk li_940_818# VDD li_940_818# li_940_818#
+ clk clk VDD VDD clk clk clk li_940_818# clk clk clk clk VSS precharge_pmos
Xlatch_nmos_pair_0 sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A li_940_3458# sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ li_940_818# sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2_0/A VSS sky130_fd_sc_hd__buf_2_1/A sky130_fd_sc_hd__buf_2_1/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A latch_nmos_pair
Xinput_diff_pair_0 ip ip ip in in VSS ip in in in in VSS li_940_3458# ip ip ip in
+ ip li_n2324_818# ip ip in ip ip ip in in in ip ip ip in ip in ip in ip in in ip
+ ip VSS ip ip in ip li_n2324_818# ip ip in in in ip ip ip in in in li_940_3458# in
+ in ip ip in ip in ip ip ip VSS ip in ip ip ip in in in ip ip in in ip in VSS ip
+ in in in in in ip in li_940_818# ip ip in ip ip li_n2324_818# in in ip ip ip in
+ ip ip ip ip in in in in in in VSS ip in in ip ip ip ip ip in in ip ip in in ip li_940_818#
+ ip ip in li_n2324_818# in in in VSS ip in in ip ip ip in ip ip ip in in ip in ip
+ in ip ip ip in in in in in VSS in ip li_n2324_818# ip ip in ip ip in ip ip in ip
+ ip li_940_3458# in in ip ip ip in in in ip ip in ip ip in in in VSS ip in VSS VSS
+ in in ip ip in in ip ip ip in in ip ip li_940_3458# in ip in ip ip in li_n2324_818#
+ ip in in in in in in ip ip in in ip ip ip ip VSS ip ip ip in in in in ip ip in ip
+ ip ip in in ip ip in in ip in in li_n2324_818# in in in in ip in in ip in ip li_940_818#
+ VSS ip ip ip ip in in ip ip VSS in in in ip in in ip ip ip in in ip in in VSS in
+ in li_n2324_818# ip in in in ip ip ip ip in in ip ip li_940_818# in ip ip in in
+ in ip in ip in ip ip ip in in in ip ip ip ip in in in ip ip in in in in ip VSS VSS
+ in in ip ip in in in input_diff_pair
C0 sky130_fd_sc_hd__buf_2_0/A li_940_818# 9.11fF
C1 ip li_940_3458# 13.70fF
C2 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_0/A 0.10fF
C3 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.02fF
C4 outp sky130_fd_sc_hd__buf_2_1/X 0.03fF
C5 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.00fF
C6 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_1/A 0.09fF
C7 clk li_n2324_818# 6.65fF
C8 sky130_fd_sc_hd__buf_2_1/a_27_47# outn 0.04fF
C9 sky130_fd_sc_hd__buf_2_0/a_27_47# VDD 0.07fF
C10 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_1/X 0.11fF
C11 outp sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.09fF
C12 ip sky130_fd_sc_hd__buf_2_0/A 2.05fF
C13 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.00fF
C14 outn sky130_fd_sc_hd__buf_2_0/A 0.05fF
C15 clk li_940_3458# 2.08fF
C16 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.05fF
C17 in sky130_fd_sc_hd__buf_2_1/A 0.67fF
C18 li_n2324_818# VDD 0.09fF
C19 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.03fF
C20 in li_940_818# 12.98fF
C21 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.03fF
C22 outn sky130_fd_sc_hd__buf_2_1/X 0.23fF
C23 VDD li_940_3458# 2.17fF
C24 outp VSS 0.44fF
C25 sky130_fd_sc_hd__buf_2_1/A VSS 1.57fF
C26 li_940_818# VSS 0.96fF
C27 clk sky130_fd_sc_hd__buf_2_0/A 3.32fF
C28 outn sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.06fF
C29 sky130_fd_sc_hd__buf_2_0/X VSS 0.04fF
C30 sky130_fd_sc_hd__buf_2_1/a_27_47# VDD 0.09fF
C31 in ip 30.51fF
C32 sky130_fd_sc_hd__nand2_4_0/a_27_47# VSS 0.28fF
C33 VDD sky130_fd_sc_hd__buf_2_0/A 30.94fF
C34 ip VSS 2.78fF
C35 outn VSS 0.56fF
C36 VDD sky130_fd_sc_hd__buf_2_1/X 0.24fF
C37 in clk 0.47fF
C38 VDD sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.02fF
C39 in VDD 0.01fF
C40 outp sky130_fd_sc_hd__buf_2_1/A 0.05fF
C41 li_n2324_818# li_940_3458# 4.64fF
C42 clk VSS 1.71fF
C43 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_1/a_27_47# 0.06fF
C44 li_940_818# sky130_fd_sc_hd__buf_2_1/A 21.09fF
C45 outp sky130_fd_sc_hd__buf_2_0/X 0.20fF
C46 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.01fF
C47 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_1/A 0.04fF
C48 outp sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.08fF
C49 VDD VSS 0.85fF
C50 sky130_fd_sc_hd__nand2_4_0/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.00fF
C51 li_n2324_818# sky130_fd_sc_hd__buf_2_0/A 1.31fF
C52 sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.01fF
C53 outn outp 1.34fF
C54 ip sky130_fd_sc_hd__buf_2_1/A 1.73fF
C55 sky130_fd_sc_hd__buf_2_0/A li_940_3458# 18.81fF
C56 outn sky130_fd_sc_hd__buf_2_1/A 0.03fF
C57 ip li_940_818# 35.81fF
C58 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.02fF
C59 outn sky130_fd_sc_hd__buf_2_0/X 0.03fF
C60 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.02fF
C61 outn sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.18fF
C62 in li_n2324_818# 49.83fF
C63 clk sky130_fd_sc_hd__buf_2_1/A 3.02fF
C64 clk li_940_818# 4.03fF
C65 sky130_fd_sc_hd__buf_2_0/a_27_47# VSS 0.03fF
C66 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.11fF
C67 in li_940_3458# 37.79fF
C68 VDD outp 0.83fF
C69 sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_0/A 0.06fF
C70 VDD sky130_fd_sc_hd__buf_2_1/A 26.23fF
C71 li_n2324_818# VSS 3.07fF
C72 VDD li_940_818# 2.08fF
C73 VDD sky130_fd_sc_hd__buf_2_0/X 0.20fF
C74 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_0/A 0.00fF
C75 li_940_3458# VSS 1.22fF
C76 clk ip 0.62fF
C77 VDD sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.01fF
C78 in sky130_fd_sc_hd__buf_2_0/A 1.07fF
C79 sky130_fd_sc_hd__buf_2_1/a_27_47# VSS 0.04fF
C80 sky130_fd_sc_hd__nand2_4_1/a_27_47# sky130_fd_sc_hd__buf_2_1/X 0.01fF
C81 VDD ip 0.03fF
C82 outn VDD 0.93fF
C83 sky130_fd_sc_hd__buf_2_0/A VSS 2.10fF
C84 sky130_fd_sc_hd__buf_2_0/a_27_47# outp 0.04fF
C85 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.02fF
C86 sky130_fd_sc_hd__buf_2_1/X VSS 0.05fF
C87 sky130_fd_sc_hd__buf_2_0/a_27_47# sky130_fd_sc_hd__buf_2_0/X 0.11fF
C88 clk VDD 14.94fF
C89 li_n2324_818# sky130_fd_sc_hd__buf_2_1/A 0.95fF
C90 li_n2324_818# li_940_818# 2.99fF
C91 sky130_fd_sc_hd__nand2_4_1/a_27_47# VSS 0.24fF
C92 sky130_fd_sc_hd__buf_2_1/A li_940_3458# 9.09fF
C93 in VSS 1.52fF
C94 li_940_818# li_940_3458# 4.44fF
C95 sky130_fd_sc_hd__buf_2_0/a_27_47# outn 0.02fF
C96 sky130_fd_sc_hd__buf_2_1/a_27_47# outp 0.02fF
C97 sky130_fd_sc_hd__buf_2_1/a_27_47# sky130_fd_sc_hd__buf_2_1/A 0.03fF
C98 li_n2324_818# ip 48.05fF
C99 outp sky130_fd_sc_hd__buf_2_0/A 0.04fF
C100 sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__buf_2_1/A 76.01fF
C101 li_940_3458# 0 -1592.65fF
C102 li_940_818# 0 -2262.83fF
C103 outn 0 21.71fF
C104 in 0 -297.33fF
C105 li_n2324_818# 0 -3722.01fF
C106 ip 0 -420.77fF
C107 VSS 0 -70.10fF
C108 sky130_fd_sc_hd__buf_2_0/A 0 -127.11fF
C109 sky130_fd_sc_hd__buf_2_1/A 0 -211.82fF
C110 VDD 0 -582.64fF
C111 clk 0 68.21fF
C112 sky130_fd_sc_hd__buf_2_1/a_27_47# 0 0.15fF
C113 sky130_fd_sc_hd__buf_2_0/a_27_47# 0 0.15fF
C114 outp 0 26.35fF
C115 sky130_fd_sc_hd__buf_2_0/X 0 43.25fF
C116 sky130_fd_sc_hd__nand2_4_1/a_27_47# 0 0.06fF
C117 sky130_fd_sc_hd__buf_2_1/X 0 23.78fF
C118 sky130_fd_sc_hd__nand2_4_0/a_27_47# 0 0.06fF
.ends

.subckt sky130_fd_pr__nfet_01v8_CFEPS5 a_n275_n238# a_n129_n152# a_n173_n64#
X0 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=8.32e+11p pd=7.76e+06u as=0p ps=0u w=650000u l=150000u
X1 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_n173_n64# a_n129_n152# a_n173_n64# a_n275_n238# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 a_n129_n152# a_n173_n64# 0.38fF
C1 a_n173_n64# a_n275_n238# 0.40fF
C2 a_n129_n152# a_n275_n238# 0.60fF
.ends

.subckt analog_top ip in rst_n i_bias_1 i_bias_2 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1
+ debug op a_probe_0 a_probe_1 a_probe_2 a_probe_3 clk d_probe_0 d_probe_1 d_probe_2
+ d_probe_3 d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1
+ VDD VSS
Xesd_cell_5 a_probe_0 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_2 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_18 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_29 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_20 ota_1/p1 VDD transmission_gate_20/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_21/in ota_1/cm VSS ota_1/p1_b transmission_gate
Xtransmission_gate_31 clock_v2_0/p1d VDD transmission_gate_31/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ip transmission_gate_31/out VSS clock_v2_0/p1d_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_70 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_19 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_21 ota_1/p2 VDD transmission_gate_21/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_21/in ota_1/in VSS ota_1/p2_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_3 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_10 transmission_gate_26/en VDD transmission_gate_10/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_w_test_0/cm transmission_gate_5/in VSS rst_n transmission_gate
Xesd_cell_6 a_probe_3 VSS VDD esd_cell
Xtransmission_gate_32 clock_v2_0/p1d VDD transmission_gate_32/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in transmission_gate_32/out VSS clock_v2_0/p1d_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_71 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_60 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_4 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_22 ota_1/p2 VDD transmission_gate_22/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_23/in ota_1/ip VSS ota_1/p2_b transmission_gate
Xtransmission_gate_11 transmission_gate_26/en VDD transmission_gate_11/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_w_test_0/cm transmission_gate_6/in VSS rst_n transmission_gate
Xota_w_test_0 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# ota_w_test_0/m1_12118_n9704#
+ ota_w_test_0/m1_12410_n9718# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580#
+ ota_w_test_0/m1_11356_n10481# ota_w_test_0/m1_11063_n10490# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_w_test_0/m1_11940_n10482#
+ ota_w_test_0/m1_12232_n10488# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580#
+ ota_w_test_0/m1_11825_n9711# ota_w_test_0/m1_11534_n9706# ota_w_test_0/m1_11242_n9716#
+ ota_w_test_0/m1_n6302_n3889# ota_w_test_0/on ota_w_test_0/sc_cmfb_0/transmission_gate_8/in
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# ota_1/p2_b ota_w_test_0/m1_11648_n10486#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# ota_w_test_0/sc_cmfb_0/transmission_gate_6/in
+ ota_w_test_0/ip ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580#
+ ota_w_test_0/m1_2462_n3318# ota_w_test_0/m1_n208_n2883# ota_w_test_0/cm ota_w_test_0/in
+ ota_w_test_0/m1_2463_n5585# ota_w_test_0/sc_cmfb_0/transmission_gate_3/out ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# ota_w_test_0/m1_n1659_n11581#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# ota_w_test_0/m1_6690_n8907#
+ ota_w_test_0/sc_cmfb_0/transmission_gate_9/in ota_1/p1_b ota_w_test_0/sc_cmfb_0/transmission_gate_4/out
+ ota_w_test_0/m1_n2176_n12171# i_bias_1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480#
+ ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# a_mux4_en_1/in1 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in
+ VDD a_mux4_en_0/in0 ota_w_test_0/m1_1038_n2886# ota_w_test_0/op ota_1/p2 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580#
+ ota_w_test_0/m1_n5574_n13620# ota_w_test_0/m1_n947_n12836# ota_1/p1 a_mux4_en_1/in2
+ a_mux4_en_0/in1 a_mux4_en_0/in2 ota_w_test
Xesd_cell_7 a_probe_2 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_50 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_61 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_23 ota_1/p1 VDD transmission_gate_23/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_23/in ota_1/cm VSS ota_1/p1_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_5 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_12 clock_v2_0/Ad VDD transmission_gate_12/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_w_test_0/op transmission_gate_17/in VSS clock_v2_0/Ad_b transmission_gate
Xsky130_fd_sc_hd__clkinv_16_0 sky130_fd_sc_hd__clkinv_4_1/Y VSS VDD d_probe_3 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_51 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_62 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_40 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_6 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_24 transmission_gate_26/en VDD transmission_gate_24/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_1/cm ota_1/ip VSS rst_n transmission_gate
Xtransmission_gate_13 clock_v2_0/Bd VDD transmission_gate_13/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_w_test_0/op transmission_gate_18/in VSS clock_v2_0/Bd_b transmission_gate
Xsky130_fd_sc_hd__clkinv_16_1 sky130_fd_sc_hd__clkinv_4_2/Y VSS VDD d_probe_2 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_52 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_63 transmission_gate_21/in transmission_gate_19/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_30 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_41 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_25 transmission_gate_26/en VDD transmission_gate_25/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_1/cm ota_1/in VSS rst_n transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_7 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_14 clock_v2_0/Bd VDD transmission_gate_14/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_w_test_0/on transmission_gate_17/in VSS clock_v2_0/Bd_b transmission_gate
Xsky130_fd_sc_hd__clkinv_16_2 sky130_fd_sc_hd__clkinv_4_3/Y VSS VDD d_probe_1 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_20 transmission_gate_23/in transmission_gate_32/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_64 transmission_gate_21/in transmission_gate_31/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_31 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_42 sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_53 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_0 rst_n VSS VDD transmission_gate_26/en sky130_fd_sc_hd__clkinv_4_0/w_82_21#
+ VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_26 transmission_gate_26/en VDD transmission_gate_26/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_1/on ota_1/op VSS rst_n transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_8 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_15 clock_v2_0/Ad VDD transmission_gate_15/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ota_w_test_0/on transmission_gate_18/in VSS clock_v2_0/Ad_b transmission_gate
Xsky130_fd_sc_hd__clkinv_16_3 sky130_fd_sc_hd__clkinv_4_4/Y VSS VDD d_probe_0 VSS
+ VDD sky130_fd_sc_hd__clkinv_16
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_65 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_21 transmission_gate_23/in transmission_gate_19/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_43 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_10 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_32 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_54 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_1 sky130_fd_sc_hd__mux4_1_0/X VSS VDD sky130_fd_sc_hd__clkinv_4_1/Y
+ sky130_fd_sc_hd__clkinv_4_1/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_9 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_27 clock_v2_0/p2_b VDD transmission_gate_27/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ onebit_dac_1/out transmission_gate_31/out VSS clock_v2_0/p2 transmission_gate
Xtransmission_gate_16 transmission_gate_26/en VDD transmission_gate_16/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_18/in transmission_gate_17/in VSS rst_n transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_22 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_11 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_66 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_44 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_55 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_33 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_2 sky130_fd_sc_hd__mux4_1_1/X VSS VDD sky130_fd_sc_hd__clkinv_4_2/Y
+ sky130_fd_sc_hd__clkinv_4_2/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_28 clock_v2_0/p2_b VDD transmission_gate_28/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ onebit_dac_1/out transmission_gate_0/out VSS clock_v2_0/p2 transmission_gate
Xtransmission_gate_17 clock_v2_0/p1d VDD transmission_gate_17/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_17/in transmission_gate_19/out VSS clock_v2_0/p1d_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_67 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_12 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_45 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_34 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_23 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_56 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xonebit_dac_0 VDD op onebit_dac_1/v_b onebit_dac_0/out VDD VSS VSS onebit_dac
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_0 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__clkinv_4_3 sky130_fd_sc_hd__mux4_1_2/X VSS VDD sky130_fd_sc_hd__clkinv_4_3/Y
+ sky130_fd_sc_hd__clkinv_4_3/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_29 clock_v2_0/p2_b VDD transmission_gate_29/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ onebit_dac_0/out transmission_gate_32/out VSS clock_v2_0/p2 transmission_gate
Xtransmission_gate_18 clock_v2_0/p1d VDD transmission_gate_18/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_18/in transmission_gate_19/in VSS clock_v2_0/p1d_b transmission_gate
Xota_1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480#
+ ota_1/m1_11825_n9711# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# ota_1/m1_12118_n9704# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# ota_1/m1_12410_n9718# ota_1/m1_n6302_n3889#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480#
+ ota_1/sc_cmfb_0/transmission_gate_9/in ota_1/m1_2463_n5585# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580#
+ ota_1/m1_n947_n12836# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480# ota_1/m1_11534_n9706#
+ ota_1/m1_11242_n9716# ota_1/m1_n2176_n12171# ota_1/sc_cmfb_0/transmission_gate_8/in
+ ota_1/sc_cmfb_0/transmission_gate_4/out ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580#
+ ota_1/p2_b ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# ota_1/sc_cmfb_0/transmission_gate_6/in
+ ota_1/ip ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_1/m1_2462_n3318# ota_1/cm
+ ota_1/m1_n208_n2883# ota_1/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580#
+ VSS ota_1/m1_6690_n8907# ota_1/p1_b i_bias_2 ota_1/m1_n5574_n13620# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480#
+ ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# ota_1/sc_cmfb_0/transmission_gate_7/in
+ ota_1/bias_a ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/bias_b ota_1/bias_d ota_1/op
+ ota_1/p2 ota_1/m1_1038_n2886# VDD ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580#
+ ota_1/cmc ota_1/bias_c ota_1/p1 ota_1/on ota_1/m1_n1659_n11581# ota
Xa_mux2_en_0 a_mux2_en_0/transmission_gate_1/en_b a_mux2_en_0/switch_5t_0/in a_mux2_en_0/switch_5t_1/transmission_gate_1/in
+ VDD a_mux2_en_0/switch_5t_0/transmission_gate_1/in ota_w_test_0/op a_mod_grp_ctrl_0
+ a_probe_0 debug a_mux2_en_0/switch_5t_1/in VSS ota_w_test_0/on a_mux2_en_0/switch_5t_1/en
+ a_mux2_en
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_13 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_68 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_46 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_57 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_24 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xonebit_dac_1 VDD op onebit_dac_1/v_b onebit_dac_1/out VSS VDD VSS onebit_dac
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_35 sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__clkinv_4_4 sky130_fd_sc_hd__mux4_1_3/X VSS VDD sky130_fd_sc_hd__clkinv_4_4/Y
+ sky130_fd_sc_hd__clkinv_4_4/w_82_21# VSS VDD sky130_fd_sc_hd__clkinv_4
Xtransmission_gate_19 clock_v2_0/p2_b VDD transmission_gate_19/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_19/in transmission_gate_19/out VSS clock_v2_0/p2 transmission_gate
Xa_mux2_en_1 a_mux2_en_1/transmission_gate_1/en_b a_mux2_en_1/switch_5t_0/in a_mux2_en_1/switch_5t_1/transmission_gate_1/in
+ VDD a_mux2_en_1/switch_5t_0/transmission_gate_1/in ota_1/op a_mod_grp_ctrl_0 a_probe_1
+ debug a_mux2_en_1/switch_5t_1/in VSS ota_1/on a_mux2_en_1/switch_5t_1/en a_mux2_en
Xsky130_fd_sc_hd__mux4_1_0 ota_1/p2_b clock_v2_0/Bd ota_1/p2 clock_v2_0/Bd_b d_clk_grp_2_ctrl_0
+ d_clk_grp_2_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_27_413#
+ sky130_fd_sc_hd__mux4_1_0/a_923_363# sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__mux4_1_0/a_834_97#
+ sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_193_413#
+ sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_69 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_47 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_58 transmission_gate_21/in transmission_gate_19/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_14 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_25 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__pfet_01v8_hvt_XAYTAL_0 onebit_dac_1/v_b VDD VDD VSS sky130_fd_pr__pfet_01v8_hvt_XAYTAL
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_36 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_2 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__mux4_1_1 clock_v2_0/p1d clock_v2_0/Ad clock_v2_0/p1d_b clock_v2_0/Ad_b
+ d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_1/X sky130_fd_sc_hd__mux4_1_1/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_1/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_27_413#
+ sky130_fd_sc_hd__mux4_1_1/a_923_363# sky130_fd_sc_hd__mux4_1_1/a_193_47# sky130_fd_sc_hd__mux4_1_1/a_834_97#
+ sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_193_413#
+ sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_26 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_48 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_15 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_59 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_3 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_37 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_sc_hd__mux4_1_2 clock_v2_0/p2 clock_v2_0/B clock_v2_0/p2_b clock_v2_0/B_b
+ d_clk_grp_1_ctrl_0 d_clk_grp_1_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_27_413#
+ sky130_fd_sc_hd__mux4_1_2/a_923_363# sky130_fd_sc_hd__mux4_1_2/a_193_47# sky130_fd_sc_hd__mux4_1_2/a_834_97#
+ sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_193_413#
+ sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_27 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_49 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_16 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_38 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_4 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_0 clock_v2_0/p1d VDD transmission_gate_0/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ ip transmission_gate_0/out VSS clock_v2_0/p1d_b transmission_gate
Xsky130_fd_sc_hd__mux4_1_3 ota_1/p1 clock_v2_0/A ota_1/p1_b clock_v2_0/A_b d_clk_grp_1_ctrl_0
+ d_clk_grp_1_ctrl_1 VSS VDD sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_277_47#
+ VSS VDD sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_27_413#
+ sky130_fd_sc_hd__mux4_1_3/a_923_363# sky130_fd_sc_hd__mux4_1_3/a_193_47# sky130_fd_sc_hd__mux4_1_3/a_834_97#
+ sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_193_413#
+ sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_17 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_28 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_39 ota_1/op ota_1/in VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_5 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_18 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_29 ota_1/on ota_1/ip VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_1 ota_1/p2 VDD transmission_gate_1/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_8/in transmission_gate_5/in VSS ota_1/p2_b transmission_gate
Xclock_v2_0 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/A clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_439_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_561_413# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X clock_v2_0/sky130_fd_sc_hd__mux2_1_0/X
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# clock_v2_0/p2_b clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_14/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_10/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315#
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X clock_v2_0/sky130_fd_sc_hd__clkbuf_16_8/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47#
+ clock_v2_0/Ad_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_4/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47#
+ clock_v2_0/A_b clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A clock_v2_0/sky130_fd_sc_hd__clkbuf_16_0/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_15/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/A
+ clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_11/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X clock_v2_0/Bd clock_v2_0/p1d_b
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1017_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_1/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_9/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_193_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkbuf_16_5/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_891_413#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B clock_v2_0/sky130_fd_sc_hd__clkbuf_16_1/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# ota_1/p2_b clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S
+ clock_v2_0/Ad clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_592_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_975_413# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_12/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_381_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y
+ clock_v2_0/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_466_413# clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y
+ clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/X
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X clock_v2_0/sky130_fd_sc_hd__nand2_1_4/a_113_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# ota_1/p1 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47#
+ ota_1/p1_b clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/X clock_v2_0/sky130_fd_sc_hd__clkbuf_16_6/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkbuf_16_2/a_110_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/A clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# clock_v2_0/B clock_v2_0/p1d
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_13/a_110_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_381_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/A
+ clk clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/X clock_v2_0/sky130_fd_sc_hd__nand2_1_0/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/A
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/X
+ ota_1/p2 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X clock_v2_0/B_b clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_634_159#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_2/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A
+ clock_v2_0/p2 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47#
+ clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/A
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47#
+ clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/X
+ clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A
+ clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/A
+ VDD VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y
+ clock_v2
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_6 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_2 clock_v2_0/p1d VDD transmission_gate_2/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ in transmission_gate_2/out VSS clock_v2_0/p1d_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_19 transmission_gate_23/in transmission_gate_19/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_7 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_3 clock_v2_0/A VDD transmission_gate_3/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_5/in ota_w_test_0/in VSS clock_v2_0/A_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_8 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_4 clock_v2_0/B VDD transmission_gate_4/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_6/in ota_w_test_0/in VSS clock_v2_0/B_b transmission_gate
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_9 sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xtransmission_gate_5 clock_v2_0/B VDD transmission_gate_5/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_5/in ota_w_test_0/ip VSS clock_v2_0/B_b transmission_gate
Xtransmission_gate_6 clock_v2_0/A VDD transmission_gate_6/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_6/in ota_w_test_0/ip VSS clock_v2_0/A_b transmission_gate
Xtransmission_gate_7 ota_1/p2 VDD transmission_gate_7/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_9/in transmission_gate_6/in VSS ota_1/p2_b transmission_gate
Xtransmission_gate_8 ota_1/p1 VDD transmission_gate_8/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_8/in ota_w_test_0/cm VSS ota_1/p1_b transmission_gate
Xtransmission_gate_9 ota_1/p1 VDD transmission_gate_9/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ transmission_gate_9/in ota_w_test_0/cm VSS ota_1/p1_b transmission_gate
Xa_mux4_en_0 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_2/a_113_47# a_mux4_en_0/switch_5t_1/transmission_gate_1/in
+ a_mux4_en_0/switch_5t_3/en a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y a_mux4_en_0/switch_5t_2/en_b
+ a_mux4_en_0/switch_5t_0/en a_mux4_en_0/sky130_fd_sc_hd__nand2_1_3/a_113_47# a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y
+ a_mux4_en_0/switch_5t_2/in a_mux4_en_0/switch_5t_0/transmission_gate_1/in a_mux4_en_0/switch_5t_2/transmission_gate_1/in
+ a_mux4_en_0/switch_5t_3/transmission_gate_1/in a_mux4_en_0/sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ a_mux4_en_0/transmission_gate_3/en_b a_mux4_en_0/switch_5t_1/en_b a_mux4_en_0/in3
+ a_mux4_en_0/switch_5t_2/en a_mux4_en_0/switch_5t_3/in a_mux4_en_0/in2 debug a_mod_grp_ctrl_1
+ a_mux4_en_0/in0 a_mux4_en_0/switch_5t_0/en_b a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_0/in
+ a_mux4_en_0/switch_5t_1/in a_probe_3 a_mux4_en_0/in1 VDD a_mux4_en_0/switch_5t_3/en_b
+ a_mux4_en_0/sky130_fd_sc_hd__nand2_1_1/a_113_47# a_mux4_en_0/switch_5t_1/en VSS
+ a_mux4_en
Xa_mux4_en_1 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_2/a_113_47# a_mux4_en_1/switch_5t_1/transmission_gate_1/in
+ a_mux4_en_1/switch_5t_3/en a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y a_mux4_en_1/switch_5t_2/en_b
+ a_mux4_en_1/switch_5t_0/en a_mux4_en_1/sky130_fd_sc_hd__nand2_1_3/a_113_47# a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y
+ a_mux4_en_1/switch_5t_2/in a_mux4_en_1/switch_5t_0/transmission_gate_1/in a_mux4_en_1/switch_5t_2/transmission_gate_1/in
+ a_mux4_en_1/switch_5t_3/transmission_gate_1/in a_mux4_en_1/sky130_fd_sc_hd__nand2_1_0/a_113_47#
+ a_mux4_en_1/transmission_gate_3/en_b a_mux4_en_1/switch_5t_1/en_b a_mux4_en_1/in3
+ a_mux4_en_1/switch_5t_2/en a_mux4_en_1/switch_5t_3/in a_mux4_en_1/in2 debug a_mod_grp_ctrl_1
+ ota_w_test_0/cm a_mux4_en_1/switch_5t_0/en_b a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_0/in
+ a_mux4_en_1/switch_5t_1/in a_probe_2 a_mux4_en_1/in1 VDD a_mux4_en_1/switch_5t_3/en_b
+ a_mux4_en_1/sky130_fd_sc_hd__nand2_1_1/a_113_47# a_mux4_en_1/switch_5t_1/en VSS
+ a_mux4_en
Xsky130_fd_sc_hd__decap_4_0 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_40 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_1 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_30 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_41 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_2 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_42 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_20 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_31 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_32 transmission_gate_9/in transmission_gate_2/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_10 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_21 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_43 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_4 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_44 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_33 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_11 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_22 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_5 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_45 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_34 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_12 transmission_gate_8/in transmission_gate_0/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_23 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_TABSMU_0 ota_1/on VSS VSS sky130_fd_pr__cap_mim_m3_1_TABSMU
Xcomparator_v2_0 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# op onebit_dac_1/v_b
+ comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X comparator_v2_0/li_n2324_818# comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47#
+ comparator_v2_0/li_940_818# comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# VSS
+ comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X VDD ota_1/p1_b comparator_v2_0/li_940_3458#
+ ota_1/on comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47#
+ ota_1/op comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A comparator_v2
Xsky130_fd_sc_hd__decap_4_6 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_46 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_35 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_13 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_24 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_0 in VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_TABSMU_1 ota_1/op VSS VSS sky130_fd_pr__cap_mim_m3_1_TABSMU
Xsky130_fd_sc_hd__decap_4_7 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_47 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_36 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_25 sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_1 ip VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_14 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_sc_hd__decap_4_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_37 transmission_gate_9/in transmission_gate_2/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_15 transmission_gate_6/in transmission_gate_18/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_26 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__nfet_01v8_CFEPS5_0 VSS onebit_dac_1/v_b VSS sky130_fd_pr__nfet_01v8_CFEPS5
Xesd_cell_2 i_bias_2 VSS VDD esd_cell
Xsky130_fd_sc_hd__decap_4_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_0 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_38 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_16 transmission_gate_5/in transmission_gate_17/in
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_27 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_3 i_bias_1 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_17 transmission_gate_8/in transmission_gate_0/out
+ VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_28 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xsky130_fd_pr__cap_mim_m3_1_CGPBWM_39 sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980#
+ sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM
Xesd_cell_4 a_probe_1 VSS VDD esd_cell
Xsky130_fd_pr__cap_mim_m3_1_CEWQ64_1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210#
+ sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64
Xtransmission_gate_30 clock_v2_0/p2_b VDD transmission_gate_30/sky130_fd_pr__nfet_01v8_6J4AMR_0/w_n646_n262#
+ onebit_dac_0/out transmission_gate_2/out VSS clock_v2_0/p2 transmission_gate
C0 clock_v2_0/Ad_b ota_w_test_0/on 0.34fF
C1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# ota_1/p1_b 0.03fF
C2 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/B 0.01fF
C3 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.09fF
C4 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y -0.00fF
C5 transmission_gate_8/in VDD 0.11fF
C6 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# -0.00fF
C7 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.35fF
C8 ota_1/ip ota_1/on 1.75fF
C9 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.12fF
C10 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C11 sky130_fd_sc_hd__mux4_1_3/a_27_47# clock_v2_0/p2 0.00fF
C12 VSS sky130_fd_sc_hd__mux4_1_1/X 0.58fF
C13 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/X 0.02fF
C14 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# -0.26fF
C15 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.08fF
C16 VSS sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.01fF
C17 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.01fF
C18 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# -0.00fF
C19 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# VDD 0.00fF
C20 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0.03fF
C21 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0.08fF
C22 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# -0.00fF
C23 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# ota_1/on 0.03fF
C24 transmission_gate_9/in VSS 0.98fF
C25 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# VDD 0.08fF
C26 clock_v2_0/Ad clock_v2_0/p2_b 0.04fF
C27 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clk 0.00fF
C28 sky130_fd_sc_hd__mux4_1_3/a_750_97# ota_1/p1_b 0.11fF
C29 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.02fF
C30 ota_w_test_0/cm transmission_gate_6/in 0.37fF
C31 a_mux4_en_0/switch_5t_0/en a_mux4_en_0/switch_5t_0/transmission_gate_1/in 0.00fF
C32 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.01fF
C33 rst_n clock_v2_0/p1d 0.22fF
C34 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_2/in -0.00fF
C35 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/A -0.05fF
C36 sky130_fd_sc_hd__mux4_1_0/a_247_21# d_clk_grp_2_ctrl_0 0.09fF
C37 sky130_fd_sc_hd__mux4_1_3/a_834_97# clock_v2_0/A_b 0.01fF
C38 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# 0.67fF
C39 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/c1_n260_n210# -0.09fF
C40 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# VDD 0.00fF
C41 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.05fF
C42 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0.06fF
C43 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.00fF
C44 VSS sky130_fd_sc_hd__mux4_1_0/a_277_47# -0.65fF
C45 a_mux4_en_0/switch_5t_1/transmission_gate_1/in VDD -0.23fF
C46 a_mux4_en_0/in0 clock_v2_0/A 0.04fF
C47 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# -0.00fF
C48 VDD a_mux4_en_0/switch_5t_3/in 0.38fF
C49 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.00fF
C50 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0.05fF
C51 ota_w_test_0/cm ota_1/p2_b 0.12fF
C52 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# -0.00fF
C53 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C54 transmission_gate_19/in ota_1/p2_b 0.29fF
C55 clock_v2_0/A ota_w_test_0/in 0.25fF
C56 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.05fF
C57 ota_w_test_0/m1_2463_n5585# ota_w_test_0/m1_2462_n3318# 0.01fF
C58 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.00fF
C59 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# transmission_gate_19/in 0.03fF
C60 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# 0.03fF
C61 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0.09fF
C62 ota_1/p1 ota_1/sc_cmfb_0/transmission_gate_4/out -0.00fF
C63 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 1.70fF
C64 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_1/op 0.07fF
C65 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VDD 0.00fF
C66 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# 0.00fF
C67 transmission_gate_9/in transmission_gate_6/in 2.41fF
C68 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480# ota_1/p1_b 0.04fF
C69 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# -0.14fF
C70 i_bias_2 ota_1/m1_1038_n2886# -0.01fF
C71 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# -0.21fF
C72 comparator_v2_0/li_n2324_818# ota_1/p1_b -0.01fF
C73 transmission_gate_19/in ota_1/in 0.05fF
C74 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0.00fF
C75 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0.00fF
C76 VDD a_mod_grp_ctrl_1 5.27fF
C77 clock_v2_0/Bd_b clock_v2_0/Ad 14.60fF
C78 ota_w_test_0/cm ota_1/p2 0.14fF
C79 transmission_gate_19/in ota_1/p2 0.22fF
C80 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0.05fF
C81 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0.00fF
C82 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.00fF
C83 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_13/a_110_47# VDD 0.14fF
C84 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_1/X 0.01fF
C85 VSS ota_1/m1_n208_n2883# 0.15fF
C86 transmission_gate_9/in ota_1/p2_b 0.07fF
C87 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.00fF
C88 VSS clk 8.65fF
C89 clock_v2_0/Ad a_mod_grp_ctrl_0 0.05fF
C90 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.09fF
C91 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.06fF
C92 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C93 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# clock_v2_0/p1d 0.04fF
C94 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y VDD 0.08fF
C95 a_mux4_en_1/in1 clock_v2_0/B_b 0.04fF
C96 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.03fF
C97 i_bias_1 clock_v2_0/B_b 1.65fF
C98 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C99 sky130_fd_sc_hd__mux4_1_2/a_1478_413# d_probe_1 0.00fF
C100 clock_v2_0/Ad_b a_mod_grp_ctrl_1 0.06fF
C101 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C102 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.03fF
C103 sky130_fd_sc_hd__mux4_1_0/a_277_47# ota_1/p2_b 0.01fF
C104 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/c1_n260_n210# 0.03fF
C105 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# 0.27fF
C106 clock_v2_0/A_b transmission_gate_5/in 0.44fF
C107 transmission_gate_9/in ota_1/p2 0.01fF
C108 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# 0.09fF
C109 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.03fF
C110 d_probe_2 d_probe_3 0.40fF
C111 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.00fF
C112 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.00fF
C113 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_14/a_110_47# -0.00fF
C114 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.06fF
C115 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.01fF
C116 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# -0.00fF
C117 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0.21fF
C118 rst_n ota_w_test_0/in 0.00fF
C119 transmission_gate_26/en clock_v2_0/A 0.19fF
C120 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# -0.00fF
C121 a_probe_0 a_mod_grp_ctrl_0 0.00fF
C122 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/X -0.00fF
C123 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# VSS 0.41fF
C124 sky130_fd_sc_hd__mux4_1_0/a_277_47# ota_1/p2 0.03fF
C125 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.02fF
C126 ota_w_test_0/op clock_v2_0/Ad 1.32fF
C127 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# 0.22fF
C128 i_bias_2 debug 0.20fF
C129 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0.12fF
C130 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.00fF
C131 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0.09fF
C132 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# clock_v2_0/p1d_b 0.01fF
C133 ota_1/ip ota_1/cm 0.44fF
C134 clock_v2_0/Bd ota_1/p1_b 0.46fF
C135 clock_v2_0/A_b clock_v2_0/B 12.56fF
C136 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.10fF
C137 clock_v2_0/p1d_b a_mod_grp_ctrl_1 0.07fF
C138 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/X -0.00fF
C139 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.00fF
C140 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# -0.00fF
C141 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# ota_1/p1_b 0.09fF
C142 ota_1/m1_n208_n2883# ota_1/in 0.00fF
C143 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.06fF
C144 ota_w_test_0/cm VDD 5.05fF
C145 sky130_fd_sc_hd__mux4_1_3/a_757_363# d_clk_grp_1_ctrl_0 0.00fF
C146 transmission_gate_19/in VDD 0.23fF
C147 VSS clock_v2_0/A_b 1.37fF
C148 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# -0.00fF
C149 a_mux4_en_0/switch_5t_0/in a_mod_grp_ctrl_1 -0.00fF
C150 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# ota_1/p1_b 0.01fF
C151 comparator_v2_0/li_n2324_818# comparator_v2_0/li_940_818# 0.00fF
C152 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0.00fF
C153 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/c1_n260_n210# 0.03fF
C154 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.00fF
C155 ota_1/p2_b sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C156 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0.00fF
C157 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0.00fF
C158 sky130_fd_sc_hd__mux4_1_0/a_757_363# d_clk_grp_2_ctrl_0 -0.00fF
C159 clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y 0.00fF
C160 sky130_fd_sc_hd__mux4_1_1/X VDD 0.71fF
C161 ota_w_test_0/m1_2462_n3318# ota_w_test_0/in 0.00fF
C162 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0.05fF
C163 transmission_gate_26/en rst_n 10.08fF
C164 sky130_fd_sc_hd__mux4_1_2/a_27_413# VDD 0.07fF
C165 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0.08fF
C166 VSS a_mux4_en_1/switch_5t_0/en 0.54fF
C167 ota_w_test_0/cm clock_v2_0/Ad_b 0.06fF
C168 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# -0.00fF
C169 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X -0.01fF
C170 transmission_gate_9/in VDD -0.09fF
C171 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# 0.04fF
C172 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X -0.00fF
C173 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_757_363# 0.01fF
C174 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A -0.01fF
C175 ip clock_v2_0/p1d 0.19fF
C176 ota_1/bias_a ota_1/cm 0.00fF
C177 sky130_fd_sc_hd__mux4_1_1/X clock_v2_0/Ad_b 0.00fF
C178 transmission_gate_6/in clock_v2_0/A_b 0.55fF
C179 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0.00fF
C180 onebit_dac_1/v_b transmission_gate_2/out 0.03fF
C181 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# -0.00fF
C182 sky130_fd_sc_hd__mux4_1_0/a_277_47# VDD 0.11fF
C183 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0.14fF
C184 VSS sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.13fF
C185 VSS a_mux4_en_0/sky130_fd_sc_hd__nand2_1_3/a_113_47# 0.00fF
C186 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# VDD -0.00fF
C187 transmission_gate_2/out in 0.01fF
C188 VSS a_mux4_en_1/sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C189 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# -0.00fF
C190 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.08fF
C191 ota_1/p2_b clock_v2_0/A_b 0.05fF
C192 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# -0.00fF
C193 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C194 ota_1/p1_b clock_v2_0/p1d 3.85fF
C195 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# -0.12fF
C196 VSS sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.01fF
C197 a_mod_grp_ctrl_0 a_mux2_en_0/transmission_gate_1/en_b 0.07fF
C198 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.02fF
C199 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# ota_w_test_0/on -0.00fF
C200 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X -0.00fF
C201 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# VSS 0.38fF
C202 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_1/X 0.05fF
C203 sky130_fd_sc_hd__mux4_1_0/a_277_47# clock_v2_0/Ad_b 0.00fF
C204 a_mux4_en_0/switch_5t_3/en a_mux4_en_0/switch_5t_3/in 0.00fF
C205 transmission_gate_19/in clock_v2_0/p1d_b 0.11fF
C206 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# -0.38fF
C207 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0.59fF
C208 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/A -0.00fF
C209 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C210 ota_1/p2 clock_v2_0/A_b 0.06fF
C211 ota_1/m1_n208_n2883# VDD 3.75fF
C212 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# 0.04fF
C213 VDD clk 2.53fF
C214 a_mux4_en_1/in1 clock_v2_0/B 0.04fF
C215 d_clk_grp_1_ctrl_1 ota_1/p1_b 0.11fF
C216 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# 0.11fF
C217 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# 0.00fF
C218 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0.04fF
C219 i_bias_1 clock_v2_0/B 0.11fF
C220 sky130_fd_sc_hd__mux4_1_1/X clock_v2_0/p1d_b 0.01fF
C221 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0.05fF
C222 a_mux4_en_1/in2 clock_v2_0/Ad 0.03fF
C223 ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# 0.24fF
C224 transmission_gate_32/out clock_v2_0/p2_b 0.21fF
C225 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.03fF
C226 transmission_gate_18/in clock_v2_0/Ad 0.37fF
C227 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n930_n880# 0.11fF
C228 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_0/A 0.01fF
C229 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# 0.42fF
C230 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C231 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_193_47# 0.00fF
C232 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A -0.01fF
C233 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# -0.00fF
C234 VSS a_mux4_en_1/in1 2.68fF
C235 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0.12fF
C236 VSS i_bias_1 2.83fF
C237 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/X 0.01fF
C238 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_2/a_113_47# a_mod_grp_ctrl_1 0.00fF
C239 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# -0.00fF
C240 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.00fF
C241 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/sc_cmfb_0/transmission_gate_6/in 0.00fF
C242 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0.00fF
C243 ota_w_test_0/op a_mux2_en_0/transmission_gate_1/en_b 0.00fF
C244 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_14/a_110_47# VDD 0.12fF
C245 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# -0.34fF
C246 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.05fF
C247 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C248 sky130_fd_sc_hd__mux4_1_1/a_193_413# VDD 0.06fF
C249 debug a_mux4_en_0/switch_5t_3/en_b -0.00fF
C250 ota_w_test_0/op ota_w_test_0/m1_n1659_n11581# 0.00fF
C251 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.01fF
C252 transmission_gate_23/in transmission_gate_21/in 0.06fF
C253 a_mod_grp_ctrl_0 a_mux2_en_0/switch_5t_1/en 0.06fF
C254 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# clock_v2_0/p1d_b 0.33fF
C255 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# 0.19fF
C256 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y 0.00fF
C257 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C258 sky130_fd_sc_hd__mux4_1_0/a_277_47# clock_v2_0/p1d_b 0.00fF
C259 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0.00fF
C260 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# -0.00fF
C261 ota_1/p1 clock_v2_0/B_b 0.47fF
C262 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# 0.21fF
C263 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.12fF
C264 a_mux4_en_0/in0 ota_1/p1_b 0.04fF
C265 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C266 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.10fF
C267 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# 0.03fF
C268 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A -0.00fF
C269 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.00fF
C270 ota_1/p2 sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.03fF
C271 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# 0.00fF
C272 VSS a_mux4_en_0/switch_5t_3/transmission_gate_1/in 0.33fF
C273 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# VDD -0.00fF
C274 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y -0.00fF
C275 d_clk_grp_1_ctrl_0 clock_v2_0/B_b 0.02fF
C276 clock_v2_0/p1d in 0.43fF
C277 VSS a_mux4_en_0/switch_5t_0/en_b 0.30fF
C278 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.05fF
C279 clock_v2_0/p2 transmission_gate_2/out 0.04fF
C280 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0.00fF
C281 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# -0.34fF
C282 ota_1/bias_b ota_1/cm 0.36fF
C283 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# 0.09fF
C284 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# -0.00fF
C285 sky130_fd_sc_hd__mux4_1_2/a_668_97# clock_v2_0/B_b -0.02fF
C286 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C287 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# VDD 0.73fF
C288 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0.04fF
C289 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# 1.58fF
C290 clock_v2_0/Ad sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.01fF
C291 VSS sky130_fd_sc_hd__mux4_1_1/a_193_47# -0.00fF
C292 VDD clock_v2_0/A_b 2.65fF
C293 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# clock_v2_0/p1d_b 0.01fF
C294 sky130_fd_sc_hd__mux4_1_3/a_277_47# ota_1/p1_b 0.04fF
C295 ota_1/ip transmission_gate_32/out 0.75fF
C296 clock_v2_0/Bd clock_v2_0/p2 0.04fF
C297 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# 0.05fF
C298 clock_v2_0/Ad ota_w_test_0/on 0.32fF
C299 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# 0.12fF
C300 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in ota_w_test_0/sc_cmfb_0/transmission_gate_8/in -0.04fF
C301 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# -0.00fF
C302 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# VDD -0.00fF
C303 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/c1_n260_n210# 0.03fF
C304 ota_1/p1 ota_1/m1_n2176_n12171# 0.16fF
C305 VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# 0.23fF
C306 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.03fF
C307 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0.00fF
C308 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0.00fF
C309 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# ota_1/ip 0.03fF
C310 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n930_n880# transmission_gate_17/in 0.11fF
C311 sky130_fd_sc_hd__mux4_1_2/a_757_363# clock_v2_0/B_b 0.00fF
C312 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# -0.00fF
C313 ota_1/m1_n1659_n11581# ota_1/p1_b 0.08fF
C314 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# -0.00fF
C315 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0.09fF
C316 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# 0.03fF
C317 transmission_gate_19/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# 0.04fF
C318 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_1/in 0.01fF
C319 a_mux4_en_1/switch_5t_0/en VDD -0.59fF
C320 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/Bd 0.00fF
C321 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# 0.11fF
C322 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A 0.10fF
C323 debug a_mux4_en_1/switch_5t_2/in 0.01fF
C324 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# 0.09fF
C325 a_mux4_en_1/switch_5t_1/en_b a_mux4_en_1/switch_5t_0/en_b 0.00fF
C326 clock_v2_0/Ad_b clock_v2_0/A_b 0.58fF
C327 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# 0.03fF
C328 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C329 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C330 sky130_fd_sc_hd__mux4_1_1/a_193_413# clock_v2_0/p1d_b 0.06fF
C331 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0.01fF
C332 VSS a_mux4_en_0/sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C333 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# -0.00fF
C334 ota_1/bias_c ota_1/cm 0.10fF
C335 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# 0.03fF
C336 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_1/bias_a 0.08fF
C337 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0.30fF
C338 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 0.30fF
C339 clock_v2_0/Bd_b clock_v2_0/p2_b 0.07fF
C340 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0.08fF
C341 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.31fF
C342 transmission_gate_26/en ota_1/p1_b 0.67fF
C343 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_2/B 0.01fF
C344 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# 0.03fF
C345 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# transmission_gate_5/in 0.80fF
C346 a_mod_grp_ctrl_0 clock_v2_0/p2_b 0.04fF
C347 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210# 0.03fF
C348 sky130_fd_sc_hd__mux4_1_2/a_1290_413# clock_v2_0/p2 0.00fF
C349 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.00fF
C350 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.00fF
C351 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# -0.00fF
C352 sky130_fd_sc_hd__mux4_1_3/a_1478_413# VDD 0.20fF
C353 a_mod_grp_ctrl_0 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C354 VSS ota_1/sc_cmfb_0/transmission_gate_7/in 2.44fF
C355 a_mux2_en_0/switch_5t_0/in a_mux2_en_0/switch_5t_1/en 0.00fF
C356 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0.05fF
C357 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C358 a_mux4_en_0/switch_5t_2/in a_mod_grp_ctrl_1 -0.00fF
C359 transmission_gate_0/out onebit_dac_1/out 0.12fF
C360 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C361 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# -0.00fF
C362 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.00fF
C363 sky130_fd_sc_hd__mux4_1_0/a_193_413# VDD 0.02fF
C364 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.01fF
C365 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0.00fF
C366 a_mux4_en_0/switch_5t_0/en a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C367 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/c1_n260_n210# -0.08fF
C368 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# -0.09fF
C369 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.05fF
C370 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# 0.11fF
C371 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# -0.65fF
C372 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.07fF
C373 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# -0.38fF
C374 clock_v2_0/p1d_b clock_v2_0/A_b 0.07fF
C375 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# -0.00fF
C376 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# -0.00fF
C377 ota_1/p1 transmission_gate_5/in 0.07fF
C378 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# 0.06fF
C379 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y 0.07fF
C380 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C381 VSS ota_1/cmc 3.03fF
C382 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C383 clock_v2_0/p1d clock_v2_0/p2 1.44fF
C384 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# VDD 0.00fF
C385 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# 0.07fF
C386 clock_v2_0/Bd_b a_mod_grp_ctrl_0 0.04fF
C387 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.25fF
C388 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# -0.00fF
C389 VSS sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.08fF
C390 transmission_gate_19/in ota_1/on 0.01fF
C391 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_0/A 0.08fF
C392 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# VDD 0.18fF
C393 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# VDD 0.07fF
C394 ota_1/cmc ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.00fF
C395 a_mux4_en_1/in1 VDD 1.53fF
C396 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0.06fF
C397 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/p1d 0.01fF
C398 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210# ota_1/op 0.04fF
C399 clock_v2_0/Ad a_mod_grp_ctrl_1 0.06fF
C400 i_bias_1 VDD 3.61fF
C401 ota_1/sc_cmfb_0/transmission_gate_4/out ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.12fF
C402 ota_w_test_0/op ota_w_test_0/sc_cmfb_0/transmission_gate_6/in 0.01fF
C403 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# -0.00fF
C404 a_mux4_en_1/in2 a_mux4_en_1/in3 0.00fF
C405 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0.08fF
C406 VSS a_mux4_en_1/switch_5t_3/in 0.04fF
C407 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/p2_b -0.00fF
C408 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.07fF
C409 VSS onebit_dac_0/out 0.81fF
C410 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0.00fF
C411 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# clock_v2_0/p1d 0.27fF
C412 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# -0.00fF
C413 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/X 0.00fF
C414 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# VDD 0.03fF
C415 ota_1/p1 clock_v2_0/B 0.64fF
C416 clock_v2_0/Ad_b a_mux4_en_1/in1 0.04fF
C417 i_bias_1 clock_v2_0/Ad_b 0.08fF
C418 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0.00fF
C419 debug a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C420 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0.00fF
C421 VSS d_probe_2 1.87fF
C422 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C423 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/p2 0.00fF
C424 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0.01fF
C425 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# -0.00fF
C426 clock_v2_0/Bd_b ota_w_test_0/op 3.10fF
C427 ota_w_test_0/op ota_w_test_0/m1_6690_n8907# 0.04fF
C428 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C429 VSS ota_1/p1 10.67fF
C430 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# -0.00fF
C431 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_1/p1 0.09fF
C432 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0.10fF
C433 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480# -0.09fF
C434 ota_w_test_0/m1_n2176_n12171# ota_w_test_0/m1_n1659_n11581# 0.03fF
C435 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.08fF
C436 d_clk_grp_1_ctrl_0 clock_v2_0/B 0.01fF
C437 d_clk_grp_2_ctrl_1 sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.01fF
C438 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0.01fF
C439 VDD a_mux4_en_0/switch_5t_3/transmission_gate_1/in -1.31fF
C440 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0.00fF
C441 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.12fF
C442 a_probe_2 a_mux4_en_1/switch_5t_3/en -0.00fF
C443 ota_w_test_0/on a_mux2_en_0/transmission_gate_1/en_b 0.00fF
C444 ota_1/p2_b ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.01fF
C445 a_mux4_en_0/switch_5t_0/en_b VDD 0.17fF
C446 a_mux4_en_0/in1 debug 0.02fF
C447 ota_w_test_0/m1_n1659_n11581# ota_w_test_0/on 0.00fF
C448 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0.08fF
C449 sky130_fd_sc_hd__mux4_1_0/a_27_47# ota_1/p2_b -0.00fF
C450 VSS d_clk_grp_1_ctrl_0 1.63fF
C451 transmission_gate_18/in transmission_gate_32/out 0.01fF
C452 transmission_gate_17/in transmission_gate_5/in -2.67fF
C453 ota_1/cmc ota_1/p2 0.02fF
C454 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C455 a_mux4_en_1/switch_5t_0/in a_mux4_en_1/transmission_gate_3/en_b 0.00fF
C456 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0.06fF
C457 VSS sky130_fd_sc_hd__mux4_1_2/a_668_97# -0.23fF
C458 VSS d_clk_grp_2_ctrl_1 1.33fF
C459 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.04fF
C460 a_mux4_en_0/switch_5t_3/en_b a_mux4_en_0/switch_5t_2/en_b 0.00fF
C461 ota_1/p2 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.01fF
C462 a_mux4_en_1/switch_5t_3/en_b a_mux4_en_1/switch_5t_2/en_b 0.00fF
C463 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# 0.00fF
C464 transmission_gate_21/in ota_1/p1_b 0.09fF
C465 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0.12fF
C466 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C467 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# -0.00fF
C468 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A 0.09fF
C469 ota_1/sc_cmfb_0/transmission_gate_9/in ota_1/p1_b -0.00fF
C470 sky130_fd_sc_hd__mux4_1_2/a_757_363# VSS -0.00fF
C471 ota_w_test_0/cm clock_v2_0/Ad 1.62fF
C472 sky130_fd_sc_hd__mux4_1_1/a_193_47# clock_v2_0/Ad_b 0.00fF
C473 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0.17fF
C474 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.03fF
C475 ota_1/p1 ota_1/p2_b 2.51fF
C476 a_mod_grp_ctrl_0 a_mux2_en_0/switch_5t_0/in 0.02fF
C477 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# transmission_gate_17/in 0.11fF
C478 d_clk_grp_2_ctrl_0 clock_v2_0/B_b 0.03fF
C479 d_probe_2 sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.00fF
C480 i_bias_2 ota_1/p1_b 0.10fF
C481 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0.00fF
C482 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_2/B -0.04fF
C483 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# 0.11fF
C484 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480# 0.54fF
C485 a_mux4_en_0/in2 debug 0.02fF
C486 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# -0.13fF
C487 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# -0.00fF
C488 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# -0.00fF
C489 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_193_47# -0.00fF
C490 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/A_b 0.00fF
C491 ota_1/p1 ota_1/in 0.16fF
C492 ota_1/sc_cmfb_0/transmission_gate_7/in VDD 1.14fF
C493 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0.07fF
C494 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.00fF
C495 ota_1/p1 ota_1/p2 3.71fF
C496 VSS transmission_gate_17/in 3.89fF
C497 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0.08fF
C498 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# -0.00fF
C499 transmission_gate_26/en clock_v2_0/p2 0.07fF
C500 a_mux2_en_1/switch_5t_1/in debug -0.00fF
C501 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in a_mux4_en_1/in2 0.00fF
C502 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# -0.00fF
C503 ota_1/m1_n5574_n13620# ota_1/p1_b 0.12fF
C504 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0.00fF
C505 sky130_fd_sc_hd__mux4_1_1/a_1478_413# d_clk_grp_2_ctrl_1 0.00fF
C506 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0.08fF
C507 a_mux4_en_0/switch_5t_0/en_b a_mux4_en_0/switch_5t_0/in -0.00fF
C508 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# -0.00fF
C509 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.04fF
C510 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_381_47# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C511 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.01fF
C512 ota_1/cmc VDD 2.35fF
C513 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A -0.01fF
C514 ota_1/p2 d_clk_grp_2_ctrl_1 0.11fF
C515 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/op -0.01fF
C516 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# VDD 0.15fF
C517 sky130_fd_sc_hd__mux4_1_3/a_1290_413# clock_v2_0/A_b 0.01fF
C518 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/c1_n260_n210# ota_1/on 0.06fF
C519 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.09fF
C520 clock_v2_0/Bd_b a_mux4_en_1/in2 0.03fF
C521 a_mux4_en_1/in2 ota_w_test_0/m1_6690_n8907# 1.37fF
C522 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y -0.00fF
C523 sky130_fd_sc_hd__mux4_1_0/a_27_47# VDD 0.00fF
C524 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C525 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# ota_1/on 0.03fF
C526 clock_v2_0/Bd_b transmission_gate_18/in 0.09fF
C527 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C528 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.01fF
C529 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.03fF
C530 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# -0.09fF
C531 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/X 0.00fF
C532 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.09fF
C533 a_mux4_en_1/switch_5t_3/en a_mod_grp_ctrl_1 0.03fF
C534 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# -0.00fF
C535 a_mux4_en_0/in0 ota_w_test_0/m1_n947_n12836# 0.02fF
C536 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0.06fF
C537 VDD a_mux4_en_1/switch_5t_3/in 0.38fF
C538 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# -0.00fF
C539 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0.18fF
C540 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__clkinv_4_4/Y 0.00fF
C541 onebit_dac_0/out VDD 0.10fF
C542 transmission_gate_17/in ota_1/p2_b 0.12fF
C543 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# -0.00fF
C544 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# -0.31fF
C545 ota_1/cmc ota_1/op -0.09fF
C546 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X -0.00fF
C547 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# 0.32fF
C548 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210# 0.03fF
C549 VSS a_mux4_en_1/switch_5t_1/en 0.56fF
C550 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# VDD -0.00fF
C551 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.09fF
C552 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.03fF
C553 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.02fF
C554 a_mux4_en_0/in1 clock_v2_0/A 0.04fF
C555 a_mux2_en_1/switch_5t_1/en debug 0.00fF
C556 sky130_fd_sc_hd__mux4_1_3/a_247_21# ota_1/p1_b 0.06fF
C557 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0.01fF
C558 d_probe_2 VDD 2.50fF
C559 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.02fF
C560 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.20fF
C561 sky130_fd_sc_hd__mux4_1_2/a_834_97# clock_v2_0/A_b 0.00fF
C562 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.01fF
C563 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# 0.79fF
C564 ota_1/p2 transmission_gate_17/in 0.09fF
C565 transmission_gate_31/out onebit_dac_0/out 0.12fF
C566 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# 0.21fF
C567 ota_1/p1 VDD 16.36fF
C568 a_mux2_en_0/switch_5t_1/en a_mod_grp_ctrl_1 0.06fF
C569 ota_1/p1 sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C570 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in ota_w_test_0/on 0.03fF
C571 clock_v2_0/A ota_w_test_0/ip 0.44fF
C572 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0.00fF
C573 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0.00fF
C574 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.01fF
C575 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0.07fF
C576 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# ota_1/p1_b 0.02fF
C577 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.02fF
C578 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/p2_b 0.00fF
C579 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# -0.00fF
C580 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# 0.06fF
C581 ota_1/m1_n208_n2883# ota_1/cm 0.06fF
C582 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/c1_n260_n210# 0.03fF
C583 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# clock_v2_0/p2 0.03fF
C584 ota_w_test_0/op a_mux4_en_1/in2 -0.03fF
C585 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# ota_1/p1 0.02fF
C586 VSS comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X 0.00fF
C587 transmission_gate_18/in ota_w_test_0/op 0.03fF
C588 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# -0.00fF
C589 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.00fF
C590 d_clk_grp_1_ctrl_0 VDD 1.54fF
C591 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_193_413# -0.00fF
C592 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# -0.00fF
C593 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.03fF
C594 ota_1/p1 clock_v2_0/Ad_b 0.99fF
C595 debug clock_v2_0/B_b 0.07fF
C596 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# -0.00fF
C597 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# 0.00fF
C598 sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980# -0.38fF
C599 sky130_fd_sc_hd__mux4_1_2/a_668_97# VDD 0.01fF
C600 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C601 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# ota_1/on 0.06fF
C602 d_clk_grp_2_ctrl_1 VDD 3.48fF
C603 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# ota_1/p1_b 0.06fF
C604 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C605 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/X 0.00fF
C606 clock_v2_0/Bd_b ota_w_test_0/on 0.10fF
C607 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/p2 0.00fF
C608 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# 0.14fF
C609 ota_w_test_0/m1_6690_n8907# ota_w_test_0/on -0.01fF
C610 ota_1/p1 ota_1/op 0.44fF
C611 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y -0.00fF
C612 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# -0.00fF
C613 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C614 sky130_fd_sc_hd__mux4_1_2/a_757_363# VDD 0.04fF
C615 a_mux4_en_0/in2 clock_v2_0/A 0.04fF
C616 onebit_dac_0/out clock_v2_0/p1d_b 0.53fF
C617 a_mux4_en_0/transmission_gate_3/en_b a_mux4_en_0/switch_5t_2/en_b -0.00fF
C618 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.00fF
C619 clock_v2_0/Ad clock_v2_0/A_b 1.10fF
C620 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/A -0.72fF
C621 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C622 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# VDD -0.05fF
C623 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B 0.00fF
C624 clock_v2_0/Ad_b d_clk_grp_2_ctrl_1 0.05fF
C625 a_mux4_en_1/switch_5t_0/in a_mux4_en_1/switch_5t_0/en_b -0.00fF
C626 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# -0.00fF
C627 a_mod_grp_ctrl_1 a_mux4_en_1/switch_5t_1/in 0.01fF
C628 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.00fF
C629 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C630 rst_n ota_w_test_0/ip 0.01fF
C631 VSS d_clk_grp_2_ctrl_0 1.60fF
C632 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S -0.00fF
C633 ota_1/p1 clock_v2_0/p1d_b 0.94fF
C634 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/c1_n260_n210# -0.07fF
C635 ota_w_test_0/op ota_w_test_0/m1_n2176_n12171# 0.00fF
C636 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0.04fF
C637 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C638 sky130_fd_sc_hd__clkinv_4_2/Y d_probe_3 0.08fF
C639 transmission_gate_17/in VDD 13.42fF
C640 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# 0.03fF
C641 a_mux4_en_1/switch_5t_3/en_b a_mux4_en_1/switch_5t_2/in -0.00fF
C642 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# 0.05fF
C643 clock_v2_0/p2_b a_mod_grp_ctrl_1 0.05fF
C644 sky130_fd_sc_hd__mux4_1_0/X d_clk_grp_2_ctrl_1 0.02fF
C645 ota_w_test_0/op ota_w_test_0/on 1.51fF
C646 a_mux4_en_1/in2 ota_w_test_0/m1_11534_n9706# 0.05fF
C647 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.00fF
C648 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0.00fF
C649 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# -0.00fF
C650 a_mod_grp_ctrl_1 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C651 sky130_fd_sc_hd__mux4_1_3/a_27_413# ota_1/p1 0.01fF
C652 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# -0.00fF
C653 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C654 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# 0.11fF
C655 sky130_fd_sc_hd__clkinv_4_3/Y clock_v2_0/B_b 0.00fF
C656 VSS ota_w_test_0/sc_cmfb_0/transmission_gate_3/out -0.29fF
C657 ota_1/bias_d ota_1/m1_n2176_n12171# 0.01fF
C658 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# -0.13fF
C659 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.00fF
C660 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0.04fF
C661 d_clk_grp_2_ctrl_1 clock_v2_0/p1d_b 0.11fF
C662 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# ota_1/in 0.04fF
C663 transmission_gate_17/in clock_v2_0/Ad_b 0.74fF
C664 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C665 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.00fF
C666 transmission_gate_19/in transmission_gate_32/out 0.80fF
C667 ota_w_test_0/m1_2462_n3318# a_mux4_en_0/in1 0.01fF
C668 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.15fF
C669 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# ota_1/p1 0.03fF
C670 sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/c1_n260_n210# ota_1/op 0.06fF
C671 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# transmission_gate_6/in 0.30fF
C672 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# VDD 0.14fF
C673 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_2/X 0.03fF
C674 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# VDD 0.14fF
C675 VSS d_probe_0 1.87fF
C676 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# ota_1/p2_b 0.19fF
C677 d_clk_grp_2_ctrl_0 ota_1/p2_b 0.00fF
C678 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.12fF
C679 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.04fF
C680 sky130_fd_sc_hd__mux4_1_3/a_668_97# clock_v2_0/A_b 0.02fF
C681 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0.05fF
C682 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0.00fF
C683 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.11fF
C684 clock_v2_0/Bd_b a_mod_grp_ctrl_1 0.06fF
C685 sky130_fd_sc_hd__mux4_1_1/a_1478_413# d_clk_grp_2_ctrl_0 -0.00fF
C686 VSS sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.01fF
C687 VSS a_mux4_en_0/switch_5t_0/en 0.55fF
C688 VSS ota_1/m1_1038_n2886# 0.19fF
C689 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# -0.00fF
C690 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.02fF
C691 a_mux2_en_0/switch_5t_0/in ota_w_test_0/on 0.02fF
C692 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# ota_1/p1_b 0.01fF
C693 a_mod_grp_ctrl_0 a_mod_grp_ctrl_1 11.47fF
C694 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# VDD 0.20fF
C695 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# ota_1/in 0.17fF
C696 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# clock_v2_0/p1d 0.15fF
C697 VDD a_mux4_en_1/switch_5t_1/en -0.85fF
C698 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C699 d_clk_grp_2_ctrl_0 ota_1/p2 0.10fF
C700 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0.00fF
C701 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# ota_1/ip 0.14fF
C702 clock_v2_0/Ad a_mux4_en_1/in1 0.04fF
C703 clock_v2_0/Ad i_bias_1 0.05fF
C704 a_mod_grp_ctrl_0 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C705 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# -0.38fF
C706 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0.06fF
C707 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C708 transmission_gate_17/in clock_v2_0/p1d_b 0.20fF
C709 a_mux4_en_0/switch_5t_1/en_b a_mux4_en_0/switch_5t_1/en 0.00fF
C710 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413# -0.00fF
C711 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# -0.00fF
C712 sky130_fd_sc_hd__mux4_1_3/a_193_47# VSS -0.00fF
C713 VSS sky130_fd_sc_hd__mux4_1_1/a_1290_413# -0.01fF
C714 clock_v2_0/A clock_v2_0/B_b 3.11fF
C715 ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0.03fF
C716 onebit_dac_1/v_b onebit_dac_1/out 0.05fF
C717 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0.06fF
C718 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C719 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C720 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0.10fF
C721 transmission_gate_19/in clock_v2_0/p2_b 0.08fF
C722 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# -0.00fF
C723 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.00fF
C724 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00fF
C725 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/on 0.00fF
C726 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_2/X 0.02fF
C727 VDD comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X 0.00fF
C728 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/B_b 0.03fF
C729 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# VDD -0.00fF
C730 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/sc_cmfb_0/transmission_gate_7/in -0.09fF
C731 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0.08fF
C732 a_mux2_en_0/switch_5t_1/in a_mux2_en_0/switch_5t_1/transmission_gate_1/in -0.00fF
C733 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/X -0.00fF
C734 ota_1/sc_cmfb_0/transmission_gate_4/out ota_1/p1_b 0.01fF
C735 debug clock_v2_0/B 0.06fF
C736 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# -0.00fF
C737 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# -0.38fF
C738 a_mux4_en_1/switch_5t_0/transmission_gate_1/in a_probe_2 0.00fF
C739 ota_1/p2_b sky130_fd_sc_hd__mux4_1_0/a_27_413# -0.00fF
C740 clock_v2_0/p1d transmission_gate_2/out 0.23fF
C741 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.04fF
C742 transmission_gate_0/out transmission_gate_5/in 0.88fF
C743 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/p2_b 0.02fF
C744 a_mux4_en_0/switch_5t_1/en_b a_mux4_en_0/switch_5t_1/in 0.00fF
C745 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0.00fF
C746 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# -0.00fF
C747 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/X 0.01fF
C748 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# 0.11fF
C749 VSS debug 4.32fF
C750 a_mux4_en_1/transmission_gate_3/en_b a_mux4_en_1/switch_5t_0/en_b -0.00fF
C751 ota_w_test_0/cm ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.01fF
C752 clock_v2_0/Bd clock_v2_0/p1d 0.62fF
C753 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.06fF
C754 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# ota_1/in 0.03fF
C755 ota_1/cmc ota_1/on -0.10fF
C756 a_mux4_en_1/in2 ota_w_test_0/on -0.10fF
C757 ota_1/cmc ota_1/sc_cmfb_0/transmission_gate_8/in -0.00fF
C758 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0.00fF
C759 ota_1/in ota_1/m1_1038_n2886# 0.00fF
C760 ota_1/p2 sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.01fF
C761 transmission_gate_9/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# 0.41fF
C762 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0.09fF
C763 ota_w_test_0/cm ota_w_test_0/m1_6690_n8907# 0.00fF
C764 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.00fF
C765 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C766 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# -0.00fF
C767 clock_v2_0/Bd_b ota_w_test_0/cm 0.10fF
C768 transmission_gate_18/in ota_w_test_0/on 0.06fF
C769 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n930_n880# 0.11fF
C770 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B VDD 0.07fF
C771 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.00fF
C772 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C773 transmission_gate_19/out clock_v2_0/p2 0.97fF
C774 ota_1/bias_b ota_1/bias_c 0.00fF
C775 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.01fF
C776 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0.09fF
C777 op onebit_dac_0/out 0.03fF
C778 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0.10fF
C779 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y -0.00fF
C780 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0.07fF
C781 rst_n clock_v2_0/B_b 0.08fF
C782 VSS ota_1/bias_d 2.73fF
C783 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y 0.00fF
C784 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C785 ota_1/p1_b comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A -0.04fF
C786 d_clk_grp_2_ctrl_0 VDD 1.39fF
C787 sky130_fd_sc_hd__mux4_1_3/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C788 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_1/p1_b 0.06fF
C789 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.05fF
C790 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.03fF
C791 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.08fF
C792 a_mux2_en_0/switch_5t_0/in a_mod_grp_ctrl_1 0.04fF
C793 ota_1/p1_b sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.03fF
C794 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# 0.30fF
C795 ota_1/ip transmission_gate_19/in 1.40fF
C796 sky130_fd_sc_hd__mux4_1_2/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C797 VSS sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.04fF
C798 transmission_gate_18/in transmission_gate_8/in 0.13fF
C799 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# clock_v2_0/p2 0.00fF
C800 VSS transmission_gate_0/out 2.06fF
C801 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_1/p2_b 0.06fF
C802 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0.08fF
C803 ota_1/p1 sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.00fF
C804 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# 0.03fF
C805 sky130_fd_sc_hd__mux4_1_2/a_1478_413# d_clk_grp_1_ctrl_0 -0.00fF
C806 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0.03fF
C807 d_clk_grp_2_ctrl_0 clock_v2_0/Ad_b 0.11fF
C808 ota_1/p2_b debug 0.31fF
C809 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0.00fF
C810 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# -0.00fF
C811 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# -0.24fF
C812 ota_1/p2_b ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.00fF
C813 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0.04fF
C814 ota_1/p1 ota_1/on 0.50fF
C815 ota_w_test_0/sc_cmfb_0/transmission_gate_3/out VDD -0.49fF
C816 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# 0.30fF
C817 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0.26fF
C818 VSS clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S -0.00fF
C819 sky130_fd_sc_hd__mux4_1_3/a_757_363# ota_1/p1_b 0.08fF
C820 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# ota_1/in 0.03fF
C821 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.10fF
C822 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.01fF
C823 ota_w_test_0/op ota_w_test_0/cm 0.00fF
C824 a_probe_2 a_mux4_en_1/switch_5t_3/transmission_gate_1/in 0.00fF
C825 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# -0.09fF
C826 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/A VDD 0.00fF
C827 VSS sky130_fd_sc_hd__clkinv_4_3/Y 0.45fF
C828 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_1/p2 0.03fF
C829 clock_v2_0/Bd a_mux4_en_0/in0 0.04fF
C830 ota_w_test_0/m1_n2176_n12171# ota_w_test_0/on 0.00fF
C831 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# 0.02fF
C832 onebit_dac_1/out clock_v2_0/p2 0.54fF
C833 VSS ota_1/m1_6690_n8907# 0.17fF
C834 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.01fF
C835 ota_1/p2 debug 0.26fF
C836 clock_v2_0/Bd ota_w_test_0/in 0.04fF
C837 clock_v2_0/A transmission_gate_5/in 0.11fF
C838 d_probe_0 VDD 2.48fF
C839 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0.00fF
C840 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210# VDD 0.00fF
C841 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A 1.56fF
C842 ota_1/p2 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.00fF
C843 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# clock_v2_0/p2 0.03fF
C844 sky130_fd_sc_hd__mux4_1_0/X d_clk_grp_2_ctrl_0 0.00fF
C845 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/A VDD -0.00fF
C846 VSS comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# 0.00fF
C847 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# -0.00fF
C848 VSS sky130_fd_sc_hd__clkinv_4_4/Y 0.39fF
C849 sky130_fd_sc_hd__mux4_1_0/a_27_413# VDD 0.07fF
C850 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0.06fF
C851 VDD a_mux4_en_0/switch_5t_0/en -0.71fF
C852 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# -0.00fF
C853 ota_1/m1_1038_n2886# VDD 2.68fF
C854 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C855 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0.07fF
C856 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0.00fF
C857 VSS comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A 0.00fF
C858 a_mux4_en_1/switch_5t_0/en_b a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y -0.00fF
C859 d_clk_grp_2_ctrl_0 clock_v2_0/p1d_b 0.16fF
C860 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# -0.00fF
C861 a_mod_grp_ctrl_0 clk 0.18fF
C862 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C863 clock_v2_0/Ad sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C864 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0.00fF
C865 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.13fF
C866 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.00fF
C867 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# -0.00fF
C868 sky130_fd_sc_hd__mux4_1_2/a_247_21# clock_v2_0/B_b 0.06fF
C869 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210# ota_1/op 0.06fF
C870 ota_w_test_0/m1_2463_n5585# ota_w_test_0/in 0.00fF
C871 clock_v2_0/A clock_v2_0/B 6.65fF
C872 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0.03fF
C873 ota_1/ip ota_1/m1_n208_n2883# 0.00fF
C874 sky130_fd_sc_hd__mux4_1_1/a_1290_413# VDD 0.10fF
C875 sky130_fd_sc_hd__mux4_1_0/a_750_97# ota_1/p2 0.09fF
C876 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# ota_1/p2_b 0.05fF
C877 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980# 0.30fF
C878 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.00fF
C879 clock_v2_0/p2_b clock_v2_0/A_b 1.54fF
C880 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/B 0.00fF
C881 VSS clock_v2_0/A 2.15fF
C882 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# transmission_gate_5/in 0.30fF
C883 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# VDD 0.82fF
C884 rst_n transmission_gate_5/in 0.09fF
C885 ota_w_test_0/cm ota_w_test_0/m1_11534_n9706# -0.01fF
C886 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C887 transmission_gate_26/en clock_v2_0/Bd 0.39fF
C888 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# ota_1/in 0.13fF
C889 VSS sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.04fF
C890 clock_v2_0/Ad ota_1/p1 0.96fF
C891 sky130_fd_sc_hd__mux4_1_1/a_1290_413# clock_v2_0/Ad_b 0.01fF
C892 VSS sky130_fd_sc_hd__mux4_1_3/X 0.60fF
C893 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0.34fF
C894 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0.00fF
C895 a_mux4_en_0/switch_5t_1/en a_probe_3 0.00fF
C896 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# -0.00fF
C897 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# VDD 0.09fF
C898 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B 0.03fF
C899 VDD debug 5.47fF
C900 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# VDD 0.00fF
C901 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# 1.05fF
C902 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# VDD 0.14fF
C903 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.00fF
C904 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0.71fF
C905 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.12fF
C906 VSS comparator_v2_0/li_940_3458# 1.72fF
C907 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.00fF
C908 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C909 VSS transmission_gate_23/in 0.37fF
C910 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0.09fF
C911 transmission_gate_6/in clock_v2_0/A 0.20fF
C912 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0.06fF
C913 clock_v2_0/Bd_b clock_v2_0/A_b 0.14fF
C914 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# 0.10fF
C915 clock_v2_0/Ad d_clk_grp_2_ctrl_1 0.00fF
C916 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0.06fF
C917 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# -0.00fF
C918 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# -0.09fF
C919 rst_n clock_v2_0/B 0.13fF
C920 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# 0.75fF
C921 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0.07fF
C922 clock_v2_0/Ad_b debug 0.07fF
C923 a_mux4_en_0/switch_5t_0/in a_mux4_en_0/switch_5t_0/en -0.00fF
C924 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/B_b 0.04fF
C925 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A VDD 0.09fF
C926 ota_1/bias_d VDD 0.39fF
C927 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.00fF
C928 ota_w_test_0/m1_n6302_n3889# VDD 0.15fF
C929 a_mod_grp_ctrl_0 clock_v2_0/A_b 0.04fF
C930 ota_w_test_0/cm a_mux4_en_1/in2 0.83fF
C931 ota_w_test_0/cm ota_w_test_0/m1_n208_n2883# 0.05fF
C932 ota_1/p1 ota_1/cm 0.17fF
C933 ota_1/p2_b clock_v2_0/A 0.36fF
C934 debug ota_1/op 0.00fF
C935 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# 0.11fF
C936 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0.05fF
C937 transmission_gate_18/in transmission_gate_19/in 0.00fF
C938 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# -0.00fF
C939 VSS rst_n 3.49fF
C940 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.00fF
C941 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# -0.00fF
C942 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# 0.19fF
C943 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.08fF
C944 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.01fF
C945 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0.00fF
C946 sky130_fd_sc_hd__mux4_1_0/a_750_97# VDD 0.10fF
C947 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_0/en 0.00fF
C948 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.01fF
C949 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# -0.09fF
C950 a_mux4_en_1/in1 a_mux4_en_1/switch_5t_1/in 0.00fF
C951 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C952 transmission_gate_0/out VDD 0.88fF
C953 ota_1/p1_b clock_v2_0/B_b 0.11fF
C954 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# -0.00fF
C955 VSS a_mux4_en_0/switch_5t_2/en_b 0.28fF
C956 ota_1/p2 clock_v2_0/A 0.16fF
C957 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.08fF
C958 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0.00fF
C959 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n930_n880# -0.31fF
C960 ota_1/bias_d ota_1/op 0.03fF
C961 transmission_gate_26/en clock_v2_0/p1d 0.11fF
C962 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210# -0.08fF
C963 sky130_fd_sc_hd__clkinv_4_2/Y VSS 0.38fF
C964 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# 0.22fF
C965 clock_v2_0/Ad_b clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# -0.00fF
C966 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S 0.07fF
C967 transmission_gate_9/in transmission_gate_18/in 0.03fF
C968 transmission_gate_23/in ota_1/p2_b 0.01fF
C969 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0.07fF
C970 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0.03fF
C971 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# 0.11fF
C972 sky130_fd_sc_hd__clkinv_4_3/Y VDD -0.54fF
C973 clock_v2_0/Ad transmission_gate_17/in 0.85fF
C974 VSS sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.02fF
C975 sky130_fd_sc_hd__mux4_1_0/a_750_97# clock_v2_0/Ad_b 0.00fF
C976 ota_w_test_0/op clock_v2_0/A_b 0.04fF
C977 transmission_gate_31/out transmission_gate_0/out 0.26fF
C978 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.03fF
C979 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# transmission_gate_5/in 0.22fF
C980 clock_v2_0/p1d_b debug 0.08fF
C981 a_mux4_en_0/switch_5t_1/in a_mux4_en_0/transmission_gate_3/en_b -0.00fF
C982 ota_1/m1_6690_n8907# VDD 1.46fF
C983 rst_n transmission_gate_6/in 0.16fF
C984 a_mux4_en_1/transmission_gate_3/en_b a_mux4_en_1/switch_5t_2/en_b -0.00fF
C985 sky130_fd_sc_hd__mux4_1_3/a_668_97# d_clk_grp_1_ctrl_0 0.03fF
C986 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B 0.00fF
C987 transmission_gate_23/in ota_1/in 0.03fF
C988 transmission_gate_17/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# 0.11fF
C989 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.00fF
C990 transmission_gate_23/in ota_1/p2 0.05fF
C991 VSS a_mux2_en_0/switch_5t_1/in 0.05fF
C992 debug a_mux4_en_0/switch_5t_0/in 0.00fF
C993 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# ota_1/p1_b 0.25fF
C994 a_mux4_en_0/switch_5t_3/en_b a_mux4_en_0/switch_5t_2/en -0.00fF
C995 a_mux4_en_0/switch_5t_2/transmission_gate_1/in a_probe_3 0.00fF
C996 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.01fF
C997 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C998 transmission_gate_31/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# 0.04fF
C999 rst_n ota_1/p2_b 1.21fF
C1000 ota_1/m1_n2176_n12171# ota_1/p1_b 0.16fF
C1001 sky130_fd_sc_hd__clkinv_4_4/Y VDD -0.05fF
C1002 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/A -0.00fF
C1003 ota_w_test_0/m1_2462_n3318# VSS 0.09fF
C1004 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n930_n880# 0.11fF
C1005 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# VDD 0.32fF
C1006 sky130_fd_sc_hd__mux4_1_3/a_834_97# ota_1/p1_b 0.01fF
C1007 VDD comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A 1.19fF
C1008 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C1009 ota_w_test_0/cm ota_w_test_0/on 0.00fF
C1010 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# 0.00fF
C1011 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_1/p1_b 0.06fF
C1012 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# ota_w_test_0/sc_cmfb_0/transmission_gate_9/in 0.06fF
C1013 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_668_97# 0.01fF
C1014 ota_1/m1_6690_n8907# ota_1/op -0.00fF
C1015 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/p2_b 0.04fF
C1016 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.03fF
C1017 rst_n ota_1/in 0.08fF
C1018 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# -0.00fF
C1019 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 7.24fF
C1020 rst_n ota_1/p2 1.17fF
C1021 clock_v2_0/Bd_b a_mux4_en_1/in1 0.04fF
C1022 ota_w_test_0/m1_6690_n8907# a_mux4_en_1/in1 0.36fF
C1023 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C1024 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.02fF
C1025 clock_v2_0/Bd_b i_bias_1 -0.20fF
C1026 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A 0.42fF
C1027 sky130_fd_sc_hd__mux4_1_1/a_834_97# VSS -0.05fF
C1028 sky130_fd_sc_hd__mux4_1_0/a_750_97# clock_v2_0/p1d_b 0.00fF
C1029 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/c1_n260_n210# ota_1/on 0.03fF
C1030 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.08fF
C1031 a_mux4_en_1/switch_5t_3/in a_mux4_en_1/switch_5t_3/en 0.00fF
C1032 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A -0.00fF
C1033 transmission_gate_0/out clock_v2_0/p1d_b 0.42fF
C1034 VSS sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.06fF
C1035 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# 0.11fF
C1036 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.03fF
C1037 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# -0.10fF
C1038 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# 0.22fF
C1039 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# 0.68fF
C1040 ota_1/cmc ota_1/sc_cmfb_0/transmission_gate_3/out -0.02fF
C1041 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# clock_v2_0/p1d_b 0.33fF
C1042 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0.09fF
C1043 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_193_47# -0.00fF
C1044 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y a_mod_grp_ctrl_1 0.00fF
C1045 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/p2 0.03fF
C1046 sky130_fd_sc_hd__mux4_1_1/a_757_363# d_clk_grp_2_ctrl_0 0.00fF
C1047 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# ota_1/on 0.03fF
C1048 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.01fF
C1049 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.00fF
C1050 VDD clock_v2_0/A 7.89fF
C1051 ota_1/bias_b ota_1/m1_n208_n2883# 0.02fF
C1052 ota_w_test_0/cm transmission_gate_8/in 0.17fF
C1053 transmission_gate_26/en ota_w_test_0/in 0.00fF
C1054 clock_v2_0/Ad_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_5/a_110_47# -0.00fF
C1055 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/cm 0.08fF
C1056 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.01fF
C1057 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.00fF
C1058 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_2/a_110_47# -0.00fF
C1059 sky130_fd_sc_hd__mux4_1_2/a_750_97# VDD 0.10fF
C1060 sky130_fd_sc_hd__mux4_1_1/a_750_97# ota_1/p2 0.00fF
C1061 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# VSS 2.06fF
C1062 sky130_fd_sc_hd__mux4_1_3/X VDD 0.71fF
C1063 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/X -0.12fF
C1064 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.15fF
C1065 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# -0.00fF
C1066 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B 0.07fF
C1067 clock_v2_0/Ad_b clock_v2_0/A 0.41fF
C1068 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# 0.00fF
C1069 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0.09fF
C1070 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0.32fF
C1071 ota_1/p1_b transmission_gate_5/in 0.16fF
C1072 a_mux4_en_0/in1 ota_w_test_0/m1_n947_n12836# 0.92fF
C1073 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# VDD 0.15fF
C1074 VSS ota_1/m1_2463_n5585# 0.05fF
C1075 transmission_gate_23/in VDD 0.37fF
C1076 ota_w_test_0/op a_mux4_en_1/in1 0.20fF
C1077 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0.04fF
C1078 ota_1/m1_n208_n2883# ota_1/bias_c -0.00fF
C1079 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_0/en_b 0.00fF
C1080 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/B -0.00fF
C1081 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# -0.14fF
C1082 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# 0.09fF
C1083 ota_1/p1 ota_1/sc_cmfb_0/transmission_gate_3/out 0.00fF
C1084 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# transmission_gate_23/in 0.00fF
C1085 onebit_dac_0/out transmission_gate_32/out 0.17fF
C1086 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.00fF
C1087 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0.09fF
C1088 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0.15fF
C1089 ota_w_test_0/cm ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# -0.02fF
C1090 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# -0.00fF
C1091 a_mux4_en_1/in2 clock_v2_0/A_b 0.03fF
C1092 VSS sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.09fF
C1093 VSS ip 1.07fF
C1094 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0.00fF
C1095 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# -0.00fF
C1096 VSS a_mux4_en_1/switch_5t_3/en_b 0.17fF
C1097 rst_n VDD 14.10fF
C1098 sky130_fd_sc_hd__mux4_1_1/a_834_97# ota_1/p2 0.00fF
C1099 ota_1/op comparator_v2_0/li_940_3458# 0.00fF
C1100 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# VDD 0.03fF
C1101 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# -0.08fF
C1102 ota_1/p1_b clock_v2_0/B 0.47fF
C1103 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 0.30fF
C1104 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# 2.72fF
C1105 clock_v2_0/p1d_b clock_v2_0/A 0.08fF
C1106 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# -0.00fF
C1107 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# VDD 0.08fF
C1108 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# 0.25fF
C1109 VDD a_mux4_en_0/switch_5t_2/en_b 0.13fF
C1110 a_mux4_en_1/switch_5t_0/en a_mux4_en_1/switch_5t_0/transmission_gate_1/in 0.00fF
C1111 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0.04fF
C1112 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# 0.13fF
C1113 clock_v2_0/Ad d_clk_grp_2_ctrl_0 0.01fF
C1114 VSS ota_1/p1_b 10.48fF
C1115 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# ota_1/p1 0.10fF
C1116 transmission_gate_31/out rst_n 0.05fF
C1117 a_probe_3 a_mux4_en_0/switch_5t_2/en 0.00fF
C1118 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_1/p1_b 0.04fF
C1119 sky130_fd_sc_hd__clkinv_4_2/Y VDD -0.21fF
C1120 rst_n clock_v2_0/Ad_b 0.12fF
C1121 a_mux4_en_0/in2 ota_w_test_0/m1_n947_n12836# 0.04fF
C1122 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# -0.00fF
C1123 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C1124 rst_n ota_1/op 0.16fF
C1125 sky130_fd_sc_hd__mux4_1_1/a_750_97# VDD 0.19fF
C1126 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# clock_v2_0/p2 0.03fF
C1127 sky130_fd_sc_hd__mux4_1_3/a_27_413# clock_v2_0/A 0.02fF
C1128 clock_v2_0/p2 clock_v2_0/B_b 4.81fF
C1129 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0.00fF
C1130 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0.06fF
C1131 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# ota_1/p1_b 0.09fF
C1132 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# 2.08fF
C1133 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.00fF
C1134 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C1135 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980# 0.29fF
C1136 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0.01fF
C1137 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B 0.09fF
C1138 onebit_dac_0/out clock_v2_0/p2_b 0.64fF
C1139 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0.05fF
C1140 sky130_fd_sc_hd__clkinv_4_2/Y clock_v2_0/Ad_b 0.00fF
C1141 a_mux2_en_0/switch_5t_1/in VDD 0.59fF
C1142 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/op -0.00fF
C1143 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A -0.00fF
C1144 a_mux4_en_1/switch_5t_3/en_b a_mux4_en_1/switch_5t_2/en -0.00fF
C1145 a_mux4_en_1/switch_5t_0/en_b a_mux4_en_1/sky130_fd_sc_hd__nand2_1_3/a_113_47# -0.00fF
C1146 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/X -0.00fF
C1147 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/Ad_b 0.03fF
C1148 debug ota_1/on 0.00fF
C1149 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0.01fF
C1150 ota_w_test_0/m1_2462_n3318# VDD 0.85fF
C1151 ota_w_test_0/on clock_v2_0/A_b 0.04fF
C1152 a_mux4_en_0/switch_5t_2/en a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C1153 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# clock_v2_0/p1d 0.15fF
C1154 ota_1/p1 clock_v2_0/p2_b 2.05fF
C1155 rst_n clock_v2_0/p1d_b 0.20fF
C1156 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0.00fF
C1157 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# transmission_gate_0/out 0.30fF
C1158 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# -0.00fF
C1159 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.04fF
C1160 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0.09fF
C1161 ota_1/p2_b ota_1/p1_b 3.35fF
C1162 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A -0.00fF
C1163 sky130_fd_sc_hd__mux4_1_1/a_247_21# d_clk_grp_2_ctrl_0 0.19fF
C1164 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_0/X 0.02fF
C1165 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.12fF
C1166 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A 0.33fF
C1167 VSS ota_1/m1_2462_n3318# 0.02fF
C1168 sky130_fd_sc_hd__mux4_1_1/a_834_97# VDD 0.01fF
C1169 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.02fF
C1170 clock_v2_0/Ad sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C1171 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0.16fF
C1172 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C1173 ota_w_test_0/m1_12118_n9704# a_mux4_en_1/in2 0.04fF
C1174 clock_v2_0/sky130_fd_sc_hd__nand2_1_0/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# -0.00fF
C1175 ota_1/bias_d ota_1/on 0.04fF
C1176 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0.05fF
C1177 sky130_fd_sc_hd__mux4_1_2/a_247_21# VDD 0.03fF
C1178 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_193_413# -0.00fF
C1179 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.13fF
C1180 a_mux4_en_1/transmission_gate_3/en_b a_mux4_en_1/switch_5t_2/in -0.00fF
C1181 VSS a_mux4_en_1/switch_5t_1/en_b 0.27fF
C1182 d_clk_grp_1_ctrl_0 clock_v2_0/p2_b 0.11fF
C1183 a_mux4_en_1/in2 a_mux4_en_1/in1 2.01fF
C1184 ota_w_test_0/m1_n208_n2883# a_mux4_en_1/in1 0.08fF
C1185 VSS onebit_dac_1/v_b 4.03fF
C1186 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_3/in 0.01fF
C1187 i_bias_1 ota_w_test_0/m1_n208_n2883# -0.02fF
C1188 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0.09fF
C1189 ota_1/in ota_1/p1_b 0.14fF
C1190 sky130_fd_sc_hd__clkinv_4_2/Y clock_v2_0/p1d_b 0.00fF
C1191 ota_1/p2 ota_1/p1_b 8.18fF
C1192 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# 0.12fF
C1193 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.01fF
C1194 a_mux4_en_0/switch_5t_2/in debug -0.00fF
C1195 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__clkinv_4_3/Y 0.03fF
C1196 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/c1_n260_n210# 0.03fF
C1197 VSS a_mux2_en_0/switch_5t_0/transmission_gate_1/in 0.09fF
C1198 VSS in 3.26fF
C1199 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/Ad_b 0.01fF
C1200 sky130_fd_sc_hd__mux4_1_1/a_750_97# clock_v2_0/p1d_b 0.11fF
C1201 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# -0.00fF
C1202 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0.14fF
C1203 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1204 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# -0.00fF
C1205 sky130_fd_sc_hd__mux4_1_1/a_277_47# d_clk_grp_2_ctrl_1 0.08fF
C1206 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out a_mux4_en_1/in1 0.02fF
C1207 clock_v2_0/Bd_b ota_1/p1 0.49fF
C1208 transmission_gate_9/in ota_w_test_0/cm 0.14fF
C1209 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0.06fF
C1210 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# -0.00fF
C1211 VSS comparator_v2_0/li_940_818# 1.49fF
C1212 ota_1/p1 ota_w_test_0/m1_6690_n8907# 0.07fF
C1213 sky130_fd_sc_hd__mux4_1_2/a_757_363# clock_v2_0/p2_b 0.06fF
C1214 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# clock_v2_0/p1d_b 0.02fF
C1215 VSS sky130_fd_sc_hd__mux4_1_1/a_668_97# -0.24fF
C1216 ota_1/p1 a_mod_grp_ctrl_0 0.05fF
C1217 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0.06fF
C1218 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.01fF
C1219 ota_1/m1_n6302_n3889# VDD 1.25fF
C1220 ota_1/m1_1038_n2886# ota_1/cm 0.08fF
C1221 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0.00fF
C1222 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0.05fF
C1223 ota_1/m1_2463_n5585# VDD 1.38fF
C1224 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# -0.00fF
C1225 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# -0.12fF
C1226 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y 0.36fF
C1227 ota_1/m1_6690_n8907# ota_1/on -0.01fF
C1228 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_27_47# -0.00fF
C1229 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0.01fF
C1230 ota_1/ip ota_1/p1 0.08fF
C1231 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# 0.06fF
C1232 VSS ota_w_test_0/sc_cmfb_0/transmission_gate_7/in 0.37fF
C1233 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.08fF
C1234 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# ota_1/p1_b 0.03fF
C1235 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C1236 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.02fF
C1237 clock_v2_0/Bd_b d_clk_grp_2_ctrl_1 0.00fF
C1238 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A VDD 0.00fF
C1239 clock_v2_0/Ad debug 0.07fF
C1240 transmission_gate_19/out clock_v2_0/p1d 0.45fF
C1241 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# 0.02fF
C1242 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980# 0.69fF
C1243 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A 0.00fF
C1244 sky130_fd_sc_hd__mux4_1_2/a_27_47# VDD 0.01fF
C1245 sky130_fd_sc_hd__mux4_1_1/a_834_97# clock_v2_0/p1d_b 0.01fF
C1246 ip VDD 2.39fF
C1247 VDD a_mux4_en_1/switch_5t_3/en_b -0.21fF
C1248 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# ota_1/on 0.00fF
C1249 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# -0.00fF
C1250 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# 0.11fF
C1251 a_mux4_en_1/in2 ota_w_test_0/m1_11825_n9711# 0.04fF
C1252 sky130_fd_sc_hd__mux4_1_2/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C1253 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C1254 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# 0.08fF
C1255 clock_v2_0/A_b a_mod_grp_ctrl_1 0.06fF
C1256 a_mux4_en_1/switch_5t_1/transmission_gate_1/in a_mux4_en_1/switch_5t_1/en_b 0.00fF
C1257 ota_w_test_0/on a_mux4_en_1/in1 0.05fF
C1258 ota_w_test_0/op ota_1/p1 0.27fF
C1259 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# -0.00fF
C1260 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y 0.09fF
C1261 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C1262 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# VDD 0.00fF
C1263 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C1264 transmission_gate_31/out ip 0.02fF
C1265 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.00fF
C1266 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# ota_1/p1 0.23fF
C1267 ota_1/p1_b VDD 21.01fF
C1268 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C1269 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.07fF
C1270 a_mux4_en_1/switch_5t_0/en a_mod_grp_ctrl_1 0.16fF
C1271 clock_v2_0/p2 clock_v2_0/B 4.21fF
C1272 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.02fF
C1273 a_mux4_en_1/switch_5t_1/en a_mux4_en_1/switch_5t_1/in -0.00fF
C1274 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980# 0.22fF
C1275 ota_1/cm ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.08fF
C1276 ota_1/p1 ota_1/bias_a 4.13fF
C1277 d_probe_3 sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C1278 clock_v2_0/Bd_b transmission_gate_17/in 0.36fF
C1279 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.01fF
C1280 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0.12fF
C1281 sky130_fd_sc_hd__mux4_1_3/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C1282 ota_1/m1_n947_n12836# VSS 0.56fF
C1283 VSS a_mux4_en_0/switch_5t_1/en 0.54fF
C1284 VSS clock_v2_0/p2 3.49fF
C1285 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.00fF
C1286 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.03fF
C1287 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# -0.13fF
C1288 clock_v2_0/Ad_b ota_1/p1_b 0.60fF
C1289 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/c1_n530_n480# -0.16fF
C1290 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.03fF
C1291 sky130_fd_sc_hd__mux4_1_3/a_193_413# d_clk_grp_1_ctrl_0 0.00fF
C1292 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# ota_1/p1_b 0.00fF
C1293 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0.02fF
C1294 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y 0.00fF
C1295 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.00fF
C1296 ota_1/p1_b ota_1/op 0.34fF
C1297 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# clock_v2_0/p1d 0.27fF
C1298 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.92fF
C1299 a_mod_grp_ctrl_1 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_1/a_113_47# 0.00fF
C1300 VSS sky130_fd_sc_hd__mux4_1_1/a_27_413# 0.00fF
C1301 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# -0.00fF
C1302 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_1/a_193_47# 0.01fF
C1303 comparator_v2_0/li_940_3458# ota_1/on 0.00fF
C1304 transmission_gate_23/in ota_1/on 0.46fF
C1305 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980# ota_1/p1_b 0.01fF
C1306 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# -0.00fF
C1307 ota_w_test_0/m1_2463_n5585# ota_w_test_0/m1_1038_n2886# 0.01fF
C1308 ip clock_v2_0/p1d_b 0.00fF
C1309 VSS a_mux4_en_0/switch_5t_1/in 0.03fF
C1310 ota_1/m1_2462_n3318# VDD 0.74fF
C1311 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0.05fF
C1312 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.06fF
C1313 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# -0.00fF
C1314 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# -0.00fF
C1315 ota_w_test_0/op transmission_gate_17/in 0.14fF
C1316 ota_w_test_0/cm clock_v2_0/A_b 0.12fF
C1317 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C1318 VDD a_mux4_en_1/switch_5t_1/en_b 0.16fF
C1319 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0.04fF
C1320 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.01fF
C1321 sky130_fd_sc_hd__clkinv_4_1/Y d_probe_3 1.63fF
C1322 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0.05fF
C1323 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C1324 onebit_dac_1/v_b VDD 2.92fF
C1325 rst_n ota_1/on 0.22fF
C1326 clock_v2_0/p1d_b ota_1/p1_b 3.75fF
C1327 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y 0.32fF
C1328 ota_1/p2_b clock_v2_0/p2 1.02fF
C1329 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.01fF
C1330 a_mux2_en_0/switch_5t_0/transmission_gate_1/in VDD 0.27fF
C1331 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.00fF
C1332 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# ota_1/p1_b 0.02fF
C1333 VDD in 2.42fF
C1334 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S -0.00fF
C1335 ota_1/m1_6690_n8907# ota_1/cm -0.00fF
C1336 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0.11fF
C1337 ota_1/p2_b ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.01fF
C1338 a_mux4_en_0/in1 clock_v2_0/Bd 0.04fF
C1339 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A 0.00fF
C1340 ota_1/m1_2462_n3318# ota_1/op -0.00fF
C1341 sky130_fd_sc_hd__mux4_1_1/a_27_413# ota_1/p2_b 0.00fF
C1342 sky130_fd_sc_hd__mux4_1_3/a_27_413# ota_1/p1_b 0.03fF
C1343 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# ota_1/in 0.17fF
C1344 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C1345 ota_1/p2 clock_v2_0/p2 0.68fF
C1346 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y 0.26fF
C1347 d_probe_1 d_clk_grp_2_ctrl_1 0.38fF
C1348 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# VDD -0.00fF
C1349 sky130_fd_sc_hd__mux4_1_1/a_668_97# VDD 0.01fF
C1350 a_mux4_en_0/switch_5t_3/in a_mux4_en_0/switch_5t_3/transmission_gate_1/in 0.00fF
C1351 clock_v2_0/Ad clock_v2_0/A 0.54fF
C1352 clock_v2_0/Bd ota_w_test_0/ip 0.02fF
C1353 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.00fF
C1354 a_mux2_en_0/transmission_gate_1/en_b debug 0.02fF
C1355 clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y -0.00fF
C1356 a_mux4_en_1/in2 ota_1/p1 0.02fF
C1357 sky130_fd_sc_hd__mux4_1_3/a_27_47# clock_v2_0/B 0.00fF
C1358 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y -0.00fF
C1359 ota_1/p2 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.05fF
C1360 transmission_gate_18/in ota_1/p1 0.16fF
C1361 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0.00fF
C1362 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# ota_1/p1_b 0.02fF
C1363 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_277_47# -0.01fF
C1364 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.02fF
C1365 d_clk_grp_2_ctrl_0 clock_v2_0/p2_b 0.02fF
C1366 VSS a_mux4_en_0/switch_5t_2/transmission_gate_1/in 0.44fF
C1367 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C1368 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in VDD 0.31fF
C1369 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0.05fF
C1370 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.16fF
C1371 VSS sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.10fF
C1372 comparator_v2_0/li_940_818# ota_1/op 0.00fF
C1373 sky130_fd_sc_hd__mux4_1_1/a_668_97# clock_v2_0/Ad_b 0.00fF
C1374 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/c1_n930_n880# -0.78fF
C1375 ota_w_test_0/m1_2463_n5585# a_mux4_en_0/in1 0.01fF
C1376 sky130_fd_sc_hd__mux4_1_1/a_277_47# d_clk_grp_2_ctrl_0 0.08fF
C1377 VSS ota_w_test_0/m1_n947_n12836# 0.40fF
C1378 ota_1/bias_b ota_1/p1 0.16fF
C1379 a_mux4_en_0/switch_5t_0/en_b a_mod_grp_ctrl_1 0.01fF
C1380 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# 0.21fF
C1381 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A 0.35fF
C1382 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.00fF
C1383 a_mux4_en_0/switch_5t_2/in a_mux4_en_0/switch_5t_2/en_b -0.00fF
C1384 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C1385 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# 0.30fF
C1386 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.13fF
C1387 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y a_mux4_en_0/switch_5t_0/en_b -0.00fF
C1388 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C1389 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y -0.00fF
C1390 clock_v2_0/Bd a_mux4_en_0/in2 0.04fF
C1391 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# transmission_gate_2/out 1.54fF
C1392 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.06fF
C1393 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_w_test_0/sc_cmfb_0/transmission_gate_8/in 0.01fF
C1394 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0.00fF
C1395 sky130_fd_sc_hd__mux4_1_3/a_750_97# clock_v2_0/B_b 0.00fF
C1396 ota_w_test_0/m1_12118_n9704# ota_w_test_0/cm -0.01fF
C1397 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# -0.00fF
C1398 i_bias_2 ota_1/m1_n5574_n13620# -0.02fF
C1399 clock_v2_0/p1d_b in 0.04fF
C1400 clock_v2_0/Bd_b d_clk_grp_2_ctrl_0 0.02fF
C1401 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in ota_w_test_0/sc_cmfb_0/transmission_gate_3/out -0.00fF
C1402 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0.00fF
C1403 clock_v2_0/Ad rst_n 0.11fF
C1404 ota_w_test_0/cm a_mux4_en_1/in1 2.25fF
C1405 transmission_gate_17/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n930_n880# 0.11fF
C1406 ota_1/p1 ota_1/bias_c 0.23fF
C1407 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# -0.15fF
C1408 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0.10fF
C1409 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# -0.13fF
C1410 sky130_fd_sc_hd__mux4_1_3/a_923_363# ota_1/p1_b -0.50fF
C1411 transmission_gate_23/in ota_1/cm 0.02fF
C1412 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C1413 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480# 0.09fF
C1414 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C1415 ota_1/m1_n947_n12836# VDD 0.29fF
C1416 a_mux4_en_0/switch_5t_1/en VDD -0.59fF
C1417 VDD clock_v2_0/p2 4.28fF
C1418 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0.10fF
C1419 ota_1/p1 ota_w_test_0/on 1.53fF
C1420 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C1421 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0.00fF
C1422 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C1423 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0.00fF
C1424 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# -0.00fF
C1425 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00fF
C1426 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0.08fF
C1427 transmission_gate_18/in transmission_gate_17/in -0.66fF
C1428 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# VDD 0.00fF
C1429 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y 0.00fF
C1430 sky130_fd_sc_hd__mux4_1_1/a_27_413# VDD 0.11fF
C1431 clock_v2_0/Ad sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.00fF
C1432 VSS ota_1/m1_12410_n9718# 0.00fF
C1433 transmission_gate_31/out clock_v2_0/p2 0.20fF
C1434 clock_v2_0/Ad_b clock_v2_0/p2 0.05fF
C1435 rst_n ota_1/cm 0.55fF
C1436 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# -0.00fF
C1437 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# 0.11fF
C1438 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0.23fF
C1439 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X -0.01fF
C1440 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# 0.11fF
C1441 sky130_fd_sc_hd__mux4_1_2/a_277_47# ota_1/p1_b 0.00fF
C1442 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# -0.00fF
C1443 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# ota_1/in 0.26fF
C1444 ota_1/m1_n947_n12836# ota_1/op 0.00fF
C1445 ota_1/p1 transmission_gate_8/in 0.12fF
C1446 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y VSS 0.66fF
C1447 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.13fF
C1448 VDD a_mux4_en_0/switch_5t_1/in 0.38fF
C1449 sky130_fd_sc_hd__mux4_1_2/X clock_v2_0/B_b 0.00fF
C1450 sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# -0.09fF
C1451 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/A -0.00fF
C1452 a_mux4_en_0/in0 a_mux4_en_0/transmission_gate_3/en_b 0.02fF
C1453 debug a_mux4_en_1/switch_5t_1/in 0.00fF
C1454 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0.00fF
C1455 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_1290_413# 0.03fF
C1456 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# transmission_gate_2/out 0.03fF
C1457 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.41fF
C1458 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.00fF
C1459 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# -0.00fF
C1460 ota_w_test_0/cm ota_w_test_0/m1_11825_n9711# -0.01fF
C1461 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n930_n880# 0.01fF
C1462 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# -0.00fF
C1463 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.00fF
C1464 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# VDD 0.05fF
C1465 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# -0.09fF
C1466 VSS a_mux4_en_1/switch_5t_0/in 0.03fF
C1467 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.00fF
C1468 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y VDD 1.52fF
C1469 transmission_gate_19/out transmission_gate_21/in 0.09fF
C1470 transmission_gate_0/out transmission_gate_32/out 0.53fF
C1471 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# -0.42fF
C1472 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# a_mux4_en_0/in0 -0.02fF
C1473 a_mux4_en_0/in1 a_mux4_en_0/in0 3.82fF
C1474 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0.05fF
C1475 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# clock_v2_0/p1d 0.15fF
C1476 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/X -0.00fF
C1477 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/c1_n930_n880# transmission_gate_17/in -0.10fF
C1478 sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.01fF
C1479 a_mux4_en_0/in1 ota_w_test_0/in 0.00fF
C1480 debug clock_v2_0/p2_b 0.06fF
C1481 VSS a_mux4_en_0/switch_5t_2/en 0.48fF
C1482 a_mux4_en_1/switch_5t_3/in a_mod_grp_ctrl_1 0.01fF
C1483 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# 0.03fF
C1484 clock_v2_0/p1d_b clock_v2_0/p2 1.95fF
C1485 ota_1/p1_b ota_1/on 0.50fF
C1486 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.02fF
C1487 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# 0.03fF
C1488 ota_w_test_0/ip ota_w_test_0/in 0.37fF
C1489 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y VDD 0.16fF
C1490 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0.00fF
C1491 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y -0.00fF
C1492 transmission_gate_17/in ota_w_test_0/on 0.04fF
C1493 clock_v2_0/Bd clock_v2_0/B_b 6.94fF
C1494 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0.00fF
C1495 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# -0.00fF
C1496 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/p1d_b 0.03fF
C1497 VDD a_mux4_en_0/switch_5t_2/transmission_gate_1/in -0.22fF
C1498 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.00fF
C1499 sky130_fd_sc_hd__mux4_1_3/a_27_413# clock_v2_0/p2 0.00fF
C1500 ota_1/p1 a_mod_grp_ctrl_1 0.06fF
C1501 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0.05fF
C1502 sky130_fd_sc_hd__mux4_1_3/a_1478_413# clock_v2_0/A_b -0.00fF
C1503 ota_w_test_0/m1_n5574_n13620# a_mux4_en_0/in0 -0.00fF
C1504 sky130_fd_sc_hd__mux4_1_3/a_27_47# VDD 0.02fF
C1505 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0.13fF
C1506 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# -0.00fF
C1507 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.01fF
C1508 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.13fF
C1509 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/c1_n260_n210# 0.03fF
C1510 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# clock_v2_0/p1d_b 0.08fF
C1511 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# 0.32fF
C1512 clock_v2_0/Bd_b debug 0.07fF
C1513 ota_w_test_0/m1_n947_n12836# VDD -0.15fF
C1514 VSS a_mux2_en_1/transmission_gate_1/en_b -0.11fF
C1515 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A 0.14fF
C1516 sky130_fd_sc_hd__mux4_1_2/a_834_97# ota_1/p1_b 0.00fF
C1517 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0.09fF
C1518 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# 0.09fF
C1519 transmission_gate_8/in transmission_gate_17/in 0.03fF
C1520 transmission_gate_0/out clock_v2_0/p2_b 0.17fF
C1521 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/c1_n260_n210# 0.03fF
C1522 d_clk_grp_2_ctrl_0 d_probe_1 0.84fF
C1523 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# VDD 0.00fF
C1524 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.00fF
C1525 ota_w_test_0/cm ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# -0.01fF
C1526 a_mux4_en_0/in0 a_mux4_en_0/in2 -0.10fF
C1527 a_mod_grp_ctrl_0 debug 17.55fF
C1528 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0.07fF
C1529 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.03fF
C1530 sky130_fd_sc_hd__mux4_1_2/a_1290_413# clock_v2_0/B_b 0.01fF
C1531 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# -0.00fF
C1532 transmission_gate_19/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.03fF
C1533 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# 0.01fF
C1534 ota_1/m1_2462_n3318# ota_1/on -0.00fF
C1535 sky130_fd_sc_hd__clkinv_4_3/Y clock_v2_0/p2_b 0.00fF
C1536 transmission_gate_19/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0.04fF
C1537 op onebit_dac_1/v_b 1.88fF
C1538 transmission_gate_26/en ota_w_test_0/ip 0.01fF
C1539 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# 0.11fF
C1540 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C1541 a_mux4_en_0/switch_5t_3/en_b a_mux4_en_0/sky130_fd_sc_hd__nand2_1_0/a_113_47# -0.00fF
C1542 VSS sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.02fF
C1543 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0.00fF
C1544 a_mux4_en_1/in1 clock_v2_0/A_b 0.03fF
C1545 VSS a_mux2_en_1/switch_5t_1/transmission_gate_1/in 0.04fF
C1546 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0.00fF
C1547 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_1290_413# -0.00fF
C1548 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0.00fF
C1549 i_bias_1 clock_v2_0/A_b 0.08fF
C1550 a_mux4_en_1/switch_5t_2/en_b a_mux4_en_1/switch_5t_2/in -0.00fF
C1551 ota_1/cm ota_1/m1_2463_n5585# 0.01fF
C1552 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.03fF
C1553 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# 0.13fF
C1554 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.32fF
C1555 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C1556 clock_v2_0/p1d clock_v2_0/B_b 0.05fF
C1557 ota_w_test_0/op debug 0.00fF
C1558 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# 0.13fF
C1559 clock_v2_0/Ad ota_1/p1_b 0.07fF
C1560 d_probe_0 d_probe_1 0.89fF
C1561 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C1562 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.09fF
C1563 comparator_v2_0/li_940_818# ota_1/on 0.00fF
C1564 clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y VDD 0.03fF
C1565 VSS sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.20fF
C1566 transmission_gate_23/in transmission_gate_32/out 0.06fF
C1567 ota_w_test_0/cm ota_1/p1 0.22fF
C1568 a_mux2_en_1/switch_5t_1/in a_mux2_en_1/switch_5t_0/in 0.00fF
C1569 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0.00fF
C1570 VSS comparator_v2_0/li_n2324_818# 7.21fF
C1571 transmission_gate_2/out transmission_gate_5/in 3.06fF
C1572 a_probe_3 a_mux4_en_0/switch_5t_0/transmission_gate_1/in 0.00fF
C1573 d_clk_grp_1_ctrl_1 clock_v2_0/B_b 0.00fF
C1574 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.00fF
C1575 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.11fF
C1576 a_mux4_en_1/in2 ota_w_test_0/sc_cmfb_0/transmission_gate_3/out -0.00fF
C1577 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.00fF
C1578 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# 0.11fF
C1579 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0.25fF
C1580 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00fF
C1581 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C1582 d_probe_2 sky130_fd_sc_hd__mux4_1_1/X 0.02fF
C1583 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y VDD -0.35fF
C1584 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# 0.65fF
C1585 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.01fF
C1586 ota_1/sc_cmfb_0/transmission_gate_6/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# 0.12fF
C1587 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# VDD 0.15fF
C1588 VSS a_mux4_en_1/transmission_gate_3/en_b 0.29fF
C1589 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.05fF
C1590 clock_v2_0/A clock_v2_0/p2_b 0.92fF
C1591 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0.08fF
C1592 rst_n transmission_gate_32/out 0.05fF
C1593 ota_1/p1 sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.00fF
C1594 VSS sky130_fd_sc_hd__mux4_1_2/X 0.70fF
C1595 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# ota_1/p1_b 0.01fF
C1596 ota_1/cm ota_1/p1_b 0.12fF
C1597 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.02fF
C1598 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_4/a_113_47# 0.00fF
C1599 transmission_gate_9/in ota_1/p1 0.09fF
C1600 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/p2 0.01fF
C1601 a_mux2_en_0/switch_5t_0/in debug 0.02fF
C1602 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/p2_b 0.10fF
C1603 a_mux4_en_1/switch_5t_0/in VDD 0.42fF
C1604 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0.10fF
C1605 ota_1/bias_a ota_1/bias_d 0.01fF
C1606 ota_1/sc_cmfb_0/transmission_gate_9/in ota_1/sc_cmfb_0/transmission_gate_4/out -0.11fF
C1607 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0.05fF
C1608 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.05fF
C1609 sky130_fd_sc_hd__mux4_1_1/a_27_47# d_clk_grp_2_ctrl_0 0.01fF
C1610 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0.00fF
C1611 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# 0.05fF
C1612 VDD a_mux4_en_0/switch_5t_2/en -0.18fF
C1613 sky130_fd_sc_hd__mux4_1_1/X d_clk_grp_2_ctrl_1 0.02fF
C1614 VSS sky130_fd_sc_hd__mux4_1_2/a_923_363# -0.11fF
C1615 ota_1/p2_b sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C1616 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.13fF
C1617 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A -0.00fF
C1618 sky130_fd_sc_hd__mux4_1_2/a_1478_413# clock_v2_0/p2 0.00fF
C1619 sky130_fd_sc_hd__clkinv_4_1/Y VSS 0.43fF
C1620 a_mux4_en_0/in0 clock_v2_0/B_b 0.04fF
C1621 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# -0.00fF
C1622 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.02fF
C1623 clock_v2_0/Bd clock_v2_0/B 3.18fF
C1624 VSS transmission_gate_2/out 2.17fF
C1625 clock_v2_0/B_b ota_w_test_0/in 0.17fF
C1626 a_mux4_en_1/switch_5t_1/en a_mod_grp_ctrl_1 0.03fF
C1627 a_mux2_en_1/switch_5t_1/en a_mux2_en_1/switch_5t_0/in 0.00fF
C1628 ota_1/bias_b ota_1/m1_1038_n2886# 0.01fF
C1629 clock_v2_0/Bd_b clock_v2_0/A 0.32fF
C1630 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.03fF
C1631 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_3/a_113_47# a_mux4_en_0/switch_5t_0/en_b -0.00fF
C1632 VSS sky130_fd_sc_hd__mux4_1_0/a_834_97# -0.06fF
C1633 a_mux4_en_1/transmission_gate_3/en_b a_mux4_en_1/switch_5t_2/en 0.00fF
C1634 ota_1/p2 sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C1635 VSS clock_v2_0/Bd 5.36fF
C1636 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0.09fF
C1637 a_mod_grp_ctrl_0 clock_v2_0/A 0.05fF
C1638 ota_1/m1_n947_n12836# ota_1/on 0.03fF
C1639 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C1640 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# -0.00fF
C1641 VSS comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# 0.00fF
C1642 sky130_fd_sc_hd__mux4_1_3/a_277_47# clock_v2_0/B_b 0.00fF
C1643 sky130_fd_sc_hd__mux4_1_0/a_277_47# d_clk_grp_2_ctrl_1 0.04fF
C1644 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.02fF
C1645 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# -0.00fF
C1646 rst_n clock_v2_0/p2_b 0.05fF
C1647 ota_1/p1 ota_1/m1_n208_n2883# 0.09fF
C1648 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# ota_1/on 0.03fF
C1649 a_mux2_en_1/transmission_gate_1/en_b VDD 0.26fF
C1650 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# -0.00fF
C1651 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0.02fF
C1652 VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# 0.40fF
C1653 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# -0.00fF
C1654 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0.03fF
C1655 transmission_gate_6/in transmission_gate_2/out 0.93fF
C1656 a_mux2_en_0/switch_5t_0/transmission_gate_1/in a_probe_0 0.00fF
C1657 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X -0.01fF
C1658 ota_1/bias_c ota_1/m1_1038_n2886# -0.00fF
C1659 a_mux4_en_1/in2 debug 0.02fF
C1660 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# -0.06fF
C1661 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.01fF
C1662 ota_w_test_0/m1_2463_n5585# VSS 0.44fF
C1663 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C1664 VSS sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0.01fF
C1665 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# 0.11fF
C1666 VSS a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.15fF
C1667 ota_w_test_0/op clock_v2_0/A 0.05fF
C1668 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.02fF
C1669 transmission_gate_26/en clock_v2_0/B_b 0.06fF
C1670 sky130_fd_sc_hd__mux4_1_3/a_750_97# VDD 0.19fF
C1671 ota_1/ip transmission_gate_23/in 0.21fF
C1672 a_mux4_en_1/switch_5t_3/en_b a_mux4_en_1/switch_5t_3/en -0.00fF
C1673 a_mux2_en_1/transmission_gate_1/en_b ota_1/op 0.00fF
C1674 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0.34fF
C1675 a_mux2_en_1/switch_5t_1/transmission_gate_1/in VDD 0.17fF
C1676 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# 0.31fF
C1677 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.04fF
C1678 clock_v2_0/Bd_b rst_n 0.18fF
C1679 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# -0.00fF
C1680 clock_v2_0/Bd ota_1/p2_b 4.69fF
C1681 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0.00fF
C1682 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_561_413# 0.00fF
C1683 sky130_fd_sc_hd__clkinv_4_1/Y ota_1/p2 0.00fF
C1684 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# -0.00fF
C1685 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C1686 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.06fF
C1687 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C1688 sky130_fd_sc_hd__clkinv_4_3/Y d_probe_1 1.63fF
C1689 clock_v2_0/p1d clock_v2_0/B 0.06fF
C1690 VSS ota_w_test_0/sc_cmfb_0/transmission_gate_8/in -0.75fF
C1691 ota_1/m1_n2176_n12171# ota_1/m1_n1659_n11581# 0.02fF
C1692 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0.00fF
C1693 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# -0.12fF
C1694 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C1695 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C1696 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# ota_1/p1 0.06fF
C1697 sky130_fd_sc_hd__mux4_1_0/a_834_97# ota_1/p2 0.00fF
C1698 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0.02fF
C1699 VSS clock_v2_0/p1d 2.98fF
C1700 clock_v2_0/Bd ota_1/p2 4.85fF
C1701 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0.01fF
C1702 ota_1/ip rst_n 0.00fF
C1703 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_2/en_b 0.00fF
C1704 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VDD 0.14fF
C1705 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.00fF
C1706 ota_w_test_0/cm ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# 0.01fF
C1707 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# ota_1/in 0.14fF
C1708 transmission_gate_18/in transmission_gate_0/out 0.05fF
C1709 d_clk_grp_1_ctrl_1 clock_v2_0/B 0.00fF
C1710 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A -0.04fF
C1711 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.00fF
C1712 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# 0.01fF
C1713 sky130_fd_sc_hd__clkinv_4_4/Y d_probe_1 0.09fF
C1714 comparator_v2_0/li_n2324_818# VDD 0.30fF
C1715 ota_1/p1 clock_v2_0/A_b 6.78fF
C1716 ota_w_test_0/sc_cmfb_0/transmission_gate_3/out ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# 0.00fF
C1717 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.05fF
C1718 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# 0.02fF
C1719 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# 0.82fF
C1720 clock_v2_0/Ad clock_v2_0/p2 0.04fF
C1721 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0.04fF
C1722 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# transmission_gate_17/in 0.11fF
C1723 sky130_fd_sc_hd__mux4_1_2/a_247_21# clock_v2_0/p2_b 0.04fF
C1724 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# -0.00fF
C1725 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# -0.14fF
C1726 transmission_gate_5/in ota_w_test_0/in 0.08fF
C1727 VSS d_clk_grp_1_ctrl_1 1.29fF
C1728 VDD a_mux4_en_1/transmission_gate_3/en_b 0.80fF
C1729 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0.00fF
C1730 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_1/a_277_47# 0.06fF
C1731 ota_w_test_0/on debug 0.00fF
C1732 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# -0.00fF
C1733 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# 0.03fF
C1734 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0.07fF
C1735 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/p1_b -0.00fF
C1736 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_1/p1_b 0.00fF
C1737 d_clk_grp_1_ctrl_0 clock_v2_0/A_b 0.12fF
C1738 sky130_fd_sc_hd__mux4_1_1/a_27_413# clock_v2_0/Ad 0.02fF
C1739 sky130_fd_sc_hd__mux4_1_2/X VDD 0.60fF
C1740 a_mod_grp_ctrl_0 a_mux2_en_0/switch_5t_1/in 0.02fF
C1741 ota_w_test_0/m1_2462_n3318# ota_w_test_0/m1_6690_n8907# 0.00fF
C1742 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# -0.14fF
C1743 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/c1_n260_n210# -0.09fF
C1744 sky130_fd_sc_hd__mux4_1_2/a_668_97# clock_v2_0/A_b 0.00fF
C1745 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A -0.00fF
C1746 comparator_v2_0/li_n2324_818# ota_1/op -0.00fF
C1747 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C1748 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.03fF
C1749 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0.00fF
C1750 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0.13fF
C1751 VSS a_mux4_en_1/switch_5t_0/en_b 0.30fF
C1752 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# ota_1/sc_cmfb_0/transmission_gate_4/out 0.00fF
C1753 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.12fF
C1754 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0.07fF
C1755 ota_1/p2_b clock_v2_0/p1d 1.38fF
C1756 a_mux4_en_0/in0 clock_v2_0/B 0.04fF
C1757 sky130_fd_sc_hd__mux4_1_2/a_923_363# VDD -0.02fF
C1758 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_1/a_834_97# 0.00fF
C1759 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C1760 a_mux4_en_0/switch_5t_0/en a_mod_grp_ctrl_1 0.02fF
C1761 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0.10fF
C1762 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# -0.00fF
C1763 sky130_fd_sc_hd__mux4_1_2/a_757_363# clock_v2_0/A_b 0.00fF
C1764 sky130_fd_sc_hd__mux4_1_3/a_1478_413# ota_1/p1 0.00fF
C1765 sky130_fd_sc_hd__clkinv_4_1/Y VDD -0.56fF
C1766 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# 0.03fF
C1767 clock_v2_0/B ota_w_test_0/in 0.00fF
C1768 sky130_fd_sc_hd__mux4_1_1/a_1478_413# clock_v2_0/p1d 0.00fF
C1769 a_mux4_en_0/switch_5t_2/in a_mux4_en_0/switch_5t_2/transmission_gate_1/in -0.00fF
C1770 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C1771 VDD transmission_gate_2/out 0.41fF
C1772 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0.07fF
C1773 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0.00fF
C1774 VSS a_mux4_en_0/in0 3.44fF
C1775 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0.00fF
C1776 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# 0.11fF
C1777 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# 0.32fF
C1778 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# 0.11fF
C1779 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# ota_1/op 0.06fF
C1780 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X -0.01fF
C1781 sky130_fd_sc_hd__mux4_1_0/a_834_97# VDD 0.00fF
C1782 VSS ota_w_test_0/in 0.52fF
C1783 clock_v2_0/Ad_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_6/a_110_47# -0.00fF
C1784 ota_1/p2 clock_v2_0/p1d 2.20fF
C1785 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# 0.02fF
C1786 ota_w_test_0/op a_mux2_en_0/switch_5t_1/in 0.02fF
C1787 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# -0.00fF
C1788 clock_v2_0/Bd VDD 5.73fF
C1789 a_mod_grp_ctrl_0 a_mux4_en_0/sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C1790 transmission_gate_26/en transmission_gate_5/in 1.84fF
C1791 a_mux4_en_1/in2 ota_w_test_0/m1_12232_n10488# 0.28fF
C1792 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.01fF
C1793 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n930_n880# 0.11fF
C1794 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# VDD 0.07fF
C1795 ota_1/m1_6690_n8907# ota_1/bias_c -0.00fF
C1796 ota_w_test_0/m1_2462_n3318# ota_w_test_0/op -0.00fF
C1797 a_mux4_en_1/in2 clock_v2_0/A 0.03fF
C1798 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0.00fF
C1799 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# VDD 0.40fF
C1800 transmission_gate_31/out transmission_gate_2/out 0.27fF
C1801 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n930_n880# 0.11fF
C1802 sky130_fd_sc_hd__mux4_1_1/X d_clk_grp_2_ctrl_0 0.00fF
C1803 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0.00fF
C1804 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/c1_n530_n480# 0.79fF
C1805 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# clock_v2_0/p1d_b 0.44fF
C1806 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# -0.00fF
C1807 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.00fF
C1808 VSS sky130_fd_sc_hd__mux4_1_3/a_277_47# -0.64fF
C1809 debug a_mux4_en_0/switch_5t_3/in 0.00fF
C1810 sky130_fd_sc_hd__mux4_1_0/a_834_97# clock_v2_0/Ad_b 0.00fF
C1811 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0.07fF
C1812 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.03fF
C1813 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n930_n880# 2.09fF
C1814 clock_v2_0/Bd clock_v2_0/Ad_b 4.65fF
C1815 a_mux2_en_0/switch_5t_0/transmission_gate_1/in a_mux2_en_0/switch_5t_1/en -0.00fF
C1816 transmission_gate_0/out transmission_gate_8/in -0.54fF
C1817 ota_1/p1 a_mux4_en_1/in1 0.09fF
C1818 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.00fF
C1819 sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# -0.14fF
C1820 VSS ota_1/m1_n1659_n11581# 0.89fF
C1821 ota_1/p1_b clock_v2_0/p2_b 3.19fF
C1822 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/X 0.25fF
C1823 transmission_gate_6/in ota_w_test_0/in 0.04fF
C1824 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/A -0.00fF
C1825 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# 0.13fF
C1826 ota_w_test_0/m1_2463_n5585# VDD 1.05fF
C1827 VSS a_mux2_en_1/switch_5t_0/in -2.37fF
C1828 VSS ota_1/m1_12118_n9704# 0.00fF
C1829 sky130_fd_sc_hd__mux4_1_2/a_1290_413# VDD 0.08fF
C1830 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# ota_1/p1 0.00fF
C1831 debug a_mod_grp_ctrl_1 5.00fF
C1832 transmission_gate_26/en clock_v2_0/B 0.08fF
C1833 sky130_fd_sc_hd__mux4_1_0/a_277_47# d_clk_grp_2_ctrl_0 0.03fF
C1834 VDD a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.08fF
C1835 a_mux4_en_0/in0 ota_1/p2_b 0.02fF
C1836 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X -0.01fF
C1837 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# -0.00fF
C1838 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# 0.07fF
C1839 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0.10fF
C1840 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.03fF
C1841 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# VDD 0.03fF
C1842 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C1843 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A -0.00fF
C1844 transmission_gate_32/out in 0.03fF
C1845 ota_w_test_0/m1_11940_n10482# a_mux4_en_1/in2 0.04fF
C1846 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X -0.01fF
C1847 VSS transmission_gate_26/en 2.18fF
C1848 clock_v2_0/p1d_b transmission_gate_2/out 0.45fF
C1849 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_3/en_b -0.00fF
C1850 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/A -0.00fF
C1851 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# 0.03fF
C1852 ota_w_test_0/sc_cmfb_0/transmission_gate_8/in VDD 0.07fF
C1853 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.00fF
C1854 a_mux4_en_0/in0 ota_1/p2 0.04fF
C1855 sky130_fd_sc_hd__mux4_1_0/a_834_97# clock_v2_0/p1d_b 0.00fF
C1856 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/c1_n260_n210# 0.03fF
C1857 clock_v2_0/Bd clock_v2_0/p1d_b 0.47fF
C1858 transmission_gate_18/in rst_n 0.11fF
C1859 clock_v2_0/Bd_b ota_1/p1_b 0.09fF
C1860 a_mux4_en_1/switch_5t_1/en_b a_mux4_en_1/switch_5t_1/in 0.00fF
C1861 VDD clock_v2_0/p1d 6.30fF
C1862 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X -0.00fF
C1863 ota_w_test_0/on clock_v2_0/A 0.05fF
C1864 sky130_fd_sc_hd__mux4_1_2/a_193_47# clock_v2_0/B_b 0.00fF
C1865 a_mod_grp_ctrl_0 ota_1/p1_b 0.06fF
C1866 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_1/sc_cmfb_0/transmission_gate_9/in 0.01fF
C1867 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C1868 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# -0.17fF
C1869 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0.00fF
C1870 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# ota_1/p1_b 0.04fF
C1871 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C1872 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# -0.00fF
C1873 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# 0.20fF
C1874 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y -0.00fF
C1875 transmission_gate_26/en transmission_gate_6/in 0.09fF
C1876 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/c1_n260_n210# ota_1/op 0.03fF
C1877 d_clk_grp_1_ctrl_1 VDD 3.52fF
C1878 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# 0.11fF
C1879 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.02fF
C1880 ota_1/ip ota_1/p1_b 0.09fF
C1881 transmission_gate_31/out clock_v2_0/p1d 0.20fF
C1882 clock_v2_0/Ad_b clock_v2_0/p1d 6.21fF
C1883 onebit_dac_1/v_b clock_v2_0/p2_b 0.01fF
C1884 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/X 0.03fF
C1885 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# -0.13fF
C1886 transmission_gate_17/in a_mux4_en_1/in1 0.00fF
C1887 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# -0.00fF
C1888 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_634_159# -0.00fF
C1889 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C1890 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_0/a_113_47# a_mod_grp_ctrl_1 0.00fF
C1891 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/c1_n260_n210# 0.03fF
C1892 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0.07fF
C1893 transmission_gate_26/en ota_1/p2_b 0.44fF
C1894 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# ota_1/p1_b 0.03fF
C1895 a_mux4_en_0/switch_5t_2/in a_mux4_en_0/switch_5t_2/en 0.00fF
C1896 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980# 0.29fF
C1897 a_mux2_en_1/transmission_gate_1/en_b ota_1/on 0.00fF
C1898 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C1899 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# ota_1/on 0.03fF
C1900 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# VDD 0.00fF
C1901 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C1902 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C1903 ota_w_test_0/cm debug 0.02fF
C1904 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.00fF
C1905 a_mux4_en_0/in1 ota_w_test_0/m1_1038_n2886# 0.03fF
C1906 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A -0.01fF
C1907 VSS ota_w_test_0/sc_cmfb_0/transmission_gate_9/in -0.68fF
C1908 VSS ota_1/sc_cmfb_0/transmission_gate_6/in 0.26fF
C1909 ota_w_test_0/op ota_1/p1_b 0.23fF
C1910 VDD a_mux4_en_1/switch_5t_0/en_b 0.17fF
C1911 transmission_gate_26/en ota_1/in 0.02fF
C1912 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980# -0.43fF
C1913 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.08fF
C1914 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n930_n880# 0.01fF
C1915 transmission_gate_26/en ota_1/p2 0.66fF
C1916 VSS a_probe_1 -1.12fF
C1917 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# 0.13fF
C1918 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.27fF
C1919 a_mux2_en_1/switch_5t_0/transmission_gate_1/in a_mux2_en_1/switch_5t_1/transmission_gate_1/in -0.00fF
C1920 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.01fF
C1921 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.03fF
C1922 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# ota_1/p1_b 0.09fF
C1923 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0.06fF
C1924 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C1925 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/c1_n260_n210# 0.03fF
C1926 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/A -0.09fF
C1927 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# -0.00fF
C1928 sky130_fd_sc_hd__mux4_1_3/a_193_413# ota_1/p1_b 0.06fF
C1929 a_mux4_en_0/in0 VDD -1.07fF
C1930 clock_v2_0/p1d_b clock_v2_0/p1d 19.79fF
C1931 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_1/en_b 0.00fF
C1932 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0.08fF
C1933 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C1934 transmission_gate_32/out clock_v2_0/p2 0.28fF
C1935 VDD ota_w_test_0/in 1.25fF
C1936 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0.01fF
C1937 ota_1/bias_a ota_1/p1_b 2.14fF
C1938 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.00fF
C1939 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y 0.28fF
C1940 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C1941 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.00fF
C1942 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.00fF
C1943 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y 0.26fF
C1944 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.42fF
C1945 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# -0.14fF
C1946 ota_1/cmc ota_1/p1 0.36fF
C1947 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C1948 a_mux4_en_0/in0 clock_v2_0/Ad_b 0.05fF
C1949 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0.03fF
C1950 sky130_fd_sc_hd__mux4_1_3/a_277_47# VDD 0.17fF
C1951 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.00fF
C1952 clock_v2_0/A a_mod_grp_ctrl_1 0.06fF
C1953 VSS a_mux4_en_0/switch_5t_0/transmission_gate_1/in 0.37fF
C1954 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.01fF
C1955 clock_v2_0/Ad_b ota_w_test_0/in 1.65fF
C1956 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0.03fF
C1957 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C1958 a_mux4_en_0/in1 a_mux4_en_0/transmission_gate_3/en_b 0.02fF
C1959 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/X 0.01fF
C1960 VSS transmission_gate_21/in 0.50fF
C1961 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# VDD -0.00fF
C1962 ota_1/sc_cmfb_0/transmission_gate_6/in ota_1/p2_b 0.02fF
C1963 comparator_v2_0/li_n2324_818# ota_1/on 0.00fF
C1964 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/c1_n260_n210# 0.03fF
C1965 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# 0.12fF
C1966 ota_w_test_0/m1_n947_n12836# ota_w_test_0/m1_n1659_n11581# 0.01fF
C1967 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n930_n880# 2.09fF
C1968 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0.09fF
C1969 ota_1/m1_n1659_n11581# VDD 0.27fF
C1970 VSS a_mux4_en_1/sky130_fd_sc_hd__nand2_1_3/a_113_47# 0.00fF
C1971 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.00fF
C1972 a_mux2_en_1/switch_5t_0/in VDD 0.00fF
C1973 VSS sky130_fd_sc_hd__mux4_1_1/a_923_363# -0.11fF
C1974 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A -0.01fF
C1975 VSS ota_1/sc_cmfb_0/transmission_gate_9/in -1.63fF
C1976 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C1977 a_mux4_en_1/in2 ota_w_test_0/m1_11242_n9716# 0.05fF
C1978 ota_w_test_0/m1_2462_n3318# ota_w_test_0/on 0.01fF
C1979 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.09fF
C1980 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# -0.00fF
C1981 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0.09fF
C1982 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.07fF
C1983 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# -0.31fF
C1984 ota_1/sc_cmfb_0/transmission_gate_6/in ota_1/p2 0.00fF
C1985 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# transmission_gate_5/in 0.18fF
C1986 VSS a_mux4_en_1/switch_5t_2/en_b 0.28fF
C1987 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n930_n880# 2.04fF
C1988 debug clk 0.20fF
C1989 VSS i_bias_2 4.38fF
C1990 ota_1/sc_cmfb_0/transmission_gate_9/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0.01fF
C1991 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y -0.01fF
C1992 clock_v2_0/p2 clock_v2_0/p2_b 12.88fF
C1993 ota_1/bias_a ota_1/m1_2462_n3318# 0.00fF
C1994 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0.08fF
C1995 transmission_gate_26/en VDD 3.34fF
C1996 ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.03fF
C1997 ota_1/bias_b ota_1/m1_n6302_n3889# 0.01fF
C1998 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# -0.00fF
C1999 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0.00fF
C2000 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C2001 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_193_413# -0.00fF
C2002 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# transmission_gate_0/out 1.54fF
C2003 ota_1/bias_b ota_1/m1_2463_n5585# 0.01fF
C2004 ota_1/m1_n1659_n11581# ota_1/op 0.00fF
C2005 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0.00fF
C2006 clock_v2_0/p1d sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 0.15fF
C2007 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# -0.00fF
C2008 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# 0.14fF
C2009 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# 0.11fF
C2010 a_mux4_en_0/in0 a_mux4_en_0/switch_5t_0/in 0.00fF
C2011 transmission_gate_21/in ota_1/p2_b 0.02fF
C2012 transmission_gate_31/out transmission_gate_26/en 0.05fF
C2013 a_mux4_en_0/in2 a_mux4_en_0/transmission_gate_3/en_b 0.02fF
C2014 a_mux4_en_0/in1 ota_w_test_0/m1_n5574_n13620# 1.39fF
C2015 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C2016 VSS ota_1/m1_n5574_n13620# 3.43fF
C2017 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C2018 ota_1/p1 d_clk_grp_1_ctrl_0 0.00fF
C2019 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# VDD 0.10fF
C2020 VSS sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.06fF
C2021 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# VDD 0.53fF
C2022 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0.00fF
C2023 d_probe_2 d_clk_grp_2_ctrl_1 0.52fF
C2024 transmission_gate_26/en ota_1/op 0.30fF
C2025 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C2026 a_mux4_en_1/in2 ota_1/p1_b 0.03fF
C2027 sky130_fd_sc_hd__mux4_1_3/a_193_47# clock_v2_0/A_b 0.01fF
C2028 VSS sky130_fd_sc_hd__mux4_1_2/a_193_47# -0.00fF
C2029 clock_v2_0/Bd_b clock_v2_0/p2 0.06fF
C2030 a_mod_grp_ctrl_1 a_mux4_en_0/switch_5t_2/en_b -0.00fF
C2031 transmission_gate_18/in ota_1/p1_b 0.19fF
C2032 d_probe_0 sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.00fF
C2033 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# 0.09fF
C2034 ota_1/bias_c ota_1/m1_2463_n5585# 0.00fF
C2035 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.01fF
C2036 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# 0.21fF
C2037 ota_w_test_0/cm clock_v2_0/A 0.31fF
C2038 a_mux4_en_0/in1 a_mux4_en_0/in2 2.80fF
C2039 transmission_gate_21/in ota_1/in 0.30fF
C2040 a_mux2_en_0/switch_5t_0/transmission_gate_1/in a_mux2_en_0/switch_5t_0/in 0.00fF
C2041 a_mux4_en_1/switch_5t_2/en a_mux4_en_1/switch_5t_2/en_b 0.00fF
C2042 transmission_gate_21/in ota_1/p2 0.62fF
C2043 a_mod_grp_ctrl_0 clock_v2_0/p2 0.04fF
C2044 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# transmission_gate_17/in -1.08fF
C2045 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_1290_413# -0.00fF
C2046 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/c1_n260_n210# -0.12fF
C2047 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_975_413# 0.00fF
C2048 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0.00fF
C2049 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/A VDD -0.00fF
C2050 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C2051 ota_1/bias_b ota_1/p1_b 0.02fF
C2052 sky130_fd_sc_hd__mux4_1_2/a_668_97# d_clk_grp_1_ctrl_0 0.00fF
C2053 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# -0.12fF
C2054 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# -0.00fF
C2055 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B 0.95fF
C2056 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# ota_1/op 0.03fF
C2057 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/A 0.00fF
C2058 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0.09fF
C2059 i_bias_2 ota_1/in 0.17fF
C2060 VSS a_mux4_en_0/switch_5t_1/en_b 0.28fF
C2061 debug clock_v2_0/A_b 0.06fF
C2062 ota_w_test_0/sc_cmfb_0/transmission_gate_9/in VDD -1.38fF
C2063 a_mux2_en_0/switch_5t_1/in a_mod_grp_ctrl_1 0.02fF
C2064 ota_1/sc_cmfb_0/transmission_gate_6/in VDD 0.16fF
C2065 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.02fF
C2066 transmission_gate_26/en clock_v2_0/p1d_b 0.17fF
C2067 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.00fF
C2068 sky130_fd_sc_hd__mux4_1_2/a_757_363# d_clk_grp_1_ctrl_0 -0.00fF
C2069 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0.05fF
C2070 transmission_gate_23/in transmission_gate_19/in 0.09fF
C2071 a_probe_1 VDD 2.27fF
C2072 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D 0.07fF
C2073 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_1/in 0.00fF
C2074 VSS sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.06fF
C2075 sky130_fd_sc_hd__mux4_1_0/a_247_21# ota_1/p2_b 0.01fF
C2076 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0.03fF
C2077 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# VDD 0.01fF
C2078 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# VDD 0.00fF
C2079 ota_1/p1 transmission_gate_17/in 0.19fF
C2080 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.07fF
C2081 ota_w_test_0/sc_cmfb_0/transmission_gate_3/out ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# 0.06fF
C2082 a_mux4_en_1/switch_5t_3/en_b a_mux4_en_1/switch_5t_3/transmission_gate_1/in -0.00fF
C2083 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0.04fF
C2084 ota_1/bias_c ota_1/p1_b 1.03fF
C2085 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.04fF
C2086 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0.06fF
C2087 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y 0.00fF
C2088 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# 0.74fF
C2089 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0.00fF
C2090 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480# ota_1/p1_b 0.04fF
C2091 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0.03fF
C2092 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0.18fF
C2093 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y -0.26fF
C2094 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# VDD 0.52fF
C2095 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# 0.03fF
C2096 ota_w_test_0/cm rst_n 0.03fF
C2097 ota_1/sc_cmfb_0/transmission_gate_6/in ota_1/op 0.01fF
C2098 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0.07fF
C2099 sky130_fd_sc_hd__mux4_1_0/a_247_21# ota_1/p2 0.03fF
C2100 ota_w_test_0/on ota_1/p1_b 0.18fF
C2101 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0.08fF
C2102 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X -0.00fF
C2103 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y VDD 0.40fF
C2104 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.01fF
C2105 sky130_fd_sc_hd__mux4_1_3/a_193_413# clock_v2_0/p2 0.00fF
C2106 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0.05fF
C2107 sky130_fd_sc_hd__mux4_1_2/a_1478_413# d_clk_grp_1_ctrl_1 -0.00fF
C2108 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# -0.02fF
C2109 ota_1/bias_b ota_1/m1_2462_n3318# 0.01fF
C2110 VDD a_mux4_en_0/switch_5t_0/transmission_gate_1/in -0.87fF
C2111 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# 0.09fF
C2112 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# -0.00fF
C2113 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980# -0.34fF
C2114 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# 0.17fF
C2115 ota_1/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0.13fF
C2116 transmission_gate_21/in VDD 2.75fF
C2117 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# 0.11fF
C2118 clock_v2_0/Ad clock_v2_0/Bd 7.70fF
C2119 VSS transmission_gate_19/out 0.08fF
C2120 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C2121 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0.06fF
C2122 VSS a_mux4_en_0/switch_5t_3/en_b 0.17fF
C2123 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.03fF
C2124 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# 0.03fF
C2125 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0.04fF
C2126 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.01fF
C2127 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0.14fF
C2128 sky130_fd_sc_hd__mux4_1_1/a_923_363# VDD -0.01fF
C2129 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0.00fF
C2130 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0.09fF
C2131 transmission_gate_8/in ota_1/p1_b 0.10fF
C2132 ota_1/sc_cmfb_0/transmission_gate_9/in VDD 0.62fF
C2133 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0.00fF
C2134 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_1/X 0.32fF
C2135 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0.08fF
C2136 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0.00fF
C2137 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# 0.14fF
C2138 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0.00fF
C2139 a_mux4_en_1/switch_5t_2/transmission_gate_1/in a_mux4_en_1/switch_5t_2/en_b 0.00fF
C2140 VDD a_mux4_en_1/switch_5t_2/en_b 0.08fF
C2141 transmission_gate_31/out transmission_gate_21/in 0.06fF
C2142 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# 0.02fF
C2143 i_bias_2 VDD 7.45fF
C2144 ota_1/bias_c ota_1/m1_2462_n3318# 0.01fF
C2145 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in a_mux4_en_1/in2 -0.00fF
C2146 a_mux4_en_0/switch_5t_0/en_b a_mux4_en_0/switch_5t_0/en -0.00fF
C2147 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# -0.01fF
C2148 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y 0.00fF
C2149 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_1/X 0.01fF
C2150 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0.08fF
C2151 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_1/p1_b 0.06fF
C2152 a_mux4_en_0/in1 clock_v2_0/B_b 0.04fF
C2153 VSS sky130_fd_sc_hd__mux4_1_0/a_757_363# -0.01fF
C2154 transmission_gate_21/in ota_1/op 0.46fF
C2155 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.01fF
C2156 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# -0.28fF
C2157 sky130_fd_sc_hd__clkinv_4_4/Y clock_v2_0/A_b 0.00fF
C2158 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# 0.02fF
C2159 sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# 0.03fF
C2160 a_mux4_en_1/in1 debug 0.02fF
C2161 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# -0.00fF
C2162 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.06fF
C2163 ota_w_test_0/ip clock_v2_0/B_b 0.19fF
C2164 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y -0.00fF
C2165 ota_1/sc_cmfb_0/transmission_gate_9/in ota_1/op 0.00fF
C2166 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# -0.00fF
C2167 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X -0.00fF
C2168 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# ota_1/in 0.26fF
C2169 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0.16fF
C2170 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.07fF
C2171 a_mux4_en_1/switch_5t_3/en_b a_mod_grp_ctrl_1 0.39fF
C2172 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# 0.03fF
C2173 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.03fF
C2174 ota_1/m1_n5574_n13620# VDD 0.77fF
C2175 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C2176 transmission_gate_19/out ota_1/p2_b 0.27fF
C2177 sky130_fd_sc_hd__mux4_1_3/a_757_363# clock_v2_0/B_b 0.00fF
C2178 VSS onebit_dac_1/out 1.06fF
C2179 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.00fF
C2180 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.02fF
C2181 sky130_fd_sc_hd__mux4_1_0/a_247_21# VDD 0.03fF
C2182 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/c1_n260_n210# 0.03fF
C2183 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y VSS 0.06fF
C2184 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.00fF
C2185 VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.23fF
C2186 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# -0.07fF
C2187 clock_v2_0/sky130_fd_sc_hd__nand2_1_2/B clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A -0.00fF
C2188 sky130_fd_sc_hd__mux4_1_0/a_27_47# d_clk_grp_2_ctrl_0 -0.00fF
C2189 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# ota_1/in 0.03fF
C2190 VSS a_mux4_en_1/switch_5t_2/in 0.05fF
C2191 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.00fF
C2192 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# 0.11fF
C2193 ota_w_test_0/op ota_w_test_0/m1_n947_n12836# 0.01fF
C2194 transmission_gate_19/out ota_1/in 1.45fF
C2195 ota_1/p1_b a_mod_grp_ctrl_1 0.07fF
C2196 transmission_gate_19/out ota_1/p2 0.21fF
C2197 clock_v2_0/A clock_v2_0/A_b 18.36fF
C2198 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# VDD 0.95fF
C2199 clock_v2_0/Ad clock_v2_0/p1d 5.92fF
C2200 a_mux4_en_0/switch_5t_0/in a_mux4_en_0/switch_5t_0/transmission_gate_1/in -0.00fF
C2201 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.03fF
C2202 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# clock_v2_0/p1d 0.04fF
C2203 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.03fF
C2204 sky130_fd_sc_hd__mux4_1_1/a_923_363# clock_v2_0/p1d_b -0.50fF
C2205 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/A -0.00fF
C2206 a_mux4_en_0/in2 clock_v2_0/B_b 0.04fF
C2207 a_mux4_en_0/switch_5t_0/en_b debug 0.00fF
C2208 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47# VDD -0.00fF
C2209 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.07fF
C2210 sky130_fd_sc_hd__mux4_1_2/a_750_97# clock_v2_0/A_b 0.00fF
C2211 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B 0.05fF
C2212 sky130_fd_sc_hd__mux4_1_3/X clock_v2_0/A_b 0.00fF
C2213 sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/c1_n260_n210# ota_1/op 0.03fF
C2214 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# transmission_gate_19/in 0.03fF
C2215 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in ota_w_test_0/on -0.00fF
C2216 d_probe_2 d_clk_grp_2_ctrl_0 0.30fF
C2217 a_mux4_en_0/switch_5t_1/en_b VDD 0.17fF
C2218 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/X -0.00fF
C2219 ota_1/m1_n1659_n11581# ota_1/on 0.00fF
C2220 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# 0.11fF
C2221 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# ota_1/in 0.03fF
C2222 ota_w_test_0/cm ota_w_test_0/m1_11242_n9716# -0.01fF
C2223 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0.03fF
C2224 sky130_fd_sc_hd__mux4_1_0/a_757_363# ota_1/p2 0.06fF
C2225 a_mux4_en_1/in2 ota_w_test_0/m1_11356_n10481# 0.05fF
C2226 ota_1/p2_b onebit_dac_1/out 0.00fF
C2227 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# 0.02fF
C2228 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C2229 sky130_fd_sc_hd__mux4_1_3/a_247_21# VDD 0.07fF
C2230 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C2231 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C2232 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0.08fF
C2233 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.00fF
C2234 VSS ota_w_test_0/m1_1038_n2886# 0.41fF
C2235 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# -0.00fF
C2236 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X -0.00fF
C2237 d_clk_grp_1_ctrl_0 d_clk_grp_2_ctrl_0 0.00fF
C2238 a_mux4_en_1/switch_5t_2/en a_mux4_en_1/switch_5t_2/in 0.00fF
C2239 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A VDD 0.05fF
C2240 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# -0.00fF
C2241 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0.01fF
C2242 transmission_gate_26/en ota_1/on 0.15fF
C2243 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0.00fF
C2244 ota_1/p2 onebit_dac_1/out 0.00fF
C2245 VSS a_probe_3 2.76fF
C2246 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_0/in 0.01fF
C2247 d_clk_grp_2_ctrl_0 d_clk_grp_2_ctrl_1 2.29fF
C2248 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# -0.13fF
C2249 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_466_413# -0.00fF
C2250 sky130_fd_sc_hd__mux4_1_1/a_247_21# clock_v2_0/p1d 0.01fF
C2251 rst_n clock_v2_0/A_b 0.25fF
C2252 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C2253 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.01fF
C2254 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0.07fF
C2255 a_mux4_en_1/switch_5t_1/en_b a_mod_grp_ctrl_1 0.08fF
C2256 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.00fF
C2257 VSS ota_1/sc_cmfb_0/transmission_gate_4/out 0.55fF
C2258 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# 0.92fF
C2259 clock_v2_0/Ad a_mux4_en_0/in0 0.04fF
C2260 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# clock_v2_0/p1d_b 0.33fF
C2261 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# -0.00fF
C2262 ota_w_test_0/ip transmission_gate_5/in 0.04fF
C2263 clock_v2_0/Ad ota_w_test_0/in 0.02fF
C2264 ota_w_test_0/cm ota_1/p1_b 0.26fF
C2265 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.07fF
C2266 transmission_gate_19/out VDD 0.82fF
C2267 VDD a_mux4_en_0/switch_5t_3/en_b -0.20fF
C2268 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0.13fF
C2269 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.05fF
C2270 sky130_fd_sc_hd__mux4_1_3/a_750_97# clock_v2_0/p2_b 0.00fF
C2271 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0.04fF
C2272 ota_1/p1 ota_1/m1_1038_n2886# 0.08fF
C2273 a_mux4_en_1/in1 clock_v2_0/A 0.04fF
C2274 d_probe_0 d_clk_grp_1_ctrl_0 0.29fF
C2275 i_bias_1 clock_v2_0/A 0.12fF
C2276 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# VDD 0.08fF
C2277 ota_1/cmc ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0.00fF
C2278 VSS a_mux4_en_0/transmission_gate_3/en_b 0.29fF
C2279 transmission_gate_31/out transmission_gate_19/out 0.84fF
C2280 a_mux4_en_0/in1 clock_v2_0/B 0.04fF
C2281 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y 0.09fF
C2282 ota_1/m1_n208_n2883# ota_1/m1_n6302_n3889# 0.01fF
C2283 transmission_gate_9/in ota_1/p1_b 0.02fF
C2284 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/X VDD 0.05fF
C2285 ota_1/m1_n208_n2883# ota_1/m1_2463_n5585# 0.02fF
C2286 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.06fF
C2287 sky130_fd_sc_hd__mux4_1_0/a_757_363# VDD 0.04fF
C2288 VSS comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A 0.00fF
C2289 transmission_gate_19/out ota_1/op 0.01fF
C2290 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.00fF
C2291 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0.05fF
C2292 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# -0.08fF
C2293 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# -0.24fF
C2294 ota_w_test_0/ip clock_v2_0/B 0.11fF
C2295 a_mux4_en_1/transmission_gate_3/en_b a_mux4_en_1/switch_5t_1/in -0.00fF
C2296 VSS a_mux4_en_0/in1 5.18fF
C2297 VSS d_probe_3 1.95fF
C2298 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0.09fF
C2299 debug a_mux4_en_1/switch_5t_3/in 0.01fF
C2300 transmission_gate_32/out transmission_gate_2/out 0.26fF
C2301 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0.01fF
C2302 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C2303 VSS ota_w_test_0/ip 0.76fF
C2304 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0.00fF
C2305 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# 0.03fF
C2306 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# VDD 0.00fF
C2307 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# transmission_gate_5/in 0.18fF
C2308 sky130_fd_sc_hd__mux4_1_0/a_757_363# clock_v2_0/Ad_b 0.00fF
C2309 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y -0.00fF
C2310 onebit_dac_1/out VDD 0.36fF
C2311 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0.06fF
C2312 transmission_gate_26/en clock_v2_0/Ad 0.06fF
C2313 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# VDD 0.05fF
C2314 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y -0.00fF
C2315 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.00fF
C2316 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# 0.03fF
C2317 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y VDD 0.02fF
C2318 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# 0.03fF
C2319 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# ota_1/p1 0.23fF
C2320 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# 0.03fF
C2321 sky130_fd_sc_hd__mux4_1_3/a_757_363# VSS -0.01fF
C2322 a_mod_grp_ctrl_0 a_mux2_en_1/switch_5t_1/transmission_gate_1/in -0.00fF
C2323 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C2324 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0.00fF
C2325 a_mux4_en_1/switch_5t_2/transmission_gate_1/in a_mux4_en_1/switch_5t_2/in -0.00fF
C2326 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A -0.00fF
C2327 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_8/a_110_47# -0.00fF
C2328 VDD a_mux4_en_1/switch_5t_2/in 0.28fF
C2329 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0.41fF
C2330 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0.05fF
C2331 sky130_fd_sc_hd__mux4_1_2/X clock_v2_0/p2_b 0.01fF
C2332 sky130_fd_sc_hd__mux4_1_1/a_1290_413# d_clk_grp_2_ctrl_1 0.03fF
C2333 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# 0.00fF
C2334 transmission_gate_19/out clock_v2_0/p1d_b 0.58fF
C2335 ota_1/p1 debug 0.07fF
C2336 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# -0.00fF
C2337 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A -0.00fF
C2338 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.00fF
C2339 VSS ota_w_test_0/m1_n5574_n13620# 1.00fF
C2340 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# 0.03fF
C2341 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.09fF
C2342 transmission_gate_31/out onebit_dac_1/out 0.13fF
C2343 ota_1/m1_n208_n2883# ota_1/p1_b 0.09fF
C2344 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# -0.16fF
C2345 a_mux4_en_0/in2 clock_v2_0/B 0.04fF
C2346 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y -0.00fF
C2347 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C2348 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C2349 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# clock_v2_0/p2 0.03fF
C2350 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C2351 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0.16fF
C2352 transmission_gate_6/in ota_w_test_0/ip 0.08fF
C2353 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0.00fF
C2354 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# -0.12fF
C2355 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# -0.37fF
C2356 sky130_fd_sc_hd__mux4_1_3/a_834_97# clock_v2_0/B_b 0.00fF
C2357 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# 0.18fF
C2358 clock_v2_0/p2 a_mod_grp_ctrl_1 0.05fF
C2359 transmission_gate_21/in ota_1/on 0.13fF
C2360 sky130_fd_sc_hd__mux4_1_2/a_923_363# clock_v2_0/p2_b -0.50fF
C2361 VSS a_mux4_en_0/in2 -2.18fF
C2362 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.08fF
C2363 transmission_gate_26/en ota_1/cm 0.49fF
C2364 ota_w_test_0/m1_n2176_n12171# ota_w_test_0/m1_n947_n12836# 0.01fF
C2365 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# -0.00fF
C2366 onebit_dac_0/out transmission_gate_0/out 0.04fF
C2367 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# 0.12fF
C2368 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# VDD 0.46fF
C2369 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0.00fF
C2370 sky130_fd_sc_hd__mux4_1_0/a_757_363# clock_v2_0/p1d_b 0.00fF
C2371 a_mux4_en_0/switch_5t_1/transmission_gate_1/in a_mux4_en_0/switch_5t_1/in -0.00fF
C2372 clock_v2_0/p2_b transmission_gate_2/out 0.13fF
C2373 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/c1_n260_n210# 0.03fF
C2374 ota_w_test_0/m1_n947_n12836# ota_w_test_0/on 0.06fF
C2375 VSS a_mux2_en_1/switch_5t_1/in 0.04fF
C2376 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/sc_cmfb_0/transmission_gate_9/in -0.00fF
C2377 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_923_363# 0.01fF
C2378 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# -0.00fF
C2379 a_mod_grp_ctrl_0 a_mux4_en_1/transmission_gate_3/en_b 0.01fF
C2380 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0.03fF
C2381 VSS a_mux2_en_0/switch_5t_1/transmission_gate_1/in -0.17fF
C2382 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0.00fF
C2383 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X -0.01fF
C2384 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# ota_1/p2_b 0.49fF
C2385 clock_v2_0/Bd clock_v2_0/p2_b 0.05fF
C2386 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0.05fF
C2387 ota_w_test_0/m1_1038_n2886# VDD 1.22fF
C2388 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# 0.04fF
C2389 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0.00fF
C2390 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# VDD -0.00fF
C2391 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/c1_n930_n880# 0.11fF
C2392 a_mux4_en_0/switch_5t_1/in a_mod_grp_ctrl_1 0.00fF
C2393 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S -0.00fF
C2394 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# ota_1/p1 0.10fF
C2395 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/X -0.00fF
C2396 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_6/a_110_47# -0.00fF
C2397 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# 0.12fF
C2398 VDD a_probe_3 -4.20fF
C2399 a_mux4_en_0/in0 ota_w_test_0/m1_n1659_n11581# 0.02fF
C2400 ota_w_test_0/m1_2462_n3318# a_mux4_en_1/in1 0.01fF
C2401 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# -0.00fF
C2402 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# clock_v2_0/p1d_b 0.08fF
C2403 transmission_gate_32/out clock_v2_0/p1d 0.21fF
C2404 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B 0.00fF
C2405 ota_1/m1_n208_n2883# ota_1/m1_2462_n3318# 0.01fF
C2406 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_592_47# 0.00fF
C2407 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0.00fF
C2408 a_mux4_en_1/switch_5t_0/in a_mux4_en_1/switch_5t_0/transmission_gate_1/in -0.00fF
C2409 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# -0.00fF
C2410 clock_v2_0/Bd_b sky130_fd_sc_hd__clkinv_4_1/Y 0.00fF
C2411 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0.28fF
C2412 ota_1/sc_cmfb_0/transmission_gate_4/out VDD 1.20fF
C2413 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.09fF
C2414 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_668_97# -0.00fF
C2415 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# -0.00fF
C2416 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# VDD 0.00fF
C2417 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A 0.37fF
C2418 ota_1/p1 ota_1/m1_6690_n8907# 0.26fF
C2419 sky130_fd_sc_hd__mux4_1_0/a_750_97# d_clk_grp_2_ctrl_1 0.12fF
C2420 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0.08fF
C2421 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_1/p2_b 0.04fF
C2422 clock_v2_0/B_b transmission_gate_5/in 0.06fF
C2423 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# ota_1/p1_b 0.01fF
C2424 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0.14fF
C2425 ota_w_test_0/op ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.01fF
C2426 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_834_97# -0.01fF
C2427 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.00fF
C2428 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.03fF
C2429 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0.08fF
C2430 ota_1/p1_b clock_v2_0/A_b 1.87fF
C2431 clock_v2_0/Bd_b clock_v2_0/Bd 20.61fF
C2432 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C2433 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C2434 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y 0.00fF
C2435 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C2436 VSS ota_1/m1_11825_n9711# 0.00fF
C2437 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# VDD 0.00fF
C2438 a_mod_grp_ctrl_0 clock_v2_0/Bd 0.04fF
C2439 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0.06fF
C2440 VSS a_mux2_en_1/switch_5t_1/en 0.49fF
C2441 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.03fF
C2442 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.05fF
C2443 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n930_n880# 2.04fF
C2444 transmission_gate_19/in clock_v2_0/p2 0.33fF
C2445 VDD a_mux4_en_0/transmission_gate_3/en_b 0.77fF
C2446 ota_1/sc_cmfb_0/transmission_gate_4/out ota_1/op 0.00fF
C2447 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.00fF
C2448 a_mux4_en_0/switch_5t_3/en a_mux4_en_0/switch_5t_3/en_b -0.00fF
C2449 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/p2 0.00fF
C2450 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# 2.08fF
C2451 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0.14fF
C2452 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0.05fF
C2453 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0.08fF
C2454 ota_w_test_0/cm ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# 0.01fF
C2455 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.00fF
C2456 VDD comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A 2.33fF
C2457 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0.06fF
C2458 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C2459 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# VDD 0.14fF
C2460 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# transmission_gate_5/in 0.30fF
C2461 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0.00fF
C2462 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in ota_w_test_0/sc_cmfb_0/transmission_gate_8/in -0.07fF
C2463 clock_v2_0/B clock_v2_0/B_b 15.54fF
C2464 clock_v2_0/p1d clock_v2_0/p2_b 1.38fF
C2465 a_mux4_en_0/in1 VDD 1.47fF
C2466 ota_w_test_0/m1_2463_n5585# ota_w_test_0/m1_6690_n8907# 0.01fF
C2467 d_probe_3 VDD 2.06fF
C2468 sky130_fd_sc_hd__mux4_1_2/a_27_413# clock_v2_0/p2 -0.00fF
C2469 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0.14fF
C2470 transmission_gate_0/out transmission_gate_17/in 1.01fF
C2471 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# -0.00fF
C2472 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/p1d 0.01fF
C2473 sky130_fd_sc_hd__mux4_1_3/a_1478_413# ota_1/p1_b -0.00fF
C2474 VDD ota_w_test_0/ip 0.86fF
C2475 ota_1/p1 clock_v2_0/A 6.44fF
C2476 ota_w_test_0/sc_cmfb_0/transmission_gate_8/in ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.00fF
C2477 VSS clock_v2_0/B_b 1.98fF
C2478 ota_w_test_0/op clock_v2_0/Bd 0.08fF
C2479 a_mod_grp_ctrl_0 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0.07fF
C2480 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0.06fF
C2481 d_clk_grp_1_ctrl_1 clock_v2_0/p2_b 0.11fF
C2482 a_mux4_en_0/in1 clock_v2_0/Ad_b 0.04fF
C2483 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# -0.00fF
C2484 sky130_fd_sc_hd__mux4_1_3/a_757_363# VDD 0.08fF
C2485 transmission_gate_21/in ota_1/cm 0.03fF
C2486 a_mux4_en_1/in2 ota_w_test_0/m1_12410_n9718# 0.04fF
C2487 a_mux4_en_1/switch_5t_0/en_b a_mux4_en_1/switch_5t_1/in -0.00fF
C2488 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X -0.00fF
C2489 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# -0.35fF
C2490 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0.12fF
C2491 d_clk_grp_1_ctrl_0 clock_v2_0/A 0.01fF
C2492 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# VDD 0.06fF
C2493 clock_v2_0/Ad_b ota_w_test_0/ip 0.02fF
C2494 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0.10fF
C2495 ota_w_test_0/m1_n5574_n13620# VDD 1.18fF
C2496 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0.08fF
C2497 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# 0.04fF
C2498 clock_v2_0/Bd_b clock_v2_0/p1d 0.50fF
C2499 d_clk_grp_1_ctrl_0 sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.00fF
C2500 sky130_fd_sc_hd__mux4_1_1/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.00fF
C2501 transmission_gate_23/in ota_1/p1 0.12fF
C2502 sky130_fd_sc_hd__mux4_1_3/X d_clk_grp_1_ctrl_0 0.00fF
C2503 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C2504 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C2505 a_mod_grp_ctrl_0 clock_v2_0/p1d 0.05fF
C2506 i_bias_2 ota_1/cm 0.07fF
C2507 transmission_gate_6/in clock_v2_0/B_b 0.06fF
C2508 sky130_fd_sc_hd__mux4_1_2/X d_probe_1 0.02fF
C2509 d_probe_3 sky130_fd_sc_hd__mux4_1_0/X 0.02fF
C2510 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.06fF
C2511 VSS ota_1/m1_n2176_n12171# 0.63fF
C2512 a_mux4_en_0/in2 VDD -0.12fF
C2513 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0.00fF
C2514 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0.09fF
C2515 VSS sky130_fd_sc_hd__mux4_1_3/a_834_97# -0.05fF
C2516 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# -0.00fF
C2517 ota_1/ip clock_v2_0/p1d 0.04fF
C2518 ota_1/p2_b clock_v2_0/B_b 0.05fF
C2519 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.06fF
C2520 a_mux4_en_0/switch_5t_0/in a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C2521 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.03fF
C2522 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# 0.12fF
C2523 ota_w_test_0/m1_11063_n10490# a_mux4_en_1/in2 0.05fF
C2524 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.09fF
C2525 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# 0.12fF
C2526 a_mux2_en_1/switch_5t_1/in VDD 0.04fF
C2527 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_750_97# -0.01fF
C2528 ota_1/p1 rst_n 1.53fF
C2529 a_mux2_en_0/switch_5t_1/transmission_gate_1/in VDD 0.71fF
C2530 transmission_gate_26/en transmission_gate_32/out 0.05fF
C2531 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# 0.06fF
C2532 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# ota_1/p1_b 0.00fF
C2533 ota_w_test_0/op ota_w_test_0/sc_cmfb_0/transmission_gate_8/in 0.00fF
C2534 a_mux4_en_0/in2 clock_v2_0/Ad_b 0.03fF
C2535 a_mux4_en_1/in2 a_mux4_en_1/transmission_gate_3/en_b 0.02fF
C2536 ota_1/cm ota_1/m1_n5574_n13620# 0.01fF
C2537 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.00fF
C2538 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# ota_1/in 0.14fF
C2539 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0.05fF
C2540 ota_1/p2 clock_v2_0/B_b 0.05fF
C2541 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.03fF
C2542 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# 0.02fF
C2543 sky130_fd_sc_hd__clkinv_4_2/Y d_probe_2 1.86fF
C2544 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.01fF
C2545 sky130_fd_sc_hd__mux4_1_3/a_277_47# clock_v2_0/p2_b 0.00fF
C2546 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C2547 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B 0.92fF
C2548 a_mux4_en_0/switch_5t_2/in a_mux4_en_0/switch_5t_3/en_b -0.00fF
C2549 sky130_fd_sc_hd__mux4_1_3/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.01fF
C2550 op onebit_dac_1/out 0.05fF
C2551 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_0/en_b 0.00fF
C2552 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0.00fF
C2553 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.02fF
C2554 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A VDD 0.31fF
C2555 clock_v2_0/B transmission_gate_5/in 0.21fF
C2556 a_mux4_en_1/switch_5t_0/in a_mod_grp_ctrl_1 0.01fF
C2557 clock_v2_0/Bd_b a_mux4_en_0/in0 0.04fF
C2558 ota_w_test_0/m1_6690_n8907# a_mux4_en_0/in0 -0.10fF
C2559 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X -0.01fF
C2560 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y 1.28fF
C2561 a_mux4_en_0/switch_5t_3/en a_probe_3 -0.00fF
C2562 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A 0.41fF
C2563 clock_v2_0/Bd_b ota_w_test_0/in 0.17fF
C2564 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A -0.15fF
C2565 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.00fF
C2566 a_mux4_en_0/switch_5t_2/en a_mod_grp_ctrl_1 0.00fF
C2567 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_1/p2_b 0.00fF
C2568 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# -0.00fF
C2569 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y 0.03fF
C2570 VSS transmission_gate_5/in 1.00fF
C2571 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980# 0.71fF
C2572 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C2573 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.06fF
C2574 sky130_fd_sc_hd__clkinv_4_2/Y d_clk_grp_2_ctrl_1 0.00fF
C2575 transmission_gate_18/in transmission_gate_2/out 1.01fF
C2576 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# 0.07fF
C2577 a_mux2_en_1/switch_5t_1/en VDD 0.22fF
C2578 transmission_gate_26/en clock_v2_0/p2_b 0.05fF
C2579 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0.00fF
C2580 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0.00fF
C2581 sky130_fd_sc_hd__mux4_1_1/a_750_97# d_clk_grp_2_ctrl_1 0.15fF
C2582 a_mux4_en_1/in2 clock_v2_0/Bd 0.03fF
C2583 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0.03fF
C2584 a_mux4_en_0/in0 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.00fF
C2585 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0.14fF
C2586 clock_v2_0/p2 clock_v2_0/A_b 0.86fF
C2587 transmission_gate_18/in clock_v2_0/Bd 0.22fF
C2588 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# -0.00fF
C2589 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0.00fF
C2590 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# clock_v2_0/p1d_b 0.33fF
C2591 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_1/p2 0.00fF
C2592 sky130_fd_sc_hd__mux4_1_0/a_750_97# d_clk_grp_2_ctrl_0 0.00fF
C2593 clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C2594 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# -0.14fF
C2595 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0.05fF
C2596 rst_n transmission_gate_17/in 0.15fF
C2597 VSS sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.05fF
C2598 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_1/B 0.02fF
C2599 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.05fF
C2600 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# 0.01fF
C2601 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# 0.11fF
C2602 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# ota_1/on 0.06fF
C2603 transmission_gate_17/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# 0.11fF
C2604 transmission_gate_6/in transmission_gate_5/in 1.83fF
C2605 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980# 0.22fF
C2606 ota_w_test_0/op a_mux4_en_0/in0 -0.00fF
C2607 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# -0.00fF
C2608 VSS clock_v2_0/B 1.58fF
C2609 a_mod_grp_ctrl_0 a_mux2_en_1/switch_5t_0/in 0.02fF
C2610 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# -0.05fF
C2611 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# -0.00fF
C2612 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# 0.04fF
C2613 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# VDD 0.33fF
C2614 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0.00fF
C2615 VDD clock_v2_0/B_b 3.26fF
C2616 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C2617 ota_w_test_0/m1_2463_n5585# ota_w_test_0/m1_n208_n2883# 0.01fF
C2618 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# 0.04fF
C2619 sky130_fd_sc_hd__mux4_1_2/a_247_21# d_clk_grp_1_ctrl_0 0.09fF
C2620 clock_v2_0/Bd_b transmission_gate_26/en 0.21fF
C2621 ota_1/p2_b transmission_gate_5/in 0.31fF
C2622 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.00fF
C2623 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_668_97# -0.00fF
C2624 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/sc_cmfb_0/transmission_gate_9/in 0.00fF
C2625 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/c1_n930_n880# 0.11fF
C2626 ota_w_test_0/cm a_mux4_en_1/switch_5t_0/in 0.00fF
C2627 clock_v2_0/Ad_b clock_v2_0/B_b 0.31fF
C2628 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0.01fF
C2629 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# 0.03fF
C2630 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A VDD -0.01fF
C2631 ota_1/p1 ota_1/m1_n6302_n3889# 0.02fF
C2632 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_923_363# 0.01fF
C2633 a_mux4_en_1/in2 ota_w_test_0/sc_cmfb_0/transmission_gate_8/in -0.00fF
C2634 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/A -0.00fF
C2635 ota_1/p1 ota_1/m1_2463_n5585# 0.09fF
C2636 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210# VDD 0.01fF
C2637 a_mux4_en_1/switch_5t_3/en_b a_mux4_en_1/switch_5t_3/in 0.00fF
C2638 ota_1/cmc ota_1/p1_b 0.71fF
C2639 ota_1/p2 transmission_gate_5/in 0.61fF
C2640 ota_1/ip transmission_gate_26/en 0.32fF
C2641 transmission_gate_6/in clock_v2_0/B 0.36fF
C2642 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/sc_cmfb_0/transmission_gate_4/out -0.00fF
C2643 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# -0.29fF
C2644 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/Bd 0.00fF
C2645 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0.05fF
C2646 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# -0.00fF
C2647 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_247_21# -0.00fF
C2648 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0.03fF
C2649 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C2650 clock_v2_0/Bd ota_w_test_0/on 0.11fF
C2651 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.00fF
C2652 ota_1/p2_b sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.00fF
C2653 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0.08fF
C2654 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.11fF
C2655 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0.05fF
C2656 ota_1/m1_n2176_n12171# VDD 0.40fF
C2657 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# ota_1/p1_b 0.25fF
C2658 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# -0.12fF
C2659 sky130_fd_sc_hd__mux4_1_1/a_1478_413# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.00fF
C2660 sky130_fd_sc_hd__mux4_1_1/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00fF
C2661 VSS transmission_gate_6/in 1.37fF
C2662 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0.09fF
C2663 transmission_gate_18/in clock_v2_0/p1d 0.24fF
C2664 d_probe_0 sky130_fd_sc_hd__clkinv_4_3/Y 0.07fF
C2665 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C2666 ota_1/p2_b clock_v2_0/B 0.06fF
C2667 sky130_fd_sc_hd__mux4_1_3/a_834_97# VDD 0.01fF
C2668 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# VDD 0.00fF
C2669 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0.00fF
C2670 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# VDD 0.14fF
C2671 ota_1/p1 sky130_fd_sc_hd__mux4_1_2/a_27_47# 0.00fF
C2672 transmission_gate_8/in transmission_gate_2/out 1.52fF
C2673 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# 0.75fF
C2674 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# -0.00fF
C2675 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# VDD 0.05fF
C2676 ota_1/bias_a ota_1/m1_n1659_n11581# 0.02fF
C2677 VSS a_mux4_en_1/switch_5t_2/en 0.67fF
C2678 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C2679 VSS ota_1/p2_b 3.41fF
C2680 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0.00fF
C2681 sky130_fd_sc_hd__mux4_1_3/a_27_47# clock_v2_0/A_b 0.09fF
C2682 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01fF
C2683 VSS sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.10fF
C2684 ota_1/p2 clock_v2_0/B 0.06fF
C2685 clock_v2_0/p1d_b clock_v2_0/B_b 0.06fF
C2686 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0.06fF
C2687 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# -0.00fF
C2688 d_probe_0 sky130_fd_sc_hd__clkinv_4_4/Y 1.85fF
C2689 sky130_fd_sc_hd__mux4_1_2/a_27_47# d_clk_grp_1_ctrl_0 -0.00fF
C2690 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0.00fF
C2691 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# 0.03fF
C2692 a_mux4_en_1/transmission_gate_3/en_b a_mod_grp_ctrl_1 0.00fF
C2693 ota_1/p1 ota_1/p1_b 35.62fF
C2694 VSS a_mux4_en_1/switch_5t_1/transmission_gate_1/in 0.43fF
C2695 VSS ota_1/in 0.66fF
C2696 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0.13fF
C2697 VSS ota_1/p2 8.85fF
C2698 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0.09fF
C2699 a_mux4_en_1/switch_5t_0/transmission_gate_1/in a_mux4_en_1/switch_5t_0/en_b 0.00fF
C2700 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.00fF
C2701 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y 0.09fF
C2702 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# 0.03fF
C2703 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/c1_n260_n210# ota_1/op 0.03fF
C2704 d_clk_grp_1_ctrl_0 ota_1/p1_b 0.16fF
C2705 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A VDD 0.30fF
C2706 ota_1/p2_b transmission_gate_6/in 0.13fF
C2707 ota_w_test_0/sc_cmfb_0/transmission_gate_9/in ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.00fF
C2708 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.00fF
C2709 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# 0.00fF
C2710 a_mux4_en_0/switch_5t_2/in a_mux4_en_0/transmission_gate_3/en_b -0.00fF
C2711 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0.03fF
C2712 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/p1d 0.01fF
C2713 VDD transmission_gate_5/in 5.66fF
C2714 transmission_gate_21/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# 0.01fF
C2715 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_1/p2_b 0.00fF
C2716 a_mux4_en_0/switch_5t_0/en_b a_mux4_en_0/switch_5t_1/en 0.00fF
C2717 a_mux4_en_1/in2 a_mux4_en_0/in0 0.85fF
C2718 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0.06fF
C2719 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# -0.00fF
C2720 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# 0.08fF
C2721 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# ota_1/cm 0.08fF
C2722 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# -0.00fF
C2723 ota_w_test_0/m1_n208_n2883# ota_w_test_0/in 0.01fF
C2724 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0.05fF
C2725 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# ota_1/p2_b 0.45fF
C2726 ota_1/p2 transmission_gate_6/in 0.37fF
C2727 a_mux4_en_0/in2 a_mux4_en_0/in3 0.00fF
C2728 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0.00fF
C2729 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A -0.00fF
C2730 sky130_fd_sc_hd__mux4_1_2/a_757_363# ota_1/p1_b 0.00fF
C2731 onebit_dac_0/out onebit_dac_1/v_b 0.04fF
C2732 sky130_fd_sc_hd__mux4_1_3/X d_probe_0 0.02fF
C2733 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0.00fF
C2734 ota_w_test_0/op ota_w_test_0/sc_cmfb_0/transmission_gate_9/in -0.00fF
C2735 clock_v2_0/Bd a_mod_grp_ctrl_1 0.05fF
C2736 ota_1/p2 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# 0.05fF
C2737 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# ota_1/on 0.01fF
C2738 ota_1/in ota_1/p2_b 1.64fF
C2739 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# 0.00fF
C2740 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/A VDD 0.00fF
C2741 ota_1/p1 ota_1/m1_2462_n3318# 0.03fF
C2742 ota_1/p2 ota_1/p2_b 28.79fF
C2743 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VDD 0.08fF
C2744 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0.04fF
C2745 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_1/B 0.11fF
C2746 sky130_fd_sc_hd__mux4_1_3/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.01fF
C2747 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0.05fF
C2748 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# -0.00fF
C2749 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0.00fF
C2750 a_mux4_en_0/switch_5t_0/en_b a_mux4_en_0/switch_5t_1/in -0.00fF
C2751 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.07fF
C2752 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.08fF
C2753 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/c1_n260_n210# 0.03fF
C2754 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# 0.47fF
C2755 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# -0.00fF
C2756 VDD clock_v2_0/B 1.89fF
C2757 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VDD 0.10fF
C2758 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0.13fF
C2759 sky130_fd_sc_hd__mux4_1_1/a_750_97# d_clk_grp_2_ctrl_0 0.01fF
C2760 ota_w_test_0/cm a_mux4_en_1/transmission_gate_3/en_b 0.02fF
C2761 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0.00fF
C2762 ota_1/ip transmission_gate_21/in 0.03fF
C2763 ota_1/p2 ota_1/in 0.53fF
C2764 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/c1_n260_n210# ota_1/op 0.06fF
C2765 transmission_gate_17/in ota_1/p1_b 0.17fF
C2766 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.01fF
C2767 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# -0.00fF
C2768 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_2/en_b 0.00fF
C2769 VSS a_mux4_en_1/switch_5t_2/transmission_gate_1/in 0.45fF
C2770 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C2771 VSS VDD 316.81fF
C2772 VSS sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.01fF
C2773 a_mod_grp_ctrl_0 i_bias_2 0.18fF
C2774 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# VDD 0.16fF
C2775 a_mux4_en_0/in1 clock_v2_0/Ad 0.04fF
C2776 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0.25fF
C2777 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# VDD 0.00fF
C2778 transmission_gate_17/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# 0.11fF
C2779 clock_v2_0/Ad_b clock_v2_0/B 0.06fF
C2780 a_mux4_en_0/in0 ota_w_test_0/m1_n2176_n12171# -0.03fF
C2781 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.05fF
C2782 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# 0.01fF
C2783 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y a_mod_grp_ctrl_1 0.05fF
C2784 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.00fF
C2785 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# VDD 0.08fF
C2786 clock_v2_0/Ad ota_w_test_0/ip 0.02fF
C2787 a_mux4_en_0/switch_5t_2/in a_mux4_en_0/in2 0.00fF
C2788 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# VDD -0.00fF
C2789 ota_1/ip i_bias_2 0.01fF
C2790 transmission_gate_18/in transmission_gate_26/en 0.07fF
C2791 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C2792 a_mux4_en_0/in0 ota_w_test_0/on 0.01fF
C2793 transmission_gate_19/out transmission_gate_32/out 0.15fF
C2794 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1017_47# -0.00fF
C2795 VSS transmission_gate_31/out 1.14fF
C2796 VSS clock_v2_0/Ad_b 3.27fF
C2797 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0.09fF
C2798 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# -0.00fF
C2799 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0.03fF
C2800 debug clock_v2_0/A 0.07fF
C2801 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/p1_b 0.06fF
C2802 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# 0.32fF
C2803 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.06fF
C2804 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# -0.00fF
C2805 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_1/p1_b 0.04fF
C2806 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C2807 sky130_fd_sc_hd__mux4_1_0/X sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.03fF
C2808 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.12fF
C2809 VSS ota_1/op 8.36fF
C2810 a_mux4_en_1/switch_5t_0/en a_mux4_en_1/switch_5t_0/in -0.00fF
C2811 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# clock_v2_0/p1d 0.25fF
C2812 a_mux2_en_1/switch_5t_0/transmission_gate_1/in a_mux2_en_1/switch_5t_1/en -0.00fF
C2813 VDD transmission_gate_6/in 6.52fF
C2814 ota_1/cm ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# 0.08fF
C2815 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X VDD 0.00fF
C2816 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# -0.00fF
C2817 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/c1_n260_n210# -0.14fF
C2818 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/B_b 0.10fF
C2819 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# VDD 0.00fF
C2820 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0.00fF
C2821 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# -0.10fF
C2822 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.03fF
C2823 clock_v2_0/p1d a_mod_grp_ctrl_1 0.06fF
C2824 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_1/X 0.02fF
C2825 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# VDD 0.15fF
C2826 ota_1/ip ota_1/m1_n5574_n13620# 0.00fF
C2827 ota_w_test_0/cm clock_v2_0/Bd 0.11fF
C2828 VSS clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0.92fF
C2829 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A 0.00fF
C2830 VDD a_mux4_en_1/switch_5t_2/en -0.36fF
C2831 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/c1_n260_n210# 0.03fF
C2832 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# 0.00fF
C2833 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__clkinv_4_3/Y 0.19fF
C2834 ota_1/p2_b VDD 7.69fF
C2835 VSS sky130_fd_sc_hd__mux4_1_0/X 0.57fF
C2836 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0.00fF
C2837 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# 0.17fF
C2838 clock_v2_0/p1d_b clock_v2_0/B 0.07fF
C2839 clock_v2_0/Ad a_mux4_en_0/in2 0.04fF
C2840 sky130_fd_sc_hd__mux4_1_2/a_1478_413# clock_v2_0/B_b -0.00fF
C2841 sky130_fd_sc_hd__mux4_1_1/a_1478_413# VDD 0.19fF
C2842 transmission_gate_9/in transmission_gate_2/out -0.55fF
C2843 onebit_dac_0/out clock_v2_0/p2 0.25fF
C2844 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# VDD -0.00fF
C2845 sky130_fd_sc_hd__mux4_1_1/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.01fF
C2846 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# ota_1/p1_b 0.01fF
C2847 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.10fF
C2848 VSS clock_v2_0/p1d_b 2.54fF
C2849 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# 0.03fF
C2850 a_mux4_en_1/switch_5t_1/transmission_gate_1/in VDD -0.19fF
C2851 ota_1/in VDD 2.28fF
C2852 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_1/en_b 0.00fF
C2853 ota_1/p2 VDD 9.56fF
C2854 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_1/a_1290_413# 0.02fF
C2855 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/a_277_47# 0.02fF
C2856 transmission_gate_31/out ota_1/p2_b 0.68fF
C2857 ota_1/p2_b clock_v2_0/Ad_b 0.72fF
C2858 sky130_fd_sc_hd__mux4_1_3/a_27_413# clock_v2_0/B 0.00fF
C2859 transmission_gate_32/out onebit_dac_1/out 0.04fF
C2860 transmission_gate_19/out clock_v2_0/p2_b 0.06fF
C2861 ota_w_test_0/m1_2463_n5585# ota_w_test_0/cm 0.00fF
C2862 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980# transmission_gate_6/in 0.30fF
C2863 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.00fF
C2864 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.03fF
C2865 sky130_fd_sc_hd__mux4_1_1/a_1478_413# clock_v2_0/Ad_b -0.00fF
C2866 VSS a_mux4_en_0/switch_5t_0/in 0.03fF
C2867 ota_1/p2_b ota_1/op 0.49fF
C2868 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0.10fF
C2869 ota_1/m1_n947_n12836# ota_1/p1 0.05fF
C2870 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_834_97# -0.01fF
C2871 VSS sky130_fd_sc_hd__mux4_1_3/a_27_413# 0.01fF
C2872 ota_1/p1 clock_v2_0/p2 1.36fF
C2873 sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# transmission_gate_5/in 0.18fF
C2874 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0.14fF
C2875 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/c1_n930_n880# 0.11fF
C2876 VSS ota_1/m1_11534_n9706# 0.00fF
C2877 transmission_gate_31/out ota_1/in 0.37fF
C2878 a_mux4_en_1/switch_5t_0/en_b a_mod_grp_ctrl_1 0.26fF
C2879 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0.00fF
C2880 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# -0.00fF
C2881 transmission_gate_31/out ota_1/p2 0.19fF
C2882 ota_1/p2 clock_v2_0/Ad_b 1.18fF
C2883 sky130_fd_sc_hd__mux4_1_3/a_750_97# clock_v2_0/A_b 0.03fF
C2884 transmission_gate_19/out sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# 0.04fF
C2885 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out ota_w_test_0/sc_cmfb_0/transmission_gate_9/in 0.03fF
C2886 ota_1/in ota_1/op 1.60fF
C2887 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.02fF
C2888 ota_1/p2 ota_1/op 0.62fF
C2889 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C2890 d_clk_grp_1_ctrl_0 clock_v2_0/p2 0.00fF
C2891 a_probe_0 a_mux2_en_0/switch_5t_1/transmission_gate_1/in 0.00fF
C2892 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# 0.73fF
C2893 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# -0.25fF
C2894 sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# -0.35fF
C2895 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# -0.00fF
C2896 sky130_fd_sc_hd__mux4_1_2/a_834_97# clock_v2_0/B_b -0.01fF
C2897 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.06fF
C2898 a_mux4_en_1/switch_5t_1/en_b a_mux4_en_1/switch_5t_1/en 0.00fF
C2899 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# 0.03fF
C2900 transmission_gate_19/in clock_v2_0/p1d 0.10fF
C2901 ota_1/p2_b clock_v2_0/p1d_b 1.49fF
C2902 sky130_fd_sc_hd__mux4_1_0/X ota_1/p2 0.01fF
C2903 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# -0.09fF
C2904 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__clkinv_4_4/Y 0.32fF
C2905 sky130_fd_sc_hd__mux4_1_1/a_1478_413# clock_v2_0/p1d_b -0.00fF
C2906 a_mux2_en_0/switch_5t_1/in debug 0.02fF
C2907 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_3/en_b -0.00fF
C2908 onebit_dac_1/out clock_v2_0/p2_b 0.44fF
C2909 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0.08fF
C2910 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0.05fF
C2911 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.07fF
C2912 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/c1_n260_n210# 0.03fF
C2913 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/sc_cmfb_0/transmission_gate_4/out -0.00fF
C2914 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# VDD 0.09fF
C2915 a_mux4_en_0/in1 ota_w_test_0/m1_n1659_n11581# 0.83fF
C2916 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C2917 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n930_n880# 0.11fF
C2918 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C2919 ota_1/p2 clock_v2_0/p1d_b 2.70fF
C2920 ota_1/ip transmission_gate_19/out 0.05fF
C2921 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C2922 ota_1/m1_1038_n2886# ota_1/m1_2463_n5585# 0.01fF
C2923 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# ota_1/in 0.22fF
C2924 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# 0.21fF
C2925 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C2926 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_757_363# 0.00fF
C2927 VDD a_mux4_en_1/switch_5t_2/transmission_gate_1/in -0.08fF
C2928 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.00fF
C2929 sky130_fd_sc_hd__mux4_1_2/a_193_413# VDD 0.02fF
C2930 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C2931 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.06fF
C2932 onebit_dac_1/v_b comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X 0.00fF
C2933 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# VDD -0.00fF
C2934 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# transmission_gate_5/in 0.22fF
C2935 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/c1_n260_n210# 0.03fF
C2936 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.03fF
C2937 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/c1_n930_n880# 0.11fF
C2938 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0.00fF
C2939 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/c1_n260_n210# ota_1/op 0.03fF
C2940 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# VDD 0.59fF
C2941 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0.06fF
C2942 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0.07fF
C2943 sky130_fd_sc_hd__mux4_1_2/a_834_97# sky130_fd_sc_hd__mux4_1_3/a_834_97# 0.01fF
C2944 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# clock_v2_0/p1d 0.15fF
C2945 VSS sky130_fd_sc_hd__mux4_1_3/a_923_363# -0.11fF
C2946 clock_v2_0/Ad clock_v2_0/B_b 0.44fF
C2947 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# 0.80fF
C2948 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# -0.00fF
C2949 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0.00fF
C2950 VSS a_mux4_en_0/switch_5t_3/en 0.29fF
C2951 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/c1_n530_n480# -0.24fF
C2952 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0.24fF
C2953 transmission_gate_31/out VDD 1.62fF
C2954 clock_v2_0/Ad_b VDD 5.15fF
C2955 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0.02fF
C2956 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# VDD 0.78fF
C2957 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# ota_1/in 0.04fF
C2958 VDD ota_1/op 8.30fF
C2959 ota_1/p1 sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.01fF
C2960 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y a_mod_grp_ctrl_0 0.06fF
C2961 ota_w_test_0/cm a_mux4_en_0/in0 0.10fF
C2962 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# -0.00fF
C2963 ota_w_test_0/cm ota_w_test_0/in 1.16fF
C2964 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0.00fF
C2965 a_mux4_en_0/in2 ota_w_test_0/m1_n1659_n11581# 0.19fF
C2966 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0.08fF
C2967 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# VDD 0.52fF
C2968 ota_1/m1_1038_n2886# ota_1/p1_b 0.06fF
C2969 a_mod_grp_ctrl_0 a_mux4_en_1/switch_5t_2/in 0.02fF
C2970 VDD clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 2.79fF
C2971 VSS sky130_fd_sc_hd__mux4_1_2/a_277_47# -0.64fF
C2972 clock_v2_0/Bd clock_v2_0/A_b 0.49fF
C2973 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A -0.01fF
C2974 sky130_fd_sc_hd__mux4_1_0/X VDD 0.60fF
C2975 sky130_fd_sc_hd__mux4_1_3/a_27_47# d_clk_grp_1_ctrl_0 0.02fF
C2976 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C2977 transmission_gate_31/out ota_1/op 0.09fF
C2978 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.03fF
C2979 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# 0.71fF
C2980 rst_n clock_v2_0/A 0.42fF
C2981 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/X -0.00fF
C2982 i_bias_2 ota_1/bias_c 0.07fF
C2983 sky130_fd_sc_hd__mux4_1_2/a_1478_413# VSS 0.16fF
C2984 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0.10fF
C2985 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_1/p2_b 0.06fF
C2986 clock_v2_0/p1d_b VDD 6.09fF
C2987 clock_v2_0/Ad_b clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C2988 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.03fF
C2989 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/c1_n260_n210# ota_1/op 0.03fF
C2990 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0.05fF
C2991 VSS a_mux4_en_0/in3 -0.21fF
C2992 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47# -0.00fF
C2993 VSS a_mux2_en_1/switch_5t_0/transmission_gate_1/in -0.44fF
C2994 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0.15fF
C2995 a_mux4_en_1/switch_5t_3/en_b debug 0.00fF
C2996 VSS sky130_fd_sc_hd__mux4_1_0/a_668_97# -0.23fF
C2997 op VSS 2.16fF
C2998 VDD a_mux4_en_0/switch_5t_0/in 0.43fF
C2999 VSS sky130_fd_sc_hd__mux4_1_3/a_1290_413# -0.01fF
C3000 sky130_fd_sc_hd__mux4_1_3/a_668_97# clock_v2_0/B_b 0.00fF
C3001 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# 0.11fF
C3002 sky130_fd_sc_hd__mux4_1_3/a_277_47# sky130_fd_sc_hd__mux4_1_2/a_27_413# 0.00fF
C3003 a_mux4_en_1/in1 a_mux4_en_1/transmission_gate_3/en_b 0.02fF
C3004 sky130_fd_sc_hd__mux4_1_3/a_27_413# VDD 0.11fF
C3005 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.00fF
C3006 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_1/p2 0.04fF
C3007 VSS ota_1/on 17.81fF
C3008 transmission_gate_31/out clock_v2_0/p1d_b 0.79fF
C3009 clock_v2_0/Ad_b clock_v2_0/p1d_b 1.74fF
C3010 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# ota_1/p1_b 0.09fF
C3011 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y -0.00fF
C3012 VSS ota_1/sc_cmfb_0/transmission_gate_8/in 0.69fF
C3013 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.03fF
C3014 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0.10fF
C3015 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# 0.00fF
C3016 VSS sky130_fd_sc_hd__mux4_1_1/a_757_363# -0.02fF
C3017 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# VDD 0.07fF
C3018 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# ota_1/p1_b 0.04fF
C3019 transmission_gate_26/en ota_w_test_0/cm 0.02fF
C3020 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/X -0.00fF
C3021 ota_1/p1_b debug 0.08fF
C3022 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.05fF
C3023 sky130_fd_sc_hd__mux4_1_1/a_27_47# sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.00fF
C3024 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# ota_1/p1_b 0.06fF
C3025 a_mux2_en_0/switch_5t_1/transmission_gate_1/in a_mux2_en_0/switch_5t_1/en 0.00fF
C3026 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VSS 0.00fF
C3027 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# -0.00fF
C3028 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0.00fF
C3029 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# 0.09fF
C3030 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# -0.00fF
C3031 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# 0.27fF
C3032 clock_v2_0/p1d clock_v2_0/A_b 0.05fF
C3033 VSS sky130_fd_sc_hd__mux4_1_2/a_834_97# -0.06fF
C3034 ip transmission_gate_0/out 0.01fF
C3035 VSS a_mux4_en_0/switch_5t_2/in 0.05fF
C3036 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0.00fF
C3037 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# 0.09fF
C3038 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0.00fF
C3039 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.00fF
C3040 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X -0.01fF
C3041 sky130_fd_sc_hd__mux4_1_3/a_757_363# clock_v2_0/p2_b 0.00fF
C3042 clock_v2_0/Bd a_mux4_en_1/in1 0.04fF
C3043 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 0.54fF
C3044 clock_v2_0/Bd i_bias_1 0.11fF
C3045 ota_1/p2_b ota_1/on 0.32fF
C3046 d_clk_grp_1_ctrl_1 clock_v2_0/A_b 0.05fF
C3047 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.07fF
C3048 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# -0.12fF
C3049 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_0/a_113_47# a_mux4_en_1/switch_5t_3/en_b -0.00fF
C3050 a_mod_grp_ctrl_0 a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C3051 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/p2_b -0.00fF
C3052 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# 0.12fF
C3053 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0.25fF
C3054 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0.08fF
C3055 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# -0.00fF
C3056 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y 0.72fF
C3057 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C3058 clock_v2_0/Bd_b a_mux4_en_0/in1 0.04fF
C3059 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# ota_1/p1_b 0.25fF
C3060 a_mux4_en_0/in1 ota_w_test_0/m1_6690_n8907# 0.01fF
C3061 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0.05fF
C3062 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# 0.22fF
C3063 clock_v2_0/Ad clock_v2_0/B 0.06fF
C3064 ota_1/in ota_1/on 0.15fF
C3065 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# 0.11fF
C3066 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0.00fF
C3067 ota_1/p2 ota_1/on 0.37fF
C3068 transmission_gate_0/out sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/c1_n930_n880# 0.03fF
C3069 a_mod_grp_ctrl_1 a_mux4_en_1/switch_5t_2/en_b 0.08fF
C3070 sky130_fd_sc_hd__mux4_1_3/a_923_363# VDD -0.01fF
C3071 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0.00fF
C3072 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A -0.01fF
C3073 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/p2 0.00fF
C3074 a_mux4_en_0/switch_5t_3/en VDD -0.69fF
C3075 clock_v2_0/Bd_b ota_w_test_0/ip 0.77fF
C3076 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# -0.13fF
C3077 sky130_fd_sc_hd__mux4_1_1/a_757_363# ota_1/p2 0.00fF
C3078 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210# 0.03fF
C3079 sky130_fd_sc_hd__clkinv_4_2/Y sky130_fd_sc_hd__mux4_1_1/a_750_97# 0.02fF
C3080 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_1/p2_b 0.01fF
C3081 VSS clock_v2_0/Ad 2.10fF
C3082 ota_1/m1_6690_n8907# ota_1/p1_b 0.02fF
C3083 ota_w_test_0/m1_2463_n5585# a_mux4_en_1/in1 0.01fF
C3084 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C3085 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0.06fF
C3086 VSS sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# 0.28fF
C3087 sky130_fd_sc_hd__mux4_1_0/a_193_413# clock_v2_0/p1d 0.00fF
C3088 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0.00fF
C3089 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A -0.01fF
C3090 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# 0.13fF
C3091 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# -0.00fF
C3092 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0.00fF
C3093 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0.04fF
C3094 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0.00fF
C3095 a_mux4_en_0/in0 clock_v2_0/A_b 0.03fF
C3096 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# -0.00fF
C3097 sky130_fd_sc_hd__clkinv_4_4/Y ota_1/p1_b 0.00fF
C3098 a_mux4_en_1/switch_5t_0/en a_mux4_en_1/switch_5t_0/en_b -0.00fF
C3099 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/c1_n260_n210# 0.03fF
C3100 ota_1/p2 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# 0.05fF
C3101 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X VDD 0.00fF
C3102 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.00fF
C3103 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/c1_n260_n210# 0.02fF
C3104 clock_v2_0/A_b ota_w_test_0/in 0.06fF
C3105 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# ota_1/p1_b -0.06fF
C3106 sky130_fd_sc_hd__mux4_1_2/a_277_47# VDD 0.12fF
C3107 ota_1/p1_b comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A -0.04fF
C3108 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# -0.00fF
C3109 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0.08fF
C3110 ota_w_test_0/sc_cmfb_0/transmission_gate_8/in a_mux4_en_1/in1 0.00fF
C3111 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_923_363# 0.00fF
C3112 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# transmission_gate_23/in 0.01fF
C3113 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# -0.26fF
C3114 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980# -0.38fF
C3115 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# VDD 0.00fF
C3116 a_mux4_en_1/in2 a_mux4_en_1/switch_5t_2/in -0.00fF
C3117 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# ota_1/ip 0.15fF
C3118 ota_w_test_0/op a_mux4_en_0/in1 0.93fF
C3119 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/A 0.00fF
C3120 VSS a_probe_0 1.41fF
C3121 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# clock_v2_0/p2 0.03fF
C3122 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n930_n880# transmission_gate_17/in 0.11fF
C3123 clock_v2_0/Bd_b a_mux4_en_0/in2 0.04fF
C3124 clock_v2_0/p1d_b sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 0.33fF
C3125 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# VSS 0.39fF
C3126 a_mux4_en_0/switch_5t_1/en_b a_mux4_en_0/switch_5t_1/transmission_gate_1/in 0.00fF
C3127 VSS ota_1/cm 3.14fF
C3128 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/c1_n260_n210# -0.12fF
C3129 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.00fF
C3130 sky130_fd_sc_hd__mux4_1_3/a_277_47# clock_v2_0/A_b 0.11fF
C3131 sky130_fd_sc_hd__mux4_1_2/a_1478_413# VDD 0.14fF
C3132 sky130_fd_sc_hd__mux4_1_1/a_834_97# sky130_fd_sc_hd__clkinv_4_2/Y 0.00fF
C3133 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# VDD -0.00fF
C3134 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0.00fF
C3135 clock_v2_0/Ad ota_1/p2_b 0.57fF
C3136 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# -0.13fF
C3137 sky130_fd_sc_hd__mux4_1_1/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.01fF
C3138 VDD a_mux4_en_0/in3 -0.63fF
C3139 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0.00fF
C3140 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0.00fF
C3141 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47# VDD -0.00fF
C3142 a_mux2_en_1/switch_5t_0/transmission_gate_1/in VDD 0.20fF
C3143 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0.00fF
C3144 ota_1/m1_6690_n8907# ota_1/m1_2462_n3318# -0.00fF
C3145 VSS sky130_fd_sc_hd__mux4_1_1/a_247_21# 0.06fF
C3146 sky130_fd_sc_hd__mux4_1_0/a_668_97# VDD 0.00fF
C3147 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# 0.14fF
C3148 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# -0.00fF
C3149 ota_1/p1_b clock_v2_0/A 6.73fF
C3150 op VDD 2.54fF
C3151 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/c1_n930_n880# 0.11fF
C3152 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# -0.15fF
C3153 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VDD 0.00fF
C3154 a_mux2_en_1/switch_5t_1/in a_mod_grp_ctrl_0 0.02fF
C3155 sky130_fd_sc_hd__mux4_1_3/a_1290_413# VDD 0.10fF
C3156 a_mux4_en_0/switch_5t_1/en_b a_mod_grp_ctrl_1 0.00fF
C3157 a_mod_grp_ctrl_0 a_mux2_en_0/switch_5t_1/transmission_gate_1/in 0.00fF
C3158 VDD ota_1/on 5.12fF
C3159 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# -0.00fF
C3160 sky130_fd_sc_hd__mux4_1_3/a_750_97# d_clk_grp_1_ctrl_0 0.01fF
C3161 VSS sky130_fd_sc_hd__mux4_1_3/a_668_97# -0.31fF
C3162 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_1/a_668_97# 0.01fF
C3163 ota_1/sc_cmfb_0/transmission_gate_8/in VDD 0.90fF
C3164 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y 0.02fF
C3165 sky130_fd_sc_hd__mux4_1_2/a_750_97# ota_1/p1_b 0.00fF
C3166 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# -0.16fF
C3167 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0.00fF
C3168 sky130_fd_sc_hd__mux4_1_3/X ota_1/p1_b 0.01fF
C3169 sky130_fd_sc_hd__mux4_1_1/a_757_363# VDD 0.08fF
C3170 ota_w_test_0/m1_1038_n2886# ota_w_test_0/m1_n208_n2883# 0.00fF
C3171 clock_v2_0/Ad ota_1/p2 0.74fF
C3172 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.00fF
C3173 ota_1/p1 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/c1_n530_n480# 0.17fF
C3174 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.06fF
C3175 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0.00fF
C3176 transmission_gate_26/en clock_v2_0/A_b 0.11fF
C3177 sky130_fd_sc_hd__mux4_1_0/a_668_97# clock_v2_0/Ad_b 0.00fF
C3178 comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# onebit_dac_1/v_b 0.00fF
C3179 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/c1_n260_n210# ota_1/on 0.03fF
C3180 ota_1/p1_b comparator_v2_0/li_940_3458# 0.00fF
C3181 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# VDD 0.30fF
C3182 ota_w_test_0/op a_mux4_en_0/in2 0.10fF
C3183 transmission_gate_23/in ota_1/p1_b 0.07fF
C3184 sky130_fd_sc_hd__mux4_1_3/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C3185 ota_1/p2_b ota_1/cm 0.28fF
C3186 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C3187 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# VDD -0.00fF
C3188 ota_w_test_0/op ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0.00fF
C3189 sky130_fd_sc_hd__mux4_1_1/a_757_363# clock_v2_0/Ad_b 0.01fF
C3190 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# VDD 0.02fF
C3191 ota_1/op ota_1/on 1.81fF
C3192 debug clock_v2_0/p2 0.06fF
C3193 sky130_fd_sc_hd__mux4_1_2/a_834_97# VDD 0.01fF
C3194 a_mux4_en_0/switch_5t_3/en_b a_mux4_en_0/switch_5t_3/in 0.00fF
C3195 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/op -0.00fF
C3196 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# clock_v2_0/p2_b 0.02fF
C3197 clock_v2_0/p2_b clock_v2_0/B_b 1.39fF
C3198 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# VDD -0.00fF
C3199 d_clk_grp_2_ctrl_1 sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C3200 VSS comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X -0.00fF
C3201 a_mux4_en_0/switch_5t_2/in VDD 0.28fF
C3202 a_mux4_en_0/in0 a_mux4_en_1/in1 2.09fF
C3203 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.00fF
C3204 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# 0.93fF
C3205 ota_1/in ota_1/cm 0.76fF
C3206 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# ota_1/p1_b 0.25fF
C3207 sky130_fd_sc_hd__mux4_1_3/a_27_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C3208 ota_1/p2 ota_1/cm 0.68fF
C3209 clock_v2_0/Bd sky130_fd_sc_hd__mux4_1_0/a_27_47# -0.00fF
C3210 rst_n ota_1/p1_b 0.73fF
C3211 onebit_dac_0/out transmission_gate_2/out 0.04fF
C3212 i_bias_1 ota_w_test_0/in 0.10fF
C3213 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0.09fF
C3214 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/c1_n930_n880# 0.11fF
C3215 a_mod_grp_ctrl_0 a_mux2_en_1/switch_5t_1/en 1.03fF
C3216 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0.23fF
C3217 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0.00fF
C3218 a_mux4_en_0/switch_5t_3/en_b a_mod_grp_ctrl_1 0.00fF
C3219 ota_1/m1_n947_n12836# ota_1/bias_d 0.03fF
C3220 sky130_fd_sc_hd__mux4_1_2/X d_clk_grp_1_ctrl_0 0.00fF
C3221 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0.30fF
C3222 sky130_fd_sc_hd__clkinv_4_1/Y d_probe_2 0.07fF
C3223 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C3224 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# ota_1/p1_b 0.04fF
C3225 VSS a_mux2_en_0/transmission_gate_1/en_b 0.01fF
C3226 clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A -0.00fF
C3227 debug a_mux4_en_0/switch_5t_1/in -0.01fF
C3228 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# 0.04fF
C3229 VSS ota_w_test_0/m1_n1659_n11581# 0.57fF
C3230 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# -0.00fF
C3231 sky130_fd_sc_hd__mux4_1_1/a_757_363# clock_v2_0/p1d_b 0.08fF
C3232 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0.09fF
C3233 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0.07fF
C3234 clock_v2_0/Bd_b clock_v2_0/B_b 3.32fF
C3235 transmission_gate_0/out clock_v2_0/p2 0.18fF
C3236 a_mux4_en_0/in1 a_mux4_en_1/in2 1.34fF
C3237 a_mux4_en_0/in1 ota_w_test_0/m1_n208_n2883# 0.01fF
C3238 i_bias_2 ota_1/m1_n208_n2883# -0.02fF
C3239 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.06fF
C3240 clock_v2_0/Ad VDD 18.79fF
C3241 sky130_fd_sc_hd__mux4_1_0/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0.01fF
C3242 ota_1/p1 clock_v2_0/Bd 0.69fF
C3243 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_2/X 0.00fF
C3244 VSS a_mux4_en_1/switch_5t_3/en 0.29fF
C3245 sky130_fd_sc_hd__mux4_1_3/a_834_97# clock_v2_0/p2_b 0.00fF
C3246 a_mod_grp_ctrl_0 clock_v2_0/B_b 0.05fF
C3247 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# 0.22fF
C3248 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0.08fF
C3249 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0.00fF
C3250 sky130_fd_sc_hd__clkinv_4_1/Y d_clk_grp_2_ctrl_1 0.00fF
C3251 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# ota_1/p1 0.23fF
C3252 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0.00fF
C3253 sky130_fd_sc_hd__mux4_1_3/a_193_47# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.01fF
C3254 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# 0.03fF
C3255 VSS a_mux4_en_1/in3 -0.21fF
C3256 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# 1.05fF
C3257 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980# transmission_gate_5/in 0.22fF
C3258 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0.08fF
C3259 comparator_v2_0/li_940_818# comparator_v2_0/li_940_3458# 0.00fF
C3260 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0.11fF
C3261 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/c1_n260_n210# -0.09fF
C3262 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.43fF
C3263 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_2/a_247_21# -0.00fF
C3264 VSS sky130_fd_sc_hd__mux4_1_0/a_193_47# -0.00fF
C3265 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0.12fF
C3266 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0.07fF
C3267 clock_v2_0/Ad clock_v2_0/Ad_b 19.81fF
C3268 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_2/a_923_363# 0.00fF
C3269 ota_1/sc_cmfb_0/transmission_gate_4/out ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# -0.02fF
C3270 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y a_mod_grp_ctrl_1 0.00fF
C3271 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C3272 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0.07fF
C3273 clock_v2_0/Bd d_clk_grp_2_ctrl_1 0.00fF
C3274 VSS ota_1/sc_cmfb_0/transmission_gate_3/out 0.43fF
C3275 a_probe_0 VDD 2.28fF
C3276 VSS a_mux2_en_0/switch_5t_1/en 0.65fF
C3277 a_mux4_en_1/in2 ota_w_test_0/m1_n5574_n13620# 0.00fF
C3278 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0.00fF
C3279 a_mod_grp_ctrl_1 a_mux4_en_1/switch_5t_2/in 0.01fF
C3280 sky130_fd_sc_hd__mux4_1_0/a_27_47# clock_v2_0/p1d 0.00fF
C3281 ota_1/cm VDD 3.37fF
C3282 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# clock_v2_0/p2 0.03fF
C3283 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0.06fF
C3284 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A -0.00fF
C3285 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0.00fF
C3286 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# -0.00fF
C3287 ota_w_test_0/op clock_v2_0/B_b 0.05fF
C3288 transmission_gate_19/out transmission_gate_19/in 0.00fF
C3289 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0.00fF
C3290 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_439_47# -0.00fF
C3291 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0.01fF
C3292 a_mux4_en_1/in2 a_mux4_en_0/in2 0.66fF
C3293 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.28fF
C3294 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/c1_n530_n480# 0.06fF
C3295 a_mux4_en_0/in1 ota_w_test_0/m1_n2176_n12171# 1.38fF
C3296 sky130_fd_sc_hd__mux4_1_1/a_247_21# VDD 0.07fF
C3297 VSS ota_1/m1_11242_n9716# 0.00fF
C3298 VSS transmission_gate_32/out 0.79fF
C3299 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# 0.31fF
C3300 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_193_413# 0.00fF
C3301 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# ota_1/sc_cmfb_0/transmission_gate_4/out -0.00fF
C3302 a_mux4_en_0/in1 ota_w_test_0/on 0.93fF
C3303 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y 0.02fF
C3304 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980# 0.75fF
C3305 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0.05fF
C3306 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47# -0.00fF
C3307 sky130_fd_sc_hd__mux4_1_3/a_668_97# VDD 0.01fF
C3308 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0.00fF
C3309 ota_1/cm ota_1/op 0.01fF
C3310 clock_v2_0/Ad clock_v2_0/p1d_b 6.17fF
C3311 a_mux4_en_0/switch_5t_1/transmission_gate_1/in a_probe_3 0.00fF
C3312 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_15/a_110_47# VDD 0.13fF
C3313 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_11/a_110_47# 0.00fF
C3314 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A -0.01fF
C3315 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# clock_v2_0/p1d_b 0.02fF
C3316 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/c1_n260_n210# 0.03fF
C3317 ota_1/p1 clock_v2_0/p1d 1.61fF
C3318 ota_1/p1 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# -0.00fF
C3319 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980# 0.29fF
C3320 clock_v2_0/Bd transmission_gate_17/in 1.49fF
C3321 clock_v2_0/A clock_v2_0/p2 0.68fF
C3322 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0.18fF
C3323 sky130_fd_sc_hd__mux4_1_1/a_247_21# clock_v2_0/Ad_b 0.06fF
C3324 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X -0.01fF
C3325 ota_1/m1_n6302_n3889# ota_1/p1_b 0.02fF
C3326 ota_1/m1_2463_n5585# ota_1/p1_b 0.09fF
C3327 VSS a_mux4_en_1/switch_5t_1/in 0.03fF
C3328 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.00fF
C3329 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# VSS 0.33fF
C3330 d_clk_grp_1_ctrl_1 ota_1/p1 0.00fF
C3331 transmission_gate_9/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/c1_n930_n880# 0.03fF
C3332 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0.35fF
C3333 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.01fF
C3334 clock_v2_0/p2_b clock_v2_0/B 4.34fF
C3335 d_clk_grp_2_ctrl_1 clock_v2_0/p1d 0.00fF
C3336 VSS clock_v2_0/sky130_fd_sc_hd__mux2_1_0/X 0.15fF
C3337 VDD comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X 0.00fF
C3338 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0.07fF
C3339 sky130_fd_sc_hd__mux4_1_3/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_277_47# 0.01fF
C3340 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/c1_n530_n480# VDD 0.00fF
C3341 ota_1/p2_b transmission_gate_32/out 0.49fF
C3342 a_mux4_en_0/in2 ota_w_test_0/m1_n2176_n12171# 0.04fF
C3343 ota_1/bias_a ota_1/m1_n2176_n12171# 0.01fF
C3344 transmission_gate_21/in sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/c1_n260_n210# 0.00fF
C3345 VSS clock_v2_0/p2_b 3.20fF
C3346 d_clk_grp_1_ctrl_1 d_clk_grp_1_ctrl_0 1.84fF
C3347 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# transmission_gate_32/out 0.03fF
C3348 a_mux4_en_0/in2 ota_w_test_0/on 0.05fF
C3349 VSS a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.06fF
C3350 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A VDD 0.24fF
C3351 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0.05fF
C3352 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_1/bias_a 0.02fF
C3353 VSS sky130_fd_sc_hd__mux4_1_1/a_277_47# -0.65fF
C3354 d_clk_grp_1_ctrl_1 d_clk_grp_2_ctrl_1 0.00fF
C3355 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# 0.02fF
C3356 VSS ota_w_test_0/sc_cmfb_0/transmission_gate_6/in -0.54fF
C3357 sky130_fd_sc_hd__mux4_1_2/a_1478_413# sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0.00fF
C3358 sky130_fd_sc_hd__mux4_1_1/a_247_21# clock_v2_0/p1d_b 0.06fF
C3359 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0.05fF
C3360 ota_1/in transmission_gate_32/out 0.03fF
C3361 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.01fF
C3362 ota_1/p2 transmission_gate_32/out 0.45fF
C3363 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.08fF
C3364 a_mux2_en_0/transmission_gate_1/en_b VDD 0.54fF
C3365 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/c1_n530_n480# -0.13fF
C3366 rst_n clock_v2_0/p2 0.06fF
C3367 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.06fF
C3368 ota_w_test_0/m1_n1659_n11581# VDD 0.02fF
C3369 a_mux4_en_0/transmission_gate_3/en_b a_mod_grp_ctrl_1 0.00fF
C3370 transmission_gate_18/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/c1_n930_n880# 0.11fF
C3371 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# -0.00fF
C3372 d_clk_grp_2_ctrl_0 sky130_fd_sc_hd__mux4_1_0/a_1478_413# -0.00fF
C3373 clock_v2_0/Bd_b clock_v2_0/B 0.79fF
C3374 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# -0.14fF
C3375 ota_1/p1 a_mux4_en_0/in0 0.04fF
C3376 ota_1/m1_2463_n5585# ota_1/m1_2462_n3318# 0.01fF
C3377 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/c1_n930_n880# -0.21fF
C3378 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# -0.00fF
C3379 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# VDD 0.15fF
C3380 sky130_fd_sc_hd__mux4_1_2/a_834_97# sky130_fd_sc_hd__mux4_1_2/a_277_47# -0.01fF
C3381 a_mod_grp_ctrl_0 clock_v2_0/B 0.04fF
C3382 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0.00fF
C3383 transmission_gate_17/in clock_v2_0/p1d 0.25fF
C3384 a_mux4_en_1/switch_5t_0/in debug 0.01fF
C3385 VDD a_mux4_en_1/switch_5t_3/en -0.70fF
C3386 VSS ota_w_test_0/m1_6690_n8907# 0.46fF
C3387 clock_v2_0/Bd_b VSS 2.31fF
C3388 sky130_fd_sc_hd__mux4_1_1/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C3389 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X -0.00fF
C3390 sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# -0.31fF
C3391 sky130_fd_sc_hd__mux4_1_3/a_247_21# clock_v2_0/A_b 0.07fF
C3392 a_mux4_en_1/in2 clock_v2_0/B_b 0.03fF
C3393 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# clock_v2_0/p2 0.05fF
C3394 ota_w_test_0/cm ota_w_test_0/m1_1038_n2886# 0.07fF
C3395 a_mux4_en_1/switch_5t_1/transmission_gate_1/in a_mux4_en_1/switch_5t_1/in -0.00fF
C3396 transmission_gate_6/in sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# 0.30fF
C3397 VSS a_mod_grp_ctrl_0 6.83fF
C3398 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0.00fF
C3399 VDD a_mux4_en_1/in3 -0.63fF
C3400 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.30fF
C3401 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# -0.00fF
C3402 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.25fF
C3403 ota_1/p2_b clock_v2_0/p2_b 2.30fF
C3404 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_193_413# -0.00fF
C3405 ota_1/p1 sky130_fd_sc_hd__mux4_1_3/a_277_47# 0.01fF
C3406 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# -0.12fF
C3407 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0.00fF
C3408 sky130_fd_sc_hd__mux4_1_3/a_27_47# clock_v2_0/A 0.01fF
C3409 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X 0.00fF
C3410 ota_1/ip VSS 2.32fF
C3411 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.67fF
C3412 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A -0.00fF
C3413 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# -0.24fF
C3414 a_mux4_en_0/switch_5t_0/en_b a_mux4_en_0/switch_5t_0/transmission_gate_1/in 0.00fF
C3415 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0.03fF
C3416 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A -0.01fF
C3417 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# -0.00fF
C3418 ota_1/p1 ota_1/m1_n1659_n11581# 0.06fF
C3419 ota_1/sc_cmfb_0/transmission_gate_3/out VDD 0.81fF
C3420 a_mux2_en_0/switch_5t_1/en VDD 0.89fF
C3421 sky130_fd_sc_hd__mux4_1_1/a_277_47# sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0.01fF
C3422 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# -0.00fF
C3423 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# VDD 0.14fF
C3424 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B 0.09fF
C3425 sky130_fd_sc_hd__mux4_1_3/a_277_47# d_clk_grp_1_ctrl_0 0.08fF
C3426 ota_1/p2 clock_v2_0/p2_b 1.19fF
C3427 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/X clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# -0.00fF
C3428 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0.00fF
C3429 ip in 0.40fF
C3430 ota_w_test_0/op clock_v2_0/B 0.05fF
C3431 ota_1/m1_2462_n3318# ota_1/p1_b 0.02fF
C3432 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/sc_cmfb_0/transmission_gate_6/in -0.00fF
C3433 sky130_fd_sc_hd__mux4_1_1/a_277_47# ota_1/p2 0.00fF
C3434 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.03fF
C3435 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# -0.13fF
C3436 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0.00fF
C3437 a_mux2_en_1/transmission_gate_1/en_b debug -0.00fF
C3438 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# ota_1/in 0.13fF
C3439 VSS ota_w_test_0/op 1.69fF
C3440 transmission_gate_26/en ota_1/p1 0.98fF
C3441 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_10/a_110_47# -0.00fF
C3442 clock_v2_0/Bd_b ota_1/p2_b 5.40fF
C3443 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0.11fF
C3444 transmission_gate_32/out VDD 1.29fF
C3445 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0.00fF
C3446 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# -0.00fF
C3447 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# -0.09fF
C3448 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/op 0.00fF
C3449 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/c1_n260_n210# 0.03fF
C3450 clock_v2_0/Bd d_clk_grp_2_ctrl_0 0.01fF
C3451 a_mod_grp_ctrl_0 ota_1/p2_b 0.04fF
C3452 VDD clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y 0.09fF
C3453 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0.11fF
C3454 sky130_fd_sc_hd__mux4_1_2/a_247_21# clock_v2_0/p2 0.01fF
C3455 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# -0.00fF
C3456 ota_1/p2_b ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0.05fF
C3457 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0.24fF
C3458 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_11/a_110_47# VDD 0.08fF
C3459 comparator_v2_0/li_940_818# ota_1/p1_b 1.36fF
C3460 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0.09fF
C3461 VSS sky130_fd_sc_hd__mux4_1_3/a_193_413# 0.01fF
C3462 ota_1/cmc ota_1/sc_cmfb_0/transmission_gate_6/in -0.03fF
C3463 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_21/c1_n530_n480# 0.13fF
C3464 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# -0.00fF
C3465 clock_v2_0/Bd_b ota_1/p2 1.54fF
C3466 ota_w_test_0/on clock_v2_0/B_b 0.05fF
C3467 VSS ota_1/bias_a 4.67fF
C3468 transmission_gate_31/out transmission_gate_32/out 1.12fF
C3469 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_1/bias_a 0.02fF
C3470 sky130_fd_sc_hd__mux4_1_1/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00fF
C3471 ota_1/ip ota_1/p2_b 1.48fF
C3472 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0.08fF
C3473 a_mux4_en_0/in1 ota_w_test_0/cm 0.09fF
C3474 ota_1/ip sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# 0.13fF
C3475 a_mod_grp_ctrl_0 ota_1/p2 0.04fF
C3476 clock_v2_0/Bd clock_v2_0/sky130_fd_sc_hd__clkbuf_16_1/a_110_47# -0.00fF
C3477 ota_1/p2 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0.02fF
C3478 a_mux4_en_0/switch_5t_2/transmission_gate_1/in a_mux4_en_0/switch_5t_2/en_b 0.00fF
C3479 VDD a_mux4_en_1/switch_5t_1/in 0.37fF
C3480 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# ota_1/p1 0.09fF
C3481 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# -0.00fF
C3482 ota_w_test_0/cm ota_w_test_0/ip 0.55fF
C3483 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/A -0.01fF
C3484 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/c1_n930_n880# transmission_gate_17/in 0.11fF
C3485 ota_1/ip ota_1/in 1.16fF
C3486 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# VDD 0.00fF
C3487 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0.03fF
C3488 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# ota_1/p2 0.00fF
C3489 ota_1/ip ota_1/p2 0.29fF
C3490 VSS a_mux2_en_0/switch_5t_0/in 0.01fF
C3491 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.01fF
C3492 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# -0.00fF
C3493 VDD clock_v2_0/sky130_fd_sc_hd__mux2_1_0/X -0.00fF
C3494 ota_w_test_0/op ota_1/p2_b 0.13fF
C3495 a_mux4_en_1/switch_5t_1/en a_mux4_en_1/switch_5t_0/en_b 0.00fF
C3496 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0.00fF
C3497 VDD clock_v2_0/p2_b 3.24fF
C3498 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0.04fF
C3499 sky130_fd_sc_hd__mux4_1_2/a_193_413# clock_v2_0/p2_b 0.04fF
C3500 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_12/a_110_47# -0.00fF
C3501 ota_w_test_0/cm ota_w_test_0/m1_n5574_n13620# 0.01fF
C3502 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/c1_n530_n480# ota_1/p1_b 0.04fF
C3503 transmission_gate_18/in transmission_gate_5/in 5.42fF
C3504 VDD a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0.02fF
C3505 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# -0.15fF
C3506 sky130_fd_sc_hd__mux4_1_1/a_277_47# VDD 0.16fF
C3507 clock_v2_0/Bd sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.01fF
C3508 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in VDD -1.17fF
C3509 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# -0.00fF
C3510 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# -0.00fF
C3511 ota_w_test_0/op ota_1/p2 1.42fF
C3512 transmission_gate_32/out clock_v2_0/p1d_b 5.94fF
C3513 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.00fF
C3514 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# ota_1/on 0.06fF
C3515 ota_1/bias_a ota_1/p2_b 0.02fF
C3516 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0.00fF
C3517 ota_1/cm ota_1/on 0.01fF
C3518 sky130_fd_sc_hd__mux4_1_2/a_27_47# clock_v2_0/p2 -0.00fF
C3519 transmission_gate_26/en transmission_gate_17/in 0.08fF
C3520 a_mux4_en_0/switch_5t_1/en_b a_mux4_en_0/switch_5t_0/en_b 0.00fF
C3521 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y 0.01fF
C3522 VSS d_probe_1 1.91fF
C3523 debug a_mux4_en_1/transmission_gate_3/en_b 0.07fF
C3524 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0.00fF
C3525 transmission_gate_31/out clock_v2_0/p2_b 0.16fF
C3526 clock_v2_0/Ad_b clock_v2_0/p2_b 0.05fF
C3527 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00fF
C3528 d_clk_grp_2_ctrl_0 clock_v2_0/p1d 0.00fF
C3529 ota_1/cmc ota_1/sc_cmfb_0/transmission_gate_9/in -0.00fF
C3530 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_11/a_110_47# clock_v2_0/p1d_b -0.00fF
C3531 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/c1_n530_n480# -0.08fF
C3532 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# VDD -0.00fF
C3533 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# transmission_gate_8/in 0.40fF
C3534 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/Ad_b 0.11fF
C3535 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/c1_n930_n880# 1.58fF
C3536 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/A clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C3537 ota_1/p2 ota_1/bias_a 0.06fF
C3538 clock_v2_0/Bd_b VDD 13.69fF
C3539 ota_1/m1_n947_n12836# ota_1/p1_b 0.08fF
C3540 sky130_fd_sc_hd__mux4_1_1/a_247_21# sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.00fF
C3541 ota_w_test_0/m1_6690_n8907# VDD 0.79fF
C3542 a_mux4_en_1/in2 clock_v2_0/B 0.03fF
C3543 ota_1/p1_b clock_v2_0/p2 3.37fF
C3544 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C3545 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A -0.00fF
C3546 a_mod_grp_ctrl_0 VDD 5.62fF
C3547 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.00fF
C3548 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0.00fF
C3549 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# 0.07fF
C3550 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# ota_1/op 0.34fF
C3551 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# VDD 0.07fF
C3552 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/A clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A -0.00fF
C3553 VSS a_mux4_en_1/in2 1.49fF
C3554 VSS ota_w_test_0/m1_n208_n2883# 1.05fF
C3555 VSS a_mux4_en_1/switch_5t_0/transmission_gate_1/in 0.37fF
C3556 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# 0.29fF
C3557 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# 0.14fF
C3558 a_mod_grp_ctrl_1 clock_v2_0/B_b 0.06fF
C3559 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.02fF
C3560 transmission_gate_18/in VSS 4.08fF
C3561 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0.00fF
C3562 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0.00fF
C3563 transmission_gate_21/in ota_1/p1 0.17fF
C3564 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# -0.35fF
C3565 clock_v2_0/Bd_b clock_v2_0/Ad_b 7.79fF
C3566 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# -0.00fF
C3567 ota_1/ip VDD 1.21fF
C3568 op comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.00fF
C3569 ota_1/cmc ota_1/m1_n5574_n13620# 0.06fF
C3570 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X -0.01fF
C3571 clock_v2_0/p1d_b clock_v2_0/p2_b 2.20fF
C3572 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# 0.09fF
C3573 clock_v2_0/Bd debug 0.06fF
C3574 a_mod_grp_ctrl_0 clock_v2_0/Ad_b 0.04fF
C3575 a_mux4_en_0/switch_5t_3/en_b a_mux4_en_0/switch_5t_3/transmission_gate_1/in -0.00fF
C3576 VSS ota_w_test_0/sc_cmfb_0/transmission_gate_4/out 0.61fF
C3577 ota_1/p1 ota_1/sc_cmfb_0/transmission_gate_9/in 0.00fF
C3578 VSS ota_1/bias_b 1.11fF
C3579 op comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X 0.00fF
C3580 ota_w_test_0/sc_cmfb_0/transmission_gate_9/in ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0.00fF
C3581 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.00fF
C3582 sky130_fd_sc_hd__mux4_1_3/a_668_97# sky130_fd_sc_hd__mux4_1_2/a_834_97# 0.00fF
C3583 sky130_fd_sc_hd__mux4_1_1/a_277_47# clock_v2_0/p1d_b 0.04fF
C3584 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0.00fF
C3585 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# 0.30fF
C3586 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__mux4_1_0/a_27_47# -0.00fF
C3587 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0.02fF
C3588 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/c1_n930_n880# 0.11fF
C3589 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0.00fF
C3590 sky130_fd_sc_hd__mux4_1_0/a_27_413# clock_v2_0/p1d 0.00fF
C3591 ota_1/p1 i_bias_2 0.10fF
C3592 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.04fF
C3593 ota_1/ip transmission_gate_31/out 0.03fF
C3594 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A -0.00fF
C3595 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# -0.00fF
C3596 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/c1_n260_n210# 0.03fF
C3597 ota_w_test_0/op VDD 2.69fF
C3598 d_clk_grp_1_ctrl_1 d_probe_0 0.69fF
C3599 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/c1_n530_n480# -0.08fF
C3600 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/X 0.00fF
C3601 VSS sky130_fd_sc_hd__mux4_1_0/a_923_363# -0.11fF
C3602 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0.14fF
C3603 sky130_fd_sc_hd__clkinv_4_3/Y sky130_fd_sc_hd__mux4_1_2/X 0.25fF
C3604 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# -0.00fF
C3605 transmission_gate_18/in transmission_gate_6/in -3.48fF
C3606 sky130_fd_sc_hd__mux4_1_3/a_750_97# clock_v2_0/A 0.00fF
C3607 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.02fF
C3608 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0.00fF
C3609 a_mux4_en_0/switch_5t_2/en a_mux4_en_0/switch_5t_2/en_b 0.00fF
C3610 transmission_gate_8/in transmission_gate_5/in 2.22fF
C3611 VSS a_probe_2 2.75fF
C3612 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# -0.01fF
C3613 transmission_gate_0/out transmission_gate_2/out 0.19fF
C3614 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# VDD 0.00fF
C3615 clock_v2_0/Bd_b clock_v2_0/p1d_b 0.13fF
C3616 ota_w_test_0/on clock_v2_0/B 0.05fF
C3617 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480# ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# -0.19fF
C3618 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0.03fF
C3619 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.04fF
C3620 sky130_fd_sc_hd__mux4_1_3/a_193_413# VDD 0.06fF
C3621 sky130_fd_sc_hd__mux4_1_3/a_193_413# sky130_fd_sc_hd__mux4_1_2/a_193_413# 0.01fF
C3622 VSS ota_1/bias_c 1.52fF
C3623 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/c1_n260_n210# 0.03fF
C3624 transmission_gate_18/in ota_1/p2_b 0.08fF
C3625 a_mux4_en_1/in2 ota_w_test_0/m1_11648_n10486# 0.05fF
C3626 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# VDD 0.05fF
C3627 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_3/a_750_97# 0.01fF
C3628 sky130_fd_sc_hd__mux4_1_2/a_27_47# sky130_fd_sc_hd__mux4_1_3/a_27_47# 0.01fF
C3629 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0.00fF
C3630 sky130_fd_sc_hd__mux4_1_1/a_1290_413# clock_v2_0/p1d 0.00fF
C3631 ota_w_test_0/op clock_v2_0/Ad_b 0.44fF
C3632 VSS ota_w_test_0/m1_n2176_n12171# 0.73fF
C3633 ota_1/bias_a VDD 3.33fF
C3634 ota_1/p1 ota_1/m1_n5574_n13620# 0.23fF
C3635 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413# clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D -0.00fF
C3636 sky130_fd_sc_hd__clkinv_4_4/Y sky130_fd_sc_hd__mux4_1_2/X 0.02fF
C3637 clock_v2_0/Bd sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.00fF
C3638 VSS clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.00fF
C3639 a_mod_grp_ctrl_0 clock_v2_0/p1d_b 0.06fF
C3640 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/c1_n530_n480# ota_1/sc_cmfb_0/transmission_gate_6/in 0.02fF
C3641 VSS sky130_fd_sc_hd__mux4_1_1/a_27_47# 0.09fF
C3642 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480# -0.10fF
C3643 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/c1_n930_n880# -0.44fF
C3644 a_mux4_en_0/in1 clock_v2_0/A_b 0.03fF
C3645 VSS ota_w_test_0/on 1.90fF
C3646 VSS clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y 0.37fF
C3647 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# 0.04fF
C3648 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0.09fF
C3649 a_mux4_en_1/in2 ota_1/p2 -0.00fF
C3650 VSS a_mux4_en_1/switch_5t_3/transmission_gate_1/in 0.34fF
C3651 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0.00fF
C3652 transmission_gate_18/in ota_1/p2 0.08fF
C3653 a_mod_grp_ctrl_0 a_mux4_en_0/switch_5t_0/in 0.00fF
C3654 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0.01fF
C3655 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/c1_n930_n880# transmission_gate_8/in 0.03fF
C3656 ota_w_test_0/cm clock_v2_0/B_b 0.18fF
C3657 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# 0.31fF
C3658 ota_1/ip clock_v2_0/p1d_b 0.00fF
C3659 clock_v2_0/A_b ota_w_test_0/ip 0.09fF
C3660 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# -0.00fF
C3661 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0.00fF
C3662 a_mux2_en_0/switch_5t_0/in VDD 0.48fF
C3663 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y -0.00fF
C3664 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# -0.00fF
C3665 ota_w_test_0/m1_1038_n2886# a_mux4_en_1/in1 0.06fF
C3666 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 1.18fF
C3667 ota_w_test_0/m1_1038_n2886# i_bias_1 -0.01fF
C3668 VDD comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# 0.08fF
C3669 debug clock_v2_0/p1d 0.07fF
C3670 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0.00fF
C3671 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# transmission_gate_6/in 0.21fF
C3672 sky130_fd_sc_hd__mux4_1_3/a_757_363# clock_v2_0/A_b 0.01fF
C3673 VSS sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/c1_n930_n880# 2.06fF
C3674 a_mux4_en_1/switch_5t_2/en a_probe_2 0.00fF
C3675 VSS transmission_gate_8/in 0.66fF
C3676 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_12/a_110_47# VDD -1.38fF
C3677 ota_1/sc_cmfb_0/transmission_gate_3/out ota_1/on 0.00fF
C3678 comparator_v2_0/li_n2324_818# comparator_v2_0/li_940_3458# 0.00fF
C3679 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980# 0.30fF
C3680 VDD sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/c1_n930_n880# 2.72fF
C3681 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0.09fF
C3682 ota_1/sc_cmfb_0/transmission_gate_8/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0.12fF
C3683 VSS clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# 0.00fF
C3684 sky130_fd_sc_hd__mux4_1_0/a_923_363# ota_1/p2 -0.50fF
C3685 sky130_fd_sc_hd__mux4_1_2/X sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C3686 clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y VDD 0.08fF
C3687 d_probe_1 VDD 2.15fF
C3688 VSS ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0.31fF
C3689 sky130_fd_sc_hd__mux4_1_3/X sky130_fd_sc_hd__mux4_1_2/X 0.06fF
C3690 ota_1/p1 sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.01fF
C3691 sky130_fd_sc_hd__mux4_1_1/a_27_47# ota_1/p2_b 0.00fF
C3692 a_mux4_en_1/switch_5t_1/transmission_gate_1/in a_probe_2 0.00fF
C3693 ota_1/p2_b ota_w_test_0/on 1.30fF
C3694 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__clkinv_4_3/Y 0.02fF
C3695 a_mux4_en_0/in2 clock_v2_0/A_b 0.03fF
C3696 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0.00fF
C3697 transmission_gate_32/out ota_1/on 0.10fF
C3698 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0.06fF
C3699 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# ota_1/p1 0.03fF
C3700 VSS a_mux4_en_0/switch_5t_1/transmission_gate_1/in 0.43fF
C3701 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0.02fF
C3702 sky130_fd_sc_hd__mux4_1_3/a_247_21# d_clk_grp_1_ctrl_0 0.19fF
C3703 transmission_gate_0/out clock_v2_0/p1d 2.73fF
C3704 VSS a_mux4_en_0/switch_5t_3/in 0.04fF
C3705 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# -0.00fF
C3706 a_probe_3 a_mux4_en_0/switch_5t_3/transmission_gate_1/in 0.00fF
C3707 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0.06fF
C3708 sky130_fd_sc_hd__mux4_1_2/a_277_47# clock_v2_0/p2_b 0.04fF
C3709 ota_1/p2 ota_w_test_0/on 0.10fF
C3710 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0.02fF
C3711 sky130_fd_sc_hd__mux4_1_3/a_247_21# sky130_fd_sc_hd__mux4_1_2/a_668_97# 0.00fF
C3712 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# clock_v2_0/p1d 0.15fF
C3713 clock_v2_0/Bd clock_v2_0/A 0.23fF
C3714 a_mod_grp_ctrl_1 clock_v2_0/B 0.05fF
C3715 VSS ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# -0.27fF
C3716 a_mux4_en_1/in2 VDD -0.44fF
C3717 ota_w_test_0/m1_n208_n2883# VDD 1.10fF
C3718 VDD a_mux4_en_1/switch_5t_0/transmission_gate_1/in -0.87fF
C3719 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# VDD 0.10fF
C3720 transmission_gate_8/in ota_1/p2_b 0.07fF
C3721 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# -0.13fF
C3722 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# 0.11fF
C3723 ota_1/p1 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0.23fF
C3724 transmission_gate_18/in VDD 13.65fF
C3725 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X -0.77fF
C3726 a_mux4_en_0/in0 debug 0.02fF
C3727 VDD clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0.13fF
C3728 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.01fF
C3729 VSS a_mod_grp_ctrl_1 3.74fF
C3730 a_mux4_en_0/in1 a_mux4_en_1/in1 0.14fF
C3731 sky130_fd_sc_hd__mux4_1_2/a_757_363# sky130_fd_sc_hd__mux4_1_3/a_247_21# 0.00fF
C3732 sky130_fd_sc_hd__mux4_1_2/a_1478_413# clock_v2_0/p2_b -0.00fF
C3733 a_mux4_en_0/in1 i_bias_1 0.08fF
C3734 VSS clock_v2_0/sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0.00fF
C3735 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0.24fF
C3736 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0.03fF
C3737 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0.04fF
C3738 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# VDD 0.00fF
C3739 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out VDD 0.12fF
C3740 a_mod_grp_ctrl_0 a_mux4_en_1/sky130_fd_sc_hd__nand2_1_2/a_113_47# 0.00fF
C3741 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0.00fF
C3742 ota_1/bias_b VDD 2.17fF
C3743 transmission_gate_8/in ota_1/p2 0.03fF
C3744 a_mux4_en_1/in2 clock_v2_0/Ad_b 0.04fF
C3745 VSS a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0.15fF
C3746 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0.10fF
C3747 i_bias_1 ota_w_test_0/ip -0.01fF
C3748 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/c1_n530_n480# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# -0.00fF
C3749 transmission_gate_18/in transmission_gate_31/out 0.00fF
C3750 ota_1/sc_cmfb_0/transmission_gate_7/in ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0.12fF
C3751 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__clkinv_4_3/Y 0.00fF
C3752 op clock_v2_0/p2_b 0.01fF
C3753 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# transmission_gate_2/out 0.30fF
C3754 transmission_gate_18/in clock_v2_0/Ad_b 0.47fF
C3755 sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/c1_n260_n210# 0.03fF
C3756 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0.00fF
C3757 sky130_fd_sc_hd__mux4_1_3/a_750_97# sky130_fd_sc_hd__mux4_1_2/a_247_21# 0.00fF
C3758 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/c1_n530_n480# ota_1/p1_b 0.04fF
C3759 clock_v2_0/Ad_b clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# -0.00fF
C3760 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# clock_v2_0/p2 0.03fF
C3761 ota_w_test_0/cm transmission_gate_5/in 0.27fF
C3762 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0.04fF
C3763 sky130_fd_sc_hd__mux4_1_0/a_923_363# VDD -0.02fF
C3764 onebit_dac_0/out onebit_dac_1/out 0.26fF
C3765 a_mux4_en_0/switch_5t_0/en_b a_mux4_en_0/transmission_gate_3/en_b 0.00fF
C3766 a_mux4_en_0/switch_5t_1/en a_mux4_en_0/switch_5t_1/in -0.00fF
C3767 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# 0.05fF
C3768 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0.00fF
C3769 sky130_fd_sc_hd__mux4_1_2/a_1290_413# sky130_fd_sc_hd__mux4_1_2/a_750_97# 0.01fF
C3770 ota_w_test_0/sc_cmfb_0/transmission_gate_3/out ota_w_test_0/sc_cmfb_0/transmission_gate_9/in -0.01fF
C3771 a_mux4_en_1/switch_5t_2/transmission_gate_1/in a_probe_2 0.00fF
C3772 VDD a_probe_2 -4.01fF
C3773 ota_w_test_0/m1_n5574_n13620# a_mux4_en_1/in1 1.43fF
C3774 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0.00fF
C3775 i_bias_1 ota_w_test_0/m1_n5574_n13620# -0.01fF
C3776 d_clk_grp_1_ctrl_1 sky130_fd_sc_hd__clkinv_4_4/Y 0.00fF
C3777 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/c1_n260_n210# sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# -0.04fF
C3778 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/p2_b 0.00fF
C3779 a_mux2_en_1/switch_5t_0/in debug -0.00fF
C3780 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# -0.00fF
C3781 clock_v2_0/Bd rst_n 0.23fF
C3782 ota_1/bias_c VDD 4.07fF
C3783 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# VDD 1.01fF
C3784 sky130_fd_sc_hd__clkinv_4_1/Y sky130_fd_sc_hd__clkinv_4_2/Y 0.17fF
C3785 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0.59fF
C3786 ota_w_test_0/m1_n2176_n12171# VDD -0.10fF
C3787 a_mux4_en_1/switch_5t_2/en a_mod_grp_ctrl_1 0.04fF
C3788 ota_1/p2_b a_mod_grp_ctrl_1 0.05fF
C3789 VDD clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0.06fF
C3790 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# -0.00fF
C3791 sky130_fd_sc_hd__mux4_1_1/a_27_47# VDD 0.01fF
C3792 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/c1_n530_n480# VDD 0.10fF
C3793 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# -0.00fF
C3794 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_0/a_668_97# -0.02fF
C3795 ota_w_test_0/on VDD 2.37fF
C3796 clock_v2_0/p1d clock_v2_0/A 0.07fF
C3797 sky130_fd_sc_hd__mux4_1_2/a_834_97# clock_v2_0/p2_b 0.00fF
C3798 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y VDD 0.31fF
C3799 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0.09fF
C3800 a_probe_0 a_mux2_en_0/switch_5t_1/en 0.00fF
C3801 ota_1/bias_d ota_1/m1_n1659_n11581# 0.02fF
C3802 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# ota_1/p2 0.00fF
C3803 ota_w_test_0/cm clock_v2_0/B 0.20fF
C3804 VDD a_mux4_en_1/switch_5t_3/transmission_gate_1/in -1.17fF
C3805 transmission_gate_18/in clock_v2_0/p1d_b 0.30fF
C3806 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0.22fF
C3807 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A VDD 0.08fF
C3808 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# transmission_gate_5/in 0.18fF
C3809 sky130_fd_sc_hd__mux4_1_1/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00fF
C3810 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0.07fF
C3811 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# -0.14fF
C3812 clock_v2_0/Bd_b clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y -0.00fF
C3813 clock_v2_0/A_b clock_v2_0/B_b 6.50fF
C3814 ota_1/p2 a_mod_grp_ctrl_1 0.06fF
C3815 clock_v2_0/Bd_b sky130_fd_sc_hd__mux4_1_1/a_757_363# 0.00fF
C3816 transmission_gate_19/out transmission_gate_17/in 0.00fF
C3817 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# 0.21fF
C3818 VDD clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# -0.00fF
C3819 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# 0.18fF
C3820 sky130_fd_sc_hd__mux4_1_1/a_27_47# clock_v2_0/Ad_b 0.05fF
C3821 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0.03fF
C3822 VSS ota_w_test_0/cm 0.92fF
C3823 VSS clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0.05fF
C3824 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# ota_1/on 0.00fF
C3825 VSS transmission_gate_19/in 0.50fF
C3826 VDD clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0.33fF
C3827 d_clk_grp_1_ctrl_1 clock_v2_0/A 0.00fF
C3828 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/c1_n530_n480# -0.25fF
C3829 sky130_fd_sc_hd__mux4_1_2/a_247_21# sky130_fd_sc_hd__mux4_1_2/X 0.00fF
C3830 clock_v2_0/p2_b 0 34.48fF
C3831 clock_v2_0/p2 0 64.24fF
C3832 sky130_fd_pr__cap_mim_m3_1_CEWQ64_1/m3_n360_n310# 0 0.63fF
C3833 sky130_fd_pr__cap_mim_m3_1_CGPBWM_39/m3_n1030_n980# 0 2.84fF
C3834 sky130_fd_pr__cap_mim_m3_1_CGPBWM_28/m3_n1030_n980# 0 2.84fF
C3835 sky130_fd_pr__cap_mim_m3_1_CGPBWM_27/m3_n1030_n980# 0 2.84fF
C3836 sky130_fd_pr__cap_mim_m3_1_CGPBWM_38/m3_n1030_n980# 0 2.84fF
C3837 sky130_fd_pr__cap_mim_m3_1_CEWQ64_0/m3_n360_n310# 0 0.63fF
C3838 sky130_fd_pr__cap_mim_m3_1_CGPBWM_26/m3_n1030_n980# 0 2.84fF
C3839 sky130_fd_pr__cap_mim_m3_1_CGPBWM_14/m3_n1030_n980# 0 2.84fF
C3840 sky130_fd_pr__cap_mim_m3_1_CGPBWM_25/m3_n1030_n980# 0 2.84fF
C3841 sky130_fd_pr__cap_mim_m3_1_CGPBWM_47/m3_n1030_n980# 0 2.84fF
C3842 sky130_fd_pr__cap_mim_m3_1_CGPBWM_24/m3_n1030_n980# 0 2.84fF
C3843 sky130_fd_pr__cap_mim_m3_1_CGPBWM_46/m3_n1030_n980# 0 2.84fF
C3844 comparator_v2_0/li_940_3458# 0 -1592.65fF
C3845 comparator_v2_0/li_940_818# 0 -2262.83fF
C3846 ota_1/on 0 -353.00fF
C3847 comparator_v2_0/li_n2324_818# 0 -3722.01fF
C3848 ota_1/op 0 -438.61fF
C3849 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/A 0 -127.11fF
C3850 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/A 0 -211.82fF
C3851 ota_1/p1_b 0 115.55fF
C3852 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/a_27_47# 0 0.15fF
C3853 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/a_27_47# 0 0.15fF
C3854 comparator_v2_0/sky130_fd_sc_hd__buf_2_0/X 0 43.25fF
C3855 comparator_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# 0 0.06fF
C3856 comparator_v2_0/sky130_fd_sc_hd__buf_2_1/X 0 23.78fF
C3857 comparator_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# 0 0.06fF
C3858 sky130_fd_pr__cap_mim_m3_1_CGPBWM_45/m3_n1030_n980# 0 2.84fF
C3859 sky130_fd_pr__cap_mim_m3_1_CGPBWM_44/m3_n1030_n980# 0 2.84fF
C3860 sky130_fd_pr__cap_mim_m3_1_CGPBWM_43/m3_n1030_n980# 0 2.84fF
C3861 sky130_fd_pr__cap_mim_m3_1_CGPBWM_42/m3_n1030_n980# 0 2.84fF
C3862 sky130_fd_pr__cap_mim_m3_1_CGPBWM_41/m3_n1030_n980# 0 2.84fF
C3863 sky130_fd_pr__cap_mim_m3_1_CGPBWM_40/m3_n1030_n980# 0 2.84fF
C3864 a_mux4_en_1/sky130_fd_sc_hd__inv_1_1/Y 0 23.85fF
C3865 a_mux4_en_1/sky130_fd_sc_hd__inv_1_0/Y 0 18.27fF
C3866 a_mux4_en_1/switch_5t_3/in 0 0.83fF
C3867 a_mux4_en_1/in3 0 0.42fF
C3868 a_mux4_en_1/transmission_gate_3/en_b 0 7.48fF
C3869 a_mux4_en_1/switch_5t_2/in 0 0.04fF
C3870 a_mux4_en_1/switch_5t_1/in 0 0.15fF
C3871 a_mux4_en_1/switch_5t_0/in 0 2.48fF
C3872 a_mux4_en_1/switch_5t_3/en 0 3.80fF
C3873 a_probe_2 0 4.74fF
C3874 a_mux4_en_1/switch_5t_3/en_b 0 8.52fF
C3875 a_mux4_en_1/switch_5t_3/transmission_gate_1/in 0 1.77fF
C3876 a_mux4_en_1/switch_5t_2/en 0 5.06fF
C3877 a_mux4_en_1/switch_5t_2/en_b 0 11.31fF
C3878 a_mux4_en_1/switch_5t_2/transmission_gate_1/in 0 1.77fF
C3879 a_mux4_en_1/switch_5t_1/en 0 12.94fF
C3880 a_mux4_en_1/switch_5t_1/en_b 0 -2.82fF
C3881 a_mux4_en_1/switch_5t_1/transmission_gate_1/in 0 1.77fF
C3882 a_mux4_en_1/switch_5t_0/en 0 4.30fF
C3883 a_mux4_en_1/switch_5t_0/en_b 0 8.42fF
C3884 a_mux4_en_1/switch_5t_0/transmission_gate_1/in 0 1.77fF
C3885 a_mux4_en_0/sky130_fd_sc_hd__inv_1_1/Y 0 23.85fF
C3886 a_mod_grp_ctrl_1 0 127.97fF
C3887 a_mux4_en_0/sky130_fd_sc_hd__inv_1_0/Y 0 18.27fF
C3888 debug 0 62.27fF
C3889 a_mux4_en_0/switch_5t_3/in 0 0.83fF
C3890 a_mux4_en_0/in3 0 0.42fF
C3891 a_mux4_en_0/transmission_gate_3/en_b 0 7.48fF
C3892 a_mux4_en_0/switch_5t_2/in 0 0.04fF
C3893 a_mux4_en_0/switch_5t_1/in 0 0.15fF
C3894 a_mux4_en_0/switch_5t_0/in 0 2.48fF
C3895 a_mux4_en_0/switch_5t_3/en 0 3.80fF
C3896 a_probe_3 0 4.75fF
C3897 a_mux4_en_0/switch_5t_3/en_b 0 8.52fF
C3898 a_mux4_en_0/switch_5t_3/transmission_gate_1/in 0 1.77fF
C3899 a_mux4_en_0/switch_5t_2/en 0 5.06fF
C3900 a_mux4_en_0/switch_5t_2/en_b 0 11.31fF
C3901 a_mux4_en_0/switch_5t_2/transmission_gate_1/in 0 1.77fF
C3902 a_mux4_en_0/switch_5t_1/en 0 12.94fF
C3903 a_mux4_en_0/switch_5t_1/en_b 0 -2.82fF
C3904 a_mux4_en_0/switch_5t_1/transmission_gate_1/in 0 1.77fF
C3905 a_mux4_en_0/switch_5t_0/en 0 4.30fF
C3906 a_mux4_en_0/switch_5t_0/en_b 0 8.42fF
C3907 a_mux4_en_0/switch_5t_0/transmission_gate_1/in 0 1.77fF
C3908 transmission_gate_8/in 0 4.25fF
C3909 transmission_gate_6/in 0 8.31fF
C3910 transmission_gate_9/in 0 -1.11fF
C3911 clock_v2_0/A 0 63.59fF
C3912 ota_w_test_0/ip 0 -8.61fF
C3913 clock_v2_0/A_b 0 77.74fF
C3914 clock_v2_0/B 0 39.11fF
C3915 transmission_gate_5/in 0 11.01fF
C3916 clock_v2_0/B_b 0 68.14fF
C3917 sky130_fd_pr__cap_mim_m3_1_CGPBWM_9/m3_n1030_n980# 0 2.84fF
C3918 ota_w_test_0/in 0 -8.63fF
C3919 clock_v2_0/p1d 0 -42.17fF
C3920 transmission_gate_2/out 0 17.37fF
C3921 in 0 14.88fF
C3922 clock_v2_0/p1d_b 0 11.93fF
C3923 clk 0 26.18fF
C3924 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_10/a_110_47# 0 1.28fF
C3925 clock_v2_0/sky130_fd_sc_hd__nand2_1_0/B 0 19.52fF
C3926 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/Y 0 33.52fF
C3927 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/S 0 9.62fF
C3928 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_505_21# 0 0.15fF
C3929 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/a_76_199# 0 0.11fF
C3930 clock_v2_0/sky130_fd_sc_hd__mux2_1_0/X 0 42.71fF
C3931 clock_v2_0/sky130_fd_sc_hd__clkinv_1_2/Y 0 24.38fF
C3932 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/A 0 23.06fF
C3933 clock_v2_0/sky130_fd_sc_hd__nand2_1_3/A 0 18.36fF
C3934 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/X 0 8.07fF
C3935 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_390_47# 0 0.10fF
C3936 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_283_47# 0 0.18fF
C3937 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/a_27_47# 0 0.18fF
C3938 clock_v2_0/sky130_fd_sc_hd__clkinv_1_1/Y 0 32.07fF
C3939 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/A 0 15.33fF
C3940 clock_v2_0/sky130_fd_sc_hd__nand2_1_2/A 0 12.52fF
C3941 clock_v2_0/sky130_fd_sc_hd__nand2_1_2/B 0 10.41fF
C3942 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_109/X 0 8.14fF
C3943 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_390_47# 0 0.10fF
C3944 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_283_47# 0 0.18fF
C3945 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/a_27_47# 0 0.18fF
C3946 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/A 0 24.52fF
C3947 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_390_47# 0 0.10fF
C3948 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_283_47# 0 0.18fF
C3949 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/a_27_47# 0 0.18fF
C3950 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/A 0 22.88fF
C3951 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_390_47# 0 0.10fF
C3952 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_283_47# 0 0.18fF
C3953 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_18/a_27_47# 0 0.18fF
C3954 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/Y 0 28.40fF
C3955 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_9/a_110_47# 0 1.28fF
C3956 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/A 0 22.93fF
C3957 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/B 0 12.62fF
C3958 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/X 0 19.67fF
C3959 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_390_47# 0 0.10fF
C3960 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_283_47# 0 0.18fF
C3961 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/a_27_47# 0 0.18fF
C3962 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/A 0 22.79fF
C3963 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_390_47# 0 0.10fF
C3964 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_283_47# 0 0.18fF
C3965 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/a_27_47# 0 0.18fF
C3966 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_108/X 0 11.25fF
C3967 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_390_47# 0 0.10fF
C3968 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_283_47# 0 0.18fF
C3969 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/a_27_47# 0 0.18fF
C3970 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/A 0 27.46fF
C3971 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/A 0 44.75fF
C3972 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_390_47# 0 0.10fF
C3973 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_283_47# 0 0.18fF
C3974 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_39/a_27_47# 0 0.18fF
C3975 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/X 0 14.09fF
C3976 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_390_47# 0 0.10fF
C3977 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_283_47# 0 0.18fF
C3978 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/a_27_47# 0 0.18fF
C3979 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_8/a_110_47# 0 1.28fF
C3980 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/A 0 18.86fF
C3981 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_118/A 0 20.20fF
C3982 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_390_47# 0 0.10fF
C3983 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_283_47# 0 0.18fF
C3984 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/a_27_47# 0 0.18fF
C3985 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/A 0 23.06fF
C3986 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_390_47# 0 0.10fF
C3987 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_283_47# 0 0.18fF
C3988 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/a_27_47# 0 0.18fF
C3989 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_29/A 0 20.23fF
C3990 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_390_47# 0 0.10fF
C3991 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_283_47# 0 0.18fF
C3992 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/a_27_47# 0 0.18fF
C3993 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_390_47# 0 0.10fF
C3994 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_283_47# 0 0.18fF
C3995 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_49/a_27_47# 0 0.18fF
C3996 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_7/a_110_47# 0 1.28fF
C3997 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/X 0 13.04fF
C3998 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_390_47# 0 0.10fF
C3999 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_283_47# 0 0.18fF
C4000 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/a_27_47# 0 0.18fF
C4001 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/A 0 24.50fF
C4002 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_390_47# 0 0.10fF
C4003 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_283_47# 0 0.18fF
C4004 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/a_27_47# 0 0.18fF
C4005 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_129/X 0 19.99fF
C4006 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_390_47# 0 0.10fF
C4007 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_283_47# 0 0.18fF
C4008 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/a_27_47# 0 0.18fF
C4009 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_117/A 0 14.35fF
C4010 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_390_47# 0 0.10fF
C4011 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_283_47# 0 0.18fF
C4012 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/a_27_47# 0 0.18fF
C4013 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/A 0 20.97fF
C4014 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_390_47# 0 0.10fF
C4015 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_283_47# 0 0.18fF
C4016 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_59/a_27_47# 0 0.18fF
C4017 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/A 0 23.98fF
C4018 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_390_47# 0 0.10fF
C4019 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_283_47# 0 0.18fF
C4020 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/a_27_47# 0 0.18fF
C4021 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_17/X 0 19.54fF
C4022 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_390_47# 0 0.10fF
C4023 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_283_47# 0 0.18fF
C4024 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/a_27_47# 0 0.18fF
C4025 clock_v2_0/sky130_fd_sc_hd__clkinv_4_4/Y 0 28.40fF
C4026 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_6/a_110_47# 0 1.28fF
C4027 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/A 0 42.29fF
C4028 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/X 0 23.44fF
C4029 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_390_47# 0 0.10fF
C4030 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_283_47# 0 0.18fF
C4031 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_159/a_27_47# 0 0.18fF
C4032 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/A 0 10.79fF
C4033 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_107/X 0 4.49fF
C4034 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_390_47# 0 0.10fF
C4035 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_283_47# 0 0.18fF
C4036 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_104/a_27_47# 0 0.18fF
C4037 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/X 0 14.02fF
C4038 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/X 0 24.11fF
C4039 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_390_47# 0 0.10fF
C4040 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_283_47# 0 0.18fF
C4041 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_69/a_27_47# 0 0.18fF
C4042 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_38/X 0 40.07fF
C4043 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_390_47# 0 0.10fF
C4044 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_283_47# 0 0.18fF
C4045 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/a_27_47# 0 0.18fF
C4046 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_390_47# 0 0.10fF
C4047 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_283_47# 0 0.18fF
C4048 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/a_27_47# 0 0.18fF
C4049 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/X 0 20.99fF
C4050 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_48/X 0 14.02fF
C4051 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_390_47# 0 0.10fF
C4052 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_283_47# 0 0.18fF
C4053 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_47/a_27_47# 0 0.18fF
C4054 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_27/A 0 21.65fF
C4055 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_390_47# 0 0.10fF
C4056 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_283_47# 0 0.18fF
C4057 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_25/a_27_47# 0 0.18fF
C4058 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_5/a_110_47# 0 1.28fF
C4059 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_390_47# 0 0.10fF
C4060 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_283_47# 0 0.18fF
C4061 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/a_27_47# 0 0.18fF
C4062 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/X 0 42.06fF
C4063 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_390_47# 0 0.10fF
C4064 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_283_47# 0 0.18fF
C4065 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/a_27_47# 0 0.18fF
C4066 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_138/A 0 20.22fF
C4067 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_390_47# 0 0.10fF
C4068 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_283_47# 0 0.18fF
C4069 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/a_27_47# 0 0.18fF
C4070 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_127/X 0 10.28fF
C4071 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_390_47# 0 0.10fF
C4072 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_283_47# 0 0.18fF
C4073 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/a_27_47# 0 0.18fF
C4074 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/B 0 54.46fF
C4075 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_390_47# 0 0.10fF
C4076 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_283_47# 0 0.18fF
C4077 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/a_27_47# 0 0.18fF
C4078 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_390_47# 0 0.10fF
C4079 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_283_47# 0 0.18fF
C4080 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/a_27_47# 0 0.18fF
C4081 clock_v2_0/sky130_fd_sc_hd__nand2_1_0/A 0 14.12fF
C4082 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/A 0 22.22fF
C4083 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_390_47# 0 0.10fF
C4084 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_283_47# 0 0.18fF
C4085 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_68/a_27_47# 0 0.18fF
C4086 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_15/X 0 19.84fF
C4087 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_390_47# 0 0.10fF
C4088 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_283_47# 0 0.18fF
C4089 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/a_27_47# 0 0.18fF
C4090 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_390_47# 0 0.10fF
C4091 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_283_47# 0 0.18fF
C4092 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/a_27_47# 0 0.18fF
C4093 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_4/a_110_47# 0 1.28fF
C4094 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/X 0 23.98fF
C4095 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_390_47# 0 0.10fF
C4096 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_283_47# 0 0.18fF
C4097 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_168/a_27_47# 0 0.18fF
C4098 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_149/X 0 25.12fF
C4099 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_390_47# 0 0.10fF
C4100 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_283_47# 0 0.18fF
C4101 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/a_27_47# 0 0.18fF
C4102 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_116/A 0 20.96fF
C4103 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_390_47# 0 0.10fF
C4104 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_283_47# 0 0.18fF
C4105 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_113/a_27_47# 0 0.18fF
C4106 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_103/A 0 17.65fF
C4107 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_390_47# 0 0.10fF
C4108 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_283_47# 0 0.18fF
C4109 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/a_27_47# 0 0.18fF
C4110 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/X 0 19.62fF
C4111 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_390_47# 0 0.10fF
C4112 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_283_47# 0 0.18fF
C4113 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/a_27_47# 0 0.18fF
C4114 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/A 0 10.32fF
C4115 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_390_47# 0 0.10fF
C4116 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_283_47# 0 0.18fF
C4117 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_89/a_27_47# 0 0.18fF
C4118 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/A 0 20.96fF
C4119 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_390_47# 0 0.10fF
C4120 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_283_47# 0 0.18fF
C4121 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_78/a_27_47# 0 0.18fF
C4122 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/X 0 14.05fF
C4123 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_390_47# 0 0.10fF
C4124 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_283_47# 0 0.18fF
C4125 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/a_27_47# 0 0.18fF
C4126 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_36/X 0 26.37fF
C4127 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_390_47# 0 0.10fF
C4128 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_283_47# 0 0.18fF
C4129 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/a_27_47# 0 0.18fF
C4130 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_58/X 0 20.09fF
C4131 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_390_47# 0 0.10fF
C4132 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_283_47# 0 0.18fF
C4133 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/a_27_47# 0 0.18fF
C4134 clock_v2_0/sky130_fd_sc_hd__clkinv_4_2/Y 0 38.00fF
C4135 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_3/a_110_47# 0 1.28fF
C4136 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_136/A 0 21.63fF
C4137 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_390_47# 0 0.10fF
C4138 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_283_47# 0 0.18fF
C4139 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/a_27_47# 0 0.18fF
C4140 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/A 0 14.02fF
C4141 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_125/X 0 24.11fF
C4142 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_390_47# 0 0.10fF
C4143 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_283_47# 0 0.18fF
C4144 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_123/a_27_47# 0 0.18fF
C4145 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_102/A 0 19.11fF
C4146 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_390_47# 0 0.10fF
C4147 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_283_47# 0 0.18fF
C4148 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/a_27_47# 0 0.18fF
C4149 clock_v2_0/sky130_fd_sc_hd__clkinv_4_8/Y 0 10.67fF
C4150 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_390_47# 0 0.10fF
C4151 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_283_47# 0 0.18fF
C4152 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_112/a_27_47# 0 0.18fF
C4153 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_390_47# 0 0.10fF
C4154 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_283_47# 0 0.18fF
C4155 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/a_27_47# 0 0.18fF
C4156 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/A 0 20.98fF
C4157 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/X 0 19.85fF
C4158 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_390_47# 0 0.10fF
C4159 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_283_47# 0 0.18fF
C4160 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_178/a_27_47# 0 0.18fF
C4161 clock_v2_0/sky130_fd_sc_hd__clkinv_4_3/Y 0 42.59fF
C4162 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_390_47# 0 0.10fF
C4163 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_283_47# 0 0.18fF
C4164 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/a_27_47# 0 0.18fF
C4165 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_390_47# 0 0.10fF
C4166 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_283_47# 0 0.18fF
C4167 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/a_27_47# 0 0.18fF
C4168 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_13/X 0 10.16fF
C4169 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_390_47# 0 0.10fF
C4170 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_283_47# 0 0.18fF
C4171 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_11/a_27_47# 0 0.18fF
C4172 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/X 0 35.47fF
C4173 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/A 0 20.02fF
C4174 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_390_47# 0 0.10fF
C4175 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_283_47# 0 0.18fF
C4176 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_44/a_27_47# 0 0.18fF
C4177 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_24/A 0 37.08fF
C4178 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_390_47# 0 0.10fF
C4179 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_283_47# 0 0.18fF
C4180 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/a_27_47# 0 0.18fF
C4181 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/Y 0 57.51fF
C4182 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_2/a_110_47# 0 1.28fF
C4183 clock_v2_0/sky130_fd_sc_hd__nand2_1_4/B 0 35.76fF
C4184 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/X 0 22.22fF
C4185 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_390_47# 0 0.10fF
C4186 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_283_47# 0 0.18fF
C4187 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_122/a_27_47# 0 0.18fF
C4188 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_101/A 0 6.80fF
C4189 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_390_47# 0 0.10fF
C4190 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_283_47# 0 0.18fF
C4191 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_100/a_27_47# 0 0.18fF
C4192 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/X 0 14.09fF
C4193 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_390_47# 0 0.10fF
C4194 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_283_47# 0 0.18fF
C4195 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/a_27_47# 0 0.18fF
C4196 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/B 0 72.22fF
C4197 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_390_47# 0 0.10fF
C4198 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_283_47# 0 0.18fF
C4199 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/a_27_47# 0 0.18fF
C4200 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/X 0 19.55fF
C4201 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/X 0 18.97fF
C4202 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_390_47# 0 0.10fF
C4203 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_283_47# 0 0.18fF
C4204 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_87/a_27_47# 0 0.18fF
C4205 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_67/A 0 24.50fF
C4206 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_390_47# 0 0.10fF
C4207 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_283_47# 0 0.18fF
C4208 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/a_27_47# 0 0.18fF
C4209 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_34/X 0 49.77fF
C4210 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_390_47# 0 0.10fF
C4211 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_283_47# 0 0.18fF
C4212 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_32/a_27_47# 0 0.18fF
C4213 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_56/X 0 13.06fF
C4214 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_390_47# 0 0.10fF
C4215 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_283_47# 0 0.18fF
C4216 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/a_27_47# 0 0.18fF
C4217 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/X 0 25.45fF
C4218 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_390_47# 0 0.10fF
C4219 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_283_47# 0 0.18fF
C4220 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_10/a_27_47# 0 0.18fF
C4221 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_1/a_110_47# 0 1.28fF
C4222 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/X 0 34.14fF
C4223 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_390_47# 0 0.10fF
C4224 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_283_47# 0 0.18fF
C4225 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/a_27_47# 0 0.18fF
C4226 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_134/A 0 20.97fF
C4227 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_390_47# 0 0.10fF
C4228 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_283_47# 0 0.18fF
C4229 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_132/a_27_47# 0 0.18fF
C4230 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/A 0 14.13fF
C4231 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_390_47# 0 0.10fF
C4232 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_283_47# 0 0.18fF
C4233 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_121/a_27_47# 0 0.18fF
C4234 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/X 0 13.78fF
C4235 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_390_47# 0 0.10fF
C4236 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_283_47# 0 0.18fF
C4237 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_187/a_27_47# 0 0.18fF
C4238 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_199/A 0 23.62fF
C4239 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/A 0 25.28fF
C4240 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_390_47# 0 0.10fF
C4241 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_283_47# 0 0.18fF
C4242 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_198/a_27_47# 0 0.18fF
C4243 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/B 0 72.14fF
C4244 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_390_47# 0 0.10fF
C4245 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_283_47# 0 0.18fF
C4246 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/a_27_47# 0 0.18fF
C4247 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/X 0 14.10fF
C4248 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_390_47# 0 0.10fF
C4249 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_283_47# 0 0.18fF
C4250 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/a_27_47# 0 0.18fF
C4251 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_77/X 0 19.67fF
C4252 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_390_47# 0 0.10fF
C4253 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_283_47# 0 0.18fF
C4254 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/a_27_47# 0 0.18fF
C4255 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_390_47# 0 0.10fF
C4256 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_283_47# 0 0.18fF
C4257 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_31/a_27_47# 0 0.18fF
C4258 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_22/A 0 34.83fF
C4259 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_390_47# 0 0.10fF
C4260 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_283_47# 0 0.18fF
C4261 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_20/a_27_47# 0 0.18fF
C4262 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/A 0 9.76fF
C4263 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_390_47# 0 0.10fF
C4264 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_283_47# 0 0.18fF
C4265 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_42/a_27_47# 0 0.18fF
C4266 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_0/a_110_47# 0 1.28fF
C4267 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_147/X 0 37.51fF
C4268 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_390_47# 0 0.10fF
C4269 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_283_47# 0 0.18fF
C4270 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_142/a_27_47# 0 0.18fF
C4271 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_390_47# 0 0.10fF
C4272 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_283_47# 0 0.18fF
C4273 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_131/a_27_47# 0 0.18fF
C4274 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_167/A 0 49.51fF
C4275 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_390_47# 0 0.10fF
C4276 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_283_47# 0 0.18fF
C4277 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/a_27_47# 0 0.18fF
C4278 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_390_47# 0 0.10fF
C4279 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_283_47# 0 0.18fF
C4280 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/a_27_47# 0 0.18fF
C4281 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_390_47# 0 0.10fF
C4282 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_283_47# 0 0.18fF
C4283 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/a_27_47# 0 0.18fF
C4284 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_99/X 0 39.94fF
C4285 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_390_47# 0 0.10fF
C4286 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_283_47# 0 0.18fF
C4287 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/a_27_47# 0 0.18fF
C4288 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_65/A 0 20.22fF
C4289 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_390_47# 0 0.10fF
C4290 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_283_47# 0 0.18fF
C4291 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/a_27_47# 0 0.18fF
C4292 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_54/X 0 25.14fF
C4293 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_390_47# 0 0.10fF
C4294 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_283_47# 0 0.18fF
C4295 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/a_27_47# 0 0.18fF
C4296 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_164/A 0 41.94fF
C4297 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_390_47# 0 0.10fF
C4298 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_283_47# 0 0.18fF
C4299 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/a_27_47# 0 0.18fF
C4300 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_157/X 0 19.63fF
C4301 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_390_47# 0 0.10fF
C4302 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_283_47# 0 0.18fF
C4303 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_152/a_27_47# 0 0.18fF
C4304 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_177/X 0 19.54fF
C4305 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_390_47# 0 0.10fF
C4306 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_283_47# 0 0.18fF
C4307 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/a_27_47# 0 0.18fF
C4308 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_197/A 0 10.74fF
C4309 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/Y 0 32.17fF
C4310 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_390_47# 0 0.10fF
C4311 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_283_47# 0 0.18fF
C4312 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_196/a_27_47# 0 0.18fF
C4313 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_169/A 0 22.16fF
C4314 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_146/X 0 23.14fF
C4315 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_390_47# 0 0.10fF
C4316 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_283_47# 0 0.18fF
C4317 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_141/a_27_47# 0 0.18fF
C4318 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_97/A 0 23.54fF
C4319 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_390_47# 0 0.10fF
C4320 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_283_47# 0 0.18fF
C4321 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/a_27_47# 0 0.18fF
C4322 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_86/A 0 22.79fF
C4323 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_390_47# 0 0.10fF
C4324 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_283_47# 0 0.18fF
C4325 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/a_27_47# 0 0.18fF
C4326 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_75/X 0 19.99fF
C4327 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_390_47# 0 0.10fF
C4328 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_283_47# 0 0.18fF
C4329 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/a_27_47# 0 0.18fF
C4330 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_163/A 0 43.11fF
C4331 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_390_47# 0 0.10fF
C4332 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_283_47# 0 0.18fF
C4333 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_162/a_27_47# 0 0.18fF
C4334 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_158/A 0 20.10fF
C4335 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_390_47# 0 0.10fF
C4336 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_283_47# 0 0.18fF
C4337 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_140/a_27_47# 0 0.18fF
C4338 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_174/X 0 19.84fF
C4339 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_390_47# 0 0.10fF
C4340 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_283_47# 0 0.18fF
C4341 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/a_27_47# 0 0.18fF
C4342 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_186/A 0 22.78fF
C4343 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_390_47# 0 0.10fF
C4344 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_283_47# 0 0.18fF
C4345 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/a_27_47# 0 0.18fF
C4346 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_390_47# 0 0.10fF
C4347 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_283_47# 0 0.18fF
C4348 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/a_27_47# 0 0.18fF
C4349 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/D 0 7.57fF
C4350 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_381_47# 0 0.03fF
C4351 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1490_369# 0 0.09fF
C4352 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_891_413# 0 0.12fF
C4353 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_1059_315# 0 0.24fF
C4354 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_466_413# 0 0.11fF
C4355 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_634_159# 0 0.12fF
C4356 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_193_47# 0 0.21fF
C4357 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_1/a_27_47# 0 0.31fF
C4358 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_63/A 0 21.63fF
C4359 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_390_47# 0 0.10fF
C4360 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_283_47# 0 0.18fF
C4361 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_61/a_27_47# 0 0.18fF
C4362 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_52/X 0 22.67fF
C4363 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_390_47# 0 0.10fF
C4364 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_283_47# 0 0.18fF
C4365 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_50/a_27_47# 0 0.18fF
C4366 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_154/X 0 21.74fF
C4367 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_390_47# 0 0.10fF
C4368 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_283_47# 0 0.18fF
C4369 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_150/a_27_47# 0 0.18fF
C4370 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_173/X 0 10.16fF
C4371 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_390_47# 0 0.10fF
C4372 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_283_47# 0 0.18fF
C4373 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_172/a_27_47# 0 0.18fF
C4374 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/Q_N 0 0.05fF
C4375 clock_v2_0/sky130_fd_sc_hd__nand2_1_1/A 0 44.99fF
C4376 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_381_47# 0 0.03fF
C4377 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1490_369# 0 0.09fF
C4378 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_891_413# 0 0.12fF
C4379 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_1059_315# 0 0.24fF
C4380 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_466_413# 0 0.11fF
C4381 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_634_159# 0 0.12fF
C4382 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_193_47# 0 0.21fF
C4383 clock_v2_0/sky130_fd_sc_hd__dfxbp_1_0/a_27_47# 0 0.31fF
C4384 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_95/A 0 25.21fF
C4385 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_390_47# 0 0.10fF
C4386 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_283_47# 0 0.18fF
C4387 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_93/a_27_47# 0 0.18fF
C4388 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_84/A 0 20.21fF
C4389 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_390_47# 0 0.10fF
C4390 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_283_47# 0 0.18fF
C4391 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/a_27_47# 0 0.18fF
C4392 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_73/X 0 10.28fF
C4393 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_390_47# 0 0.10fF
C4394 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_283_47# 0 0.18fF
C4395 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_71/a_27_47# 0 0.18fF
C4396 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_184/A 0 20.18fF
C4397 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_390_47# 0 0.10fF
C4398 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_283_47# 0 0.18fF
C4399 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/a_27_47# 0 0.18fF
C4400 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_195/X 0 33.91fF
C4401 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_390_47# 0 0.10fF
C4402 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_283_47# 0 0.18fF
C4403 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/a_27_47# 0 0.18fF
C4404 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/Y 0 106.51fF
C4405 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_96/X 0 40.72fF
C4406 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_390_47# 0 0.10fF
C4407 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_283_47# 0 0.18fF
C4408 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/a_27_47# 0 0.18fF
C4409 VDD 0 -38260.64fF
C4410 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_82/A 0 14.35fF
C4411 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_390_47# 0 0.10fF
C4412 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_283_47# 0 0.18fF
C4413 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_80/a_27_47# 0 0.18fF
C4414 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_182/A 0 14.37fF
C4415 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_390_47# 0 0.10fF
C4416 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_283_47# 0 0.18fF
C4417 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_180/a_27_47# 0 0.18fF
C4418 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_193/X 0 34.61fF
C4419 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_390_47# 0 0.10fF
C4420 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_283_47# 0 0.18fF
C4421 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/a_27_47# 0 0.18fF
C4422 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_92/X 0 50.29fF
C4423 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_390_47# 0 0.10fF
C4424 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_283_47# 0 0.18fF
C4425 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_90/a_27_47# 0 0.18fF
C4426 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_191/X 0 42.28fF
C4427 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_390_47# 0 0.10fF
C4428 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_283_47# 0 0.18fF
C4429 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_190/a_27_47# 0 0.18fF
C4430 clock_v2_0/sky130_fd_sc_hd__clkinv_4_7/A 0 69.53fF
C4431 clock_v2_0/sky130_fd_sc_hd__clkinv_4_5/Y 0 107.06fF
C4432 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/A 0 19.99fF
C4433 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_390_47# 0 0.10fF
C4434 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_283_47# 0 0.18fF
C4435 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_8/a_27_47# 0 0.18fF
C4436 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/Y 0 58.90fF
C4437 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/A 0 19.81fF
C4438 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_390_47# 0 0.10fF
C4439 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_283_47# 0 0.18fF
C4440 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_6/a_27_47# 0 0.18fF
C4441 clock_v2_0/sky130_fd_sc_hd__nand2_4_3/a_27_47# 0 0.06fF
C4442 clock_v2_0/sky130_fd_sc_hd__clkinv_4_1/A 0 117.01fF
C4443 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_390_47# 0 0.10fF
C4444 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_283_47# 0 0.18fF
C4445 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_5/a_27_47# 0 0.18fF
C4446 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/Y 0 58.46fF
C4447 clock_v2_0/sky130_fd_sc_hd__nand2_4_2/a_27_47# 0 0.06fF
C4448 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/Y 0 60.89fF
C4449 clock_v2_0/sky130_fd_sc_hd__nand2_4_1/a_27_47# 0 0.06fF
C4450 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/B 0 72.21fF
C4451 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_390_47# 0 0.10fF
C4452 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_283_47# 0 0.18fF
C4453 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/a_27_47# 0 0.18fF
C4454 clock_v2_0/sky130_fd_sc_hd__nand2_4_0/a_27_47# 0 0.06fF
C4455 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_3/A 0 23.61fF
C4456 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/A 0 25.28fF
C4457 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_390_47# 0 0.10fF
C4458 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_283_47# 0 0.18fF
C4459 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_2/a_27_47# 0 0.18fF
C4460 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_15/a_110_47# 0 1.28fF
C4461 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_390_47# 0 0.10fF
C4462 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_283_47# 0 0.18fF
C4463 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/a_27_47# 0 0.18fF
C4464 clock_v2_0/sky130_fd_sc_hd__clkinv_1_3/A 0 90.21fF
C4465 clock_v2_0/sky130_fd_sc_hd__clkinv_4_10/Y 0 28.47fF
C4466 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_14/a_110_47# 0 1.28fF
C4467 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_1/A 0 10.73fF
C4468 clock_v2_0/sky130_fd_sc_hd__clkinv_1_0/Y 0 32.17fF
C4469 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_390_47# 0 0.10fF
C4470 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_283_47# 0 0.18fF
C4471 clock_v2_0/sky130_fd_sc_hd__clkdlybuf4s50_1_0/a_27_47# 0 0.18fF
C4472 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_13/a_110_47# 0 1.28fF
C4473 clock_v2_0/sky130_fd_sc_hd__clkinv_4_9/Y 0 74.50fF
C4474 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_12/a_110_47# 0 1.28fF
C4475 clock_v2_0/sky130_fd_sc_hd__clkbuf_16_11/a_110_47# 0 1.28fF
C4476 sky130_fd_pr__cap_mim_m3_1_CEWQ64_18/m3_n360_n310# 0 0.63fF
C4477 sky130_fd_sc_hd__mux4_1_3/X 0 52.90fF
C4478 sky130_fd_sc_hd__mux4_1_3/a_834_97# 0 0.02fF
C4479 sky130_fd_sc_hd__mux4_1_3/a_668_97# 0 0.03fF
C4480 sky130_fd_sc_hd__mux4_1_3/a_27_47# 0 0.03fF
C4481 sky130_fd_sc_hd__mux4_1_3/a_1478_413# 0 0.11fF
C4482 sky130_fd_sc_hd__mux4_1_3/a_1290_413# 0 0.15fF
C4483 sky130_fd_sc_hd__mux4_1_3/a_750_97# 0 0.03fF
C4484 sky130_fd_sc_hd__mux4_1_3/a_277_47# 0 0.07fF
C4485 sky130_fd_sc_hd__mux4_1_3/a_247_21# 0 0.27fF
C4486 transmission_gate_0/out 0 3.97fF
C4487 ip 0 8.23fF
C4488 sky130_fd_pr__cap_mim_m3_1_CGPBWM_4/m3_n1030_n980# 0 2.84fF
C4489 sky130_fd_pr__cap_mim_m3_1_CEWQ64_38/m3_n360_n310# 0 0.63fF
C4490 sky130_fd_pr__cap_mim_m3_1_CEWQ64_49/m3_n360_n310# 0 0.63fF
C4491 sky130_fd_pr__cap_mim_m3_1_CEWQ64_27/m3_n360_n310# 0 0.63fF
C4492 sky130_fd_sc_hd__mux4_1_2/X 0 26.26fF
C4493 d_clk_grp_1_ctrl_1 0 19.38fF
C4494 d_clk_grp_1_ctrl_0 0 20.35fF
C4495 sky130_fd_sc_hd__mux4_1_2/a_834_97# 0 0.02fF
C4496 sky130_fd_sc_hd__mux4_1_2/a_668_97# 0 0.03fF
C4497 sky130_fd_sc_hd__mux4_1_2/a_27_47# 0 0.03fF
C4498 sky130_fd_sc_hd__mux4_1_2/a_1478_413# 0 0.11fF
C4499 sky130_fd_sc_hd__mux4_1_2/a_1290_413# 0 0.15fF
C4500 sky130_fd_sc_hd__mux4_1_2/a_750_97# 0 0.03fF
C4501 sky130_fd_sc_hd__mux4_1_2/a_277_47# 0 0.07fF
C4502 sky130_fd_sc_hd__mux4_1_2/a_247_21# 0 0.27fF
C4503 sky130_fd_pr__cap_mim_m3_1_CEWQ64_37/m3_n360_n310# 0 0.63fF
C4504 sky130_fd_pr__cap_mim_m3_1_CGPBWM_3/m3_n1030_n980# 0 2.84fF
C4505 sky130_fd_pr__cap_mim_m3_1_CEWQ64_15/m3_n360_n310# 0 0.63fF
C4506 sky130_fd_pr__cap_mim_m3_1_CEWQ64_26/m3_n360_n310# 0 0.63fF
C4507 sky130_fd_sc_hd__mux4_1_1/X 0 26.31fF
C4508 sky130_fd_sc_hd__mux4_1_1/a_834_97# 0 0.02fF
C4509 sky130_fd_sc_hd__mux4_1_1/a_668_97# 0 0.03fF
C4510 sky130_fd_sc_hd__mux4_1_1/a_27_47# 0 0.03fF
C4511 sky130_fd_sc_hd__mux4_1_1/a_1478_413# 0 0.11fF
C4512 sky130_fd_sc_hd__mux4_1_1/a_1290_413# 0 0.15fF
C4513 sky130_fd_sc_hd__mux4_1_1/a_750_97# 0 0.03fF
C4514 sky130_fd_sc_hd__mux4_1_1/a_277_47# 0 0.07fF
C4515 sky130_fd_sc_hd__mux4_1_1/a_247_21# 0 0.27fF
C4516 sky130_fd_pr__cap_mim_m3_1_CGPBWM_2/m3_n1030_n980# 0 2.84fF
C4517 sky130_fd_pr__cap_mim_m3_1_CEWQ64_36/m3_n360_n310# 0 0.63fF
C4518 sky130_fd_pr__cap_mim_m3_1_CEWQ64_14/m3_n360_n310# 0 0.63fF
C4519 sky130_fd_pr__cap_mim_m3_1_CEWQ64_47/m3_n360_n310# 0 0.63fF
C4520 sky130_fd_pr__cap_mim_m3_1_CEWQ64_69/m3_n360_n310# 0 0.63fF
C4521 sky130_fd_sc_hd__mux4_1_0/X 0 26.26fF
C4522 d_clk_grp_2_ctrl_1 0 17.02fF
C4523 d_clk_grp_2_ctrl_0 0 17.69fF
C4524 sky130_fd_sc_hd__mux4_1_0/a_834_97# 0 0.02fF
C4525 sky130_fd_sc_hd__mux4_1_0/a_668_97# 0 0.03fF
C4526 sky130_fd_sc_hd__mux4_1_0/a_27_47# 0 0.03fF
C4527 sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0 0.11fF
C4528 sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0 0.15fF
C4529 sky130_fd_sc_hd__mux4_1_0/a_750_97# 0 0.03fF
C4530 sky130_fd_sc_hd__mux4_1_0/a_277_47# 0 0.07fF
C4531 sky130_fd_sc_hd__mux4_1_0/a_247_21# 0 0.27fF
C4532 a_mux2_en_1/switch_5t_0/in 0 1.63fF
C4533 a_mux2_en_1/transmission_gate_1/en_b 0 0.82fF
C4534 a_mux2_en_1/switch_5t_1/in 0 0.73fF
C4535 a_mux2_en_1/switch_5t_1/en 0 7.11fF
C4536 a_probe_1 0 -6.88fF
C4537 a_mux2_en_1/switch_5t_1/transmission_gate_1/in 0 1.77fF
C4538 a_mux2_en_1/switch_5t_0/transmission_gate_1/in 0 1.77fF
C4539 sky130_fd_pr__cap_mim_m3_1_CEWQ64_35/m3_n360_n310# 0 0.63fF
C4540 onebit_dac_1/out 0 -4.96fF
C4541 sky130_fd_pr__cap_mim_m3_1_CGPBWM_1/m3_n1030_n980# 0 2.84fF
C4542 sky130_fd_pr__cap_mim_m3_1_CEWQ64_24/m3_n360_n310# 0 0.63fF
C4543 sky130_fd_pr__cap_mim_m3_1_CEWQ64_46/m3_n360_n310# 0 0.63fF
C4544 a_mux2_en_0/switch_5t_0/in 0 1.63fF
C4545 a_mux2_en_0/transmission_gate_1/en_b 0 0.82fF
C4546 a_mux2_en_0/switch_5t_1/in 0 0.73fF
C4547 a_mux2_en_0/switch_5t_1/en 0 7.11fF
C4548 a_probe_0 0 -1.47fF
C4549 a_mod_grp_ctrl_0 0 110.64fF
C4550 a_mux2_en_0/switch_5t_1/transmission_gate_1/in 0 1.77fF
C4551 a_mux2_en_0/switch_5t_0/transmission_gate_1/in 0 1.77fF
C4552 ota_1/m1_1038_n2886# 0 -76.00fF
C4553 ota_1/m1_n208_n2883# 0 -83.42fF
C4554 ota_1/m1_n6302_n3889# 0 10.46fF
C4555 ota_1/m1_2463_n5585# 0 0.31fF
C4556 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0 1.37fF
C4557 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# 0 1.37fF
C4558 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0 1.37fF
C4559 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# 0 1.37fF
C4560 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# 0 1.37fF
C4561 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0 1.37fF
C4562 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# 0 1.37fF
C4563 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# 0 1.37fF
C4564 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# 0 1.37fF
C4565 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0 1.37fF
C4566 ota_1/sc_cmfb_0/transmission_gate_9/in 0 -27.99fF
C4567 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# 0 1.37fF
C4568 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# 0 1.37fF
C4569 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# 0 1.37fF
C4570 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0 1.37fF
C4571 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0 1.37fF
C4572 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# 0 1.37fF
C4573 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0 1.37fF
C4574 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# 0 1.37fF
C4575 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0 1.37fF
C4576 ota_1/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0 1.37fF
C4577 ota_1/sc_cmfb_0/transmission_gate_8/in 0 -0.42fF
C4578 ota_1/sc_cmfb_0/transmission_gate_6/in 0 2.41fF
C4579 ota_1/sc_cmfb_0/transmission_gate_7/in 0 1.91fF
C4580 ota_1/cm 0 -36.78fF
C4581 ota_1/sc_cmfb_0/transmission_gate_4/out 0 0.84fF
C4582 ota_1/sc_cmfb_0/transmission_gate_3/out 0 -4.68fF
C4583 ota_1/m1_2462_n3318# 0 -13.18fF
C4584 ota_1/m1_12410_n11263# 0 0.16fF
C4585 ota_1/m1_12118_n11263# 0 0.30fF
C4586 ota_1/m1_11826_n11260# 0 0.32fF
C4587 ota_1/m1_11534_n11258# 0 0.23fF
C4588 ota_1/m1_11244_n11260# 0 0.24fF
C4589 ota_1/m1_12232_n10488# 0 0.22fF
C4590 ota_1/m1_11940_n10482# 0 0.34fF
C4591 ota_1/m1_11648_n10486# 0 0.25fF
C4592 ota_1/m1_11356_n10481# 0 0.26fF
C4593 ota_1/m1_11063_n10490# 0 0.26fF
C4594 ota_1/m1_12410_n9718# 0 0.16fF
C4595 ota_1/m1_12118_n9704# 0 0.27fF
C4596 ota_1/m1_11825_n9711# 0 0.29fF
C4597 ota_1/m1_11534_n9706# 0 0.22fF
C4598 ota_1/m1_11242_n9716# 0 0.23fF
C4599 ota_1/cmc 0 1.10fF
C4600 ota_1/bias_a 0 -298.49fF
C4601 ota_1/m1_n5574_n13620# 0 183.14fF
C4602 ota_1/m1_6690_n8907# 0 -73.84fF
C4603 ota_1/bias_c 0 43.28fF
C4604 i_bias_2 0 -23.49fF
C4605 ota_1/m1_n1659_n11581# 0 3.21fF
C4606 ota_1/m1_n947_n12836# 0 7.99fF
C4607 ota_1/m1_n2176_n12171# 0 12.82fF
C4608 ota_1/bias_d 0 119.38fF
C4609 ota_1/bias_b 0 12.75fF
C4610 transmission_gate_19/in 0 3.38fF
C4611 sky130_fd_pr__cap_mim_m3_1_CGPBWM_0/m3_n1030_n980# 0 2.84fF
C4612 onebit_dac_1/v_b 0 30.49fF
C4613 onebit_dac_0/out 0 -1.49fF
C4614 op 0 30.01fF
C4615 sky130_fd_pr__cap_mim_m3_1_CEWQ64_56/m3_n360_n310# 0 0.63fF
C4616 ota_1/ip 0 13.86fF
C4617 sky130_fd_pr__cap_mim_m3_1_CEWQ64_45/m3_n360_n310# 0 0.63fF
C4618 transmission_gate_19/out 0 -6.85fF
C4619 sky130_fd_pr__cap_mim_m3_1_CEWQ64_33/m3_n360_n310# 0 0.63fF
C4620 sky130_fd_pr__cap_mim_m3_1_CEWQ64_55/m3_n360_n310# 0 0.63fF
C4621 transmission_gate_17/in 0 -4.37fF
C4622 transmission_gate_18/in 0 13.53fF
C4623 sky130_fd_pr__cap_mim_m3_1_CEWQ64_9/m3_n360_n310# 0 0.63fF
C4624 sky130_fd_pr__cap_mim_m3_1_CEWQ64_32/m3_n360_n310# 0 0.63fF
C4625 sky130_fd_pr__cap_mim_m3_1_CEWQ64_65/m3_n360_n310# 0 0.63fF
C4626 d_probe_0 0 -41.93fF
C4627 sky130_fd_sc_hd__clkinv_4_4/Y 0 26.71fF
C4628 sky130_fd_pr__cap_mim_m3_1_CEWQ64_8/m3_n360_n310# 0 0.63fF
C4629 sky130_fd_pr__cap_mim_m3_1_CEWQ64_53/m3_n360_n310# 0 0.63fF
C4630 sky130_fd_pr__cap_mim_m3_1_CEWQ64_42/m3_n360_n310# 0 0.63fF
C4631 d_probe_1 0 -42.67fF
C4632 sky130_fd_sc_hd__clkinv_4_3/Y 0 13.72fF
C4633 sky130_fd_pr__cap_mim_m3_1_CEWQ64_7/m3_n360_n310# 0 0.63fF
C4634 sky130_fd_pr__cap_mim_m3_1_CEWQ64_41/m3_n360_n310# 0 0.63fF
C4635 sky130_fd_pr__cap_mim_m3_1_CEWQ64_52/m3_n360_n310# 0 0.63fF
C4636 d_probe_2 0 -39.34fF
C4637 sky130_fd_sc_hd__clkinv_4_2/Y 0 13.89fF
C4638 clock_v2_0/Bd 0 46.97fF
C4639 clock_v2_0/Bd_b 0 71.54fF
C4640 sky130_fd_pr__cap_mim_m3_1_CEWQ64_6/m3_n360_n310# 0 0.63fF
C4641 ota_1/in 0 20.14fF
C4642 sky130_fd_pr__cap_mim_m3_1_CEWQ64_51/m3_n360_n310# 0 0.63fF
C4643 d_probe_3 0 -38.10fF
C4644 sky130_fd_sc_hd__clkinv_4_1/Y 0 13.72fF
C4645 clock_v2_0/Ad 0 37.43fF
C4646 clock_v2_0/Ad_b 0 68.98fF
C4647 sky130_fd_pr__cap_mim_m3_1_CEWQ64_5/m3_n360_n310# 0 0.63fF
C4648 sky130_fd_pr__cap_mim_m3_1_CEWQ64_50/m3_n360_n310# 0 0.63fF
C4649 ota_w_test_0/m1_1038_n2886# 0 -76.00fF
C4650 ota_w_test_0/m1_n208_n2883# 0 -83.42fF
C4651 ota_w_test_0/m1_n2176_n12171# 0 12.82fF
C4652 a_mux4_en_0/in2 0 116.58fF
C4653 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_19/m3_n630_n580# 0 1.37fF
C4654 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_18/m3_n630_n580# 0 1.37fF
C4655 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_29/m3_n630_n580# 0 1.37fF
C4656 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_17/m3_n630_n580# 0 1.37fF
C4657 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_28/m3_n630_n580# 0 1.37fF
C4658 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_16/m3_n630_n580# 0 1.37fF
C4659 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_27/m3_n630_n580# 0 1.37fF
C4660 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_26/m3_n630_n580# 0 1.37fF
C4661 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_25/m3_n630_n580# 0 1.37fF
C4662 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_35/m3_n630_n580# 0 1.37fF
C4663 ota_w_test_0/sc_cmfb_0/transmission_gate_9/in 0 -27.99fF
C4664 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_24/m3_n630_n580# 0 1.37fF
C4665 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_33/m3_n630_n580# 0 1.37fF
C4666 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_34/m3_n630_n580# 0 1.37fF
C4667 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_23/m3_n630_n580# 0 1.37fF
C4668 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_22/m3_n630_n580# 0 1.37fF
C4669 ota_1/p2 0 70.38fF
C4670 ota_1/p2_b 0 16.61fF
C4671 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_32/m3_n630_n580# 0 1.37fF
C4672 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_21/m3_n630_n580# 0 1.37fF
C4673 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_31/m3_n630_n580# 0 1.37fF
C4674 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_20/m3_n630_n580# 0 1.37fF
C4675 ota_w_test_0/sc_cmfb_0/unit_cap_mim_m3m4_30/m3_n630_n580# 0 1.37fF
C4676 ota_w_test_0/sc_cmfb_0/transmission_gate_8/in 0 -0.42fF
C4677 ota_w_test_0/sc_cmfb_0/transmission_gate_6/in 0 2.41fF
C4678 ota_w_test_0/sc_cmfb_0/transmission_gate_7/in 0 1.91fF
C4679 ota_w_test_0/cm 0 -8.72fF
C4680 ota_1/p1 0 -12.50fF
C4681 ota_w_test_0/op 0 -2.79fF
C4682 ota_w_test_0/sc_cmfb_0/transmission_gate_4/out 0 0.84fF
C4683 ota_w_test_0/on 0 -63.99fF
C4684 ota_w_test_0/sc_cmfb_0/transmission_gate_3/out 0 -4.68fF
C4685 ota_w_test_0/m1_12410_n11263# 0 0.16fF
C4686 ota_w_test_0/m1_12118_n11263# 0 0.30fF
C4687 ota_w_test_0/m1_11826_n11260# 0 0.32fF
C4688 ota_w_test_0/m1_11534_n11258# 0 0.23fF
C4689 ota_w_test_0/m1_11244_n11260# 0 0.24fF
C4690 ota_w_test_0/m1_12232_n10488# 0 0.22fF
C4691 ota_w_test_0/m1_11940_n10482# 0 0.34fF
C4692 ota_w_test_0/m1_11648_n10486# 0 0.25fF
C4693 ota_w_test_0/m1_11356_n10481# 0 0.26fF
C4694 ota_w_test_0/m1_11063_n10490# 0 0.26fF
C4695 a_mux4_en_1/in1 0 12.23fF
C4696 ota_w_test_0/m1_12410_n9718# 0 0.16fF
C4697 ota_w_test_0/m1_12118_n9704# 0 0.27fF
C4698 ota_w_test_0/m1_11825_n9711# 0 0.29fF
C4699 ota_w_test_0/m1_11534_n9706# 0 0.22fF
C4700 ota_w_test_0/m1_11242_n9716# 0 0.23fF
C4701 ota_w_test_0/m1_6690_n8907# 0 -73.84fF
C4702 ota_w_test_0/m1_2462_n3318# 0 -13.18fF
C4703 a_mux4_en_0/in1 0 61.18fF
C4704 VSS 0 -37531.12fF
C4705 i_bias_1 0 -16.95fF
C4706 ota_w_test_0/m1_n5574_n13620# 0 183.14fF
C4707 a_mux4_en_0/in0 0 -291.59fF
C4708 a_mux4_en_1/in2 0 7.25fF
C4709 ota_w_test_0/m1_2463_n5585# 0 0.31fF
C4710 ota_w_test_0/m1_n1659_n11581# 0 3.21fF
C4711 ota_w_test_0/m1_n947_n12836# 0 7.99fF
C4712 ota_w_test_0/m1_n6302_n3889# 0 10.46fF
C4713 transmission_gate_26/en 0 30.18fF
C4714 rst_n 0 49.56fF
C4715 transmission_gate_23/in 0 -0.20fF
C4716 sky130_fd_pr__cap_mim_m3_1_CEWQ64_4/m3_n360_n310# 0 0.63fF
C4717 sky130_fd_pr__cap_mim_m3_1_CEWQ64_71/m3_n360_n310# 0 0.63fF
C4718 transmission_gate_32/out 0 15.70fF
C4719 sky130_fd_pr__cap_mim_m3_1_CEWQ64_3/m3_n360_n310# 0 0.63fF
C4720 sky130_fd_pr__cap_mim_m3_1_CGPBWM_19/m3_n1030_n980# 0 2.84fF
C4721 sky130_fd_pr__cap_mim_m3_1_CEWQ64_70/m3_n360_n310# 0 0.63fF
C4722 transmission_gate_31/out 0 3.48fF
C4723 transmission_gate_21/in 0 -5.23fF
C4724 sky130_fd_pr__cap_mim_m3_1_CGPBWM_29/m3_n1030_n980# 0 2.84fF
C4725 sky130_fd_pr__cap_mim_m3_1_CEWQ64_2/m3_n360_n310# 0 0.63fF
.ends

