* NGSPICE file created from transmission_gate.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_UNG2NQ a_n416_n136# a_352_n136# a_n128_n136# a_n224_n136#
+ a_64_n136# a_160_n136# a_n320_n136# w_n646_n356# a_n32_n136# a_n508_n136# a_448_n136#
+ a_n512_n234# a_256_n136# VSUBS
X0 a_n224_n136# a_n512_n234# a_n320_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X1 a_352_n136# a_n512_n234# a_256_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X2 a_n128_n136# a_n512_n234# a_n224_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X3 a_256_n136# a_n512_n234# a_160_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.488e+11p ps=3.38e+06u w=1.36e+06u l=150000u
X4 a_n416_n136# a_n512_n234# a_n508_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=4.216e+11p ps=3.34e+06u w=1.36e+06u l=150000u
X5 a_n320_n136# a_n512_n234# a_n416_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
X6 a_n32_n136# a_n512_n234# a_n128_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X7 a_448_n136# a_n512_n234# a_352_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.216e+11p pd=3.34e+06u as=0p ps=0u w=1.36e+06u l=150000u
X8 a_64_n136# a_n512_n234# a_n32_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=4.488e+11p pd=3.38e+06u as=0p ps=0u w=1.36e+06u l=150000u
X9 a_160_n136# a_n512_n234# a_64_n136# w_n646_n356# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.36e+06u l=150000u
C0 a_352_n136# a_256_n136# 0.33fF
C1 a_160_n136# a_n224_n136# 0.05fF
C2 a_352_n136# a_n32_n136# 0.05fF
C3 a_64_n136# a_160_n136# 0.33fF
C4 a_n32_n136# a_256_n136# 0.07fF
C5 a_n508_n136# w_n646_n356# 0.13fF
C6 a_n508_n136# a_n512_n234# 0.06fF
C7 a_352_n136# a_448_n136# 0.33fF
C8 a_256_n136# a_448_n136# 0.12fF
C9 a_n32_n136# a_448_n136# 0.04fF
C10 a_n320_n136# a_n508_n136# 0.12fF
C11 a_n128_n136# w_n646_n356# 0.05fF
C12 a_n128_n136# a_n512_n234# 0.06fF
C13 a_n508_n136# a_n416_n136# 0.33fF
C14 w_n646_n356# a_n224_n136# 0.06fF
C15 a_64_n136# w_n646_n356# 0.05fF
C16 a_64_n136# a_n512_n234# 0.06fF
C17 a_n128_n136# a_n320_n136# 0.12fF
C18 a_n128_n136# a_n416_n136# 0.07fF
C19 a_n320_n136# a_n224_n136# 0.33fF
C20 a_n224_n136# a_n416_n136# 0.12fF
C21 a_64_n136# a_n320_n136# 0.05fF
C22 a_352_n136# a_n508_n136# 0.02fF
C23 a_160_n136# w_n646_n356# 0.06fF
C24 a_64_n136# a_n416_n136# 0.04fF
C25 a_256_n136# a_n508_n136# 0.02fF
C26 a_n32_n136# a_n508_n136# 0.04fF
C27 a_352_n136# a_n128_n136# 0.04fF
C28 a_448_n136# a_n508_n136# 0.02fF
C29 a_160_n136# a_n320_n136# 0.04fF
C30 a_352_n136# a_n224_n136# 0.03fF
C31 a_160_n136# a_n416_n136# 0.03fF
C32 a_256_n136# a_n128_n136# 0.05fF
C33 a_256_n136# a_n224_n136# 0.04fF
C34 a_n32_n136# a_n128_n136# 0.33fF
C35 a_352_n136# a_64_n136# 0.07fF
C36 a_n32_n136# a_n224_n136# 0.12fF
C37 a_64_n136# a_256_n136# 0.12fF
C38 w_n646_n356# a_n512_n234# 1.13fF
C39 a_64_n136# a_n32_n136# 0.33fF
C40 a_448_n136# a_n128_n136# 0.03fF
C41 a_448_n136# a_n224_n136# 0.03fF
C42 a_64_n136# a_448_n136# 0.05fF
C43 a_352_n136# a_160_n136# 0.12fF
C44 a_n320_n136# w_n646_n356# 0.06fF
C45 a_n320_n136# a_n512_n234# 0.06fF
C46 a_256_n136# a_160_n136# 0.33fF
C47 w_n646_n356# a_n416_n136# 0.08fF
C48 a_n32_n136# a_160_n136# 0.12fF
C49 a_448_n136# a_160_n136# 0.07fF
C50 a_n320_n136# a_n416_n136# 0.33fF
C51 a_352_n136# w_n646_n356# 0.08fF
C52 a_n128_n136# a_n508_n136# 0.05fF
C53 a_n508_n136# a_n224_n136# 0.07fF
C54 a_256_n136# w_n646_n356# 0.06fF
C55 a_256_n136# a_n512_n234# 0.06fF
C56 a_n32_n136# w_n646_n356# 0.05fF
C57 a_64_n136# a_n508_n136# 0.03fF
C58 a_352_n136# a_n320_n136# 0.03fF
C59 a_448_n136# w_n646_n356# 0.13fF
C60 a_448_n136# a_n512_n234# 0.06fF
C61 a_352_n136# a_n416_n136# 0.02fF
C62 a_n128_n136# a_n224_n136# 0.33fF
C63 a_256_n136# a_n320_n136# 0.03fF
C64 a_256_n136# a_n416_n136# 0.03fF
C65 a_n32_n136# a_n320_n136# 0.07fF
C66 a_64_n136# a_n128_n136# 0.12fF
C67 a_n32_n136# a_n416_n136# 0.05fF
C68 a_160_n136# a_n508_n136# 0.03fF
C69 a_64_n136# a_n224_n136# 0.07fF
C70 a_448_n136# a_n320_n136# 0.02fF
C71 a_448_n136# a_n416_n136# 0.02fF
C72 a_160_n136# a_n128_n136# 0.07fF
C73 w_n646_n356# VSUBS 2.52fF
.ends

.subckt sky130_fd_pr__nfet_01v8_6J4AMR a_256_n52# a_n32_n52# a_n224_n52# a_448_n52#
+ a_n416_n52# a_160_n52# a_n610_n226# a_n128_n52# a_n512_n140# a_352_n52# a_n320_n52#
+ a_n508_n52# a_64_n52#
X0 a_n32_n52# a_n512_n140# a_n128_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X1 a_n416_n52# a_n512_n140# a_n508_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.612e+11p ps=1.66e+06u w=520000u l=150000u
X2 a_n224_n52# a_n512_n140# a_n320_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X3 a_n128_n52# a_n512_n140# a_n224_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_n320_n52# a_n512_n140# a_n416_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X5 a_160_n52# a_n512_n140# a_64_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X6 a_352_n52# a_n512_n140# a_256_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.716e+11p pd=1.7e+06u as=1.716e+11p ps=1.7e+06u w=520000u l=150000u
X7 a_256_n52# a_n512_n140# a_160_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X8 a_448_n52# a_n512_n140# a_352_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=1.612e+11p pd=1.66e+06u as=0p ps=0u w=520000u l=150000u
X9 a_64_n52# a_n512_n140# a_n32_n52# a_n610_n226# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
C0 a_n32_n52# a_448_n52# 0.02fF
C1 a_n32_n52# a_n128_n52# 0.13fF
C2 a_n512_n140# a_n508_n52# 0.09fF
C3 a_448_n52# a_160_n52# 0.03fF
C4 a_448_n52# a_64_n52# 0.02fF
C5 a_448_n52# a_352_n52# 0.13fF
C6 a_n128_n52# a_160_n52# 0.03fF
C7 a_64_n52# a_n128_n52# 0.05fF
C8 a_n128_n52# a_352_n52# 0.02fF
C9 a_448_n52# a_256_n52# 0.05fF
C10 a_n128_n52# a_256_n52# 0.02fF
C11 a_64_n52# a_n512_n140# 0.09fF
C12 a_n512_n140# a_256_n52# 0.09fF
C13 a_n224_n52# a_n320_n52# 0.13fF
C14 a_n416_n52# a_n320_n52# 0.13fF
C15 a_n508_n52# a_n320_n52# 0.05fF
C16 a_448_n52# a_n128_n52# 0.01fF
C17 a_n224_n52# a_n416_n52# 0.05fF
C18 a_n224_n52# a_n508_n52# 0.03fF
C19 a_n32_n52# a_n320_n52# 0.03fF
C20 a_n416_n52# a_n508_n52# 0.13fF
C21 a_n32_n52# a_n224_n52# 0.05fF
C22 a_n320_n52# a_160_n52# 0.02fF
C23 a_448_n52# a_n512_n140# 0.09fF
C24 a_64_n52# a_n320_n52# 0.02fF
C25 a_n320_n52# a_352_n52# 0.01fF
C26 a_n512_n140# a_n128_n52# 0.09fF
C27 a_n224_n52# a_160_n52# 0.02fF
C28 a_64_n52# a_n224_n52# 0.03fF
C29 a_n224_n52# a_352_n52# 0.01fF
C30 a_n320_n52# a_256_n52# 0.01fF
C31 a_n32_n52# a_n416_n52# 0.02fF
C32 a_n32_n52# a_n508_n52# 0.02fF
C33 a_n224_n52# a_256_n52# 0.02fF
C34 a_n416_n52# a_160_n52# 0.01fF
C35 a_n508_n52# a_160_n52# 0.01fF
C36 a_64_n52# a_n416_n52# 0.02fF
C37 a_n416_n52# a_352_n52# 0.01fF
C38 a_64_n52# a_n508_n52# 0.01fF
C39 a_n508_n52# a_352_n52# 0.01fF
C40 a_n416_n52# a_256_n52# 0.01fF
C41 a_n508_n52# a_256_n52# 0.01fF
C42 a_n32_n52# a_160_n52# 0.05fF
C43 a_n32_n52# a_64_n52# 0.13fF
C44 a_n32_n52# a_352_n52# 0.02fF
C45 a_64_n52# a_160_n52# 0.13fF
C46 a_352_n52# a_160_n52# 0.05fF
C47 a_n32_n52# a_256_n52# 0.03fF
C48 a_64_n52# a_352_n52# 0.03fF
C49 a_160_n52# a_256_n52# 0.13fF
C50 a_64_n52# a_256_n52# 0.05fF
C51 a_352_n52# a_256_n52# 0.13fF
C52 a_448_n52# a_n320_n52# 0.01fF
C53 a_n128_n52# a_n320_n52# 0.05fF
C54 a_448_n52# a_n224_n52# 0.01fF
C55 a_n224_n52# a_n128_n52# 0.13fF
C56 a_448_n52# a_n416_n52# 0.01fF
C57 a_448_n52# a_n508_n52# 0.01fF
C58 a_n512_n140# a_n320_n52# 0.09fF
C59 a_n416_n52# a_n128_n52# 0.03fF
C60 a_n508_n52# a_n128_n52# 0.02fF
C61 a_448_n52# a_n610_n226# 0.07fF
C62 a_352_n52# a_n610_n226# 0.05fF
C63 a_256_n52# a_n610_n226# 0.04fF
C64 a_160_n52# a_n610_n226# 0.04fF
C65 a_64_n52# a_n610_n226# 0.04fF
C66 a_n32_n52# a_n610_n226# 0.04fF
C67 a_n128_n52# a_n610_n226# 0.04fF
C68 a_n224_n52# a_n610_n226# 0.04fF
C69 a_n320_n52# a_n610_n226# 0.04fF
C70 a_n416_n52# a_n610_n226# 0.05fF
C71 a_n508_n52# a_n610_n226# 0.07fF
C72 a_n512_n140# a_n610_n226# 1.45fF
.ends

.subckt transmission_gate in out en en_b VDD VSS
Xsky130_fd_pr__pfet_01v8_UNG2NQ_0 in in out in out in out VDD in out out en_b out
+ VSS sky130_fd_pr__pfet_01v8_UNG2NQ
Xsky130_fd_pr__nfet_01v8_6J4AMR_0 out in in out in in VSS out en in out out out sky130_fd_pr__nfet_01v8_6J4AMR
C0 out en_b 0.03fF
C1 out VDD 0.40fF
C2 out in 0.71fF
C3 en en_b 0.14fF
C4 en VDD 0.05fF
C5 en in 1.30fF
C6 VDD en_b 0.10fF
C7 en out 0.05fF
C8 in en_b 1.18fF
C9 in VDD 0.92fF
C10 en VSS 1.66fF
C11 out VSS 1.04fF
C12 in VSS 1.15fF
C13 en_b VSS 0.24fF
C14 VDD VSS 3.18fF
.ends

