magic
tech sky130A
timestamp 1655484843
<< error_s >>
rect 129 180 158 183
rect 339 180 368 183
rect 549 180 578 183
rect 759 180 788 183
rect 969 180 998 183
rect 1179 180 1208 183
rect 1389 180 1418 183
rect 1599 180 1628 183
rect 1809 180 1838 183
rect 2019 180 2048 183
rect 2229 180 2258 183
rect 2439 180 2468 183
rect 2649 180 2678 183
rect 2859 180 2888 183
rect 3069 180 3098 183
rect 3279 180 3308 183
rect 3489 180 3518 183
rect 3699 180 3728 183
rect 3909 180 3938 183
rect 4119 180 4148 183
rect 129 163 135 180
rect 339 163 345 180
rect 549 163 555 180
rect 759 163 765 180
rect 969 163 975 180
rect 1179 163 1185 180
rect 1389 163 1395 180
rect 1599 163 1605 180
rect 1809 163 1815 180
rect 2019 163 2025 180
rect 2229 163 2235 180
rect 2439 163 2445 180
rect 2649 163 2655 180
rect 2859 163 2865 180
rect 3069 163 3075 180
rect 3279 163 3285 180
rect 3489 163 3495 180
rect 3699 163 3705 180
rect 3909 163 3915 180
rect 4119 163 4125 180
rect 129 160 158 163
rect 339 160 368 163
rect 549 160 578 163
rect 759 160 788 163
rect 969 160 998 163
rect 1179 160 1208 163
rect 1389 160 1418 163
rect 1599 160 1628 163
rect 1809 160 1838 163
rect 2019 160 2048 163
rect 2229 160 2258 163
rect 2439 160 2468 163
rect 2649 160 2678 163
rect 2859 160 2888 163
rect 3069 160 3098 163
rect 3279 160 3308 163
rect 3489 160 3518 163
rect 3699 160 3728 163
rect 3909 160 3938 163
rect 4119 160 4148 163
rect 0 44 31 144
rect 46 44 77 144
rect 105 44 136 144
rect 151 44 182 144
rect 210 44 241 144
rect 256 44 287 144
rect 315 44 346 144
rect 361 44 392 144
rect 420 44 451 144
rect 466 44 497 144
rect 525 44 556 144
rect 571 44 602 144
rect 630 44 661 144
rect 676 44 707 144
rect 735 44 766 144
rect 781 44 812 144
rect 840 44 871 144
rect 886 44 917 144
rect 945 44 976 144
rect 991 44 1022 144
rect 1050 44 1081 144
rect 1096 44 1127 144
rect 1155 44 1186 144
rect 1201 44 1232 144
rect 1260 44 1291 144
rect 1306 44 1337 144
rect 1365 44 1396 144
rect 1411 44 1442 144
rect 1470 44 1501 144
rect 1516 44 1547 144
rect 1575 44 1606 144
rect 1621 44 1652 144
rect 1680 44 1711 144
rect 1726 44 1757 144
rect 1785 44 1816 144
rect 1831 44 1862 144
rect 1890 44 1921 144
rect 1936 44 1967 144
rect 1995 44 2026 144
rect 2041 44 2072 144
rect 2100 44 2131 144
rect 2146 44 2177 144
rect 2205 44 2236 144
rect 2251 44 2282 144
rect 2310 44 2341 144
rect 2356 44 2387 144
rect 2415 44 2446 144
rect 2461 44 2492 144
rect 2520 44 2551 144
rect 2566 44 2597 144
rect 2625 44 2656 144
rect 2671 44 2702 144
rect 2730 44 2761 144
rect 2776 44 2807 144
rect 2835 44 2866 144
rect 2881 44 2912 144
rect 2940 44 2971 144
rect 2986 44 3017 144
rect 3045 44 3076 144
rect 3091 44 3122 144
rect 3150 44 3181 144
rect 3196 44 3227 144
rect 3255 44 3286 144
rect 3301 44 3332 144
rect 3360 44 3391 144
rect 3406 44 3437 144
rect 3465 44 3496 144
rect 3511 44 3542 144
rect 3570 44 3601 144
rect 3616 44 3647 144
rect 3675 44 3706 144
rect 3721 44 3752 144
rect 3780 44 3811 144
rect 3826 44 3857 144
rect 3885 44 3916 144
rect 3931 44 3962 144
rect 3990 44 4021 144
rect 4036 44 4067 144
rect 4095 44 4126 144
rect 4141 44 4172 144
rect 4200 44 4231 144
rect 4246 44 4277 144
rect 4305 44 4336 144
rect 4351 44 4382 144
rect 234 25 263 28
rect 444 25 473 28
rect 654 25 683 28
rect 864 25 893 28
rect 1074 25 1103 28
rect 1284 25 1313 28
rect 1494 25 1523 28
rect 1704 25 1733 28
rect 1914 25 1943 28
rect 2124 25 2153 28
rect 2334 25 2363 28
rect 2544 25 2573 28
rect 2754 25 2783 28
rect 2964 25 2993 28
rect 3174 25 3203 28
rect 3384 25 3413 28
rect 3594 25 3623 28
rect 3804 25 3833 28
rect 4014 25 4043 28
rect 4224 25 4253 28
rect 234 8 240 25
rect 444 8 450 25
rect 654 8 660 25
rect 864 8 870 25
rect 1074 8 1080 25
rect 1284 8 1290 25
rect 1494 8 1500 25
rect 1704 8 1710 25
rect 1914 8 1920 25
rect 2124 8 2130 25
rect 2334 8 2340 25
rect 2544 8 2550 25
rect 2754 8 2760 25
rect 2964 8 2970 25
rect 3174 8 3180 25
rect 3384 8 3390 25
rect 3594 8 3600 25
rect 3804 8 3810 25
rect 4014 8 4020 25
rect 4224 8 4230 25
rect 234 5 263 8
rect 444 5 473 8
rect 654 5 683 8
rect 864 5 893 8
rect 1074 5 1103 8
rect 1284 5 1313 8
rect 1494 5 1523 8
rect 1704 5 1733 8
rect 1914 5 1943 8
rect 2124 5 2153 8
rect 2334 5 2363 8
rect 2544 5 2573 8
rect 2754 5 2783 8
rect 2964 5 2993 8
rect 3174 5 3203 8
rect 3384 5 3413 8
rect 3594 5 3623 8
rect 3804 5 3833 8
rect 4014 5 4043 8
rect 4224 5 4253 8
rect 129 -40 158 -37
rect 339 -40 368 -37
rect 549 -40 578 -37
rect 759 -40 788 -37
rect 969 -40 998 -37
rect 1179 -40 1208 -37
rect 1389 -40 1418 -37
rect 1599 -40 1628 -37
rect 1809 -40 1838 -37
rect 2019 -40 2048 -37
rect 2229 -40 2258 -37
rect 2439 -40 2468 -37
rect 2649 -40 2678 -37
rect 2859 -40 2888 -37
rect 3069 -40 3098 -37
rect 3279 -40 3308 -37
rect 3489 -40 3518 -37
rect 3699 -40 3728 -37
rect 3909 -40 3938 -37
rect 4119 -40 4148 -37
rect 129 -57 135 -40
rect 339 -57 345 -40
rect 549 -57 555 -40
rect 759 -57 765 -40
rect 969 -57 975 -40
rect 1179 -57 1185 -40
rect 1389 -57 1395 -40
rect 1599 -57 1605 -40
rect 1809 -57 1815 -40
rect 2019 -57 2025 -40
rect 2229 -57 2235 -40
rect 2439 -57 2445 -40
rect 2649 -57 2655 -40
rect 2859 -57 2865 -40
rect 3069 -57 3075 -40
rect 3279 -57 3285 -40
rect 3489 -57 3495 -40
rect 3699 -57 3705 -40
rect 3909 -57 3915 -40
rect 4119 -57 4125 -40
rect 129 -60 158 -57
rect 339 -60 368 -57
rect 549 -60 578 -57
rect 759 -60 788 -57
rect 969 -60 998 -57
rect 1179 -60 1208 -57
rect 1389 -60 1418 -57
rect 1599 -60 1628 -57
rect 1809 -60 1838 -57
rect 2019 -60 2048 -57
rect 2229 -60 2258 -57
rect 2439 -60 2468 -57
rect 2649 -60 2678 -57
rect 2859 -60 2888 -57
rect 3069 -60 3098 -57
rect 3279 -60 3308 -57
rect 3489 -60 3518 -57
rect 3699 -60 3728 -57
rect 3909 -60 3938 -57
rect 4119 -60 4148 -57
rect 0 -176 31 -76
rect 46 -176 77 -76
rect 105 -176 136 -76
rect 151 -176 182 -76
rect 210 -176 241 -76
rect 256 -176 287 -76
rect 315 -176 346 -76
rect 361 -176 392 -76
rect 420 -176 451 -76
rect 466 -176 497 -76
rect 525 -176 556 -76
rect 571 -176 602 -76
rect 630 -176 661 -76
rect 676 -176 707 -76
rect 735 -176 766 -76
rect 781 -176 812 -76
rect 840 -176 871 -76
rect 886 -176 917 -76
rect 945 -176 976 -76
rect 991 -176 1022 -76
rect 1050 -176 1081 -76
rect 1096 -176 1127 -76
rect 1155 -176 1186 -76
rect 1201 -176 1232 -76
rect 1260 -176 1291 -76
rect 1306 -176 1337 -76
rect 1365 -176 1396 -76
rect 1411 -176 1442 -76
rect 1470 -176 1501 -76
rect 1516 -176 1547 -76
rect 1575 -176 1606 -76
rect 1621 -176 1652 -76
rect 1680 -176 1711 -76
rect 1726 -176 1757 -76
rect 1785 -176 1816 -76
rect 1831 -176 1862 -76
rect 1890 -176 1921 -76
rect 1936 -176 1967 -76
rect 1995 -176 2026 -76
rect 2041 -176 2072 -76
rect 2100 -176 2131 -76
rect 2146 -176 2177 -76
rect 2205 -176 2236 -76
rect 2251 -176 2282 -76
rect 2310 -176 2341 -76
rect 2356 -176 2387 -76
rect 2415 -176 2446 -76
rect 2461 -176 2492 -76
rect 2520 -176 2551 -76
rect 2566 -176 2597 -76
rect 2625 -176 2656 -76
rect 2671 -176 2702 -76
rect 2730 -176 2761 -76
rect 2776 -176 2807 -76
rect 2835 -176 2866 -76
rect 2881 -176 2912 -76
rect 2940 -176 2971 -76
rect 2986 -176 3017 -76
rect 3045 -176 3076 -76
rect 3091 -176 3122 -76
rect 3150 -176 3181 -76
rect 3196 -176 3227 -76
rect 3255 -176 3286 -76
rect 3301 -176 3332 -76
rect 3360 -176 3391 -76
rect 3406 -176 3437 -76
rect 3465 -176 3496 -76
rect 3511 -176 3542 -76
rect 3570 -176 3601 -76
rect 3616 -176 3647 -76
rect 3675 -176 3706 -76
rect 3721 -176 3752 -76
rect 3780 -176 3811 -76
rect 3826 -176 3857 -76
rect 3885 -176 3916 -76
rect 3931 -176 3962 -76
rect 3990 -176 4021 -76
rect 4036 -176 4067 -76
rect 4095 -176 4126 -76
rect 4141 -176 4172 -76
rect 4200 -176 4231 -76
rect 4246 -176 4277 -76
rect 4305 -176 4336 -76
rect 4351 -176 4382 -76
rect 234 -195 263 -192
rect 444 -195 473 -192
rect 654 -195 683 -192
rect 864 -195 893 -192
rect 1074 -195 1103 -192
rect 1284 -195 1313 -192
rect 1494 -195 1523 -192
rect 1704 -195 1733 -192
rect 1914 -195 1943 -192
rect 2124 -195 2153 -192
rect 2334 -195 2363 -192
rect 2544 -195 2573 -192
rect 2754 -195 2783 -192
rect 2964 -195 2993 -192
rect 3174 -195 3203 -192
rect 3384 -195 3413 -192
rect 3594 -195 3623 -192
rect 3804 -195 3833 -192
rect 4014 -195 4043 -192
rect 4224 -195 4253 -192
rect 234 -212 240 -195
rect 444 -212 450 -195
rect 654 -212 660 -195
rect 864 -212 870 -195
rect 1074 -212 1080 -195
rect 1284 -212 1290 -195
rect 1494 -212 1500 -195
rect 1704 -212 1710 -195
rect 1914 -212 1920 -195
rect 2124 -212 2130 -195
rect 2334 -212 2340 -195
rect 2544 -212 2550 -195
rect 2754 -212 2760 -195
rect 2964 -212 2970 -195
rect 3174 -212 3180 -195
rect 3384 -212 3390 -195
rect 3594 -212 3600 -195
rect 3804 -212 3810 -195
rect 4014 -212 4020 -195
rect 4224 -212 4230 -195
rect 234 -215 263 -212
rect 444 -215 473 -212
rect 654 -215 683 -212
rect 864 -215 893 -212
rect 1074 -215 1103 -212
rect 1284 -215 1313 -212
rect 1494 -215 1523 -212
rect 1704 -215 1733 -212
rect 1914 -215 1943 -212
rect 2124 -215 2153 -212
rect 2334 -215 2363 -212
rect 2544 -215 2573 -212
rect 2754 -215 2783 -212
rect 2964 -215 2993 -212
rect 3174 -215 3203 -212
rect 3384 -215 3413 -212
rect 3594 -215 3623 -212
rect 3804 -215 3833 -212
rect 4014 -215 4043 -212
rect 4224 -215 4253 -212
rect 129 -260 158 -257
rect 339 -260 368 -257
rect 549 -260 578 -257
rect 759 -260 788 -257
rect 969 -260 998 -257
rect 1179 -260 1208 -257
rect 1389 -260 1418 -257
rect 1599 -260 1628 -257
rect 1809 -260 1838 -257
rect 2019 -260 2048 -257
rect 2229 -260 2258 -257
rect 2439 -260 2468 -257
rect 2649 -260 2678 -257
rect 2859 -260 2888 -257
rect 3069 -260 3098 -257
rect 3279 -260 3308 -257
rect 3489 -260 3518 -257
rect 3699 -260 3728 -257
rect 3909 -260 3938 -257
rect 4119 -260 4148 -257
rect 129 -277 135 -260
rect 339 -277 345 -260
rect 549 -277 555 -260
rect 759 -277 765 -260
rect 969 -277 975 -260
rect 1179 -277 1185 -260
rect 1389 -277 1395 -260
rect 1599 -277 1605 -260
rect 1809 -277 1815 -260
rect 2019 -277 2025 -260
rect 2229 -277 2235 -260
rect 2439 -277 2445 -260
rect 2649 -277 2655 -260
rect 2859 -277 2865 -260
rect 3069 -277 3075 -260
rect 3279 -277 3285 -260
rect 3489 -277 3495 -260
rect 3699 -277 3705 -260
rect 3909 -277 3915 -260
rect 4119 -277 4125 -260
rect 129 -280 158 -277
rect 339 -280 368 -277
rect 549 -280 578 -277
rect 759 -280 788 -277
rect 969 -280 998 -277
rect 1179 -280 1208 -277
rect 1389 -280 1418 -277
rect 1599 -280 1628 -277
rect 1809 -280 1838 -277
rect 2019 -280 2048 -277
rect 2229 -280 2258 -277
rect 2439 -280 2468 -277
rect 2649 -280 2678 -277
rect 2859 -280 2888 -277
rect 3069 -280 3098 -277
rect 3279 -280 3308 -277
rect 3489 -280 3518 -277
rect 3699 -280 3728 -277
rect 3909 -280 3938 -277
rect 4119 -280 4148 -277
rect 0 -396 31 -296
rect 46 -396 77 -296
rect 105 -396 136 -296
rect 151 -396 182 -296
rect 210 -396 241 -296
rect 256 -396 287 -296
rect 315 -396 346 -296
rect 361 -396 392 -296
rect 420 -396 451 -296
rect 466 -396 497 -296
rect 525 -396 556 -296
rect 571 -396 602 -296
rect 630 -396 661 -296
rect 676 -396 707 -296
rect 735 -396 766 -296
rect 781 -396 812 -296
rect 840 -396 871 -296
rect 886 -396 917 -296
rect 945 -396 976 -296
rect 991 -396 1022 -296
rect 1050 -396 1081 -296
rect 1096 -396 1127 -296
rect 1155 -396 1186 -296
rect 1201 -396 1232 -296
rect 1260 -396 1291 -296
rect 1306 -396 1337 -296
rect 1365 -396 1396 -296
rect 1411 -396 1442 -296
rect 1470 -396 1501 -296
rect 1516 -396 1547 -296
rect 1575 -396 1606 -296
rect 1621 -396 1652 -296
rect 1680 -396 1711 -296
rect 1726 -396 1757 -296
rect 1785 -396 1816 -296
rect 1831 -396 1862 -296
rect 1890 -396 1921 -296
rect 1936 -396 1967 -296
rect 1995 -396 2026 -296
rect 2041 -396 2072 -296
rect 2100 -396 2131 -296
rect 2146 -396 2177 -296
rect 2205 -396 2236 -296
rect 2251 -396 2282 -296
rect 2310 -396 2341 -296
rect 2356 -396 2387 -296
rect 2415 -396 2446 -296
rect 2461 -396 2492 -296
rect 2520 -396 2551 -296
rect 2566 -396 2597 -296
rect 2625 -396 2656 -296
rect 2671 -396 2702 -296
rect 2730 -396 2761 -296
rect 2776 -396 2807 -296
rect 2835 -396 2866 -296
rect 2881 -396 2912 -296
rect 2940 -396 2971 -296
rect 2986 -396 3017 -296
rect 3045 -396 3076 -296
rect 3091 -396 3122 -296
rect 3150 -396 3181 -296
rect 3196 -396 3227 -296
rect 3255 -396 3286 -296
rect 3301 -396 3332 -296
rect 3360 -396 3391 -296
rect 3406 -396 3437 -296
rect 3465 -396 3496 -296
rect 3511 -396 3542 -296
rect 3570 -396 3601 -296
rect 3616 -396 3647 -296
rect 3675 -396 3706 -296
rect 3721 -396 3752 -296
rect 3780 -396 3811 -296
rect 3826 -396 3857 -296
rect 3885 -396 3916 -296
rect 3931 -396 3962 -296
rect 3990 -396 4021 -296
rect 4036 -396 4067 -296
rect 4095 -396 4126 -296
rect 4141 -396 4172 -296
rect 4200 -396 4231 -296
rect 4246 -396 4277 -296
rect 4305 -396 4336 -296
rect 4351 -396 4382 -296
rect 234 -415 263 -412
rect 444 -415 473 -412
rect 654 -415 683 -412
rect 864 -415 893 -412
rect 1074 -415 1103 -412
rect 1284 -415 1313 -412
rect 1494 -415 1523 -412
rect 1704 -415 1733 -412
rect 1914 -415 1943 -412
rect 2124 -415 2153 -412
rect 2334 -415 2363 -412
rect 2544 -415 2573 -412
rect 2754 -415 2783 -412
rect 2964 -415 2993 -412
rect 3174 -415 3203 -412
rect 3384 -415 3413 -412
rect 3594 -415 3623 -412
rect 3804 -415 3833 -412
rect 4014 -415 4043 -412
rect 4224 -415 4253 -412
rect 234 -432 240 -415
rect 444 -432 450 -415
rect 654 -432 660 -415
rect 864 -432 870 -415
rect 1074 -432 1080 -415
rect 1284 -432 1290 -415
rect 1494 -432 1500 -415
rect 1704 -432 1710 -415
rect 1914 -432 1920 -415
rect 2124 -432 2130 -415
rect 2334 -432 2340 -415
rect 2544 -432 2550 -415
rect 2754 -432 2760 -415
rect 2964 -432 2970 -415
rect 3174 -432 3180 -415
rect 3384 -432 3390 -415
rect 3594 -432 3600 -415
rect 3804 -432 3810 -415
rect 4014 -432 4020 -415
rect 4224 -432 4230 -415
rect 234 -435 263 -432
rect 444 -435 473 -432
rect 654 -435 683 -432
rect 864 -435 893 -432
rect 1074 -435 1103 -432
rect 1284 -435 1313 -432
rect 1494 -435 1523 -432
rect 1704 -435 1733 -432
rect 1914 -435 1943 -432
rect 2124 -435 2153 -432
rect 2334 -435 2363 -432
rect 2544 -435 2573 -432
rect 2754 -435 2783 -432
rect 2964 -435 2993 -432
rect 3174 -435 3203 -432
rect 3384 -435 3413 -432
rect 3594 -435 3623 -432
rect 3804 -435 3833 -432
rect 4014 -435 4043 -432
rect 4224 -435 4253 -432
rect 129 -480 158 -477
rect 339 -480 368 -477
rect 549 -480 578 -477
rect 759 -480 788 -477
rect 969 -480 998 -477
rect 1179 -480 1208 -477
rect 1389 -480 1418 -477
rect 1599 -480 1628 -477
rect 1809 -480 1838 -477
rect 2019 -480 2048 -477
rect 2229 -480 2258 -477
rect 2439 -480 2468 -477
rect 2649 -480 2678 -477
rect 2859 -480 2888 -477
rect 3069 -480 3098 -477
rect 3279 -480 3308 -477
rect 3489 -480 3518 -477
rect 3699 -480 3728 -477
rect 3909 -480 3938 -477
rect 4119 -480 4148 -477
rect 129 -497 135 -480
rect 339 -497 345 -480
rect 549 -497 555 -480
rect 759 -497 765 -480
rect 969 -497 975 -480
rect 1179 -497 1185 -480
rect 1389 -497 1395 -480
rect 1599 -497 1605 -480
rect 1809 -497 1815 -480
rect 2019 -497 2025 -480
rect 2229 -497 2235 -480
rect 2439 -497 2445 -480
rect 2649 -497 2655 -480
rect 2859 -497 2865 -480
rect 3069 -497 3075 -480
rect 3279 -497 3285 -480
rect 3489 -497 3495 -480
rect 3699 -497 3705 -480
rect 3909 -497 3915 -480
rect 4119 -497 4125 -480
rect 129 -500 158 -497
rect 339 -500 368 -497
rect 549 -500 578 -497
rect 759 -500 788 -497
rect 969 -500 998 -497
rect 1179 -500 1208 -497
rect 1389 -500 1418 -497
rect 1599 -500 1628 -497
rect 1809 -500 1838 -497
rect 2019 -500 2048 -497
rect 2229 -500 2258 -497
rect 2439 -500 2468 -497
rect 2649 -500 2678 -497
rect 2859 -500 2888 -497
rect 3069 -500 3098 -497
rect 3279 -500 3308 -497
rect 3489 -500 3518 -497
rect 3699 -500 3728 -497
rect 3909 -500 3938 -497
rect 4119 -500 4148 -497
rect 0 -616 31 -516
rect 46 -616 77 -516
rect 105 -616 136 -516
rect 151 -616 182 -516
rect 210 -616 241 -516
rect 256 -616 287 -516
rect 315 -616 346 -516
rect 361 -616 392 -516
rect 420 -616 451 -516
rect 466 -616 497 -516
rect 525 -616 556 -516
rect 571 -616 602 -516
rect 630 -616 661 -516
rect 676 -616 707 -516
rect 735 -616 766 -516
rect 781 -616 812 -516
rect 840 -616 871 -516
rect 886 -616 917 -516
rect 945 -616 976 -516
rect 991 -616 1022 -516
rect 1050 -616 1081 -516
rect 1096 -616 1127 -516
rect 1155 -616 1186 -516
rect 1201 -616 1232 -516
rect 1260 -616 1291 -516
rect 1306 -616 1337 -516
rect 1365 -616 1396 -516
rect 1411 -616 1442 -516
rect 1470 -616 1501 -516
rect 1516 -616 1547 -516
rect 1575 -616 1606 -516
rect 1621 -616 1652 -516
rect 1680 -616 1711 -516
rect 1726 -616 1757 -516
rect 1785 -616 1816 -516
rect 1831 -616 1862 -516
rect 1890 -616 1921 -516
rect 1936 -616 1967 -516
rect 1995 -616 2026 -516
rect 2041 -616 2072 -516
rect 2100 -616 2131 -516
rect 2146 -616 2177 -516
rect 2205 -616 2236 -516
rect 2251 -616 2282 -516
rect 2310 -616 2341 -516
rect 2356 -616 2387 -516
rect 2415 -616 2446 -516
rect 2461 -616 2492 -516
rect 2520 -616 2551 -516
rect 2566 -616 2597 -516
rect 2625 -616 2656 -516
rect 2671 -616 2702 -516
rect 2730 -616 2761 -516
rect 2776 -616 2807 -516
rect 2835 -616 2866 -516
rect 2881 -616 2912 -516
rect 2940 -616 2971 -516
rect 2986 -616 3017 -516
rect 3045 -616 3076 -516
rect 3091 -616 3122 -516
rect 3150 -616 3181 -516
rect 3196 -616 3227 -516
rect 3255 -616 3286 -516
rect 3301 -616 3332 -516
rect 3360 -616 3391 -516
rect 3406 -616 3437 -516
rect 3465 -616 3496 -516
rect 3511 -616 3542 -516
rect 3570 -616 3601 -516
rect 3616 -616 3647 -516
rect 3675 -616 3706 -516
rect 3721 -616 3752 -516
rect 3780 -616 3811 -516
rect 3826 -616 3857 -516
rect 3885 -616 3916 -516
rect 3931 -616 3962 -516
rect 3990 -616 4021 -516
rect 4036 -616 4067 -516
rect 4095 -616 4126 -516
rect 4141 -616 4172 -516
rect 4200 -616 4231 -516
rect 4246 -616 4277 -516
rect 4305 -616 4336 -516
rect 4351 -616 4382 -516
rect 234 -635 263 -632
rect 444 -635 473 -632
rect 654 -635 683 -632
rect 864 -635 893 -632
rect 1074 -635 1103 -632
rect 1284 -635 1313 -632
rect 1494 -635 1523 -632
rect 1704 -635 1733 -632
rect 1914 -635 1943 -632
rect 2124 -635 2153 -632
rect 2334 -635 2363 -632
rect 2544 -635 2573 -632
rect 2754 -635 2783 -632
rect 2964 -635 2993 -632
rect 3174 -635 3203 -632
rect 3384 -635 3413 -632
rect 3594 -635 3623 -632
rect 3804 -635 3833 -632
rect 4014 -635 4043 -632
rect 4224 -635 4253 -632
rect 234 -652 240 -635
rect 444 -652 450 -635
rect 654 -652 660 -635
rect 864 -652 870 -635
rect 1074 -652 1080 -635
rect 1284 -652 1290 -635
rect 1494 -652 1500 -635
rect 1704 -652 1710 -635
rect 1914 -652 1920 -635
rect 2124 -652 2130 -635
rect 2334 -652 2340 -635
rect 2544 -652 2550 -635
rect 2754 -652 2760 -635
rect 2964 -652 2970 -635
rect 3174 -652 3180 -635
rect 3384 -652 3390 -635
rect 3594 -652 3600 -635
rect 3804 -652 3810 -635
rect 4014 -652 4020 -635
rect 4224 -652 4230 -635
rect 234 -655 263 -652
rect 444 -655 473 -652
rect 654 -655 683 -652
rect 864 -655 893 -652
rect 1074 -655 1103 -652
rect 1284 -655 1313 -652
rect 1494 -655 1523 -652
rect 1704 -655 1733 -652
rect 1914 -655 1943 -652
rect 2124 -655 2153 -652
rect 2334 -655 2363 -652
rect 2544 -655 2573 -652
rect 2754 -655 2783 -652
rect 2964 -655 2993 -652
rect 3174 -655 3203 -652
rect 3384 -655 3413 -652
rect 3594 -655 3623 -652
rect 3804 -655 3833 -652
rect 4014 -655 4043 -652
rect 4224 -655 4253 -652
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_0
timestamp 1655484843
transform 1 0 2191 0 1 94
box -2191 -94 2191 94
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_1
timestamp 1655484843
transform 1 0 2191 0 1 -126
box -2191 -94 2191 94
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_2
timestamp 1655484843
transform 1 0 2191 0 1 -346
box -2191 -94 2191 94
use sky130_fd_pr__nfet_01v8_J3WY8C  sky130_fd_pr__nfet_01v8_J3WY8C_3
timestamp 1655484843
transform 1 0 2191 0 1 -566
box -2191 -94 2191 94
<< end >>
