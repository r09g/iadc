magic
tech sky130A
magscale 1 2
timestamp 1653693763
<< nwell >>
rect 163 464 1457 1114
rect 157 -688 1451 -38
<< pwell >>
rect 163 0 1457 462
rect 157 -1152 1451 -690
<< nmos >>
rect 363 210 393 314
rect 459 210 489 314
rect 555 210 585 314
rect 651 210 681 314
rect 747 210 777 314
rect 843 210 873 314
rect 939 210 969 314
rect 1035 210 1065 314
rect 1131 210 1161 314
rect 1227 210 1257 314
rect 357 -942 387 -838
rect 453 -942 483 -838
rect 549 -942 579 -838
rect 645 -942 675 -838
rect 741 -942 771 -838
rect 837 -942 867 -838
rect 933 -942 963 -838
rect 1029 -942 1059 -838
rect 1125 -942 1155 -838
rect 1221 -942 1251 -838
<< pmos >>
rect 363 622 393 894
rect 459 622 489 894
rect 555 622 585 894
rect 651 622 681 894
rect 747 622 777 894
rect 843 622 873 894
rect 939 622 969 894
rect 1035 622 1065 894
rect 1131 622 1161 894
rect 1227 622 1257 894
rect 357 -530 387 -258
rect 453 -530 483 -258
rect 549 -530 579 -258
rect 645 -530 675 -258
rect 741 -530 771 -258
rect 837 -530 867 -258
rect 933 -530 963 -258
rect 1029 -530 1059 -258
rect 1125 -530 1155 -258
rect 1221 -530 1251 -258
<< ndiff >>
rect 301 302 363 314
rect 301 222 313 302
rect 347 222 363 302
rect 301 210 363 222
rect 393 302 459 314
rect 393 222 409 302
rect 443 222 459 302
rect 393 210 459 222
rect 489 302 555 314
rect 489 222 505 302
rect 539 222 555 302
rect 489 210 555 222
rect 585 302 651 314
rect 585 222 601 302
rect 635 222 651 302
rect 585 210 651 222
rect 681 302 747 314
rect 681 222 697 302
rect 731 222 747 302
rect 681 210 747 222
rect 777 302 843 314
rect 777 222 793 302
rect 827 222 843 302
rect 777 210 843 222
rect 873 302 939 314
rect 873 222 889 302
rect 923 222 939 302
rect 873 210 939 222
rect 969 302 1035 314
rect 969 222 985 302
rect 1019 222 1035 302
rect 969 210 1035 222
rect 1065 302 1131 314
rect 1065 222 1081 302
rect 1115 222 1131 302
rect 1065 210 1131 222
rect 1161 302 1227 314
rect 1161 222 1177 302
rect 1211 222 1227 302
rect 1161 210 1227 222
rect 1257 302 1319 314
rect 1257 222 1273 302
rect 1307 222 1319 302
rect 1257 210 1319 222
rect 295 -850 357 -838
rect 295 -930 307 -850
rect 341 -930 357 -850
rect 295 -942 357 -930
rect 387 -850 453 -838
rect 387 -930 403 -850
rect 437 -930 453 -850
rect 387 -942 453 -930
rect 483 -850 549 -838
rect 483 -930 499 -850
rect 533 -930 549 -850
rect 483 -942 549 -930
rect 579 -850 645 -838
rect 579 -930 595 -850
rect 629 -930 645 -850
rect 579 -942 645 -930
rect 675 -850 741 -838
rect 675 -930 691 -850
rect 725 -930 741 -850
rect 675 -942 741 -930
rect 771 -850 837 -838
rect 771 -930 787 -850
rect 821 -930 837 -850
rect 771 -942 837 -930
rect 867 -850 933 -838
rect 867 -930 883 -850
rect 917 -930 933 -850
rect 867 -942 933 -930
rect 963 -850 1029 -838
rect 963 -930 979 -850
rect 1013 -930 1029 -850
rect 963 -942 1029 -930
rect 1059 -850 1125 -838
rect 1059 -930 1075 -850
rect 1109 -930 1125 -850
rect 1059 -942 1125 -930
rect 1155 -850 1221 -838
rect 1155 -930 1171 -850
rect 1205 -930 1221 -850
rect 1155 -942 1221 -930
rect 1251 -850 1313 -838
rect 1251 -930 1267 -850
rect 1301 -930 1313 -850
rect 1251 -942 1313 -930
<< pdiff >>
rect 301 882 363 894
rect 301 634 313 882
rect 347 634 363 882
rect 301 622 363 634
rect 393 882 459 894
rect 393 634 409 882
rect 443 634 459 882
rect 393 622 459 634
rect 489 882 555 894
rect 489 634 505 882
rect 539 634 555 882
rect 489 622 555 634
rect 585 882 651 894
rect 585 634 601 882
rect 635 634 651 882
rect 585 622 651 634
rect 681 882 747 894
rect 681 634 697 882
rect 731 634 747 882
rect 681 622 747 634
rect 777 882 843 894
rect 777 634 793 882
rect 827 634 843 882
rect 777 622 843 634
rect 873 882 939 894
rect 873 634 889 882
rect 923 634 939 882
rect 873 622 939 634
rect 969 882 1035 894
rect 969 634 985 882
rect 1019 634 1035 882
rect 969 622 1035 634
rect 1065 882 1131 894
rect 1065 634 1081 882
rect 1115 634 1131 882
rect 1065 622 1131 634
rect 1161 882 1227 894
rect 1161 634 1177 882
rect 1211 634 1227 882
rect 1161 622 1227 634
rect 1257 882 1319 894
rect 1257 634 1273 882
rect 1307 634 1319 882
rect 1257 622 1319 634
rect 295 -270 357 -258
rect 295 -518 307 -270
rect 341 -518 357 -270
rect 295 -530 357 -518
rect 387 -270 453 -258
rect 387 -518 403 -270
rect 437 -518 453 -270
rect 387 -530 453 -518
rect 483 -270 549 -258
rect 483 -518 499 -270
rect 533 -518 549 -270
rect 483 -530 549 -518
rect 579 -270 645 -258
rect 579 -518 595 -270
rect 629 -518 645 -270
rect 579 -530 645 -518
rect 675 -270 741 -258
rect 675 -518 691 -270
rect 725 -518 741 -270
rect 675 -530 741 -518
rect 771 -270 837 -258
rect 771 -518 787 -270
rect 821 -518 837 -270
rect 771 -530 837 -518
rect 867 -270 933 -258
rect 867 -518 883 -270
rect 917 -518 933 -270
rect 867 -530 933 -518
rect 963 -270 1029 -258
rect 963 -518 979 -270
rect 1013 -518 1029 -270
rect 963 -530 1029 -518
rect 1059 -270 1125 -258
rect 1059 -518 1075 -270
rect 1109 -518 1125 -270
rect 1059 -530 1125 -518
rect 1155 -270 1221 -258
rect 1155 -518 1171 -270
rect 1205 -518 1221 -270
rect 1155 -530 1221 -518
rect 1251 -270 1313 -258
rect 1251 -518 1267 -270
rect 1301 -518 1313 -270
rect 1251 -530 1313 -518
<< ndiffc >>
rect 313 222 347 302
rect 409 222 443 302
rect 505 222 539 302
rect 601 222 635 302
rect 697 222 731 302
rect 793 222 827 302
rect 889 222 923 302
rect 985 222 1019 302
rect 1081 222 1115 302
rect 1177 222 1211 302
rect 1273 222 1307 302
rect 307 -930 341 -850
rect 403 -930 437 -850
rect 499 -930 533 -850
rect 595 -930 629 -850
rect 691 -930 725 -850
rect 787 -930 821 -850
rect 883 -930 917 -850
rect 979 -930 1013 -850
rect 1075 -930 1109 -850
rect 1171 -930 1205 -850
rect 1267 -930 1301 -850
<< pdiffc >>
rect 313 634 347 882
rect 409 634 443 882
rect 505 634 539 882
rect 601 634 635 882
rect 697 634 731 882
rect 793 634 827 882
rect 889 634 923 882
rect 985 634 1019 882
rect 1081 634 1115 882
rect 1177 634 1211 882
rect 1273 634 1307 882
rect 307 -518 341 -270
rect 403 -518 437 -270
rect 499 -518 533 -270
rect 595 -518 629 -270
rect 691 -518 725 -270
rect 787 -518 821 -270
rect 883 -518 917 -270
rect 979 -518 1013 -270
rect 1075 -518 1109 -270
rect 1171 -518 1205 -270
rect 1267 -518 1301 -270
<< psubdiff >>
rect 199 392 295 426
rect 1325 392 1421 426
rect 199 330 233 392
rect 1387 330 1421 392
rect 199 70 233 132
rect 1387 70 1421 132
rect 199 36 295 70
rect 1325 36 1421 70
rect 193 -760 289 -726
rect 1319 -760 1415 -726
rect 193 -822 227 -760
rect 1381 -822 1415 -760
rect 193 -1082 227 -1020
rect 1381 -1082 1415 -1020
rect 193 -1116 289 -1082
rect 1319 -1116 1415 -1082
<< nsubdiff >>
rect 199 1044 295 1078
rect 1325 1044 1421 1078
rect 199 982 233 1044
rect 1387 982 1421 1044
rect 199 534 233 596
rect 1387 534 1421 596
rect 199 500 295 534
rect 1325 500 1421 534
rect 193 -108 289 -74
rect 1319 -108 1415 -74
rect 193 -170 227 -108
rect 1381 -170 1415 -108
rect 193 -618 227 -556
rect 1381 -618 1415 -556
rect 193 -652 289 -618
rect 1319 -652 1415 -618
<< psubdiffcont >>
rect 295 392 1325 426
rect 199 132 233 330
rect 1387 132 1421 330
rect 295 36 1325 70
rect 289 -760 1319 -726
rect 193 -1020 227 -822
rect 1381 -1020 1415 -822
rect 289 -1116 1319 -1082
<< nsubdiffcont >>
rect 295 1044 1325 1078
rect 199 596 233 982
rect 1387 596 1421 982
rect 295 500 1325 534
rect 289 -108 1319 -74
rect 193 -556 227 -170
rect 1381 -556 1415 -170
rect 289 -652 1319 -618
<< poly >>
rect 297 976 1323 992
rect 297 942 313 976
rect 347 942 505 976
rect 539 942 697 976
rect 731 942 889 976
rect 923 942 1081 976
rect 1115 942 1273 976
rect 1307 942 1323 976
rect 297 926 1323 942
rect 363 894 393 926
rect 459 894 489 926
rect 555 894 585 926
rect 651 894 681 926
rect 747 894 777 926
rect 843 894 873 926
rect 939 894 969 926
rect 1035 894 1065 926
rect 1131 894 1161 926
rect 1227 894 1257 926
rect 363 596 393 622
rect 459 596 489 622
rect 555 596 585 622
rect 651 596 681 622
rect 747 596 777 622
rect 843 596 873 622
rect 939 596 969 622
rect 1035 596 1065 622
rect 1131 596 1161 622
rect 1227 596 1257 622
rect 363 314 393 340
rect 459 314 489 340
rect 555 314 585 340
rect 651 314 681 340
rect 747 314 777 340
rect 843 314 873 340
rect 939 314 969 340
rect 1035 314 1065 340
rect 1131 314 1161 340
rect 1227 314 1257 340
rect 363 188 393 210
rect 459 188 489 210
rect 555 188 585 210
rect 651 188 681 210
rect 747 188 777 210
rect 843 188 873 210
rect 939 188 969 210
rect 1035 188 1065 210
rect 1131 188 1161 210
rect 1227 188 1257 210
rect 297 168 1323 188
rect 297 134 313 168
rect 347 134 505 168
rect 539 134 697 168
rect 731 134 889 168
rect 923 134 1081 168
rect 1115 134 1273 168
rect 1307 134 1323 168
rect 297 122 1323 134
rect 291 -176 1317 -160
rect 291 -210 307 -176
rect 341 -210 499 -176
rect 533 -210 691 -176
rect 725 -210 883 -176
rect 917 -210 1075 -176
rect 1109 -210 1267 -176
rect 1301 -210 1317 -176
rect 291 -226 1317 -210
rect 357 -258 387 -226
rect 453 -258 483 -226
rect 549 -258 579 -226
rect 645 -258 675 -226
rect 741 -258 771 -226
rect 837 -258 867 -226
rect 933 -258 963 -226
rect 1029 -258 1059 -226
rect 1125 -258 1155 -226
rect 1221 -258 1251 -226
rect 357 -556 387 -530
rect 453 -556 483 -530
rect 549 -556 579 -530
rect 645 -556 675 -530
rect 741 -556 771 -530
rect 837 -556 867 -530
rect 933 -556 963 -530
rect 1029 -556 1059 -530
rect 1125 -556 1155 -530
rect 1221 -556 1251 -530
rect 357 -838 387 -812
rect 453 -838 483 -812
rect 549 -838 579 -812
rect 645 -838 675 -812
rect 741 -838 771 -812
rect 837 -838 867 -812
rect 933 -838 963 -812
rect 1029 -838 1059 -812
rect 1125 -838 1155 -812
rect 1221 -838 1251 -812
rect 357 -964 387 -942
rect 453 -964 483 -942
rect 549 -964 579 -942
rect 645 -964 675 -942
rect 741 -964 771 -942
rect 837 -964 867 -942
rect 933 -964 963 -942
rect 1029 -964 1059 -942
rect 1125 -964 1155 -942
rect 1221 -964 1251 -942
rect 291 -984 1317 -964
rect 291 -1018 307 -984
rect 341 -1018 499 -984
rect 533 -1018 691 -984
rect 725 -1018 883 -984
rect 917 -1018 1075 -984
rect 1109 -1018 1267 -984
rect 1301 -1018 1317 -984
rect 291 -1030 1317 -1018
<< polycont >>
rect 313 942 347 976
rect 505 942 539 976
rect 697 942 731 976
rect 889 942 923 976
rect 1081 942 1115 976
rect 1273 942 1307 976
rect 313 134 347 168
rect 505 134 539 168
rect 697 134 731 168
rect 889 134 923 168
rect 1081 134 1115 168
rect 1273 134 1307 168
rect 307 -210 341 -176
rect 499 -210 533 -176
rect 691 -210 725 -176
rect 883 -210 917 -176
rect 1075 -210 1109 -176
rect 1267 -210 1301 -176
rect 307 -1018 341 -984
rect 499 -1018 533 -984
rect 691 -1018 725 -984
rect 883 -1018 917 -984
rect 1075 -1018 1109 -984
rect 1267 -1018 1301 -984
<< locali >>
rect 199 1044 295 1078
rect 1325 1044 1421 1078
rect 199 982 233 1044
rect 1387 982 1421 1044
rect 297 942 313 976
rect 347 942 363 976
rect 489 942 505 976
rect 539 942 555 976
rect 681 942 697 976
rect 731 942 747 976
rect 873 942 889 976
rect 923 942 939 976
rect 1065 942 1081 976
rect 1115 942 1131 976
rect 1257 942 1273 976
rect 1307 942 1323 976
rect 313 882 347 898
rect 313 618 347 634
rect 409 882 443 898
rect 409 618 443 634
rect 505 882 539 898
rect 505 618 539 634
rect 601 882 635 898
rect 601 618 635 634
rect 697 882 731 898
rect 697 618 731 634
rect 793 882 827 898
rect 793 618 827 634
rect 889 882 923 898
rect 889 618 923 634
rect 985 882 1019 898
rect 985 618 1019 634
rect 1081 882 1115 898
rect 1081 618 1115 634
rect 1177 882 1211 898
rect 1177 618 1211 634
rect 1273 882 1307 898
rect 1273 618 1307 634
rect 199 534 233 596
rect 1387 534 1421 596
rect 199 500 295 534
rect 1325 500 1421 534
rect 199 392 295 426
rect 1325 392 1421 426
rect 199 330 233 392
rect 1387 332 1421 392
rect 313 302 347 318
rect 313 206 347 222
rect 409 302 443 318
rect 409 206 443 222
rect 505 302 539 318
rect 505 206 539 222
rect 601 302 635 318
rect 601 206 635 222
rect 697 302 731 318
rect 697 206 731 222
rect 793 302 827 318
rect 793 206 827 222
rect 889 302 923 318
rect 889 206 923 222
rect 985 302 1019 318
rect 985 206 1019 222
rect 1081 302 1115 318
rect 1081 206 1115 222
rect 1177 302 1211 318
rect 1177 206 1211 222
rect 1273 302 1307 318
rect 1273 206 1307 222
rect 297 134 313 168
rect 347 134 363 168
rect 489 134 505 168
rect 539 134 555 168
rect 681 134 697 168
rect 731 134 747 168
rect 873 134 889 168
rect 923 134 939 168
rect 1065 134 1081 168
rect 1115 134 1131 168
rect 1257 134 1273 168
rect 1307 134 1323 168
rect 199 70 233 132
rect 1387 70 1421 132
rect 199 36 295 70
rect 1325 36 1421 70
rect 193 -108 289 -74
rect 1319 -108 1415 -74
rect 193 -170 227 -108
rect 1381 -170 1415 -108
rect 291 -210 307 -176
rect 341 -210 357 -176
rect 483 -210 499 -176
rect 533 -210 549 -176
rect 675 -210 691 -176
rect 725 -210 741 -176
rect 867 -210 883 -176
rect 917 -210 933 -176
rect 1059 -210 1075 -176
rect 1109 -210 1125 -176
rect 1251 -210 1267 -176
rect 1301 -210 1317 -176
rect 307 -270 341 -254
rect 307 -534 341 -518
rect 403 -270 437 -254
rect 403 -534 437 -518
rect 499 -270 533 -254
rect 499 -534 533 -518
rect 595 -270 629 -254
rect 595 -534 629 -518
rect 691 -270 725 -254
rect 691 -534 725 -518
rect 787 -270 821 -254
rect 787 -534 821 -518
rect 883 -270 917 -254
rect 883 -534 917 -518
rect 979 -270 1013 -254
rect 979 -534 1013 -518
rect 1075 -270 1109 -254
rect 1075 -534 1109 -518
rect 1171 -270 1205 -254
rect 1171 -534 1205 -518
rect 1267 -270 1301 -254
rect 1267 -534 1301 -518
rect 193 -618 227 -556
rect 1381 -618 1415 -556
rect 193 -652 289 -618
rect 1319 -652 1415 -618
rect 193 -760 289 -726
rect 1319 -760 1415 -726
rect 193 -822 227 -760
rect 1381 -820 1415 -760
rect 307 -850 341 -834
rect 307 -946 341 -930
rect 403 -850 437 -834
rect 403 -946 437 -930
rect 499 -850 533 -834
rect 499 -946 533 -930
rect 595 -850 629 -834
rect 595 -946 629 -930
rect 691 -850 725 -834
rect 691 -946 725 -930
rect 787 -850 821 -834
rect 787 -946 821 -930
rect 883 -850 917 -834
rect 883 -946 917 -930
rect 979 -850 1013 -834
rect 979 -946 1013 -930
rect 1075 -850 1109 -834
rect 1075 -946 1109 -930
rect 1171 -850 1205 -834
rect 1171 -946 1205 -930
rect 1267 -850 1301 -834
rect 1267 -946 1301 -930
rect 291 -1018 307 -984
rect 341 -1018 357 -984
rect 483 -1018 499 -984
rect 533 -1018 549 -984
rect 675 -1018 691 -984
rect 725 -1018 741 -984
rect 867 -1018 883 -984
rect 917 -1018 933 -984
rect 1059 -1018 1075 -984
rect 1109 -1018 1125 -984
rect 1251 -1018 1267 -984
rect 1301 -1018 1317 -984
rect 193 -1082 227 -1020
rect 1381 -1082 1415 -1020
rect 193 -1116 289 -1082
rect 1319 -1116 1415 -1082
<< viali >>
rect 313 942 347 976
rect 505 942 539 976
rect 697 942 731 976
rect 889 942 923 976
rect 1081 942 1115 976
rect 1273 942 1307 976
rect 313 634 347 882
rect 409 634 443 882
rect 505 634 539 882
rect 601 634 635 882
rect 697 634 731 882
rect 793 634 827 882
rect 889 634 923 882
rect 985 634 1019 882
rect 1081 634 1115 882
rect 1177 634 1211 882
rect 1273 634 1307 882
rect 1387 596 1421 982
rect 1387 330 1421 332
rect 313 222 347 302
rect 409 222 443 302
rect 505 222 539 302
rect 601 222 635 302
rect 697 222 731 302
rect 793 222 827 302
rect 889 222 923 302
rect 985 222 1019 302
rect 1081 222 1115 302
rect 1177 222 1211 302
rect 1273 222 1307 302
rect 313 134 347 168
rect 505 134 539 168
rect 697 134 731 168
rect 889 134 923 168
rect 1081 134 1115 168
rect 1273 134 1307 168
rect 1387 132 1421 330
rect 307 -210 341 -176
rect 499 -210 533 -176
rect 691 -210 725 -176
rect 883 -210 917 -176
rect 1075 -210 1109 -176
rect 1267 -210 1301 -176
rect 307 -518 341 -270
rect 403 -518 437 -270
rect 499 -518 533 -270
rect 595 -518 629 -270
rect 691 -518 725 -270
rect 787 -518 821 -270
rect 883 -518 917 -270
rect 979 -518 1013 -270
rect 1075 -518 1109 -270
rect 1171 -518 1205 -270
rect 1267 -518 1301 -270
rect 1381 -556 1415 -170
rect 1381 -822 1415 -820
rect 307 -930 341 -850
rect 403 -930 437 -850
rect 499 -930 533 -850
rect 595 -930 629 -850
rect 691 -930 725 -850
rect 787 -930 821 -850
rect 883 -930 917 -850
rect 979 -930 1013 -850
rect 1075 -930 1109 -850
rect 1171 -930 1205 -850
rect 1267 -930 1301 -850
rect 307 -1018 341 -984
rect 499 -1018 533 -984
rect 691 -1018 725 -984
rect 883 -1018 917 -984
rect 1075 -1018 1109 -984
rect 1267 -1018 1301 -984
rect 1381 -1020 1415 -822
<< metal1 >>
rect 129 1044 1211 1078
rect -133 934 27 986
rect 79 934 89 986
rect -300 438 -238 490
rect -186 438 -176 490
rect -298 -38 -236 14
rect -184 -38 -174 14
rect -133 -326 -81 934
rect -10 438 0 490
rect 52 481 62 490
rect 129 481 163 1044
rect 294 934 304 986
rect 356 934 366 986
rect 409 894 443 1044
rect 487 934 497 986
rect 549 934 559 986
rect 601 894 635 1044
rect 678 934 688 986
rect 740 934 750 986
rect 793 894 827 1044
rect 870 934 880 986
rect 932 934 942 986
rect 985 894 1019 1044
rect 1062 934 1072 986
rect 1124 934 1134 986
rect 1177 894 1211 1044
rect 1381 1062 1892 1114
rect 1254 934 1264 986
rect 1316 934 1326 986
rect 1381 982 1427 1062
rect 307 882 353 894
rect 307 634 313 882
rect 347 634 353 882
rect 307 622 353 634
rect 403 882 449 894
rect 403 634 409 882
rect 443 634 449 882
rect 403 622 449 634
rect 499 882 545 894
rect 499 634 505 882
rect 539 634 545 882
rect 499 622 545 634
rect 595 882 641 894
rect 595 634 601 882
rect 635 634 641 882
rect 595 622 641 634
rect 691 882 737 894
rect 691 634 697 882
rect 731 634 737 882
rect 691 622 737 634
rect 787 882 833 894
rect 787 634 793 882
rect 827 634 833 882
rect 787 622 833 634
rect 883 882 929 894
rect 883 634 889 882
rect 923 634 929 882
rect 883 622 929 634
rect 979 882 1025 894
rect 979 634 985 882
rect 1019 634 1025 882
rect 979 622 1025 634
rect 1075 882 1121 894
rect 1075 634 1081 882
rect 1115 634 1121 882
rect 1075 622 1121 634
rect 1171 882 1217 894
rect 1171 634 1177 882
rect 1211 634 1217 882
rect 1171 622 1217 634
rect 1267 882 1313 894
rect 1267 634 1273 882
rect 1307 634 1313 882
rect 1267 622 1313 634
rect 52 447 163 481
rect 52 438 62 447
rect -31 127 27 179
rect 79 127 89 179
rect -31 14 21 127
rect 129 70 163 447
rect 313 481 347 622
rect 505 481 539 622
rect 697 481 731 622
rect 889 481 923 622
rect 1081 481 1115 622
rect 1273 481 1307 622
rect 1381 596 1387 982
rect 1421 630 1427 982
rect 1421 596 1727 630
rect 1381 584 1427 596
rect 313 447 1530 481
rect 313 314 347 447
rect 505 314 539 447
rect 697 314 731 447
rect 889 314 923 447
rect 1081 314 1115 447
rect 1273 314 1307 447
rect 1381 333 1427 344
rect 307 302 353 314
rect 307 222 313 302
rect 347 222 353 302
rect 307 210 353 222
rect 403 302 449 314
rect 403 222 409 302
rect 443 222 449 302
rect 403 210 449 222
rect 499 302 545 314
rect 499 222 505 302
rect 539 222 545 302
rect 499 210 545 222
rect 595 302 641 314
rect 595 222 601 302
rect 635 222 641 302
rect 595 210 641 222
rect 691 302 737 314
rect 691 222 697 302
rect 731 222 737 302
rect 691 210 737 222
rect 787 302 833 314
rect 787 222 793 302
rect 827 222 833 302
rect 787 210 833 222
rect 883 302 929 314
rect 883 222 889 302
rect 923 222 929 302
rect 883 210 929 222
rect 979 302 1025 314
rect 979 222 985 302
rect 1019 222 1025 302
rect 979 210 1025 222
rect 1075 302 1121 314
rect 1075 222 1081 302
rect 1115 222 1121 302
rect 1075 210 1121 222
rect 1171 302 1217 314
rect 1171 222 1177 302
rect 1211 222 1217 302
rect 1171 210 1217 222
rect 1267 302 1313 314
rect 1267 222 1273 302
rect 1307 222 1313 302
rect 1368 281 1378 333
rect 1430 281 1440 333
rect 1267 210 1313 222
rect 297 179 363 182
rect 294 127 304 179
rect 356 127 366 179
rect 297 122 363 127
rect 409 70 443 210
rect 489 179 555 182
rect 485 127 495 179
rect 547 127 557 179
rect 489 122 555 127
rect 601 70 635 210
rect 681 179 747 182
rect 677 127 687 179
rect 739 127 749 179
rect 681 122 747 127
rect 793 70 827 210
rect 873 179 939 182
rect 869 127 879 179
rect 931 127 941 179
rect 873 122 939 127
rect 985 70 1019 210
rect 1065 178 1131 182
rect 1062 126 1072 178
rect 1124 126 1134 178
rect 1065 122 1131 126
rect 1177 70 1211 210
rect 1257 178 1323 182
rect 1254 126 1264 178
rect 1316 126 1326 178
rect 1381 132 1387 281
rect 1421 132 1427 281
rect 1257 122 1323 126
rect 129 36 1211 70
rect -41 -38 -31 14
rect 21 -38 31 14
rect 1381 0 1427 132
rect 1496 5 1530 447
rect 1571 281 1581 333
rect 1633 281 1643 333
rect -31 -218 21 -38
rect 123 -108 1205 -74
rect 73 -218 83 -166
rect -313 -378 -81 -326
rect -300 -715 -238 -663
rect -186 -715 -176 -663
rect -133 -973 -81 -378
rect -17 -715 -7 -663
rect 45 -671 55 -663
rect 123 -671 157 -108
rect 288 -218 298 -166
rect 350 -218 360 -166
rect 403 -258 437 -108
rect 481 -218 491 -166
rect 543 -218 553 -166
rect 595 -258 629 -108
rect 672 -218 682 -166
rect 734 -218 744 -166
rect 787 -258 821 -108
rect 864 -218 874 -166
rect 926 -218 936 -166
rect 979 -258 1013 -108
rect 1056 -218 1066 -166
rect 1118 -218 1128 -166
rect 1171 -258 1205 -108
rect 1248 -218 1258 -166
rect 1310 -218 1320 -166
rect 1375 -170 1421 -38
rect 1477 -47 1487 5
rect 1539 -47 1549 5
rect 301 -270 347 -258
rect 301 -518 307 -270
rect 341 -518 347 -270
rect 301 -530 347 -518
rect 397 -270 443 -258
rect 397 -518 403 -270
rect 437 -518 443 -270
rect 397 -530 443 -518
rect 493 -270 539 -258
rect 493 -518 499 -270
rect 533 -518 539 -270
rect 493 -530 539 -518
rect 589 -270 635 -258
rect 589 -518 595 -270
rect 629 -518 635 -270
rect 589 -530 635 -518
rect 685 -270 731 -258
rect 685 -518 691 -270
rect 725 -518 731 -270
rect 685 -530 731 -518
rect 781 -270 827 -258
rect 781 -518 787 -270
rect 821 -518 827 -270
rect 781 -530 827 -518
rect 877 -270 923 -258
rect 877 -518 883 -270
rect 917 -518 923 -270
rect 877 -530 923 -518
rect 973 -270 1019 -258
rect 973 -518 979 -270
rect 1013 -518 1019 -270
rect 973 -530 1019 -518
rect 1069 -270 1115 -258
rect 1069 -518 1075 -270
rect 1109 -518 1115 -270
rect 1069 -530 1115 -518
rect 1165 -270 1211 -258
rect 1165 -518 1171 -270
rect 1205 -518 1211 -270
rect 1165 -530 1211 -518
rect 1261 -270 1307 -258
rect 1261 -518 1267 -270
rect 1301 -518 1307 -270
rect 1375 -505 1381 -170
rect 1415 -505 1421 -170
rect 1261 -530 1307 -518
rect 45 -705 157 -671
rect 45 -715 55 -705
rect -133 -1025 21 -973
rect 73 -1025 83 -973
rect 123 -1082 157 -705
rect 307 -671 341 -530
rect 499 -671 533 -530
rect 691 -671 725 -530
rect 883 -671 917 -530
rect 1075 -671 1109 -530
rect 1267 -671 1301 -530
rect 1362 -557 1372 -505
rect 1424 -557 1434 -505
rect 1375 -568 1421 -557
rect 1496 -671 1530 -47
rect 307 -705 1530 -671
rect 307 -838 341 -705
rect 499 -838 533 -705
rect 691 -838 725 -705
rect 883 -838 917 -705
rect 1075 -838 1109 -705
rect 1267 -838 1301 -705
rect 1375 -820 1421 -808
rect 1590 -820 1624 281
rect 1693 -505 1727 596
rect 1782 -47 1792 5
rect 1844 -47 1895 5
rect 1674 -557 1684 -505
rect 1736 -557 1746 -505
rect 301 -850 347 -838
rect 301 -930 307 -850
rect 341 -930 347 -850
rect 301 -942 347 -930
rect 397 -850 443 -838
rect 397 -930 403 -850
rect 437 -930 443 -850
rect 397 -942 443 -930
rect 493 -850 539 -838
rect 493 -930 499 -850
rect 533 -930 539 -850
rect 493 -942 539 -930
rect 589 -850 635 -838
rect 589 -930 595 -850
rect 629 -930 635 -850
rect 589 -942 635 -930
rect 685 -850 731 -838
rect 685 -930 691 -850
rect 725 -930 731 -850
rect 685 -942 731 -930
rect 781 -850 827 -838
rect 781 -930 787 -850
rect 821 -930 827 -850
rect 781 -942 827 -930
rect 877 -850 923 -838
rect 877 -930 883 -850
rect 917 -930 923 -850
rect 877 -942 923 -930
rect 973 -850 1019 -838
rect 973 -930 979 -850
rect 1013 -930 1019 -850
rect 973 -942 1019 -930
rect 1069 -850 1115 -838
rect 1069 -930 1075 -850
rect 1109 -930 1115 -850
rect 1069 -942 1115 -930
rect 1165 -850 1211 -838
rect 1165 -930 1171 -850
rect 1205 -930 1211 -850
rect 1165 -942 1211 -930
rect 1261 -850 1307 -838
rect 1261 -930 1267 -850
rect 1301 -930 1307 -850
rect 1261 -942 1307 -930
rect 291 -973 357 -970
rect 288 -1025 298 -973
rect 350 -1025 360 -973
rect 291 -1030 357 -1025
rect 403 -1082 437 -942
rect 483 -973 549 -970
rect 479 -1025 489 -973
rect 541 -1025 551 -973
rect 483 -1030 549 -1025
rect 595 -1082 629 -942
rect 675 -973 741 -970
rect 671 -1025 681 -973
rect 733 -1025 743 -973
rect 675 -1030 741 -1025
rect 787 -1082 821 -942
rect 867 -973 933 -970
rect 863 -1025 873 -973
rect 925 -1025 935 -973
rect 867 -1030 933 -1025
rect 979 -1082 1013 -942
rect 1059 -974 1125 -970
rect 1056 -1026 1066 -974
rect 1118 -1026 1128 -974
rect 1059 -1030 1125 -1026
rect 1171 -1082 1205 -942
rect 1251 -974 1317 -970
rect 1248 -1026 1258 -974
rect 1310 -1026 1320 -974
rect 1375 -1020 1381 -820
rect 1415 -854 1624 -820
rect 1415 -1020 1421 -854
rect 1251 -1030 1317 -1026
rect 123 -1116 1205 -1082
rect 1375 -1102 1421 -1020
rect 1374 -1154 1885 -1102
<< via1 >>
rect 27 934 79 986
rect -238 438 -186 490
rect -236 -38 -184 14
rect 0 438 52 490
rect 304 976 356 986
rect 304 942 313 976
rect 313 942 347 976
rect 347 942 356 976
rect 304 934 356 942
rect 497 976 549 986
rect 497 942 505 976
rect 505 942 539 976
rect 539 942 549 976
rect 497 934 549 942
rect 688 976 740 986
rect 688 942 697 976
rect 697 942 731 976
rect 731 942 740 976
rect 688 934 740 942
rect 880 976 932 986
rect 880 942 889 976
rect 889 942 923 976
rect 923 942 932 976
rect 880 934 932 942
rect 1072 976 1124 986
rect 1072 942 1081 976
rect 1081 942 1115 976
rect 1115 942 1124 976
rect 1072 934 1124 942
rect 1264 976 1316 986
rect 1264 942 1273 976
rect 1273 942 1307 976
rect 1307 942 1316 976
rect 1264 934 1316 942
rect 27 127 79 179
rect 1378 332 1430 333
rect 1378 281 1387 332
rect 1387 281 1421 332
rect 1421 281 1430 332
rect 304 168 356 179
rect 304 134 313 168
rect 313 134 347 168
rect 347 134 356 168
rect 304 127 356 134
rect 495 168 547 179
rect 495 134 505 168
rect 505 134 539 168
rect 539 134 547 168
rect 495 127 547 134
rect 687 168 739 179
rect 687 134 697 168
rect 697 134 731 168
rect 731 134 739 168
rect 687 127 739 134
rect 879 168 931 179
rect 879 134 889 168
rect 889 134 923 168
rect 923 134 931 168
rect 879 127 931 134
rect 1072 168 1124 178
rect 1072 134 1081 168
rect 1081 134 1115 168
rect 1115 134 1124 168
rect 1072 126 1124 134
rect 1264 168 1316 178
rect 1264 134 1273 168
rect 1273 134 1307 168
rect 1307 134 1316 168
rect 1264 126 1316 134
rect -31 -38 21 14
rect 1581 281 1633 333
rect 21 -218 73 -166
rect -238 -715 -186 -663
rect -7 -715 45 -663
rect 298 -176 350 -166
rect 298 -210 307 -176
rect 307 -210 341 -176
rect 341 -210 350 -176
rect 298 -218 350 -210
rect 491 -176 543 -166
rect 491 -210 499 -176
rect 499 -210 533 -176
rect 533 -210 543 -176
rect 491 -218 543 -210
rect 682 -176 734 -166
rect 682 -210 691 -176
rect 691 -210 725 -176
rect 725 -210 734 -176
rect 682 -218 734 -210
rect 874 -176 926 -166
rect 874 -210 883 -176
rect 883 -210 917 -176
rect 917 -210 926 -176
rect 874 -218 926 -210
rect 1066 -176 1118 -166
rect 1066 -210 1075 -176
rect 1075 -210 1109 -176
rect 1109 -210 1118 -176
rect 1066 -218 1118 -210
rect 1258 -176 1310 -166
rect 1258 -210 1267 -176
rect 1267 -210 1301 -176
rect 1301 -210 1310 -176
rect 1258 -218 1310 -210
rect 1487 -47 1539 5
rect 21 -1025 73 -973
rect 1372 -556 1381 -505
rect 1381 -556 1415 -505
rect 1415 -556 1424 -505
rect 1372 -557 1424 -556
rect 1792 -47 1844 5
rect 1684 -557 1736 -505
rect 298 -984 350 -973
rect 298 -1018 307 -984
rect 307 -1018 341 -984
rect 341 -1018 350 -984
rect 298 -1025 350 -1018
rect 489 -984 541 -973
rect 489 -1018 499 -984
rect 499 -1018 533 -984
rect 533 -1018 541 -984
rect 489 -1025 541 -1018
rect 681 -984 733 -973
rect 681 -1018 691 -984
rect 691 -1018 725 -984
rect 725 -1018 733 -984
rect 681 -1025 733 -1018
rect 873 -984 925 -973
rect 873 -1018 883 -984
rect 883 -1018 917 -984
rect 917 -1018 925 -984
rect 873 -1025 925 -1018
rect 1066 -984 1118 -974
rect 1066 -1018 1075 -984
rect 1075 -1018 1109 -984
rect 1109 -1018 1118 -984
rect 1066 -1026 1118 -1018
rect 1258 -984 1310 -974
rect 1258 -1018 1267 -984
rect 1267 -1018 1301 -984
rect 1301 -1018 1310 -984
rect 1258 -1026 1310 -1018
<< metal2 >>
rect 27 986 79 996
rect 304 986 356 996
rect 497 986 549 996
rect 688 986 740 996
rect 880 986 932 996
rect 1072 986 1124 996
rect 1264 986 1316 996
rect 79 934 304 986
rect 356 934 497 986
rect 549 934 688 986
rect 740 934 880 986
rect 932 934 1072 986
rect 1124 934 1264 986
rect 1316 934 1323 986
rect 27 924 79 934
rect 304 924 356 934
rect 497 924 549 934
rect 688 924 740 934
rect 880 924 932 934
rect 1072 924 1124 934
rect 1264 924 1316 934
rect -238 490 -186 500
rect 0 490 52 500
rect -186 438 0 490
rect -238 428 -186 438
rect 0 428 52 438
rect 1378 333 1430 343
rect 1581 333 1633 343
rect 1430 281 1581 333
rect 1378 271 1430 281
rect 1581 271 1633 281
rect 27 179 79 189
rect 304 179 356 189
rect 495 179 547 189
rect 687 179 739 189
rect 879 179 931 189
rect 1072 179 1124 188
rect 1264 179 1316 188
rect 79 127 304 179
rect 356 127 495 179
rect 547 127 687 179
rect 739 127 879 179
rect 931 178 1323 179
rect 931 127 1072 178
rect 27 117 79 127
rect 304 117 356 127
rect 495 117 547 127
rect 687 117 739 127
rect 879 117 931 127
rect 1124 127 1264 178
rect 1072 116 1124 126
rect 1316 127 1323 178
rect 1264 116 1316 126
rect -236 14 -184 24
rect -31 14 21 24
rect -184 -38 -31 14
rect -236 -48 -184 -38
rect -31 -48 21 -38
rect 1487 5 1539 15
rect 1792 5 1844 15
rect 1539 -47 1792 5
rect 1487 -57 1539 -47
rect 1792 -57 1844 -47
rect 21 -166 73 -156
rect 298 -166 350 -156
rect 491 -166 543 -156
rect 682 -166 734 -156
rect 874 -166 926 -156
rect 1066 -166 1118 -156
rect 1258 -166 1310 -156
rect 73 -218 298 -166
rect 350 -218 491 -166
rect 543 -218 682 -166
rect 734 -218 874 -166
rect 926 -218 1066 -166
rect 1118 -218 1258 -166
rect 1310 -218 1317 -166
rect 21 -228 73 -218
rect 298 -228 350 -218
rect 491 -228 543 -218
rect 682 -228 734 -218
rect 874 -228 926 -218
rect 1066 -228 1118 -218
rect 1258 -228 1310 -218
rect 1372 -505 1424 -495
rect 1684 -505 1736 -495
rect 1424 -557 1684 -505
rect 1372 -567 1424 -557
rect 1684 -567 1736 -557
rect -238 -663 -186 -653
rect -7 -663 45 -653
rect -186 -715 -7 -663
rect -238 -725 -186 -715
rect -7 -725 45 -715
rect 21 -973 73 -963
rect 298 -973 350 -963
rect 489 -973 541 -963
rect 681 -973 733 -963
rect 873 -973 925 -963
rect 1066 -973 1118 -964
rect 1258 -973 1310 -964
rect 73 -1025 298 -973
rect 350 -1025 489 -973
rect 541 -1025 681 -973
rect 733 -1025 873 -973
rect 925 -974 1317 -973
rect 925 -1025 1066 -974
rect 21 -1035 73 -1025
rect 298 -1035 350 -1025
rect 489 -1035 541 -1025
rect 681 -1035 733 -1025
rect 873 -1035 925 -1025
rect 1118 -1025 1258 -974
rect 1066 -1036 1118 -1026
rect 1310 -1025 1317 -974
rect 1258 -1036 1310 -1026
<< labels >>
flabel metal1 -285 464 -285 464 1 FreeSans 400 0 0 0 v_hi
port 1 n
flabel metal1 -280 -690 -280 -690 1 FreeSans 400 0 0 0 v_lo
port 2 n
flabel metal1 -275 -14 -275 -14 1 FreeSans 400 0 0 0 v
port 3 n
flabel metal1 -286 -352 -286 -352 1 FreeSans 400 0 0 0 v_b
port 4 n
flabel metal1 1879 -24 1879 -24 1 FreeSans 400 0 0 0 out
port 5 n
flabel metal1 1868 1086 1868 1086 1 FreeSans 400 0 0 0 VDD
port 6 n power bidirectional
flabel metal1 1867 -1131 1867 -1131 1 FreeSans 400 0 0 0 VSS
port 7 n ground bidirectional
flabel metal1 -1 -192 -1 -192 3 FreeSans 400 0 0 0 transmission_gate_1/en_b
flabel metal1 -2 -688 -2 -688 3 FreeSans 400 0 0 0 transmission_gate_1/in
flabel metal1 -2 -999 -2 -999 3 FreeSans 400 0 0 0 transmission_gate_1/en
flabel metal1 1489 -689 1489 -689 7 FreeSans 400 0 0 0 transmission_gate_1/out
flabel metal1 1398 -43 1398 -43 5 FreeSans 400 0 0 0 transmission_gate_1/VDD
flabel metal1 1398 -1149 1398 -1149 1 FreeSans 400 0 0 0 transmission_gate_1/VSS
flabel metal1 5 960 5 960 3 FreeSans 400 0 0 0 transmission_gate_0/en_b
flabel metal1 4 464 4 464 3 FreeSans 400 0 0 0 transmission_gate_0/in
flabel metal1 4 153 4 153 3 FreeSans 400 0 0 0 transmission_gate_0/en
flabel metal1 1495 463 1495 463 7 FreeSans 400 0 0 0 transmission_gate_0/out
flabel metal1 1404 1109 1404 1109 5 FreeSans 400 0 0 0 transmission_gate_0/VDD
flabel metal1 1404 3 1404 3 1 FreeSans 400 0 0 0 transmission_gate_0/VSS
<< end >>
