magic
tech sky130A
timestamp 1653453365
<< metal3 >>
rect -315 -290 264 290
<< mimcap >>
rect -265 220 215 240
rect -265 -220 -245 220
rect 195 -220 215 220
rect -265 -240 215 -220
<< mimcapcontact >>
rect -245 -220 195 220
<< properties >>
string FIXED_BBOX -315 -290 265 290
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.799 l 4.799 val 49.726 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
