magic
tech sky130A
magscale 1 2
timestamp 1654644491
<< nmos >>
rect -1217 -140 -1097 140
rect -1039 -140 -919 140
rect -861 -140 -741 140
rect -683 -140 -563 140
rect -505 -140 -385 140
rect -327 -140 -207 140
rect -149 -140 -29 140
rect 29 -140 149 140
rect 207 -140 327 140
rect 385 -140 505 140
rect 563 -140 683 140
rect 741 -140 861 140
rect 919 -140 1039 140
rect 1097 -140 1217 140
<< ndiff >>
rect -1275 128 -1217 140
rect -1275 -128 -1263 128
rect -1229 -128 -1217 128
rect -1275 -140 -1217 -128
rect -1097 128 -1039 140
rect -1097 -128 -1085 128
rect -1051 -128 -1039 128
rect -1097 -140 -1039 -128
rect -919 128 -861 140
rect -919 -128 -907 128
rect -873 -128 -861 128
rect -919 -140 -861 -128
rect -741 128 -683 140
rect -741 -128 -729 128
rect -695 -128 -683 128
rect -741 -140 -683 -128
rect -563 128 -505 140
rect -563 -128 -551 128
rect -517 -128 -505 128
rect -563 -140 -505 -128
rect -385 128 -327 140
rect -385 -128 -373 128
rect -339 -128 -327 128
rect -385 -140 -327 -128
rect -207 128 -149 140
rect -207 -128 -195 128
rect -161 -128 -149 128
rect -207 -140 -149 -128
rect -29 128 29 140
rect -29 -128 -17 128
rect 17 -128 29 128
rect -29 -140 29 -128
rect 149 128 207 140
rect 149 -128 161 128
rect 195 -128 207 128
rect 149 -140 207 -128
rect 327 128 385 140
rect 327 -128 339 128
rect 373 -128 385 128
rect 327 -140 385 -128
rect 505 128 563 140
rect 505 -128 517 128
rect 551 -128 563 128
rect 505 -140 563 -128
rect 683 128 741 140
rect 683 -128 695 128
rect 729 -128 741 128
rect 683 -140 741 -128
rect 861 128 919 140
rect 861 -128 873 128
rect 907 -128 919 128
rect 861 -140 919 -128
rect 1039 128 1097 140
rect 1039 -128 1051 128
rect 1085 -128 1097 128
rect 1039 -140 1097 -128
rect 1217 128 1275 140
rect 1217 -128 1229 128
rect 1263 -128 1275 128
rect 1217 -140 1275 -128
<< ndiffc >>
rect -1263 -128 -1229 128
rect -1085 -128 -1051 128
rect -907 -128 -873 128
rect -729 -128 -695 128
rect -551 -128 -517 128
rect -373 -128 -339 128
rect -195 -128 -161 128
rect -17 -128 17 128
rect 161 -128 195 128
rect 339 -128 373 128
rect 517 -128 551 128
rect 695 -128 729 128
rect 873 -128 907 128
rect 1051 -128 1085 128
rect 1229 -128 1263 128
<< poly >>
rect -1199 212 -1115 228
rect -1199 195 -1183 212
rect -1217 178 -1183 195
rect -1131 195 -1115 212
rect -1021 212 -937 228
rect -1021 195 -1005 212
rect -1131 178 -1097 195
rect -1217 140 -1097 178
rect -1039 178 -1005 195
rect -953 195 -937 212
rect -843 212 -759 228
rect -843 195 -827 212
rect -953 178 -919 195
rect -1039 140 -919 178
rect -861 178 -827 195
rect -775 195 -759 212
rect -665 212 -581 228
rect -665 195 -649 212
rect -775 178 -741 195
rect -861 140 -741 178
rect -683 178 -649 195
rect -597 195 -581 212
rect -487 212 -403 228
rect -487 195 -471 212
rect -597 178 -563 195
rect -683 140 -563 178
rect -505 178 -471 195
rect -419 195 -403 212
rect -309 212 -225 228
rect -309 195 -293 212
rect -419 178 -385 195
rect -505 140 -385 178
rect -327 178 -293 195
rect -241 195 -225 212
rect -131 212 -47 228
rect -131 195 -115 212
rect -241 178 -207 195
rect -327 140 -207 178
rect -149 178 -115 195
rect -63 195 -47 212
rect 47 212 131 228
rect 47 195 63 212
rect -63 178 -29 195
rect -149 140 -29 178
rect 29 178 63 195
rect 115 195 131 212
rect 225 212 309 228
rect 225 195 241 212
rect 115 178 149 195
rect 29 140 149 178
rect 207 178 241 195
rect 293 195 309 212
rect 403 212 487 228
rect 403 195 419 212
rect 293 178 327 195
rect 207 140 327 178
rect 385 178 419 195
rect 471 195 487 212
rect 581 212 665 228
rect 581 195 597 212
rect 471 178 505 195
rect 385 140 505 178
rect 563 178 597 195
rect 649 195 665 212
rect 759 212 843 228
rect 759 195 775 212
rect 649 178 683 195
rect 563 140 683 178
rect 741 178 775 195
rect 827 195 843 212
rect 937 212 1021 228
rect 937 195 953 212
rect 827 178 861 195
rect 741 140 861 178
rect 919 178 953 195
rect 1005 195 1021 212
rect 1115 212 1199 228
rect 1115 195 1131 212
rect 1005 178 1039 195
rect 919 140 1039 178
rect 1097 178 1131 195
rect 1183 195 1199 212
rect 1183 178 1217 195
rect 1097 140 1217 178
rect -1217 -178 -1097 -140
rect -1217 -195 -1183 -178
rect -1199 -212 -1183 -195
rect -1131 -195 -1097 -178
rect -1039 -178 -919 -140
rect -1039 -195 -1005 -178
rect -1131 -212 -1115 -195
rect -1199 -228 -1115 -212
rect -1021 -212 -1005 -195
rect -953 -195 -919 -178
rect -861 -178 -741 -140
rect -861 -195 -827 -178
rect -953 -212 -937 -195
rect -1021 -228 -937 -212
rect -843 -212 -827 -195
rect -775 -195 -741 -178
rect -683 -178 -563 -140
rect -683 -195 -649 -178
rect -775 -212 -759 -195
rect -843 -228 -759 -212
rect -665 -212 -649 -195
rect -597 -195 -563 -178
rect -505 -178 -385 -140
rect -505 -195 -471 -178
rect -597 -212 -581 -195
rect -665 -228 -581 -212
rect -487 -212 -471 -195
rect -419 -195 -385 -178
rect -327 -178 -207 -140
rect -327 -195 -293 -178
rect -419 -212 -403 -195
rect -487 -228 -403 -212
rect -309 -212 -293 -195
rect -241 -195 -207 -178
rect -149 -178 -29 -140
rect -149 -195 -115 -178
rect -241 -212 -225 -195
rect -309 -228 -225 -212
rect -131 -212 -115 -195
rect -63 -195 -29 -178
rect 29 -178 149 -140
rect 29 -195 63 -178
rect -63 -212 -47 -195
rect -131 -228 -47 -212
rect 47 -212 63 -195
rect 115 -195 149 -178
rect 207 -178 327 -140
rect 207 -195 241 -178
rect 115 -212 131 -195
rect 47 -228 131 -212
rect 225 -212 241 -195
rect 293 -195 327 -178
rect 385 -178 505 -140
rect 385 -195 419 -178
rect 293 -212 309 -195
rect 225 -228 309 -212
rect 403 -212 419 -195
rect 471 -195 505 -178
rect 563 -178 683 -140
rect 563 -195 597 -178
rect 471 -212 487 -195
rect 403 -228 487 -212
rect 581 -212 597 -195
rect 649 -195 683 -178
rect 741 -178 861 -140
rect 741 -195 775 -178
rect 649 -212 665 -195
rect 581 -228 665 -212
rect 759 -212 775 -195
rect 827 -195 861 -178
rect 919 -178 1039 -140
rect 919 -195 953 -178
rect 827 -212 843 -195
rect 759 -228 843 -212
rect 937 -212 953 -195
rect 1005 -195 1039 -178
rect 1097 -178 1217 -140
rect 1097 -195 1131 -178
rect 1005 -212 1021 -195
rect 937 -228 1021 -212
rect 1115 -212 1131 -195
rect 1183 -195 1217 -178
rect 1183 -212 1199 -195
rect 1115 -228 1199 -212
<< polycont >>
rect -1183 178 -1131 212
rect -1005 178 -953 212
rect -827 178 -775 212
rect -649 178 -597 212
rect -471 178 -419 212
rect -293 178 -241 212
rect -115 178 -63 212
rect 63 178 115 212
rect 241 178 293 212
rect 419 178 471 212
rect 597 178 649 212
rect 775 178 827 212
rect 953 178 1005 212
rect 1131 178 1183 212
rect -1183 -212 -1131 -178
rect -1005 -212 -953 -178
rect -827 -212 -775 -178
rect -649 -212 -597 -178
rect -471 -212 -419 -178
rect -293 -212 -241 -178
rect -115 -212 -63 -178
rect 63 -212 115 -178
rect 241 -212 293 -178
rect 419 -212 471 -178
rect 597 -212 649 -178
rect 775 -212 827 -178
rect 953 -212 1005 -178
rect 1131 -212 1183 -178
<< locali >>
rect -1263 178 -1183 212
rect -1131 178 -1115 212
rect -1021 178 -1005 212
rect -953 178 -937 212
rect -843 178 -827 212
rect -775 178 -759 212
rect -665 178 -649 212
rect -597 178 -581 212
rect -487 178 -471 212
rect -419 178 -403 212
rect -309 178 -293 212
rect -241 178 -225 212
rect -131 178 -115 212
rect -63 178 -47 212
rect 47 178 63 212
rect 115 178 131 212
rect 225 178 241 212
rect 293 178 309 212
rect 403 178 419 212
rect 471 178 487 212
rect 581 178 597 212
rect 649 178 665 212
rect 759 178 775 212
rect 827 178 843 212
rect 937 178 953 212
rect 1005 178 1021 212
rect 1115 178 1131 212
rect 1183 178 1263 212
rect -1263 128 -1229 178
rect -1263 -178 -1229 -128
rect -1085 128 -1051 144
rect -1085 -144 -1051 -128
rect -907 128 -873 144
rect -907 -144 -873 -128
rect -729 128 -695 144
rect -729 -144 -695 -128
rect -551 128 -517 144
rect -551 -144 -517 -128
rect -373 128 -339 144
rect -373 -144 -339 -128
rect -195 128 -161 144
rect -195 -144 -161 -128
rect -17 128 17 144
rect -17 -144 17 -128
rect 161 128 195 144
rect 161 -144 195 -128
rect 339 128 373 144
rect 339 -144 373 -128
rect 517 128 551 144
rect 517 -144 551 -128
rect 695 128 729 144
rect 695 -144 729 -128
rect 873 128 907 144
rect 873 -144 907 -128
rect 1051 128 1085 144
rect 1051 -144 1085 -128
rect 1229 128 1263 178
rect 1229 -178 1263 -128
rect -1263 -212 -1183 -178
rect -1131 -212 -1115 -178
rect -1021 -212 -1005 -178
rect -953 -212 -937 -178
rect -843 -212 -827 -178
rect -775 -212 -759 -178
rect -665 -212 -649 -178
rect -597 -212 -581 -178
rect -487 -212 -471 -178
rect -419 -212 -403 -178
rect -309 -212 -293 -178
rect -241 -212 -225 -178
rect -131 -212 -115 -178
rect -63 -212 -47 -178
rect 47 -212 63 -178
rect 115 -212 131 -178
rect 225 -212 241 -178
rect 293 -212 309 -178
rect 403 -212 419 -178
rect 471 -212 487 -178
rect 581 -212 597 -178
rect 649 -212 665 -178
rect 759 -212 775 -178
rect 827 -212 843 -178
rect 937 -212 953 -178
rect 1005 -212 1021 -178
rect 1115 -212 1131 -178
rect 1183 -212 1263 -178
<< viali >>
rect -1005 178 -953 212
rect -827 178 -775 212
rect -649 178 -597 212
rect -471 178 -419 212
rect -293 178 -241 212
rect -115 178 -63 212
rect 63 178 115 212
rect 241 178 293 212
rect 419 178 471 212
rect 597 178 649 212
rect 775 178 827 212
rect 953 178 1005 212
rect -1005 -212 -953 -178
rect -827 -212 -775 -178
rect -649 -212 -597 -178
rect -471 -212 -419 -178
rect -293 -212 -241 -178
rect -115 -212 -63 -178
rect 63 -212 115 -178
rect 241 -212 293 -178
rect 419 -212 471 -178
rect 597 -212 649 -178
rect 775 -212 827 -178
rect 953 -212 1005 -178
<< metal1 >>
rect -1017 212 -941 218
rect -1017 178 -1005 212
rect -953 178 -941 212
rect -1017 172 -941 178
rect -839 212 -763 218
rect -839 178 -827 212
rect -775 178 -763 212
rect -839 172 -763 178
rect -661 212 -585 218
rect -661 178 -649 212
rect -597 178 -585 212
rect -661 172 -585 178
rect -483 212 -407 218
rect -483 178 -471 212
rect -419 178 -407 212
rect -483 172 -407 178
rect -305 212 -229 218
rect -305 178 -293 212
rect -241 178 -229 212
rect -305 172 -229 178
rect -127 212 -51 218
rect -127 178 -115 212
rect -63 178 -51 212
rect -127 172 -51 178
rect 51 212 127 218
rect 51 178 63 212
rect 115 178 127 212
rect 51 172 127 178
rect 229 212 305 218
rect 229 178 241 212
rect 293 178 305 212
rect 229 172 305 178
rect 407 212 483 218
rect 407 178 419 212
rect 471 178 483 212
rect 407 172 483 178
rect 585 212 661 218
rect 585 178 597 212
rect 649 178 661 212
rect 585 172 661 178
rect 763 212 839 218
rect 763 178 775 212
rect 827 178 839 212
rect 763 172 839 178
rect 941 212 1017 218
rect 941 178 953 212
rect 1005 178 1017 212
rect 941 172 1017 178
rect -1017 -178 -941 -172
rect -1017 -212 -1005 -178
rect -953 -212 -941 -178
rect -1017 -218 -941 -212
rect -839 -178 -763 -172
rect -839 -212 -827 -178
rect -775 -212 -763 -178
rect -839 -218 -763 -212
rect -661 -178 -585 -172
rect -661 -212 -649 -178
rect -597 -212 -585 -178
rect -661 -218 -585 -212
rect -483 -178 -407 -172
rect -483 -212 -471 -178
rect -419 -212 -407 -178
rect -483 -218 -407 -212
rect -305 -178 -229 -172
rect -305 -212 -293 -178
rect -241 -212 -229 -178
rect -305 -218 -229 -212
rect -127 -178 -51 -172
rect -127 -212 -115 -178
rect -63 -212 -51 -178
rect -127 -218 -51 -212
rect 51 -178 127 -172
rect 51 -212 63 -178
rect 115 -212 127 -178
rect 51 -218 127 -212
rect 229 -178 305 -172
rect 229 -212 241 -178
rect 293 -212 305 -178
rect 229 -218 305 -212
rect 407 -178 483 -172
rect 407 -212 419 -178
rect 471 -212 483 -178
rect 407 -218 483 -212
rect 585 -178 661 -172
rect 585 -212 597 -178
rect 649 -212 661 -178
rect 585 -218 661 -212
rect 763 -178 839 -172
rect 763 -212 775 -178
rect 827 -212 839 -178
rect 763 -218 839 -212
rect 941 -178 1017 -172
rect 941 -212 953 -178
rect 1005 -212 1017 -178
rect 941 -218 1017 -212
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.4 l 0.6 m 1 nf 14 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 0 viadrn 0 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
