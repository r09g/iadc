magic
tech sky130A
timestamp 1653369027
<< pwell >>
rect -370 -130 370 130
<< nmos >>
rect -270 -25 -255 25
rect -165 -25 -150 25
rect -60 -25 -45 25
rect 45 -25 60 25
rect 150 -25 165 25
rect 255 -25 270 25
<< ndiff >>
rect -301 19 -270 25
rect -301 -19 -295 19
rect -278 -19 -270 19
rect -301 -25 -270 -19
rect -255 19 -224 25
rect -255 -19 -247 19
rect -230 -19 -224 19
rect -255 -25 -224 -19
rect -196 19 -165 25
rect -196 -19 -190 19
rect -173 -19 -165 19
rect -196 -25 -165 -19
rect -150 19 -119 25
rect -150 -19 -142 19
rect -125 -19 -119 19
rect -150 -25 -119 -19
rect -91 19 -60 25
rect -91 -19 -85 19
rect -68 -19 -60 19
rect -91 -25 -60 -19
rect -45 19 -14 25
rect -45 -19 -37 19
rect -20 -19 -14 19
rect -45 -25 -14 -19
rect 14 19 45 25
rect 14 -19 20 19
rect 37 -19 45 19
rect 14 -25 45 -19
rect 60 19 91 25
rect 60 -19 68 19
rect 85 -19 91 19
rect 60 -25 91 -19
rect 119 19 150 25
rect 119 -19 125 19
rect 142 -19 150 19
rect 119 -25 150 -19
rect 165 19 196 25
rect 165 -19 173 19
rect 190 -19 196 19
rect 165 -25 196 -19
rect 224 19 255 25
rect 224 -19 230 19
rect 247 -19 255 19
rect 224 -25 255 -19
rect 270 19 301 25
rect 270 -19 278 19
rect 295 -19 301 19
rect 270 -25 301 -19
<< ndiffc >>
rect -295 -19 -278 19
rect -247 -19 -230 19
rect -190 -19 -173 19
rect -142 -19 -125 19
rect -85 -19 -68 19
rect -37 -19 -20 19
rect 20 -19 37 19
rect 68 -19 85 19
rect 125 -19 142 19
rect 173 -19 190 19
rect 230 -19 247 19
rect 278 -19 295 19
<< psubdiff >>
rect -352 95 -304 112
rect 304 95 352 112
rect -352 64 -335 95
rect 335 64 352 95
rect -352 -95 -335 -64
rect 335 -95 352 -64
rect -352 -112 -304 -95
rect 304 -112 352 -95
<< psubdiffcont >>
rect -304 95 304 112
rect -352 -64 -335 64
rect 335 -64 352 64
rect -304 -112 304 -95
<< poly >>
rect -279 61 -246 69
rect -279 44 -271 61
rect -254 44 -246 61
rect -279 36 -246 44
rect -174 61 -141 69
rect -174 44 -166 61
rect -149 44 -141 61
rect -174 36 -141 44
rect 141 61 174 69
rect 141 44 149 61
rect 166 44 174 61
rect -270 25 -255 36
rect -165 25 -150 36
rect -60 25 -45 38
rect 45 25 60 38
rect 141 36 174 44
rect 246 61 279 69
rect 246 44 254 61
rect 271 44 279 61
rect 246 36 279 44
rect 150 25 165 36
rect 255 25 270 36
rect -270 -36 -255 -25
rect -279 -44 -246 -36
rect -165 -38 -150 -25
rect -60 -36 -45 -25
rect 45 -36 60 -25
rect -279 -61 -271 -44
rect -254 -61 -246 -44
rect -279 -69 -246 -61
rect -69 -44 -36 -36
rect -69 -61 -61 -44
rect -44 -61 -36 -44
rect -69 -69 -36 -61
rect 36 -44 69 -36
rect 150 -38 165 -25
rect 255 -36 270 -25
rect 36 -61 44 -44
rect 61 -61 69 -44
rect 36 -69 69 -61
rect 246 -44 279 -36
rect 246 -61 254 -44
rect 271 -61 279 -44
rect 246 -69 279 -61
<< polycont >>
rect -271 44 -254 61
rect -166 44 -149 61
rect 149 44 166 61
rect 254 44 271 61
rect -271 -61 -254 -44
rect -61 -61 -44 -44
rect 44 -61 61 -44
rect 254 -61 271 -44
<< locali >>
rect -352 95 -304 112
rect 304 95 352 112
rect -352 64 -335 95
rect -271 61 -254 95
rect 254 61 271 95
rect 335 64 352 95
rect -295 44 -271 61
rect -254 44 -230 61
rect -174 44 -166 61
rect -149 44 149 61
rect 166 44 174 61
rect 230 44 254 61
rect 271 44 295 61
rect -295 19 -278 44
rect -295 -44 -278 -19
rect -247 19 -230 44
rect -247 -44 -230 -19
rect -190 24 -173 27
rect -190 -27 -173 -19
rect -142 24 -125 27
rect -142 -27 -125 -19
rect -85 26 -68 27
rect -85 -27 -68 -19
rect -37 19 -20 27
rect -37 -27 -20 -24
rect 20 19 37 27
rect 20 -27 37 -24
rect 68 26 85 27
rect 68 -27 85 -19
rect 125 24 142 27
rect 125 -27 142 -19
rect 173 24 190 27
rect 173 -27 190 -19
rect 230 19 247 44
rect 230 -44 247 -19
rect 278 19 295 44
rect 278 -44 295 -19
rect -295 -61 -271 -44
rect -254 -61 -230 -44
rect -69 -61 -61 -44
rect -44 -61 44 -44
rect 61 -61 69 -44
rect 230 -61 254 -44
rect 271 -61 295 -44
rect -352 -95 -335 -64
rect -271 -95 -254 -61
rect 254 -95 271 -61
rect 335 -95 352 -64
rect -352 -112 -304 -95
rect 304 -112 352 -95
<< viali >>
rect -166 44 -149 61
rect 149 44 166 61
rect -190 19 -173 24
rect -190 7 -173 19
rect -142 19 -125 24
rect -142 7 -125 19
rect -85 19 -68 26
rect -85 9 -68 19
rect -37 -19 -20 -7
rect -37 -24 -20 -19
rect 20 -19 37 -7
rect 20 -24 37 -19
rect 68 19 85 26
rect 68 9 85 19
rect 125 19 142 24
rect 125 7 142 19
rect 173 19 190 24
rect 173 7 190 19
rect -61 -61 -44 -44
rect 44 -61 61 -44
<< metal1 >>
rect -172 61 -143 64
rect 143 61 172 64
rect -172 44 -166 61
rect -149 44 149 61
rect 166 44 174 61
rect 224 44 229 70
rect 255 44 259 70
rect -172 41 -143 44
rect 143 41 172 44
rect -196 24 -167 27
rect -204 -2 -199 24
rect -173 4 -167 24
rect -148 24 -119 27
rect -91 26 -62 29
rect 62 26 91 29
rect -148 4 -142 24
rect -173 -2 -168 4
rect -147 -2 -142 4
rect -116 -2 -111 24
rect -91 9 -85 26
rect -68 10 68 26
rect -68 9 -62 10
rect -91 6 -62 9
rect 62 9 68 10
rect 85 9 91 26
rect 119 24 148 27
rect 62 1 91 9
rect -43 -7 -13 -4
rect -43 -24 -37 -7
rect -20 -24 -13 -7
rect -43 -27 -13 -24
rect -18 -30 -13 -27
rect 13 -7 43 -4
rect 13 -24 20 -7
rect 37 -24 43 -7
rect 13 -27 43 -24
rect 62 -25 68 1
rect 94 -25 97 1
rect 113 -2 116 24
rect 142 4 148 24
rect 167 24 196 27
rect 167 4 173 24
rect 142 -2 147 4
rect 168 -2 173 4
rect 199 -2 204 24
rect 13 -30 18 -27
rect -67 -44 -38 -41
rect 38 -42 67 -41
rect 35 -44 67 -42
rect -69 -61 -61 -44
rect -44 -61 44 -44
rect 61 -61 67 -44
rect -67 -64 -38 -61
rect 38 -64 67 -61
<< via1 >>
rect 229 44 255 70
rect -199 7 -190 24
rect -190 7 -173 24
rect -199 -2 -173 7
rect -142 7 -125 24
rect -125 7 -116 24
rect -142 -2 -116 7
rect -13 -30 13 -4
rect 68 -25 94 1
rect 116 7 125 24
rect 125 7 142 24
rect 116 -2 142 7
rect 173 7 190 24
rect 190 7 199 24
rect 173 -2 199 7
<< metal2 >>
rect -199 58 199 75
rect -199 24 -173 58
rect -230 -2 -199 12
rect -230 -5 -173 -2
rect -142 24 142 36
rect -116 19 116 24
rect 68 1 94 5
rect -142 -44 -116 -2
rect -272 -61 -116 -44
rect -13 -4 13 1
rect -13 -73 13 -30
rect 116 -5 142 -2
rect 173 24 199 58
rect 173 -5 199 -2
rect 229 70 255 75
rect 229 39 255 44
rect 68 -33 94 -25
rect 229 -33 247 39
rect 68 -51 247 -33
rect -13 -90 295 -73
<< properties >>
string FIXED_BBOX -343 -103 343 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
